//
// Conformal-LEC Version 15.10-d003 ( 23-Apr-2015) ( 64 bit executable)
//
module top ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 );
input  n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 ;
output n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 ;

wire  C0 , C1 , 
    RI19a859b8_2755 , 
    RI19a23510_2794 , 
    RI19a22f70_2797 , 
    RI1754a798_67 , 
    RI19a23e70_2789 , 
    RI19ad04a8_2209 , 
    RI1754c610_2 , 
    RI17465568_1242 , 
    RI19a8fd50_2684 , 
    RI1753aa78_586 , 
    RI1749f948_958 , 
    RI19ab7530_2399 , 
    RI17534808_603 , 
    RI173ba970_1846 , 
    RI17403660_1491 , 
    RI173efea8_1586 , 
    RI174741a8_1170 , 
    RI19a9a160_2611 , 
    RI174bfb80_814 , 
    RI19ac9938_2258 , 
    RI1738f1d0_2058 , 
    RI173d7ec0_1703 , 
    RI1744f998_1348 , 
    RI174cedd8_767 , 
    RI19ac4460_2297 , 
    RI1746f630_1193 , 
    RI19a8a2d8_2723 , 
    RI174b8308_838 , 
    RI19abbe50_2368 , 
    RI1738a658_2081 , 
    RI173d3348_1726 , 
    RI1744ae20_1371 , 
    RI1747e270_1121 , 
    RI19aa5560_2527 , 
    RI174cf300_766 , 
    RI19a869a8_2748 , 
    RI17398f50_2010 , 
    RI173e1c40_1655 , 
    RI17459a60_1299 , 
    RI173a7500_1940 , 
    RI1747dbe0_1123 , 
    RI19a93fe0_2654 , 
    RI174ce8b0_768 , 
    RI19ac4280_2298 , 
    RI173988c0_2012 , 
    RI173e15b0_1657 , 
    RI174593d0_1301 , 
    RI1749b118_980 , 
    RI19aa7e28_2510 , 
    RI1752d698_625 , 
    RI19a89e28_2725 , 
    RI173b5df8_1869 , 
    RI173fee30_1513 , 
    RI173c2620_1808 , 
    RI1740fb40_1431 , 
    RI174944d0_1013 , 
    RI19aaac18_2490 , 
    RI17522c70_658 , 
    RI19aa5a88_2525 , 
    RI173af1b0_1902 , 
    RI173f7ea0_1547 , 
    RI1733d8d0_2141 , 
    RI17468d30_1225 , 
    RI19a8d410_2702 , 
    RI174b1a08_870 , 
    RI19abe4c0_2347 , 
    RI17343168_2114 , 
    RI173cc6e8_1759 , 
    RI17415720_1403 , 
    RI1745d570_1281 , 
    RI17473488_1174 , 
    RI19a99698_2616 , 
    RI174be6e0_818 , 
    RI19ac90c8_2262 , 
    RI1738e4b0_2062 , 
    RI173d71a0_1707 , 
    RI1744ec78_1352 , 
    RI174909c0_1031 , 
    RI19aad468_2473 , 
    RI1751cfa0_676 , 
    RI19abe2e0_2348 , 
    RI173ab6a0_1920 , 
    RI173f4390_1565 , 
    RI1750ecc0_720 , 
    RI17497608_998 , 
    RI19aaa510_2493 , 
    RI17488d10_1069 , 
    RI19aa0970_2564 , 
    RI17510bb0_714 , 
    RI19acf680_2215 , 
    RI173a3d38_1957 , 
    RI173eca28_1602 , 
    RI17483130_1097 , 
    RI174a6590_925 , 
    RI19ab2148_2439 , 
    RI17337cf0_2169 , 
    RI173c1270_1814 , 
    RI17409f60_1459 , 
    RI17460d38_1264 , 
    RI17335c20_2179 , 
    RI17495bc8_1006 , 
    RI19aabb90_2484 , 
    RI17525088_651 , 
    RI19aaf448_2459 , 
    RI173b08a8_1895 , 
    RI173f9598_1540 , 
    RI1738bd50_2074 , 
    RI1746a428_1218 , 
    RI19a8bbb0_2713 , 
    RI174b3100_863 , 
    RI19abd188_2358 , 
    RI17344860_2107 , 
    RI173ce128_1751 , 
    RI17445c18_1396 , 
    RI17444ef8_1400 , 
    RI174a3ae8_938 , 
    RI19ab52f8_2415 , 
    RI17335590_2181 , 
    RI173beb10_1826 , 
    RI17407800_1471 , 
    RI17447ce8_1386 , 
    RI17478690_1149 , 
    RI19a97dc0_2627 , 
    RI174c62a0_794 , 
    RI19ac7b38_2272 , 
    RI17393370_2038 , 
    RI173dc060_1683 , 
    RI17453b38_1328 , 
    RI17465bf8_1240 , 
    RI19a8ffa8_2683 , 
    RI174ae8d0_885 , 
    RI19ac0680_2328 , 
    RI17340030_2129 , 
    RI173c95b0_1774 , 
    RI174125e8_1418 , 
    RI17482de8_1098 , 
    RI19aa3aa8_2540 , 
    RI17507628_743 , 
    RI19a84e00_2760 , 
    RI1739dac8_1987 , 
    RI173e6b00_1631 , 
    RI1745e5d8_1276 , 
    RI17508ff0_738 , 
    RI19a82f88_2773 , 
    RI17475210_1165 , 
    RI19a98630_2623 , 
    RI174c1548_809 , 
    RI19ac81c8_2269 , 
    RI17390238_2053 , 
    RI173d8f28_1698 , 
    RI17450a00_1343 , 
    RI17492a90_1021 , 
    RI19aac6d0_2480 , 
    RI17520330_666 , 
    RI19ab3c00_2425 , 
    RI173ad770_1910 , 
    RI173f6460_1555 , 
    RI1752f060_620 , 
    RI174c8be0_786 , 
    RI174809d0_1109 , 
    RI19aa4a98_2532 , 
    RI17501ef8_754 , 
    RI19a85e68_2753 , 
    RI1739b6b0_1998 , 
    RI173e43a0_1643 , 
    RI1745c1c0_1287 , 
    RI1749df08_966 , 
    RI19ab8d90_2389 , 
    RI17531ec8_611 , 
    RI173b8f30_1854 , 
    RI17401c20_1499 , 
    RI173dfeb8_1664 , 
    RI174a5f00_927 , 
    RI19ab4380_2422 , 
    RI174972c0_999 , 
    RI19aaa330_2494 , 
    RI175274a0_644 , 
    RI19aa12d0_2559 , 
    RI173b1fa0_1888 , 
    RI173fac90_1533 , 
    RI1739b9f8_1997 , 
    RI1746bb20_1211 , 
    RI19a8cb28_2706 , 
    RI174b47f8_856 , 
    RI19abddb8_2351 , 
    RI17345f58_2100 , 
    RI173cf820_1744 , 
    RI17447310_1389 , 
    RI174b6580_847 , 
    RI19abcdc8_2360 , 
    RI174a7fd0_917 , 
    RI19ab3138_2431 , 
    RI17339730_2161 , 
    RI173c2cb0_1806 , 
    RI1740b9a0_1451 , 
    RI173895f0_2086 , 
    RI1747c830_1129 , 
    RI19a93068_2661 , 
    RI174cc9c0_774 , 
    RI19ac3290_2305 , 
    RI17397510_2018 , 
    RI173e0200_1663 , 
    RI17458020_1307 , 
    RI1744fce0_1347 , 
    RI17465f40_1239 , 
    RI19a90188_2682 , 
    RI174aec18_884 , 
    RI19ac0860_2327 , 
    RI17340378_2128 , 
    RI173c98f8_1773 , 
    RI17412930_1417 , 
    RI17483478_1096 , 
    RI19aa3c88_2539 , 
    RI17508078_741 , 
    RI19a85058_2759 , 
    RI1739e158_1985 , 
    RI173e7190_1629 , 
    RI1745ec68_1274 , 
    RI174820c8_1102 , 
    RI19aa3238_2544 , 
    RI174737d0_1173 , 
    RI19a998f0_2615 , 
    RI174bec08_817 , 
    RI19ac92a8_2261 , 
    RI1738e7f8_2061 , 
    RI173d74e8_1706 , 
    RI1744efc0_1351 , 
    RI17491050_1029 , 
    RI19aad648_2472 , 
    RI1751d9f0_674 , 
    RI19abf690_2337 , 
    RI173abd30_1918 , 
    RI173f4a20_1563 , 
    RI17512aa0_708 , 
    RI1751ab88_683 , 
    RI19a23678_2793 , 
    RI17480688_1110 , 
    RI19aa48b8_2533 , 
    RI175019d0_755 , 
    RI19a85c10_2754 , 
    RI1739b368_1999 , 
    RI173e4058_1644 , 
    RI1745be78_1288 , 
    RI1749dbc0_967 , 
    RI19ab8b38_2390 , 
    RI175319a0_612 , 
    RI173b8be8_1855 , 
    RI174018d8_1500 , 
    RI173ddaa0_1675 , 
    RI174b8650_837 , 
    RI19acb300_2246 , 
    RI174613c8_1262 , 
    RI19a91e98_2669 , 
    RI174aa0a0_907 , 
    RI19ac21b0_2313 , 
    RI1733b800_2151 , 
    RI173c4d80_1796 , 
    RI1740da70_1441 , 
    RI1747e5b8_1120 , 
    RI19aa5740_2526 , 
    RI174cf828_765 , 
    RI19a86c00_2747 , 
    RI17399298_2009 , 
    RI173e1f88_1654 , 
    RI17459da8_1298 , 
    RI173a7848_1939 , 
    RI1747df28_1122 , 
    RI19a94238_2653 , 
    RI17398c08_2011 , 
    RI173e18f8_1656 , 
    RI17459718_1300 , 
    RI1748cb68_1050 , 
    RI19aafad8_2456 , 
    RI175172d0_694 , 
    RI19a85508_2757 , 
    RI173a7b90_1938 , 
    RI173f0880_1583 , 
    RI174a9d58_908 , 
    RI173f9c28_1538 , 
    RI17487618_1076 , 
    RI19a9fae8_2571 , 
    RI1750e798_721 , 
    RI19ace870_2221 , 
    RI173a2640_1964 , 
    RI173eb330_1609 , 
    RI17475558_1164 , 
    RI174a4b50_933 , 
    RI19ab36d8_2428 , 
    RI173365f8_2176 , 
    RI173bfb78_1821 , 
    RI17408868_1466 , 
    RI17453160_1331 , 
    RI17335f68_2178 , 
    RI17495f10_1005 , 
    RI19aa9688_2500 , 
    RI175255b0_650 , 
    RI19a981f8_2625 , 
    RI173b0bf0_1894 , 
    RI173f98e0_1539 , 
    RI1738e168_2063 , 
    RI1746a770_1217 , 
    RI19a8be08_2712 , 
    RI174b3448_862 , 
    RI19abd2f0_2357 , 
    RI17344ba8_2106 , 
    RI173ce470_1750 , 
    RI17445f60_1395 , 
    RI17340a08_2126 , 
    RI174a0668_954 , 
    RI19ab7f80_2395 , 
    RI17535ca8_599 , 
    RI173bb690_1842 , 
    RI17404380_1487 , 
    RI173f8f08_1542 , 
    RI17474ec8_1166 , 
    RI19a983d8_2624 , 
    RI174c1020_810 , 
    RI19ac7f70_2270 , 
    RI1738fef0_2054 , 
    RI173d8be0_1699 , 
    RI174506b8_1344 , 
    RI173d39d8_1724 , 
    RI17461710_1261 , 
    RI19a920f0_2668 , 
    RI174aa3e8_906 , 
    RI19ac2390_2312 , 
    RI1733bb48_2150 , 
    RI173c50c8_1795 , 
    RI1740ddb8_1440 , 
    RI1747ec48_1118 , 
    RI19aa5dd0_2524 , 
    RI174d0278_763 , 
    RI19a86fc0_2745 , 
    RI17399928_2007 , 
    RI173e2618_1652 , 
    RI1745a438_1296 , 
    RI17509518_737 , 
    RI19a831e0_2772 , 
    RI174758a0_1163 , 
    RI19a98888_2622 , 
    RI174c1f98_807 , 
    RI19ac8330_2268 , 
    RI173908c8_2051 , 
    RI173d95b8_1696 , 
    RI17451090_1341 , 
    RI17492dd8_1020 , 
    RI19aac838_2479 , 
    RI17520858_665 , 
    RI19ab54d8_2414 , 
    RI173adab8_1909 , 
    RI173f67a8_1554 , 
    RI17532918_609 , 
    RI173b1c58_1889 , 
    RI17488680_1071 , 
    RI19aa05b0_2566 , 
    RI17510160_716 , 
    RI19acf1d0_2217 , 
    RI173a36a8_1959 , 
    RI173ec398_1604 , 
    RI1747e900_1119 , 
    RI17337660_2171 , 
    RI173c0be0_1816 , 
    RI174098d0_1461 , 
    RI1745c508_1286 , 
    RI17405730_1481 , 
    RI17493468_1018 , 
    RI19aaca18_2478 , 
    RI175212a8_663 , 
    RI19ab6cc0_2403 , 
    RI173ae148_1907 , 
    RI173f6e38_1552 , 
    RI17332458_2196 , 
    RI17467980_1231 , 
    RI19a8efb8_2690 , 
    RI174b0658_876 , 
    RI19abfa50_2335 , 
    RI17341db8_2120 , 
    RI173cb338_1765 , 
    RI17414370_1409 , 
    RI174b68c8_846 , 
    RI19abaa28_2376 , 
    RI174a8318_916 , 
    RI19ab0e10_2447 , 
    RI17339a78_2160 , 
    RI173c2ff8_1805 , 
    RI1740bce8_1450 , 
    RI173a0228_1975 , 
    RI1747cb78_1128 , 
    RI19a932c0_2660 , 
    RI174ccee8_773 , 
    RI19ac34e8_2304 , 
    RI17397858_2017 , 
    RI173e0548_1662 , 
    RI17458368_1306 , 
    RI173915e8_2047 , 
    RI17468010_1229 , 
    RI19a8f210_2689 , 
    RI174b0ce8_874 , 
    RI19abfc30_2334 , 
    RI17342448_2118 , 
    RI173cb9c8_1763 , 
    RI17414a00_1407 , 
    RI17485200_1087 , 
    RI19aa2e78_2546 , 
    RI1750aee0_732 , 
    RI19a83f78_2766 , 
    RI1739fee0_1976 , 
    RI173e8f18_1620 , 
    RI174609f0_1265 , 
    RI173e9f80_1615 , 
    RI17477628_1154 , 
    RI19a976b8_2630 , 
    RI174c4e00_798 , 
    RI19ac74a8_2275 , 
    RI17392650_2042 , 
    RI173db340_1687 , 
    RI17452e18_1332 , 
    RI17494ea8_1010 , 
    RI19aab410_2487 , 
    RI17523be8_655 , 
    RI19aaa858_2492 , 
    RI173afb88_1899 , 
    RI173f8878_1544 , 
    RI17344518_2108 , 
    RI1751b0b0_682 , 
    RI19a23858_2792 , 
    RI173c39d0_1802 , 
    RI1749a3f8_984 , 
    RI19aa71f8_2515 , 
    RI1752c1f8_629 , 
    RI19a88460_2736 , 
    RI173b50d8_1873 , 
    RI173fe110_1517 , 
    RI173b95c0_1852 , 
    RI1746ec58_1196 , 
    RI19a89888_2727 , 
    RI174b7930_841 , 
    RI19abb5e0_2372 , 
    RI17389c80_2084 , 
    RI173d2970_1729 , 
    RI1744a448_1374 , 
    RI173d2cb8_1728 , 
    RI174a9380_911 , 
    RI19ab1860_2442 , 
    RI1733aae0_2155 , 
    RI173c4060_1800 , 
    RI1740cd50_1445 , 
    RI17411f58_1420 , 
    RI17491398_1028 , 
    RI19aad828_2471 , 
    RI1751df18_673 , 
    RI19ac0a40_2326 , 
    RI173ac078_1917 , 
    RI173f4d68_1562 , 
    RI17516358_697 , 
    RI1733be90_2149 , 
    RI1749baf0_977 , 
    RI19ab9a38_2383 , 
    RI1752e610_622 , 
    RI173b67d0_1866 , 
    RI173ff808_1510 , 
    RI173c9268_1775 , 
    RI17470350_1189 , 
    RI19a9c5f0_2595 , 
    RI174b9460_834 , 
    RI19acb828_2243 , 
    RI1738b378_2077 , 
    RI173d4068_1722 , 
    RI1744bb40_1367 , 
    RI173dd410_1677 , 
    RI1746b148_1214 , 
    RI19a8c498_2709 , 
    RI174b3e20_859 , 
    RI19abd890_2354 , 
    RI17345580_2103 , 
    RI173cee48_1747 , 
    RI17446938_1392 , 
    RI174a9a10_909 , 
    RI19ab1ef0_2440 , 
    RI1733b170_2153 , 
    RI173c46f0_1798 , 
    RI1740d3e0_1443 , 
    RI175361d0_598 , 
    RI1746f978_1192 , 
    RI19a9bfd8_2598 , 
    RI1738a9a0_2080 , 
    RI173d3690_1725 , 
    RI1744b168_1370 , 
    RI174c7c68_789 , 
    RI19ac6080_2284 , 
    RI1746ae00_1215 , 
    RI19a8c240_2710 , 
    RI174b3ad8_860 , 
    RI19abd6b0_2355 , 
    RI17345238_2104 , 
    RI173ceb00_1748 , 
    RI174465f0_1393 , 
    RI17488338_1072 , 
    RI19aa0358_2567 , 
    RI1750fc38_717 , 
    RI19acef78_2218 , 
    RI173a3360_1960 , 
    RI173ec050_1605 , 
    RI1747c4e8_1130 , 
    RI173a2cd0_1962 , 
    RI174793b0_1145 , 
    RI19a96038_2640 , 
    RI174c7740_790 , 
    RI19ac5e28_2285 , 
    RI17394090_2034 , 
    RI173dcd80_1679 , 
    RI17454858_1324 , 
    RI174968e8_1002 , 
    RI19aa9d90_2497 , 
    RI17526528_647 , 
    RI19a9cc08_2592 , 
    RI173b15c8_1891 , 
    RI173fa2b8_1536 , 
    RI17394db0_2030 , 
    RI17539830_589 , 
    RI17539218_590 , 
    RI175385e8_592 , 
    RI17537fd0_593 , 
    RI175379b8_594 , 
    RI17536770_597 , 
    RI17539e48_588 , 
    RI174844e0_1091 , 
    RI19aa2248_2551 , 
    RI17509a40_736 , 
    RI19a83438_2771 , 
    RI1739f1c0_1980 , 
    RI173e81f8_1624 , 
    RI1745fcd0_1269 , 
    RI174a1a18_948 , 
    RI19ab63d8_2407 , 
    RI173334c0_2191 , 
    RI173bca40_1836 , 
    RI174046c8_1486 , 
    RI174d1208_760 , 
    RI19a876c8_2742 , 
    RI174709e0_1187 , 
    RI19a9ca28_2593 , 
    RI174b9eb0_832 , 
    RI19acbc60_2241 , 
    RI1738ba08_2075 , 
    RI173d46f8_1720 , 
    RI1744c1d0_1365 , 
    RI1748df18_1044 , 
    RI19ab0870_2450 , 
    RI175191c0_688 , 
    RI19ac1d78_2315 , 
    RI173a8f40_1932 , 
    RI173f1c30_1577 , 
    RI174b75e8_842 , 
    RI173ad0e0_1912 , 
    RI17483b08_1094 , 
    RI19aa1d20_2554 , 
    RI17508ac8_739 , 
    RI19a82d30_2774 , 
    RI1739e7e8_1983 , 
    RI173e7820_1627 , 
    RI1745f2f8_1272 , 
    RI174a1040_951 , 
    RI19ab5d48_2410 , 
    RI17332ae8_2194 , 
    RI173bc068_1839 , 
    RI17404d58_1484 , 
    RI173fda80_1519 , 
    RI174a1388_950 , 
    RI19ab5f28_2409 , 
    RI174672f0_1233 , 
    RI19a8e8b0_2693 , 
    RI174affc8_878 , 
    RI19abf4b0_2338 , 
    RI17341728_2122 , 
    RI173caca8_1767 , 
    RI17413ce0_1411 , 
    RI174b1d50_869 , 
    RI19abe6a0_2346 , 
    RI174a3458_940 , 
    RI19ab4dd0_2417 , 
    RI17334f00_2183 , 
    RI173be480_1828 , 
    RI17407170_1473 , 
    RI174146b8_1408 , 
    RI17478000_1151 , 
    RI19a97820_2629 , 
    RI174c5850_796 , 
    RI19ac7700_2274 , 
    RI17392ce0_2040 , 
    RI173db9d0_1685 , 
    RI174534a8_1330 , 
    RI1738ca70_2070 , 
    RI17463150_1253 , 
    RI19a90cc8_2677 , 
    RI174abe28_898 , 
    RI19ac1148_2322 , 
    RI1733d588_2142 , 
    RI173c6b08_1787 , 
    RI1740f7f8_1432 , 
    RI1748be48_1054 , 
    RI19a9e030_2584 , 
    RI1747d898_1124 , 
    RI19a93d88_2655 , 
    RI174ce388_769 , 
    RI19ac40a0_2299 , 
    RI17398578_2013 , 
    RI173e1268_1658 , 
    RI17459088_1302 , 
    RI1749add0_981 , 
    RI19aa7c48_2511 , 
    RI1752d170_626 , 
    RI19a88e38_2732 , 
    RI173b5ab0_1870 , 
    RI173feae8_1514 , 
    RI173c0208_1819 , 
    RI1752a308_635 , 
    RI19a95048_2647 , 
    RI1748a750_1061 , 
    RI19a9f548_2574 , 
    RI17513a18_705 , 
    RI19ace168_2224 , 
    RI173a5778_1949 , 
    RI173ee468_1594 , 
    RI17493120_1019 , 
    RI173bee58_1825 , 
    RI17495880_1007 , 
    RI19aab938_2485 , 
    RI17524b60_652 , 
    RI19aadb70_2470 , 
    RI173b0560_1896 , 
    RI173f9250_1541 , 
    RI17389938_2085 , 
    RI17469d98_1220 , 
    RI19a8dfc8_2697 , 
    RI174b2a70_865 , 
    RI19abeda8_2342 , 
    RI173441d0_2109 , 
    RI173cd750_1754 , 
    RI17445588_1398 , 
    RI173a3018_1961 , 
    RI174796f8_1144 , 
    RI19a96290_2639 , 
    RI173943d8_2033 , 
    RI173dd0c8_1678 , 
    RI17454ba0_1323 , 
    RI17496c30_1001 , 
    RI19aa9f70_2496 , 
    RI17526a50_646 , 
    RI19a9e6c0_2581 , 
    RI173b1910_1890 , 
    RI173fa600_1535 , 
    RI173971c8_2019 , 
    RI173f53f8_1560 , 
    RI174a0320_955 , 
    RI19ab7da0_2396 , 
    RI17535780_600 , 
    RI173bb348_1843 , 
    RI17404038_1488 , 
    RI173f6af0_1553 , 
    RI173e4a30_1641 , 
    RI1748ffe8_1034 , 
    RI19aaf628_2458 , 
    RI1751c028_679 , 
    RI19a23150_2796 , 
    RI173aacc8_1923 , 
    RI173f39b8_1568 , 
    RI17502420_753 , 
    RI17464848_1246 , 
    RI19a919e8_2671 , 
    RI174ad520_891 , 
    RI19ac1b98_2316 , 
    RI1733ec80_2135 , 
    RI173c8200_1780 , 
    RI17410ef0_1425 , 
    RI1733c1d8_2148 , 
    RI1749be38_976 , 
    RI19ab9c18_2382 , 
    RI1752eb38_621 , 
    RI173b6b18_1865 , 
    RI173ffb50_1509 , 
    RI173cb680_1764 , 
    RI17470698_1188 , 
    RI19a9c848_2594 , 
    RI174b9988_833 , 
    RI19acba08_2242 , 
    RI1738b6c0_2076 , 
    RI173d43b0_1721 , 
    RI1744be88_1366 , 
    RI173dd758_1676 , 
    RI1746b490_1213 , 
    RI19a8c6f0_2708 , 
    RI174b4168_858 , 
    RI19abd9f8_2353 , 
    RI173458c8_2102 , 
    RI173cf190_1746 , 
    RI17446c80_1391 , 
    RI174889c8_1070 , 
    RI19aa0790_2565 , 
    RI17510688_715 , 
    RI19acf428_2216 , 
    RI173a39f0_1958 , 
    RI173ec6e0_1603 , 
    RI17480d18_1108 , 
    RI174a2dc8_942 , 
    RI173ad428_1911 , 
    RI17483e50_1093 , 
    RI19aa1f00_2553 , 
    RI1739eb30_1982 , 
    RI173e7b68_1626 , 
    RI1745f640_1271 , 
    RI17332e30_2193 , 
    RI173bc3b0_1838 , 
    RI174050a0_1483 , 
    RI173ffe98_1508 , 
    RI17400f00_1503 , 
    RI1748ec38_1040 , 
    RI19aae7a0_2465 , 
    RI1751a138_685 , 
    RI19a23330_2795 , 
    RI173a9918_1929 , 
    RI173f2608_1574 , 
    RI174be1b8_819 , 
    RI174118c8_1422 , 
    RI1749f600_959 , 
    RI19ab73c8_2400 , 
    RI175342e0_604 , 
    RI173ba628_1847 , 
    RI17403318_1492 , 
    RI173eda90_1597 , 
    RI17473e60_1171 , 
    RI19a99f80_2612 , 
    RI174bf658_815 , 
    RI19ac96e0_2259 , 
    RI1738ee88_2059 , 
    RI173d7b78_1704 , 
    RI1744f650_1349 , 
    RI1738cdb8_2069 , 
    RI174637e0_1251 , 
    RI19a90f20_2676 , 
    RI174ac4b8_896 , 
    RI19ac12b0_2321 , 
    RI1733dc18_2140 , 
    RI173c7198_1785 , 
    RI1740fe88_1430 , 
    RI173e5750_1637 , 
    RI17472df8_1176 , 
    RI19a9bd80_2599 , 
    RI174bd768_821 , 
    RI19acb120_2247 , 
    RI1738de20_2064 , 
    RI173d6b10_1709 , 
    RI1744e5e8_1354 , 
    RI17490678_1032 , 
    RI19aad300_2474 , 
    RI1751ca78_677 , 
    RI19abcfa8_2359 , 
    RI173ab358_1921 , 
    RI173f4048_1566 , 
    RI1750b408_731 , 
    RI173b2630_1886 , 
    RI1748ade0_1059 , 
    RI19a9d400_2589 , 
    RI17514468_703 , 
    RI19acc200_2238 , 
    RI173a5e08_1947 , 
    RI173eeaf8_1592 , 
    RI17497950_997 , 
    RI174a8660_915 , 
    RI19ab0ff0_2446 , 
    RI17339dc0_2159 , 
    RI173c3340_1804 , 
    RI1740c030_1449 , 
    RI173b6e60_1864 , 
    RI173bf1a0_1824 , 
    RI174a4808_934 , 
    RI19ab34f8_2429 , 
    RI173362b0_2177 , 
    RI173bf830_1822 , 
    RI17408520_1467 , 
    RI17450d48_1342 , 
    RI1744b7f8_1368 , 
    RI17461a58_1260 , 
    RI19a922d0_2667 , 
    RI174aa730_905 , 
    RI19ac25e8_2311 , 
    RI173c5410_1794 , 
    RI1740e100_1439 , 
    RI1747ef90_1117 , 
    RI19aa5fb0_2523 , 
    RI174d07a0_762 , 
    RI19a87218_2744 , 
    RI17399c70_2006 , 
    RI173e2960_1651 , 
    RI1745a780_1295 , 
    RI173acd98_1913 , 
    RI174837c0_1095 , 
    RI19aa3ee0_2538 , 
    RI175085a0_740 , 
    RI19a852b0_2758 , 
    RI1739e4a0_1984 , 
    RI173e74d8_1628 , 
    RI1745efb0_1273 , 
    RI174a0cf8_952 , 
    RI19ab5a00_2411 , 
    RI173327a0_2195 , 
    RI173bbd20_1840 , 
    RI17404a10_1485 , 
    RI173fb668_1530 , 
    RI17400870_1505 , 
    RI17462ac0_1255 , 
    RI19a92e10_2662 , 
    RI174ab798_900 , 
    RI19ac30b0_2306 , 
    RI1733cef8_2144 , 
    RI173c6478_1789 , 
    RI1740f168_1434 , 
    RI17411238_1424 , 
    RI1749ef70_961 , 
    RI19ab7008_2402 , 
    RI17533890_606 , 
    RI173b9f98_1849 , 
    RI17402c88_1494 , 
    RI173e9260_1619 , 
    RI1746aab8_1216 , 
    RI19a8bfe8_2711 , 
    RI174b3790_861 , 
    RI19abd4d0_2356 , 
    RI17344ef0_2105 , 
    RI173ce7b8_1749 , 
    RI174462a8_1394 , 
    RI17487ff0_1073 , 
    RI19aa0100_2568 , 
    RI1750f710_718 , 
    RI19aced20_2219 , 
    RI173ebd08_1606 , 
    RI1747a0d0_1141 , 
    RI17479068_1146 , 
    RI19a95de0_2641 , 
    RI174c7218_791 , 
    RI19ac5bd0_2286 , 
    RI17393d48_2035 , 
    RI173dca38_1680 , 
    RI17454510_1325 , 
    RI174965a0_1003 , 
    RI19aa9bb0_2498 , 
    RI17526000_648 , 
    RI19a9b420_2603 , 
    RI173b1280_1892 , 
    RI173f9f70_1537 , 
    RI17392998_2041 , 
    RI17482758_1100 , 
    RI19aa3580_2542 , 
    RI17506bd8_745 , 
    RI19a84950_2762 , 
    RI1739d438_1989 , 
    RI173e6470_1633 , 
    RI1745df48_1278 , 
    RI1749fc90_957 , 
    RI19ab7878_2398 , 
    RI17534d30_602 , 
    RI173bacb8_1845 , 
    RI174039a8_1490 , 
    RI173f22c0_1575 , 
    RI174ae240_887 , 
    RI19ac04a0_2329 , 
    RI1733f9a0_2131 , 
    RI173c8f20_1776 , 
    RI17411c10_1421 , 
    RI1749b7a8_978 , 
    RI19ab98d0_2384 , 
    RI1752e0e8_623 , 
    RI173b6488_1867 , 
    RI173ff4c0_1511 , 
    RI173c6e50_1786 , 
    RI17470008_1190 , 
    RI19a9c398_2596 , 
    RI174b8f38_835 , 
    RI19acb648_2244 , 
    RI1738b030_2078 , 
    RI173d3d20_1723 , 
    RI174d0cc8_761 , 
    RI19a87470_2743 , 
    RI1748dbd0_1045 , 
    RI19ab0528_2451 , 
    RI17518c98_689 , 
    RI19ab3a20_2426 , 
    RI173a8bf8_1933 , 
    RI173f18e8_1578 , 
    RI174b51d0_853 , 
    RI174a3110_941 , 
    RI19ab4bf0_2418 , 
    RI17334bb8_2184 , 
    RI173be138_1829 , 
    RI17406e28_1474 , 
    RI174122a0_1419 , 
    RI1738c728_2071 , 
    RI17462e08_1254 , 
    RI19a90a70_2678 , 
    RI174abae0_899 , 
    RI19ac0f68_2323 , 
    RI1733d240_2143 , 
    RI173c67c0_1788 , 
    RI1740f4b0_1433 , 
    RI17480340_1111 , 
    RI19aa46d8_2534 , 
    RI175014a8_756 , 
    RI1739b020_2000 , 
    RI173e3d10_1645 , 
    RI1745bb30_1289 , 
    RI173e50c0_1639 , 
    RI17472768_1178 , 
    RI19a9b8d0_2601 , 
    RI174bcd18_823 , 
    RI19acadd8_2249 , 
    RI1738d790_2066 , 
    RI173d6480_1711 , 
    RI1744df58_1356 , 
    RI17529de0_636 , 
    RI19a93518_2659 , 
    RI1748a408_1062 , 
    RI19a9f368_2575 , 
    RI175134f0_706 , 
    RI19acdf10_2225 , 
    RI173a5430_1950 , 
    RI173ee120_1595 , 
    RI17490d08_1030 , 
    RI174a7c88_918 , 
    RI19ab2f58_2432 , 
    RI173393e8_2162 , 
    RI173c2968_1807 , 
    RI1740b658_1452 , 
    RI17332110_2197 , 
    RI174951f0_1009 , 
    RI19aab5f0_2486 , 
    RI17524110_654 , 
    RI19aac388_2481 , 
    RI173afed0_1898 , 
    RI173f8bc0_1543 , 
    RI17346930_2097 , 
    RI17469a50_1221 , 
    RI19a8dd70_2698 , 
    RI174b2728_866 , 
    RI19abebc8_2343 , 
    RI17343e88_2110 , 
    RI173cd408_1755 , 
    RI17445240_1399 , 
    RI174a4178_936 , 
    RI19ab5820_2412 , 
    RI17407e90_1469 , 
    RI1744c518_1364 , 
    RI17478d20_1147 , 
    RI19a95b88_2642 , 
    RI174c6cf0_792 , 
    RI19ac5978_2287 , 
    RI17393a00_2036 , 
    RI173dc6f0_1681 , 
    RI174541c8_1326 , 
    RI173f50b0_1561 , 
    RI17482aa0_1099 , 
    RI19aa38c8_2541 , 
    RI17507100_744 , 
    RI19a84ba8_2761 , 
    RI1739d780_1988 , 
    RI173e67b8_1632 , 
    RI1745e290_1277 , 
    RI1749ffd8_956 , 
    RI19ab7a58_2397 , 
    RI17535258_601 , 
    RI173bb000_1844 , 
    RI17403cf0_1489 , 
    RI173f46d8_1564 , 
    RI173e22d0_1653 , 
    RI1748fca0_1035 , 
    RI19aaf268_2460 , 
    RI1751bb00_680 , 
    RI19a23c18_2790 , 
    RI173aa980_1924 , 
    RI173f3670_1569 , 
    RI174cfd50_764 , 
    RI17464500_1247 , 
    RI19a91808_2672 , 
    RI174ad1d8_892 , 
    RI19ac1a30_2317 , 
    RI1733e938_2136 , 
    RI173c7eb8_1781 , 
    RI17410ba8_1426 , 
    RI174a09b0_953 , 
    RI1747d550_1125 , 
    RI19a93ba8_2656 , 
    RI174cde60_770 , 
    RI19ac3d58_2300 , 
    RI17398230_2014 , 
    RI173e0f20_1659 , 
    RI17458d40_1303 , 
    RI1749aa88_982 , 
    RI19aa7a68_2512 , 
    RI1752cc48_627 , 
    RI19a88be0_2733 , 
    RI173b5768_1871 , 
    RI173fe7a0_1515 , 
    RI173bddf0_1830 , 
    RI17400bb8_1504 , 
    RI1748e260_1043 , 
    RI19ab0a50_2449 , 
    RI175196e8_687 , 
    RI19ad0238_2210 , 
    RI173a9288_1931 , 
    RI173f1f78_1576 , 
    RI174ba3d8_831 , 
    RI17411580_1423 , 
    RI1749f2b8_960 , 
    RI19ab71e8_2401 , 
    RI17533db8_605 , 
    RI173ba2e0_1848 , 
    RI17402fd0_1493 , 
    RI173eb678_1608 , 
    RI17473b18_1172 , 
    RI19a99d28_2613 , 
    RI174bf130_816 , 
    RI19ac9500_2260 , 
    RI1738eb40_2060 , 
    RI173d7830_1705 , 
    RI1744f308_1350 , 
    RI173e5408_1638 , 
    RI17472ab0_1177 , 
    RI19a9bb28_2600 , 
    RI174bd240_822 , 
    RI19acaf40_2248 , 
    RI1738dad8_2065 , 
    RI173d67c8_1710 , 
    RI1744e2a0_1355 , 
    RI17490330_1033 , 
    RI19aaf790_2457 , 
    RI1751c550_678 , 
    RI19a83b40_2768 , 
    RI173ab010_1922 , 
    RI173f3d00_1567 , 
    RI17507b50_742 , 
    RI173b0218_1897 , 
    RI1748aa98_1060 , 
    RI19a9f728_2573 , 
    RI17513f40_704 , 
    RI19ace3c0_2223 , 
    RI173a5ac0_1948 , 
    RI173ee7b0_1593 , 
    RI17495538_1008 , 
    RI174a44c0_935 , 
    RI19ab3318_2430 , 
    RI173bf4e8_1823 , 
    RI174081d8_1468 , 
    RI1744e930_1353 , 
    RI1744b4b0_1369 , 
    RI1733f310_2133 , 
    RI1746f2e8_1194 , 
    RI19a8a080_2724 , 
    RI174b7fc0_839 , 
    RI19abbc70_2369 , 
    RI1738a310_2082 , 
    RI173d3000_1727 , 
    RI1744aad8_1372 , 
    RI1748c820_1051 , 
    RI19a9e468_2582 , 
    RI17516da8_695 , 
    RI19acd100_2231 , 
    RI173f0538_1584 , 
    RI174a7940_919 , 
    RI173a6e70_1942 , 
    RI17486f88_1078 , 
    RI19aa19d8_2555 , 
    RI1750dd48_723 , 
    RI19a82b50_2775 , 
    RI173a1fb0_1966 , 
    RI173eaca0_1611 , 
    RI17470d28_1186 , 
    RI17465220_1243 , 
    RI19a8faf8_2685 , 
    RI174a6248_926 , 
    RI19ab4560_2421 , 
    RI173379a8_2170 , 
    RI173c0f28_1815 , 
    RI17409c18_1460 , 
    RI1745e920_1275 , 
    RI173358d8_2180 , 
    RI17474838_1168 , 
    RI19a9a610_2609 , 
    RI174c05d0_812 , 
    RI19ac9de8_2256 , 
    RI1738f860_2056 , 
    RI173d8550_1701 , 
    RI17450028_1346 , 
    RI17492748_1022 , 
    RI19aac040_2482 , 
    RI1751fe08_667 , 
    RI19ab2508_2437 , 
    RI173f6118_1556 , 
    RI1752b7a8_631 , 
    RI174a5870_929 , 
    RI19ab3de0_2424 , 
    RI17336fd0_2173 , 
    RI173c0550_1818 , 
    RI17409240_1463 , 
    RI17457cd8_1308 , 
    RI174a5bb8_928 , 
    RI19ab4038_2423 , 
    RI17496f78_1000 , 
    RI19aaa150_2495 , 
    RI17526f78_645 , 
    RI19a9fcc8_2570 , 
    RI173fa948_1534 , 
    RI173995e0_2008 , 
    RI1746b7d8_1212 , 
    RI19a8c948_2707 , 
    RI174b44b0_857 , 
    RI19abdbd8_2352 , 
    RI17345c10_2101 , 
    RI173cf4d8_1745 , 
    RI17446fc8_1390 , 
    RI174b6238_848 , 
    RI19abcbe8_2361 , 
    RI1747c1a0_1131 , 
    RI19a95930_2643 , 
    RI174cbf70_776 , 
    RI19ac5720_2288 , 
    RI17396e80_2020 , 
    RI173dfb70_1665 , 
    RI17457648_1310 , 
    RI17390f58_2049 , 
    RI17467638_1232 , 
    RI19a8ed60_2691 , 
    RI174b0310_877 , 
    RI19abf870_2336 , 
    RI17341a70_2121 , 
    RI173caff0_1766 , 
    RI17414028_1410 , 
    RI17484b70_1089 , 
    RI19aa27e8_2549 , 
    RI1750a490_734 , 
    RI19a838e8_2769 , 
    RI1739f850_1978 , 
    RI173e8888_1622 , 
    RI17460360_1267 , 
    RI17481d80_1103 , 
    RI19aa3058_2545 , 
    RI1751a660_684 , 
    RI1749d878_968 , 
    RI19ab8958_2391 , 
    RI17531478_613 , 
    RI173b88a0_1856 , 
    RI17401590_1501 , 
    RI173db688_1686 , 
    RI17499a20_987 , 
    RI19aa6d48_2517 , 
    RI1752b280_632 , 
    RI19a88028_2738 , 
    RI173b4700_1876 , 
    RI173fd738_1520 , 
    RI173b4a48_1875 , 
    RI1746e280_1199 , 
    RI19a894c8_2729 , 
    RI174b6f58_844 , 
    RI19abaf50_2374 , 
    RI173599e0_2088 , 
    RI173d1f98_1732 , 
    RI17449a70_1377 , 
    RI174872d0_1077 , 
    RI19a9f908_2572 , 
    RI1750e270_722 , 
    RI19ace618_2222 , 
    RI173a22f8_1965 , 
    RI173eafe8_1610 , 
    RI17473140_1175 , 
    RI173406c0_2127 , 
    RI17474b80_1167 , 
    RI19a9a868_2608 , 
    RI174c0af8_811 , 
    RI19aca040_2255 , 
    RI1738fba8_2055 , 
    RI173d8898_1700 , 
    RI17450370_1345 , 
    RI17337318_2172 , 
    RI173c0898_1817 , 
    RI17409588_1462 , 
    RI1745a0f0_1297 , 
    RI174053e8_1482 , 
    RI173912a0_2048 , 
    RI17484eb8_1088 , 
    RI19aa2c20_2547 , 
    RI1750a9b8_733 , 
    RI19a83d20_2767 , 
    RI1739fb98_1977 , 
    RI173e8bd0_1621 , 
    RI174606a8_1266 , 
    RI173e9c38_1616 , 
    RI174772e0_1155 , 
    RI19a97460_2631 , 
    RI174c48d8_799 , 
    RI19ac7250_2276 , 
    RI17392308_2043 , 
    RI173daff8_1688 , 
    RI17452ad0_1333 , 
    RI17494b60_1011 , 
    RI19aab0c8_2488 , 
    RI175236c0_656 , 
    RI19aa8f80_2503 , 
    RI173af840_1900 , 
    RI173f8530_1545 , 
    RI17342100_2119 , 
    RI173c3688_1803 , 
    RI1749a0b0_985 , 
    RI19aa7090_2516 , 
    RI1752bcd0_630 , 
    RI19a88208_2737 , 
    RI173b4d90_1874 , 
    RI173fddc8_1518 , 
    RI173b71a8_1863 , 
    RI1746e5c8_1198 , 
    RI19a89720_2728 , 
    RI174b72a0_843 , 
    RI19abb298_2373 , 
    RI173892a8_2087 , 
    RI173d22e0_1731 , 
    RI17449db8_1376 , 
    RI174a9038_912 , 
    RI19ab16f8_2443 , 
    RI1733a798_2156 , 
    RI173c3d18_1801 , 
    RI1740ca08_1446 , 
    RI173fb320_1531 , 
    RI173413e0_2123 , 
    RI17475be8_1162 , 
    RI19a98ae0_2621 , 
    RI174c24c0_806 , 
    RI19ac8510_2267 , 
    RI17390c10_2050 , 
    RI173d9900_1695 , 
    RI174513d8_1340 , 
    RI174620e8_1258 , 
    RI19a92708_2665 , 
    RI174aadc0_903 , 
    RI19ac2a98_2309 , 
    RI1733c520_2147 , 
    RI173c5aa0_1792 , 
    RI1740e790_1437 , 
    RI1747f620_1115 , 
    RI19aa62f8_2521 , 
    RI1739a300_2004 , 
    RI173e2ff0_1649 , 
    RI1745ae10_1293 , 
    RI17491a28_1026 , 
    RI19aadfa8_2468 , 
    RI1751e968_671 , 
    RI19ac36c8_2303 , 
    RI173ac708_1915 , 
    RI1751d4c8_675 , 
    RI17461da0_1259 , 
    RI19a92528_2666 , 
    RI174aaa78_904 , 
    RI19ac2840_2310 , 
    RI173c5758_1793 , 
    RI1740e448_1438 , 
    RI1747f2d8_1116 , 
    RI19aa6190_2522 , 
    RI17399fb8_2005 , 
    RI173e2ca8_1650 , 
    RI1745aac8_1294 , 
    RI1748d540_1047 , 
    RI19ab01e0_2453 , 
    RI17518248_691 , 
    RI19a94df0_2648 , 
    RI173a8568_1935 , 
    RI173f1258_1580 , 
    RI174b09a0_875 , 
    RI17336940_2175 , 
    RI17476278_1160 , 
    RI19a98f90_2619 , 
    RI174c2f10_804 , 
    RI19ac89c0_2265 , 
    RI173d9f90_1693 , 
    RI17451a68_1338 , 
    RI17493af8_1016 , 
    RI19aacdd8_2476 , 
    RI17521cf8_661 , 
    RI19ab9df8_2381 , 
    RI173ae7d8_1905 , 
    RI173f74c8_1550 , 
    RI17336c88_2174 , 
    RI173b2978_1885 , 
    RI17489058_1068 , 
    RI19a9e8a0_2580 , 
    RI175110d8_713 , 
    RI19acd358_2230 , 
    RI173a4080_1956 , 
    RI173ecd70_1601 , 
    RI17485548_1086 , 
    RI174a68d8_924 , 
    RI19ab2328_2438 , 
    RI17338038_2168 , 
    RI173c15b8_1813 , 
    RI1740a2a8_1458 , 
    RI17477970_1153 , 
    RI17406108_1478 , 
    RI17493e40_1015 , 
    RI19aad120_2475 , 
    RI17522220_660 , 
    RI19abba90_2370 , 
    RI173aeb20_1904 , 
    RI173f7810_1549 , 
    RI173390a0_2163 , 
    RI174686a0_1227 , 
    RI19a8cd80_2705 , 
    RI174b1378_872 , 
    RI19abdf98_2350 , 
    RI17342ad8_2116 , 
    RI173cc058_1761 , 
    RI17415090_1405 , 
    RI174a8cf0_913 , 
    RI19ab1518_2444 , 
    RI1733a450_2157 , 
    RI1740c6c0_1447 , 
    RI173e46e8_1642 , 
    RI17391fc0_2044 , 
    RI174689e8_1226 , 
    RI19a8cfd8_2704 , 
    RI174b16c0_871 , 
    RI19abe100_2349 , 
    RI17342e20_2115 , 
    RI173cc3a0_1760 , 
    RI174153d8_1404 , 
    RI17485f20_1083 , 
    RI19aa0f10_2561 , 
    RI1750c380_728 , 
    RI19acfd88_2212 , 
    RI173a0f48_1971 , 
    RI174658b0_1241 , 
    RI173ea958_1612 , 
    RI174816f0_1105 , 
    RI19aa5218_2529 , 
    RI17503398_750 , 
    RI19a864f8_2750 , 
    RI1739c3d0_1994 , 
    RI1745cee0_1283 , 
    RI1749ec28_962 , 
    RI19ab9498_2386 , 
    RI17533368_607 , 
    RI173b9c50_1850 , 
    RI17402940_1495 , 
    RI173e6e48_1630 , 
    RI173c43a8_1799 , 
    RI1749b460_979 , 
    RI19ab96f0_2385 , 
    RI1752dbc0_624 , 
    RI173b6140_1868 , 
    RI173ff178_1512 , 
    RI173c4a38_1797 , 
    RI1746fcc0_1191 , 
    RI19a9c1b8_2597 , 
    RI174b8a10_836 , 
    RI19acb4e0_2245 , 
    RI1738ace8_2079 , 
    RI1744a100_1375 , 
    RI17466918_1236 , 
    RI19a8e220_2696 , 
    RI17462430_1257 , 
    RI19a92960_2664 , 
    RI174ab108_902 , 
    RI19ac2cf0_2308 , 
    RI1733c868_2146 , 
    RI173c5de8_1791 , 
    RI1740ead8_1436 , 
    RI1747f968_1114 , 
    RI19aa6640_2520 , 
    RI17500530_759 , 
    RI19a87920_2741 , 
    RI1739a648_2003 , 
    RI173e3338_1648 , 
    RI1745b158_1292 , 
    RI174744f0_1169 , 
    RI19a9a3b8_2610 , 
    RI174c00a8_813 , 
    RI19ac9b90_2257 , 
    RI1738f518_2057 , 
    RI173d8208_1702 , 
    RI17491d70_1025 , 
    RI19aae110_2467 , 
    RI1751ee90_670 , 
    RI19ac4f28_2292 , 
    RI173aca50_1914 , 
    RI173f5740_1559 , 
    RI17520d80_664 , 
    RI174989b8_992 , 
    RI19aa8bc0_2505 , 
    RI1748a0c0_1063 , 
    RI19a9f188_2576 , 
    RI17512fc8_707 , 
    RI19acdcb8_2226 , 
    RI173a50e8_1951 , 
    RI173eddd8_1596 , 
    RI1748e8f0_1041 , 
    RI174a75f8_920 , 
    RI19ab2d78_2433 , 
    RI17338d58_2164 , 
    RI173c22d8_1809 , 
    RI1740afc8_1454 , 
    RI17512578_709 , 
    RI17406450_1477 , 
    RI17494188_1014 , 
    RI19aaaa38_2491 , 
    RI17522748_659 , 
    RI19aa4318_2536 , 
    RI173aee68_1903 , 
    RI173f7b58_1548 , 
    RI1733b4b8_2152 , 
    RI17466c60_1235 , 
    RI19a8e478_2695 , 
    RI174af938_880 , 
    RI19abf0f0_2340 , 
    RI17341098_2124 , 
    RI173ca618_1769 , 
    RI17413650_1413 , 
    RI17484198_1092 , 
    RI19aa2068_2552 , 
    RI1739ee78_1981 , 
    RI173e7eb0_1625 , 
    RI1745f988_1270 , 
    RI174789d8_1148 , 
    RI19a98018_2626 , 
    RI174c67c8_793 , 
    RI19ac7d90_2271 , 
    RI173936b8_2037 , 
    RI173dc3a8_1682 , 
    RI17453e80_1327 , 
    RI17503de8_748 , 
    RI19a841d0_2765 , 
    RI1739ca60_1992 , 
    RI173e5a98_1636 , 
    RI174a6f68_922 , 
    RI19ab29b8_2435 , 
    RI17498670_993 , 
    RI19aa8878_2506 , 
    RI17529390_638 , 
    RI19a90368_2681 , 
    RI173b3350_1882 , 
    RI173fc388_1526 , 
    RI173a71b8_1941 , 
    RI1746ced0_1205 , 
    RI19a8af08_2718 , 
    RI174b5ba8_850 , 
    RI19abc8a0_2363 , 
    RI17347308_2094 , 
    RI173d0bd0_1738 , 
    RI174486c0_1383 , 
    RI17466fa8_1234 , 
    RI19a8e6d0_2694 , 
    RI174afc80_879 , 
    RI19abf2d0_2339 , 
    RI173ca960_1768 , 
    RI17413998_1412 , 
    RI174920b8_1024 , 
    RI19aae458_2466 , 
    RI1751f3b8_669 , 
    RI19ac6878_2281 , 
    RI173f5a88_1558 , 
    RI17524638_653 , 
    RI1740a5f0_1457 , 
    RI17498328_994 , 
    RI19aa8530_2507 , 
    RI17528e68_639 , 
    RI19a8eb08_2692 , 
    RI173b3008_1883 , 
    RI173fc040_1527 , 
    RI173a4da0_1952 , 
    RI1746cb88_1206 , 
    RI19a8acb0_2719 , 
    RI174b5860_851 , 
    RI19abc6c0_2364 , 
    RI17346fc0_2095 , 
    RI173d0888_1739 , 
    RI17448378_1384 , 
    RI174996d8_988 , 
    RI19aa6b68_2518 , 
    RI1752ad58_633 , 
    RI19a87dd0_2739 , 
    RI173b43b8_1877 , 
    RI173fd3f0_1521 , 
    RI1746df38_1200 , 
    RI19a89270_2730 , 
    RI174b6c10_845 , 
    RI19abad70_2375 , 
    RI17359698_2089 , 
    RI173d1c50_1733 , 
    RI17449728_1378 , 
    RI1747a418_1140 , 
    RI19a96bf0_2635 , 
    RI174c9108_785 , 
    RI19ac69e0_2280 , 
    RI173950f8_2029 , 
    RI173ddde8_1674 , 
    RI174558c0_1319 , 
    RI174665d0_1237 , 
    RI19a90818_2679 , 
    RI174af2a8_882 , 
    RI19ac0d88_2324 , 
    RI173c9f88_1771 , 
    RI17412fc0_1415 , 
    RI1749c4c8_974 , 
    RI19aba050_2380 , 
    RI1752f588_619 , 
    RI173b74f0_1862 , 
    RI174001e0_1507 , 
    RI173cdde0_1752 , 
    RI173964a8_2023 , 
    RI173eee40_1591 , 
    RI1733fce8_2130 , 
    RI174adef8_888 , 
    RI19ac0338_2330 , 
    RI1733f658_2132 , 
    RI173c8bd8_1777 , 
    RI17454ee8_1322 , 
    RI174a4e98_932 , 
    RI19ab3840_2427 , 
    RI173bfec0_1820 , 
    RI17408bb0_1465 , 
    RI17455578_1320 , 
    RI17479a40_1143 , 
    RI19a964e8_2638 , 
    RI174c8190_788 , 
    RI19ac63c8_2283 , 
    RI17394720_2032 , 
    RI17496258_1004 , 
    RI19aa9868_2499 , 
    RI17525ad8_649 , 
    RI19a99ad0_2614 , 
    RI173b0f38_1893 , 
    RI17390580_2052 , 
    RI1747fcb0_1113 , 
    RI19aa6988_2519 , 
    RI17500a58_758 , 
    RI19a87b78_2740 , 
    RI1739a990_2002 , 
    RI173e3680_1647 , 
    RI1745b4a0_1291 , 
    RI1749d1e8_970 , 
    RI19ab82c8_2394 , 
    RI17530a28_615 , 
    RI173b8210_1858 , 
    RI173d6e58_1708 , 
    RI1744a790_1373 , 
    RI17511600_712 , 
    RI19acd5b0_2229 , 
    RI1747adf0_1137 , 
    RI19a946e8_2651 , 
    RI174ca080_782 , 
    RI19ac4910_2295 , 
    RI17395ad0_2026 , 
    RI173de7c0_1671 , 
    RI17456298_1316 , 
    RI17486268_1082 , 
    RI19aa10f0_2560 , 
    RI1750c8a8_727 , 
    RI19acffe0_2211 , 
    RI173a1290_1970 , 
    RI17467cc8_1230 , 
    RI174a37a0_939 , 
    RI19ab5118_2416 , 
    RI17335248_2182 , 
    RI173be7c8_1827 , 
    RI174074b8_1472 , 
    RI174458d0_1397 , 
    RI1749cb58_972 , 
    RI19aba578_2378 , 
    RI17455230_1321 , 
    RI17523198_657 , 
    RI19aa7540_2514 , 
    RI17464b90_1245 , 
    RI19a8f648_2687 , 
    RI174ad868_890 , 
    RI19abff78_2332 , 
    RI1733efc8_2134 , 
    RI173c8548_1779 , 
    RI173c8890_1778 , 
    RI174916e0_1027 , 
    RI19aadd50_2469 , 
    RI1751e440_672 , 
    RI19ac1f58_2314 , 
    RI173ac3c0_1916 , 
    RI17519c10_686 , 
    RI17515e30_698 , 
    RI19accc50_2233 , 
    RI173efb60_1587 , 
    RI174a96c8_910 , 
    RI19ab1ba8_2441 , 
    RI1733ae28_2154 , 
    RI1740d098_1444 , 
    RI17457990_1309 , 
    RI1749a740_983 , 
    RI19aa7888_2513 , 
    RI1752c720_628 , 
    RI19a88a00_2734 , 
    RI173b5420_1872 , 
    RI173fe458_1516 , 
    RI173bb9d8_1841 , 
    RI1746efa0_1195 , 
    RI19a89bd0_2726 , 
    RI174b7c78_840 , 
    RI19abb748_2371 , 
    RI17389fc8_2083 , 
    RI175279c8_643 , 
    RI19aa29c8_2548 , 
    RI173b22e8_1887 , 
    RI173fafd8_1532 , 
    RI1739de10_1986 , 
    RI173a7ed8_1937 , 
    RI17497c98_996 , 
    RI19aa8080_2509 , 
    RI17528418_641 , 
    RI19a8b958_2714 , 
    RI173fb9b0_1529 , 
    RI173a0570_1974 , 
    RI1746c1b0_1209 , 
    RI19a8a878_2721 , 
    RI174b4e88_854 , 
    RI19abc378_2366 , 
    RI173465e8_2098 , 
    RI173cfeb0_1742 , 
    RI174479a0_1387 , 
    RI174acb48_894 , 
    RI19ac1670_2319 , 
    RI17395e18_2025 , 
    RI1746c840_1207 , 
    RI19a8aad0_2720 , 
    RI174b5518_852 , 
    RI19abc4e0_2365 , 
    RI17346c78_2096 , 
    RI173d0540_1740 , 
    RI17448030_1385 , 
    RI17489a30_1065 , 
    RI19a9efa8_2577 , 
    RI17512050_710 , 
    RI19acda60_2227 , 
    RI173a4a58_1953 , 
    RI173ed748_1598 , 
    RI1748c190_1053 , 
    RI174a2738_944 , 
    RI19ab4740_2420 , 
    RI173341e0_2187 , 
    RI173bd760_1832 , 
    RI1740d728_1442 , 
    RI1748c4d8_1052 , 
    RI19a9e288_2583 , 
    RI17516880_696 , 
    RI19accea8_2232 , 
    RI173f01f0_1585 , 
    RI174a5528_930 , 
    RI17499390_989 , 
    RI19aa9430_2501 , 
    RI1752a830_634 , 
    RI19a96998_2636 , 
    RI173b4070_1878 , 
    RI173fd0a8_1522 , 
    RI1746dbf0_1201 , 
    RI19a89018_2731 , 
    RI17359350_2090 , 
    RI173d1908_1734 , 
    RI174493e0_1379 , 
    RI17466288_1238 , 
    RI19a905c0_2680 , 
    RI174aef60_883 , 
    RI19ac0ba8_2325 , 
    RI173c9c40_1772 , 
    RI17412c78_1416 , 
    RI1746e910_1197 , 
    RI1752ffd8_617 , 
    RI173b7b80_1860 , 
    RI173d2628_1730 , 
    RI17497fe0_995 , 
    RI19aa81e8_2508 , 
    RI17528940_640 , 
    RI19a8d230_2703 , 
    RI173b2cc0_1884 , 
    RI173fbcf8_1528 , 
    RI173a2988_1963 , 
    RI17485bd8_1084 , 
    RI19aa0d30_2562 , 
    RI1750be58_729 , 
    RI19acfb30_2213 , 
    RI173a0c00_1972 , 
    RI173e98f0_1617 , 
    RI17463498_1252 , 
    RI1748d888_1046 , 
    RI19ab03c0_2452 , 
    RI17518770_690 , 
    RI19aa40c0_2537 , 
    RI173a88b0_1934 , 
    RI173f15a0_1579 , 
    RI174b2db8_864 , 
    RI17484828_1090 , 
    RI19aa24a0_2550 , 
    RI17509f68_735 , 
    RI19a83690_2770 , 
    RI1739f508_1979 , 
    RI173e8540_1623 , 
    RI17460018_1268 , 
    RI174a1d60_947 , 
    RI19ab65b8_2406 , 
    RI17333808_2190 , 
    RI173bcd88_1835 , 
    RI17405a78_1480 , 
    RI17406ae0_1475 , 
    RI1749cea0_971 , 
    RI19aba8c0_2377 , 
    RI17530500_616 , 
    RI173b7ec8_1859 , 
    RI173d4a40_1719 , 
    RI17471700_1183 , 
    RI19a9aac0_2607 , 
    RI174bb350_828 , 
    RI19aca298_2254 , 
    RI173d5418_1716 , 
    RI1744cef0_1361 , 
    RI173a4710_1954 , 
    RI1747b138_1136 , 
    RI19a94940_2650 , 
    RI174ca5a8_781 , 
    RI19ac4b68_2294 , 
    RI173deb08_1670 , 
    RI174565e0_1315 , 
    RI174720d8_1180 , 
    RI19a9b1c8_2604 , 
    RI174bc2c8_825 , 
    RI19aca9a0_2251 , 
    RI1738d100_2068 , 
    RI173d5df0_1713 , 
    RI1744d8c8_1358 , 
    RI173df198_1668 , 
    RI17485890_1085 , 
    RI19aa0b50_2563 , 
    RI1750b930_730 , 
    RI19acf8d8_2214 , 
    RI173a08b8_1973 , 
    RI173e95a8_1618 , 
    RI17461080_1263 , 
    RI174a2a80_943 , 
    RI19ab48a8_2419 , 
    RI17334528_2186 , 
    RI173bdaa8_1831 , 
    RI17406798_1476 , 
    RI17464ed8_1244 , 
    RI19a8f8a0_2686 , 
    RI174adbb0_889 , 
    RI19ac0158_2331 , 
    RI17482410_1101 , 
    RI19aa3418_2543 , 
    RI175066b0_746 , 
    RI19a846f8_2763 , 
    RI1739d0f0_1990 , 
    RI173e6128_1634 , 
    RI1745dc00_1279 , 
    RI173cfb68_1743 , 
    RI1744d238_1360 , 
    RI17471a48_1182 , 
    RI19a9ad18_2606 , 
    RI174bb878_827 , 
    RI19aca4f0_2253 , 
    RI173d5760_1715 , 
    RI174caff8_779 , 
    RI19ac5108_2291 , 
    RI174865b0_1081 , 
    RI19aa1438_2558 , 
    RI1750cdd0_726 , 
    RI19a82538_2778 , 
    RI173a15d8_1969 , 
    RI173ea2c8_1614 , 
    RI1746a0e0_1219 , 
    RI174693c0_1223 , 
    RI19a8d8c0_2700 , 
    RI174b2098_868 , 
    RI19abe808_2345 , 
    RI173437f8_2112 , 
    RI173ccd78_1757 , 
    RI17444bb0_1401 , 
    RI17479d88_1142 , 
    RI19a96740_2637 , 
    RI174c86b8_787 , 
    RI19ac6620_2282 , 
    RI17394a68_2031 , 
    RI1744d580_1359 , 
    RI17471070_1185 , 
    RI19a9ce60_2591 , 
    RI174ba900_830 , 
    RI19acbe40_2240 , 
    RI1738c098_2073 , 
    RI173d4d88_1718 , 
    RI1744c860_1363 , 
    RI1753a460_587 , 
    RI175373a0_595 , 
    RI174a16d0_949 , 
    RI19ab6090_2408 , 
    RI17478348_1150 , 
    RI19a97b68_2628 , 
    RI174c5d78_795 , 
    RI19ac7958_2273 , 
    RI17393028_2039 , 
    RI173dbd18_1684 , 
    RI174537f0_1329 , 
    RI17514990_702 , 
    RI17410860_1427 , 
    RI1749e250_965 , 
    RI19ab8f70_2388 , 
    RI175323f0_610 , 
    RI173b9278_1853 , 
    RI17401f68_1498 , 
    RI173a1c68_1967 , 
    RI173d9270_1697 , 
    RI1748ef80_1039 , 
    RI19aae980_2464 , 
    RI173a9c60_1928 , 
    RI173f2950_1573 , 
    RI174c1a70_808 , 
    RI17471d90_1181 , 
    RI19a9af70_2605 , 
    RI174bbda0_826 , 
    RI19aca748_2252 , 
    RI173d5aa8_1714 , 
    RI1748f610_1037 , 
    RI19aaeea8_2462 , 
    RI173aa2f0_1926 , 
    RI173f2fe0_1571 , 
    RI174a72b0_921 , 
    RI19ab2b98_2434 , 
    RI17338a10_2165 , 
    RI173c1f90_1810 , 
    RI1740ac80_1455 , 
    RI174bdc90_820 , 
    RI17494818_1012 , 
    RI19aaad80_2489 , 
    RI173af4f8_1901 , 
    RI173f81e8_1546 , 
    RI17469078_1224 , 
    RI19a8d668_2701 , 
    RI173434b0_2113 , 
    RI173cca30_1758 , 
    RI17415a68_1402 , 
    RI1748f2c8_1038 , 
    RI19aaeb60_2463 , 
    RI173a9fa8_1927 , 
    RI173f2c98_1572 , 
    RI174c5328_797 , 
    RI17463b28_1250 , 
    RI19a91100_2675 , 
    RI174ac800_895 , 
    RI19ac1490_2320 , 
    RI1733df60_2139 , 
    RI173c74e0_1784 , 
    RI174101d0_1429 , 
    RI17499d68_986 , 
    RI17492400_1023 , 
    RI19aabcf8_2483 , 
    RI1749e8e0_963 , 
    RI19ab92b8_2387 , 
    RI17532e40_608 , 
    RI173b9908_1851 , 
    RI174025f8_1496 , 
    RI173a95d0_1930 , 
    RI174af5f0_881 , 
    RI19abef88_2341 , 
    RI17340d50_2125 , 
    RI173ca2d0_1770 , 
    RI17413308_1414 , 
    RI17476f98_1156 , 
    RI19a97208_2632 , 
    RI174c43b0_800 , 
    RI19ac6ff8_2277 , 
    RI173dacb0_1689 , 
    RI17452788_1334 , 
    RI1748b470_1057 , 
    RI19a9d9a0_2587 , 
    RI1747cec0_1127 , 
    RI19a936f8_2658 , 
    RI174cd410_772 , 
    RI19ac3920_2302 , 
    RI17397ba0_2016 , 
    RI173e0890_1661 , 
    RI174586b0_1305 , 
    RI1749c810_973 , 
    RI19aba398_2379 , 
    RI17462778_1256 , 
    RI19a92bb8_2663 , 
    RI174ab450_901 , 
    RI19ac2f48_2307 , 
    RI1733cbb0_2145 , 
    RI173c6130_1790 , 
    RI1740ee20_1435 , 
    RI1747a760_1139 , 
    RI19a96e48_2634 , 
    RI174c9630_784 , 
    RI19ac6bc0_2279 , 
    RI17395440_2028 , 
    RI173de130_1673 , 
    RI17455c08_1318 , 
    RI1752fab0_618 , 
    RI173b7838_1861 , 
    RI17400528_1506 , 
    RI173d01f8_1741 , 
    RI173967f0_2022 , 
    RI1746d218_1204 , 
    RI19a8b250_2717 , 
    RI174b5ef0_849 , 
    RI19abca80_2362 , 
    RI17347650_2093 , 
    RI173d0f18_1737 , 
    RI17448a08_1382 , 
    RI174896e8_1066 , 
    RI19a9ed50_2578 , 
    RI173bc6f8_1837 , 
    RI1748d1f8_1048 , 
    RI19ab0000_2454 , 
    RI17517d20_692 , 
    RI19a887a8_2735 , 
    RI173a8220_1936 , 
    RI173f0f10_1581 , 
    RI174ae588_886 , 
    RI1747bb10_1133 , 
    RI19a954f8_2645 , 
    RI174cb520_778 , 
    RI19ac52e8_2290 , 
    RI173df4e0_1667 , 
    RI17456fb8_1312 , 
    RI174c3e88_801 , 
    RI19ac6e18_2278 , 
    RI17487960_1075 , 
    RI174713b8_1184 , 
    RI19a9d1a8_2590 , 
    RI174bae28_829 , 
    RI19acc020_2239 , 
    RI1738c3e0_2072 , 
    RI173d50d0_1717 , 
    RI1744cba8_1362 , 
    RI17514eb8_701 , 
    RI19acc5c0_2236 , 
    RI17457300_1311 , 
    RI1746d560_1203 , 
    RI19a8b4a8_2716 , 
    RI17358cc0_2092 , 
    RI173d1278_1736 , 
    RI17448d50_1381 , 
    RI17476c50_1157 , 
    RI19a97028_2633 , 
    RI17391c78_2045 , 
    RI173da968_1690 , 
    RI17452440_1335 , 
    RI17530f50_614 , 
    RI175153e0_700 , 
    RI19acc818_2235 , 
    RI1747d208_1126 , 
    RI19a93950_2657 , 
    RI174cd938_771 , 
    RI19ac3b00_2301 , 
    RI17397ee8_2015 , 
    RI173e0bd8_1660 , 
    RI174589f8_1304 , 
    RI174a20a8_946 , 
    RI19ab6900_2405 , 
    RI17333b50_2189 , 
    RI173bd0d0_1834 , 
    RI17405dc0_1479 , 
    RI17408ef8_1464 , 
    RI17476908_1158 , 
    RI19a99440_2617 , 
    RI174c3960_802 , 
    RI19ac8e70_2263 , 
    RI17391930_2046 , 
    RI173da620_1691 , 
    RI174520f8_1336 , 
    RI174813a8_1106 , 
    RI19aa4ed0_2530 , 
    RI17502e70_751 , 
    RI19a86318_2751 , 
    RI1739c088_1995 , 
    RI1745cb98_1284 , 
    RI17469708_1222 , 
    RI19a8db18_2699 , 
    RI174b23e0_867 , 
    RI19abe9e8_2344 , 
    RI17343b40_2111 , 
    RI173cd0c0_1756 , 
    RI17486c40_1079 , 
    RI19aa17f8_2556 , 
    RI1750d820_724 , 
    RI19a82970_2776 , 
    RI17499048_990 , 
    RI19aa90e8_2502 , 
    RI173b3d28_1879 , 
    RI173fcd60_1523 , 
    RI173ade00_1908 , 
    RI173a6498_1945 , 
    RI173ef188_1590 , 
    RI1749c180_975 , 
    RI1748b7b8_1056 , 
    RI19a9dbf8_2586 , 
    RI173a67e0_1944 , 
    RI173ef4d0_1589 , 
    RI1749e598_964 , 
    RI1747be58_1132 , 
    RI19a95750_2644 , 
    RI174cba48_777 , 
    RI19ac5540_2289 , 
    RI17396b38_2021 , 
    RI173df828_1666 , 
    RI174765c0_1159 , 
    RI19a991e8_2618 , 
    RI174c3438_803 , 
    RI19ac8c18_2264 , 
    RI173da2d8_1692 , 
    RI17451db0_1337 , 
    RI1748ceb0_1049 , 
    RI19aafcb8_2455 , 
    RI175177f8_693 , 
    RI19a86de0_2746 , 
    RI173f0bc8_1582 , 
    RI174ac170_897 , 
    RI1748b128_1058 , 
    RI19a9d658_2588 , 
    RI19acc3e0_2237 , 
    RI173a6150_1946 , 
    RI174a89a8_914 , 
    RI19ab11d0_2445 , 
    RI1733a108_2158 , 
    RI1740c378_1448 , 
    RI173cda98_1753 , 
    RI174a23f0_945 , 
    RI19ab6ae0_2404 , 
    RI17333e98_2188 , 
    RI173bd418_1833 , 
    RI1740b310_1453 , 
    RI17500f80_757 , 
    RI19a85760_2756 , 
    RI174937b0_1017 , 
    RI19aacbf8_2477 , 
    RI175217d0_662 , 
    RI19ab8778_2392 , 
    RI173ae490_1906 , 
    RI173f7180_1551 , 
    RI17334870_2185 , 
    RI174a3e30_937 , 
    RI19ab5640_2413 , 
    RI17407b48_1470 , 
    RI173f5dd0_1557 , 
    RI173de478_1672 , 
    RI1746be68_1210 , 
    RI19a8a530_2722 , 
    RI174b4b40_855 , 
    RI19abc198_2367 , 
    RI173462a0_2099 , 
    RI17447658_1388 , 
    RI174893a0_1067 , 
    RI19a9eaf8_2579 , 
    RI173a43c8_1955 , 
    RI173ed0b8_1600 , 
    RI17463e70_1249 , 
    RI19a91358_2674 , 
    RI1733e2a8_2138 , 
    RI173c7828_1783 , 
    RI17410518_1428 , 
    RI174641b8_1248 , 
    RI19a915b0_2673 , 
    RI174ace90_893 , 
    RI19ac1850_2318 , 
    RI1733e5f0_2137 , 
    RI173c7b70_1782 , 
    RI17475f30_1161 , 
    RI19a98d38_2620 , 
    RI174c29e8_805 , 
    RI19ac8768_2266 , 
    RI173d9c48_1694 , 
    RI17451720_1339 , 
    RI1748f958_1036 , 
    RI19aaf088_2461 , 
    RI1751b5d8_681 , 
    RI19a23a38_2791 , 
    RI173aa638_1925 , 
    RI173f3328_1570 , 
    RI174cc498_775 , 
    RI1748bb00_1055 , 
    RI19a9de50_2585 , 
    RI17515908_699 , 
    RI19acc9f8_2234 , 
    RI173a6b28_1943 , 
    RI173ef818_1588 , 
    RI1751f8e0_668 , 
    RI19ab0c30_2448 , 
    RI17527ef0_642 , 
    RI17468358_1228 , 
    RI19a8f3f0_2688 , 
    RI174b1030_873 , 
    RI19abfd98_2333 , 
    RI17342790_2117 , 
    RI173cbd10_1762 , 
    RI17414d48_1406 , 
    RI17487ca8_1074 , 
    RI19a9ff20_2569 , 
    RI1750f1e8_719 , 
    RI19aceac8_2220 , 
    RI173eb9c0_1607 , 
    RI17477cb8_1152 , 
    RI17333178_2192 , 
    RI174022b0_1497 , 
    RI17456c70_1313 , 
    RI17472420_1179 , 
    RI19a9b678_2602 , 
    RI174bc7f0_824 , 
    RI19acabf8_2250 , 
    RI1738d448_2067 , 
    RI173d6138_1712 , 
    RI1744dc10_1357 , 
    RI1745b7e8_1290 , 
    RI173c1900_1812 , 
    RI17481a38_1104 , 
    RI19aa53f8_2528 , 
    RI175038c0_749 , 
    RI19a86750_2749 , 
    RI1739c718_1993 , 
    RI1745d228_1282 , 
    RI174c9b58_783 , 
    RI19ac46b8_2296 , 
    RI1747b480_1135 , 
    RI19a94b98_2649 , 
    RI174a6c20_923 , 
    RI19ab2670_2436 , 
    RI17338380_2167 , 
    RI1748e5a8_1042 , 
    RI174caad0_780 , 
    RI19ac4dc0_2293 , 
    RI17396160_2024 , 
    RI173dee50_1669 , 
    RI17456928_1314 , 
    RI1747aaa8_1138 , 
    RI19a94490_2652 , 
    RI17395788_2027 , 
    RI17455f50_1317 , 
    RI1747fff8_1112 , 
    RI19aa44f8_2535 , 
    RI1739acd8_2001 , 
    RI173e39c8_1646 , 
    RI1749d530_969 , 
    RI19ab8430_2393 , 
    RI173b8558_1857 , 
    RI17401248_1502 , 
    RI17481060_1107 , 
    RI19aa4cf0_2531 , 
    RI17502948_752 , 
    RI19a860c0_2752 , 
    RI1739bd40_1996 , 
    RI173e4d78_1640 , 
    RI1745c850_1285 , 
    RI17511b28_711 , 
    RI19acd808_2228 , 
    RI173ed400_1599 , 
    RI17489d78_1064 , 
    RI1747b7c8_1134 , 
    RI19a952a0_2646 , 
    RI173386c8_2166 , 
    RI173c1c48_1811 , 
    RI1740a938_1456 , 
    RI174a51e0_931 , 
    RI17359008_2091 , 
    RI175298b8_637 , 
    RI19a91c40_2670 , 
    RI173b3698_1881 , 
    RI173fc6d0_1525 , 
    RI17498d00_991 , 
    RI19aa8da0_2504 , 
    RI173b39e0_1880 , 
    RI173fca18_1524 , 
    RI173ab9e8_1919 , 
    RI173d15c0_1735 , 
    RI17506188_747 , 
    RI19a843b0_2764 , 
    RI1739cda8_1991 , 
    RI173e5de0_1635 , 
    RI1745d8b8_1280 , 
    RI1746d8a8_1202 , 
    RI19a8b700_2715 , 
    RI1750d2f8_725 , 
    RI19a82790_2777 , 
    RI174868f8_1080 , 
    RI19aa1618_2557 , 
    RI173a1920_1968 , 
    RI173ea610_1613 , 
    RI1746c4f8_1208 , 
    RI17449098_1380 , 
    RI1754bad0_26 , 
    RI1754a5b8_71 , 
    RI1754a630_70 , 
    RI1754a6a8_69 , 
    RI1754a720_68 , 
    RI17538c00_591 , 
    RI19a25298_2780 , 
    RI1754b788_33 , 
    RI1754b878_31 , 
    RI1754c430_6 , 
    RI17536d88_596 , 
    RI1754b800_32 , 
    RI1754b530_38 , 
    RI19a822e0_2779 , 
    RI19ad0700_2208 , 
    RI1754bcb0_22 , 
    RI19a24ed8_2782 , 
    RI19a250b8_2781 , 
    RI1754be18_19 , 
    RI1754b350_42 , 
    RI1754c250_10 , 
    RI1754b1e8_45 , 
    RI19a24320_2787 , 
    RI19a24578_2786 , 
    RI1754b5a8_37 , 
    RI19ad21b8_2198 , 
    RI1754c160_12 , 
    RI1754a900_64 , 
    RI19a24c80_2783 , 
    RI1754bf08_17 , 
    RI1754ac48_57 , 
    RI1754bf80_16 , 
    RI1754bc38_23 , 
    RI19a240c8_2788 , 
    RI1754c070_14 , 
    RI1754b3c8_41 , 
    RI1754af18_51 , 
    RI1754b080_48 , 
    RI1754af90_50 , 
    RI1754bda0_20 , 
    RI1754aea0_52 , 
    RI1754b260_44 , 
    RI19ad0bb0_2206 , 
    RI19a24a28_2784 , 
    RI1754ae28_53 , 
    RI1754a888_65 , 
    RI1754bbc0_24 , 
    RI19ad0e08_2205 , 
    RI1754a810_66 , 
    RI1754b440_40 , 
    RI1754adb0_54 , 
    RI1754c3b8_7 , 
    RI19ad1060_2204 , 
    RI1754ba58_27 , 
    RI1754c340_8 , 
    RI1754aa68_61 , 
    RI1754ad38_55 , 
    RI19ad12b8_2203 , 
    RI1754be90_18 , 
    RI1754c2c8_9 , 
    RI1754c1d8_11 , 
    RI19a247d0_2785 , 
    RI1754b170_46 , 
    RI1754aae0_60 , 
    RI1754acc0_56 , 
    RI1754a978_63 , 
    RI19ad1588_2202 , 
    RI1754b620_36 , 
    RI1754bd28_21 , 
    RI1754b9e0_28 , 
    RI1754bb48_25 , 
    RI1754ab58_59 , 
    RI1754abd0_58 , 
    RI1754b2d8_43 , 
    RI1754c598_3 , 
    RI19ad1858_2201 , 
    RI1754b4b8_39 , 
    RI1754b0f8_47 , 
    RI1754c0e8_13 , 
    RI1754bff8_15 , 
    RI1754b698_35 , 
    RI19ad1c18_2200 , 
    RI1754c520_4 , 
    RI1754b968_29 , 
    RI19ad1ee8_2199 , 
    RI1754b008_49 , 
    RI1754c4a8_5 , 
    RI1754b710_34 , 
    RI1754a9f0_62 , 
    RI1754b8f0_30 , 
    RI19ad0958_2207 , 
    R_147ef_11ce6748 , 
    R_5f38_10569f58 , 
    R_13287_11ce6b08 , 
    R_c94b_102f7608 , 
    R_20a_1204ce78 , 
    R_12f29_10571bb8 , 
    R_13a43_13a1dec8 , 
    R_1474d_1056fbd8 , 
    R_14493_12657988 , 
    R_11fd1_11ce17e8 , 
    R_14705_1264d248 , 
    R_105_f8cc2b8 , 
    R_13cb9_11ce3c28 , 
    R_138ee_13309fa8 , 
    R_129dc_11543018 , 
    R_10bcf_11ce1ba8 , 
    R_13b6e_13a1e648 , 
    R_14840_13a13ec8 , 
    R_13482_10563838 , 
    R_12d08_12650088 , 
    R_10303_12b42dd8 , 
    R_1437c_1056ac78 , 
    R_87e9_1056cd98 , 
    R_a30d_13320588 , 
    R_144a2_133222e8 , 
    R_1236b_13a1c8e8 , 
    R_1396e_105627f8 , 
    R_9ba7_10567258 , 
    R_1f3_13797a68 , 
    R_11c_13796528 , 
    R_7a_1331e148 , 
    R_117c9_1264ba88 , 
    R_13b3f_1153ed38 , 
    R_11abc_1264c2a8 , 
    R_20d_137962a8 , 
    R_207_1265a548 , 
    R_14828_1207a118 , 
    R_148eb_105aa7d8 , 
    R_f3a4_10568bf8 , 
    R_1b6_13799d68 , 
    R_13429_1207f4d8 , 
    R_14506_1056e878 , 
    R_159_12b3d158 , 
    R_108_105aaeb8 , 
    R_102_13794cc8 , 
    R_b1_12053638 , 
    R_54_13309d28 , 
    R_145d8_12b3ae58 , 
    R_1278a_12083718 , 
    R_13640_11cdeae8 , 
    R_f706_11542578 , 
    R_dc82_1153ebf8 , 
    R_1491b_1265ef08 , 
    R_14a05_10569738 , 
    R_13fc5_102eac28 , 
    R_1405a_115415d8 , 
    R_136b3_126461c8 , 
    R_1a0_132f9c88 , 
    R_16f_1265bee8 , 
    R_1480d_105a9dd8 , 
    R_61_13304288 , 
    R_e082_13798fa8 , 
    R_10c7d_12082bd8 , 
    R_14793_1379e188 , 
    R_11ee1_102f4688 , 
    R_128ba_12b27758 , 
    R_70_120513d8 , 
    R_129f0_12049bd8 , 
    R_117e7_102f5588 , 
    R_fee6_13309e68 , 
    R_148f7_132f3ce8 , 
    R_1362d_11ce39a8 , 
    R_10693_126510c8 , 
    R_11998_12656808 , 
    R_143ec_11537df8 , 
    R_138e8_1264afe8 , 
    R_12650_12649b48 , 
    R_137a1_105b63f8 , 
    R_13afd_120772d8 , 
    R_1490c_1264a7c8 , 
    R_105e5_13306f88 , 
    R_12e2b_132fa868 , 
    R_144e7_12b38e78 , 
    R_143e4_11cddf08 , 
    R_1324a_1264c348 , 
    R_1215a_11542ed8 , 
    R_f685_11541678 , 
    R_149ba_102ecb68 , 
    R_135dc_12646088 , 
    R_1476c_11cd7928 , 
    R_146bd_11537998 , 
    R_1df_12b39378 , 
    R_13ee8_133069e8 , 
    R_130_1265ac28 , 
    R_65_12047c98 , 
    R_13d75_1330d6a8 , 
    R_13933_12081198 , 
    R_133b5_12648388 , 
    R_125a0_13311488 , 
    R_8c_1379a808 , 
    R_eadc_1207ead8 , 
    R_134c7_126487e8 , 
    R_11df5_1056e9b8 , 
    R_144d5_102f8aa8 , 
    R_12b2a_102eed28 , 
    R_143d2_11538898 , 
    R_1462c_102f8508 , 
    R_13269_11543658 , 
    R_f4_1331e0a8 , 
    R_d7_132fde28 , 
    R_238_1204ec78 , 
    R_21b_1265e508 , 
    R_12f3d_12b38b58 , 
    R_112f1_1153c858 , 
    R_f09_f8c93d8 , 
    R_1487c_11cd99a8 , 
    R_c08f_1207cb98 , 
    R_923a_13a1ab88 , 
    R_14042_102f2108 , 
    R_143e8_102f3b48 , 
    R_c2e7_13a19e68 , 
    R_c175_12045118 , 
    R_1450f_102f8b48 , 
    R_12b14_12077238 , 
    R_149e4_13a1c528 , 
    R_12a04_11ce2968 , 
    R_145ed_13a14e68 , 
    R_13884_13796488 , 
    R_13b0b_1330a688 , 
    R_b5a4_102f4868 , 
    R_14584_1056ec38 , 
    R_13cee_12653148 , 
    R_10bed_12080ab8 , 
    R_117f0_102ef4a8 , 
    R_10a2a_133048c8 , 
    R_1be_137995e8 , 
    R_151_12b448b8 , 
    R_ef06_10563c98 , 
    R_f9d4_1056b178 , 
    R_e88a_13a13a68 , 
    R_13c67_102f38c8 , 
    R_128eb_10568dd8 , 
    R_12eaf_f8c3118 , 
    R_204_12039778 , 
    R_14951_1265ebe8 , 
    R_149c3_11ce5348 , 
    R_1ad_12b28e78 , 
    R_13f99_102f0da8 , 
    R_162_12b25e58 , 
    R_12003_11cdf628 , 
    R_10b_11539478 , 
    R_ff_1203c6f8 , 
    R_1484f_1153ea18 , 
    R_a8_12b425b8 , 
    R_5d_13312068 , 
    R_210_12043bd8 , 
    R_13d84_102f4188 , 
    R_142e1_10568658 , 
    R_10f30_11cd9ae8 , 
    R_1293d_12b43d78 , 
    R_10b34_1056da18 , 
    R_11a07_102eb4e8 , 
    R_145b1_12082db8 , 
    R_12c96_13a190a8 , 
    R_d3b0_10565958 , 
    R_13f2c_102f4b88 , 
    R_fb8a_13a18608 , 
    R_130d5_13319c88 , 
    R_13f89_102f36e8 , 
    R_146ff_13a1a4a8 , 
    R_10ccb_1264f868 , 
    R_124c3_1056f138 , 
    R_10786_102f2568 , 
    R_12a16_10568e78 , 
    R_10726_102ef408 , 
    R_137d3_12656da8 , 
    R_13863_11cddb48 , 
    R_14993_102f27e8 , 
    R_bab1_1264a2c8 , 
    R_1451e_10565818 , 
    R_12a46_126515c8 , 
    R_e7da_102f3508 , 
    R_12756_13a1f0e8 , 
    R_c4_13797ba8 , 
    R_128da_1207ec18 , 
    R_c282_12076838 , 
    R_1272e_1056cbb8 , 
    R_14a5f_120797b8 , 
    R_14448_12663648 , 
    R_c2_12048058 , 
    R_1372d_11ce2aa8 , 
    R_f878_1207c7d8 , 
    R_13a76_13797888 , 
    R_13a17_13796b68 , 
    R_1cb_12044ad8 , 
    R_14462_12b3f8b8 , 
    R_6021_1379bd48 , 
    R_144_13795128 , 
    R_1383e_105671b8 , 
    R_147ab_1056a6d8 , 
    R_c6_1330e0a8 , 
    R_249_12654368 , 
    R_1305a_13796ca8 , 
    R_12e4b_13307348 , 
    R_14a38_137a1e28 , 
    R_d1de_11cd9ea8 , 
    R_138e2_11cd83c8 , 
    R_13e62_1056dab8 , 
    R_114a7_1331d748 , 
    R_12f53_13319648 , 
    R_f8a4_11543a18 , 
    R_11ec3_13a157c8 , 
    R_12c06_11cdac68 , 
    R_12be8_12649788 , 
    R_136c6_11cdc6a8 , 
    R_1482e_13a1a228 , 
    R_10ba7_115431f8 , 
    R_89f2_11545098 , 
    R_11953_1153c538 , 
    R_9e64_11ce48a8 , 
    R_e77d_11ce3ea8 , 
    R_1091c_13a1a2c8 , 
    R_114ec_12650628 , 
    R_1286a_11cdcd88 , 
    R_10d6d_1265db08 , 
    R_1228f_1331f0e8 , 
    R_1c5_126590a8 , 
    R_14490_132f7d48 , 
    R_1a1_1264a408 , 
    R_976e_12056398 , 
    R_6845_12648ec8 , 
    R_16e_1379a3a8 , 
    R_14a_12657528 , 
    R_12718_10566fd8 , 
    R_145c9_12075438 , 
    R_c0_132fa5e8 , 
    R_9c_12655f48 , 
    R_d230_102edec8 , 
    R_69_12658888 , 
    R_13097_11ce5b68 , 
    R_11051_1264a5e8 , 
    R_145f0_11536818 , 
    R_13ccd_132f9288 , 
    R_e0_12661ac8 , 
    R_22f_1331df68 , 
    R_12a2a_11cd9f48 , 
    R_10a54_11540458 , 
    R_d027_13795628 , 
    R_144d2_105677f8 , 
    R_14638_11cd9228 , 
    R_1454b_10568338 , 
    R_147fe_1265bb28 , 
    R_e861_12650448 , 
    R_c03c_137931e8 , 
    R_13574_102f97c8 , 
    R_10e6d_102ec0c8 , 
    R_c8_1331c348 , 
    R_247_12b3bad8 , 
    R_77_126636e8 , 
    R_13a50_1056bb78 , 
    R_129a5_11543798 , 
    R_ef35_102f6d48 , 
    R_1028c_137951c8 , 
    R_1348b_12051838 , 
    R_11f8b_11cdc428 , 
    R_1452d_f8c5878 , 
    R_12a3b_12650308 , 
    R_13fd5_12079d58 , 
    R_dd89_13302de8 , 
    R_13dcc_102f7ec8 , 
    R_14822_102f5768 , 
    R_baf1_12084e38 , 
    R_1315c_11ce75a8 , 
    R_df0e_12654d68 , 
    R_efea_11cdc248 , 
    R_fe90_13a14a08 , 
    R_1453c_102ec208 , 
    R_aaa7_102edba8 , 
    R_13c4e_13a1c988 , 
    R_f758_13a13d88 , 
    R_1485e_12b38f18 , 
    R_ece9_1264c488 , 
    R_14a35_12037f18 , 
    R_1190c_102ecfc8 , 
    R_12810_12650d08 , 
    R_f016_12044df8 , 
    R_1494e_13a14f08 , 
    R_14344_1264eaa8 , 
    R_10e_1265af48 , 
    R_13f62_12075758 , 
    R_fc_133201c8 , 
    R_1378e_11cdd8c8 , 
    R_147eb_120847f8 , 
    R_13331_13308ec8 , 
    R_213_12654f48 , 
    R_146ae_1265dc48 , 
    R_201_1153b138 , 
    R_11d47_f8cc0d8 , 
    R_c820_13a19328 , 
    R_edbe_132fbd08 , 
    R_be_132f4148 , 
    R_a1_12043c78 , 
    R_131b9_102f29c8 , 
    R_12eb9_1153f738 , 
    R_146e1_1153fb98 , 
    R_1487f_13a173e8 , 
    R_13fb4_11544af8 , 
    R_1446b_10568798 , 
    R_ef60_1264cf28 , 
    R_1463b_1207bd38 , 
    R_13166_1153aff8 , 
    R_10a4b_10565bd8 , 
    R_14599_12080c98 , 
    R_10b18_12080018 , 
    R_7254_12055078 , 
    R_db04_1207b3d8 , 
    R_149f9_10570cb8 , 
    R_14a4a_1265d608 , 
    R_14796_1264b808 , 
    R_120d3_1379f3a8 , 
    R_119cb_102f2068 , 
    R_12acb_10565458 , 
    R_145b4_12083358 , 
    R_11ae9_12651528 , 
    R_13af6_f8ce6f8 , 
    R_13451_102f0128 , 
    R_ef8c_1204e098 , 
    R_ca_12b3e058 , 
    R_245_f8c5ff8 , 
    R_af_12b2a8b8 , 
    R_10e57_11544eb8 , 
    R_b243_f8c5698 , 
    R_13633_13a13248 , 
    R_11c97_10562078 , 
    R_13838_102f5e48 , 
    R_efb7_13a1bc68 , 
    R_d4db_10566038 , 
    R_10bc8_11ce66a8 , 
    R_c9c0_102eee68 , 
    R_13608_10563798 , 
    R_8f_12b299b8 , 
    R_59_133089c8 , 
    R_134f1_102ebf88 , 
    R_10499_1331e828 , 
    R_14424_102f8f08 , 
    R_1d6_133209e8 , 
    R_ebe2_13a18568 , 
    R_139_12b44ef8 , 
    R_97_13792c48 , 
    R_144ed_105660d8 , 
    R_120c8_11541d58 , 
    R_11736_11cde408 , 
    R_149a8_13317528 , 
    R_1450c_1056eff8 , 
    R_147d9_120828b8 , 
    R_11ea5_1264a9a8 , 
    R_11425_1207c918 , 
    R_d53e_1207c2d8 , 
    R_14787_12b352b8 , 
    R_13cf3_10571078 , 
    R_13f36_1330ebe8 , 
    R_d00d_102ee968 , 
    R_a1e6_11cde368 , 
    R_13f77_13a19648 , 
    R_118_132f5f48 , 
    R_13688_120832b8 , 
    R_1f7_105a9978 , 
    R_f630_1056b858 , 
    R_136a1_1153fa58 , 
    R_1b7_126577a8 , 
    R_158_12b27938 , 
    R_ec_1330a868 , 
    R_223_f8c32f8 , 
    R_133bf_11543338 , 
    R_f2a8_102f47c8 , 
    R_e112_12076e78 , 
    R_12b72_1056c6b8 , 
    R_2f00_102f3d28 , 
    R_14819_1331de28 , 
    R_e809_13313c48 , 
    R_14358_11cd8788 , 
    R_1473e_11543b58 , 
    R_139c7_102ed1a8 , 
    R_13d65_12036a78 , 
    R_12c10_102ea548 , 
    R_13870_11ce5e88 , 
    R_dede_13a16448 , 
    R_12c49_12b27438 , 
    R_1192b_12645e08 , 
    R_bd66_126533c8 , 
    R_13fa2_1379f6c8 , 
    R_13407_1056df18 , 
    R_118b0_1204acb8 , 
    R_13c3e_126496e8 , 
    R_1438a_11cda268 , 
    R_11e51_102fa268 , 
    R_102b9_132f6588 , 
    R_d9_1330dec8 , 
    R_bc_13799c28 , 
    R_236_13795f88 , 
    R_ffee_1264d568 , 
    R_10ea9_102f8788 , 
    R_14852_13a154a8 , 
    R_e696_11cdce28 , 
    R_1ae_1203c3d8 , 
    R_1457e_133027e8 , 
    R_161_12656c68 , 
    R_127_12b3cc58 , 
    R_ea26_1265a4a8 , 
    R_1e8_11539298 , 
    R_139e4_102f59e8 , 
    R_1477b_1204f218 , 
    R_1459c_12056a78 , 
    R_1336e_11545138 , 
    R_108cd_102f7ce8 , 
    R_13b4f_13305c28 , 
    R_1a2_12b423d8 , 
    R_16d_12664c28 , 
    R_14656_11ce6ce8 , 
    R_827e_1207e998 , 
    R_11ab0_1204a358 , 
    R_144ab_12b39af8 , 
    R_144c3_12080338 , 
    R_12794_102f5b28 , 
    R_13149_102f7888 , 
    R_144e4_12b28838 , 
    R_13e_12660da8 , 
    R_123_1330d888 , 
    R_e7_137956c8 , 
    R_cc_12038918 , 
    R_137c7_102f79c8 , 
    R_243_13796d48 , 
    R_13795_13795588 , 
    R_228_10570c18 , 
    R_13f01_1056e2d8 , 
    R_13d8e_11cd77e8 , 
    R_1ec_12039ef8 , 
    R_f175_13a17ca8 , 
    R_1d1_126540e8 , 
    R_14409_12b434b8 , 
    R_138b2_102f06c8 , 
    R_14653_1207e0d8 , 
    R_13044_102f7a68 , 
    R_13133_13a1ae08 , 
    R_10b8f_1265ad68 , 
    R_12e35_12b3b858 , 
    R_12df0_12050bb8 , 
    R_fc88_1207be78 , 
    R_13804_102ef548 , 
    R_13b68_137a1ba8 , 
    R_134_13312b68 , 
    R_14990_1331ae08 , 
    R_1db_12043db8 , 
    R_ccdc_102f6488 , 
    R_1494b_11ce61a8 , 
    R_12c39_10562ed8 , 
    R_131c2_11ce4b28 , 
    R_12d97_126626a8 , 
    R_12d59_12b26b78 , 
    R_1352d_13315188 , 
    R_12c4f_13321d48 , 
    R_1343e_10562d98 , 
    R_1345b_102fa088 , 
    R_1167d_115410d8 , 
    R_14008_1264dec8 , 
    R_11bc8_11544e18 , 
    R_13c9a_1207e178 , 
    R_148be_12b27f78 , 
    R_14360_105ad078 , 
    R_13aa3_12078138 , 
    R_116da_13a1a7c8 , 
    R_14732_102f5448 , 
    R_cec6_132f3608 , 
    R_133dc_13a1ea08 , 
    R_14942_f8c5058 , 
    R_13a0f_10563018 , 
    R_bd10_f8ce978 , 
    R_12da1_12647528 , 
    R_12af5_12052418 , 
    R_13cf9_13a1c0c8 , 
    R_13658_12646628 , 
    R_149bd_1204adf8 , 
    R_13233_11cde908 , 
    R_12585_1207a898 , 
    R_118e9_10564a58 , 
    R_1359a_13a18928 , 
    R_12451_13a1d568 , 
    R_dcbb_1265bf88 , 
    R_f424_13a1b948 , 
    R_1226a_11cdef48 , 
    R_14641_13a12d48 , 
    R_1257c_11ce4448 , 
    R_e309_120806f8 , 
    R_11ccc_13314be8 , 
    R_146c0_13a15908 , 
    R_14843_13a196e8 , 
    R_11d00_1207f9d8 , 
    R_14a1d_13a14c88 , 
    R_13d54_11ce00c8 , 
    R_135b5_132fdd88 , 
    R_d40b_10569058 , 
    R_145f9_102ee148 , 
    R_14882_1056d838 , 
    R_101a4_f8c2ad8 , 
    R_13abf_13a15188 , 
    R_eab3_126509e8 , 
    R_8296_13322608 , 
    R_6d_12036618 , 
    R_50_12b3c118 , 
    R_11b19_102ee508 , 
    R_de1d_13a193c8 , 
    R_14477_11cdcc48 , 
    R_1195d_12038198 , 
    R_14527_102eb6c8 , 
    R_be8c_126504e8 , 
    R_11e87_12b3c398 , 
    R_14a02_13309aa8 , 
    R_12b_1203e6d8 , 
    R_f1_13799ea8 , 
    R_21e_126608a8 , 
    R_1e4_12b28338 , 
    R_115ff_13304148 , 
    R_10d8e_1264cfc8 , 
    R_11500_12083c18 , 
    R_c4bc_137945e8 , 
    R_1465c_10568f18 , 
    R_133e6_11cd9048 , 
    R_7c4f_11ce4a88 , 
    R_11f78_12b2c118 , 
    R_1013a_132f59a8 , 
    R_149e1_105b62b8 , 
    R_150_1330cac8 , 
    R_111_12b3e238 , 
    R_f9_1204ba78 , 
    R_ba_1331bc68 , 
    R_4b_1264c028 , 
    R_216_1204a038 , 
    R_13733_f8d0098 , 
    R_1fe_120539f8 , 
    R_146de_12648748 , 
    R_1bf_1265cd48 , 
    R_74_1331da68 , 
    R_f5c3_1264d108 , 
    R_f1f7_120367f8 , 
    R_e338_13301ac8 , 
    R_1486d_1056e558 , 
    R_13e2d_12047fb8 , 
    R_12344_137a0de8 , 
    R_14729_10570178 , 
    R_13364_105717f8 , 
    R_11160_1153e298 , 
    R_10a01_11cde228 , 
    R_13c6f_12041658 , 
    R_148c4_10568978 , 
    R_11c81_132f7348 , 
    R_10ec5_11cdb028 , 
    R_14441_12659008 , 
    R_cbab_105a9a18 , 
    R_1238a_126482e8 , 
    R_a6_12660448 , 
    R_12b36_11ce6428 , 
    R_dc46_10566498 , 
    R_11f_137936e8 , 
    R_ce_12055fd8 , 
    R_241_132fd748 , 
    R_147f8_1207ccd8 , 
    R_1f0_13798a08 , 
    R_1467d_1056bcb8 , 
    R_14668_11546178 , 
    R_132cc_1153edd8 , 
    R_136ba_11ce37c8 , 
    R_12c23_102f1d48 , 
    R_106be_1264edc8 , 
    R_11bde_10564878 , 
    R_11a1a_11cd9a48 , 
    R_9548_11ce6ba8 , 
    R_f451_11542438 , 
    R_119b7_105663f8 , 
    R_142e5_102f2388 , 
    R_147e4_13a19dc8 , 
    R_d862_12661348 , 
    R_d940_13a19d28 , 
    R_eb8c_13a19288 , 
    R_1175e_11cda088 , 
    R_146f9_11ce4768 , 
    R_14551_102eae08 , 
    R_14578_12b3a6d8 , 
    R_1467a_13a13568 , 
    R_1130e_1056bfd8 , 
    R_1493f_1056d3d8 , 
    R_14948_102f76a8 , 
    R_10230_1153d1b8 , 
    R_f4d1_13a17848 , 
    R_14772_11cda8a8 , 
    R_1466e_1203e138 , 
    R_14999_120382d8 , 
    R_9d72_102f18e8 , 
    R_eeaf_10566f38 , 
    R_13083_12b3ff98 , 
    R_e288_11541fd8 , 
    R_13969_102ea408 , 
    R_13825_1264d928 , 
    R_134a8_13a13c48 , 
    R_fcde_115390b8 , 
    R_14566_102f6988 , 
    R_f5eb_11544558 , 
    R_12318_102ec348 , 
    R_d2c9_11cd9408 , 
    R_16c_132f7ca8 , 
    R_d894_1056f778 , 
    R_12323_102ec8e8 , 
    R_1a3_13303108 , 
    R_118ba_13307ac8 , 
    R_12704_10562938 , 
    R_148c7_1264d888 , 
    R_148bb_12661d48 , 
    R_1221a_13a1d248 , 
    R_135b0_12651348 , 
    R_1470e_10562898 , 
    R_efa_1207d1d8 , 
    R_ce1e_102f95e8 , 
    R_126e3_105b5c78 , 
    R_14026_102ecd48 , 
    R_11e36_102ed608 , 
    R_11515_12039318 , 
    R_108e3_1056dd38 , 
    R_128f4_1207aa78 , 
    R_147ae_1207ce18 , 
    R_12235_12650e48 , 
    R_12183_12052eb8 , 
    R_14647_102f04e8 , 
    R_13aef_11cdd968 , 
    R_1249f_102f9368 , 
    R_f34d_13a18ec8 , 
    R_12c3f_f8cfd78 , 
    R_13d5d_1153d4d8 , 
    R_12126_102ef228 , 
    R_ad_12b3b358 , 
    R_92_13312d48 , 
    R_113db_f8cb4f8 , 
    R_10d98_f8c6318 , 
    R_1481f_1264dce8 , 
    R_ad98_102f3aa8 , 
    R_55_132f50e8 , 
    R_102d5_f8ced38 , 
    R_144ae_11545ef8 , 
    R_a3e0_12655308 , 
    R_5dbf_13a15f48 , 
    R_e2_1203f858 , 
    R_22d_1379de68 , 
    R_135c4_105b5bd8 , 
    R_13cff_13a16308 , 
    R_12692_102eb8a8 , 
    R_13375_13794a48 , 
    R_12f6a_10562438 , 
    R_128c4_102ea5e8 , 
    R_122f0_12650f88 , 
    R_14855_12056f78 , 
    R_14885_13795a88 , 
    R_bb92_11ce0ca8 , 
    R_8b04_1265cf28 , 
    R_e71c_115426b8 , 
    R_14a23_120545d8 , 
    R_149_1330f408 , 
    R_b8_13305048 , 
    R_1c6_1379cce8 , 
    R_e13d_102eb448 , 
    R_14617_11ce2f08 , 
    R_13557_11545778 , 
    R_148cd_12082c78 , 
    R_11768_1264ffe8 , 
    R_12503_11cdd008 , 
    R_1239d_1330d1a8 , 
    R_1448c_105662b8 , 
    R_160_f8c0d78 , 
    R_143_13795e48 , 
    R_1252c_102f1208 , 
    R_1cc_f8cc858 , 
    R_149de_11cde7c8 , 
    R_1af_12b40678 , 
    R_a28f_11ce5708 , 
    R_f7ae_11ce57a8 , 
    R_1243d_10571118 , 
    R_d0df_126478e8 , 
    R_1498d_1153fe18 , 
    R_10350_11cda6c8 , 
    R_103a6_10569878 , 
    R_128b0_1056c118 , 
    R_14936_10561e98 , 
    R_10d1b_11cd7748 , 
    R_ed92_102eea08 , 
    R_145d2_11cdb208 , 
    R_109f6_1153ca38 , 
    R_cc46_1207b298 , 
    R_11006_126501c8 , 
    R_188_1265c348 , 
    R_187_12b25d18 , 
    R_12f_1379dbe8 , 
    R_db_12663f08 , 
    R_84_12652ce8 , 
    R_81_12042a58 , 
    R_234_12b43af8 , 
    R_1e0_133037e8 , 
    R_13ed7_1207ad98 , 
    R_189_f8c6458 , 
    R_186_126553a8 , 
    R_157_132f7a28 , 
    R_d0_105aa238 , 
    R_23f_13307848 , 
    R_11399_12b3c1b8 , 
    R_1b8_11537358 , 
    R_f82c_f8cdc58 , 
    R_d9ca_10562bb8 , 
    R_145f6_f8c3398 , 
    R_1449c_11ce71e8 , 
    R_13850_13a1fe08 , 
    R_135e3_13306da8 , 
    R_ec0b_132fa368 , 
    R_147e0_13a12fc8 , 
    R_13add_132ff728 , 
    R_f65b_12084578 , 
    R_10cb4_11cdf9e8 , 
    R_18a_133173e8 , 
    R_185_12042cd8 , 
    R_134d0_12651028 , 
    R_144f3_102f3fa8 , 
    R_12dd1_f8c52d8 , 
    R_135a9_10567938 , 
    R_11b39_102ec988 , 
    R_1386a_102ebda8 , 
    R_14747_12042b98 , 
    R_148d0_137a0a28 , 
    R_11f4d_137986e8 , 
    R_13d05_12081378 , 
    R_f56e_102f2608 , 
    R_62_12b26498 , 
    R_10e0b_1056abd8 , 
    R_ba73_1264c8e8 , 
    R_14888_12653288 , 
    R_fc34_1379c428 , 
    R_18b_12663fa8 , 
    R_184_1153acd8 , 
    R_119d5_1331dc48 , 
    R_122b5_13305688 , 
    R_e051_12649f08 , 
    R_ca0a_10567438 , 
    R_10a84_115427f8 , 
    R_668e_10563f18 , 
    R_14539_102f7108 , 
    R_c3d6_11cdb7a8 , 
    R_11703_132fa728 , 
    R_1472f_105708f8 , 
    R_1307a_11cdc1a8 , 
    R_fdae_1153d258 , 
    R_13ac5_102ee3c8 , 
    R_120bd_1153ff58 , 
    R_13f6e_12649dc8 , 
    R_1177b_1207fbb8 , 
    R_f804_1379efe8 , 
    R_111d5_13a17c08 , 
    R_14750_13304008 , 
    R_137d9_12055e98 , 
    R_87_132ffa48 , 
    R_7e_137949a8 , 
    R_f140_1056f598 , 
    R_d43f_12079678 , 
    R_11900_1056f6d8 , 
    R_18c_12660e48 , 
    R_c969_1330f9a8 , 
    R_183_126587e8 , 
    R_11093_102f60c8 , 
    R_f31e_120770f8 , 
    R_f06_1265f728 , 
    R_d5cf_102f5128 , 
    R_10874_12037838 , 
    R_11324_13a1f228 , 
    R_13621_120823b8 , 
    R_120dd_f8cdcf8 , 
    R_148d3_12049a98 , 
    R_13e42_12648888 , 
    R_144c0_12078db8 , 
    R_12978_13316d08 , 
    R_11b5e_13a1b088 , 
    R_13025_13a1ef08 , 
    R_e615_12084bb8 , 
    R_149b7_102ea4a8 , 
    R_1497e_1207ef38 , 
    R_11fee_12b2a3b8 , 
    R_11b_12b43198 , 
    R_5e_126647c8 , 
    R_1f4_1265d108 , 
    R_1445f_13792888 , 
    R_13981_13798aa8 , 
    R_14569_11cdbfc8 , 
    R_114_12b3e4b8 , 
    R_f6_12664188 , 
    R_9f_12054d58 , 
    R_66_13308068 , 
    R_219_1203c338 , 
    R_132a5_12654868 , 
    R_f9aa_11cdd5a8 , 
    R_1fb_126610c8 , 
    R_1a4_13798648 , 
    R_16b_1331a2c8 , 
    R_9a_12658568 , 
    R_13c54_102f6e88 , 
    R_14933_1207e5d8 , 
    R_a6b7_1264b588 , 
    R_10fad_13a15548 , 
    R_18d_13321a28 , 
    R_182_13315cc8 , 
    R_14a58_102f65c8 , 
    R_c8f6_132f4a08 , 
    R_1458d_13a17ac8 , 
    R_126d9_11545598 , 
    R_10942_102f85a8 , 
    R_14a32_12654ea8 , 
    R_b7bc_12b28798 , 
    R_1389f_11cda3a8 , 
    R_14602_102ed7e8 , 
    R_100bf_1330b9e8 , 
    R_112eb_115386b8 , 
    R_146d5_105b59f8 , 
    R_1206a_1207c878 , 
    R_e2de_1264ce88 , 
    R_13b3a_11cddaa8 , 
    R_13739_10563bf8 , 
    R_148d6_11cd86e8 , 
    R_1319d_11544918 , 
    R_12f7f_12077eb8 , 
    R_1242c_f8cda78 , 
    R_14483_12054fd8 , 
    R_14456_102ea728 , 
    R_6b42_120790d8 , 
    R_1186d_f8cbb38 , 
    R_147d3_12648e28 , 
    R_11add_1056c4d8 , 
    R_13c18_1264df68 , 
    R_13e19_132f7c08 , 
    R_b6_1265e148 , 
    R_13bb8_1265edc8 , 
    R_146a8_12050118 , 
    R_18e_12043ef8 , 
    R_181_12647a28 , 
    R_b677_12083178 , 
    R_1176f_1379f8a8 , 
    R_11d7b_102f2d88 , 
    R_145bd_1207cff8 , 
    R_13bae_105700d8 , 
    R_10fed_1330ad68 , 
    R_1479f_11cde4a8 , 
    R_71_1265e8c8 , 
    R_3ca5_102eebe8 , 
    R_14769_1056b718 , 
    R_139ba_11ce35e8 , 
    R_ccf5_13a128e8 , 
    R_13964_1207def8 , 
    R_13920_133128e8 , 
    R_13b74_11cd8dc8 , 
    R_13e6d_11cd90e8 , 
    R_13ae8_11545db8 , 
    R_e946_13796668 , 
    R_12db3_10562b18 , 
    R_7b5f_1264bc68 , 
    R_139f5_132fc348 , 
    R_cd6e_10562a78 , 
    R_13626_12077cd8 , 
    R_148dc_102f3c88 , 
    R_11db0_13302748 , 
    R_1470b_115413f8 , 
    R_fd8e_120835d8 , 
    R_142aa_102f2a68 , 
    R_1267b_1056b538 , 
    R_10df7_1264ae08 , 
    R_b753_102ebe48 , 
    R_14a47_102eeb48 , 
    R_12f94_1379c068 , 
    R_f3d0_1264e3c8 , 
    R_13cd6_10565638 , 
    R_123b1_12b3e378 , 
    R_144cf_f8c96f8 , 
    R_13d0c_102f6168 , 
    R_13c61_12081d78 , 
    R_134f6_11ce6608 , 
    R_112c2_12b294b8 , 
    R_11922_1056c898 , 
    R_11971_1207dbd8 , 
    R_138_1265b308 , 
    R_d2_12654c28 , 
    R_23d_12656088 , 
    R_8a_1379cba8 , 
    R_38ad_12048418 , 
    R_7b_12651de8 , 
    R_13889_10564918 , 
    R_13188_12079c18 , 
    R_13b8c_13a15728 , 
    R_947f_1056eaf8 , 
    R_1d7_12649648 , 
    R_149db_102f1668 , 
    R_ac1d_120826d8 , 
    R_13a06_105668f8 , 
    R_18f_132fc988 , 
    R_180_1265fea8 , 
    R_10e36_11ce6d88 , 
    R_136a7_12035cb8 , 
    R_148df_13a1d608 , 
    R_1380f_12080838 , 
    R_1485b_1265a688 , 
    R_14930_102f1a28 , 
    R_10044_102f1c08 , 
    R_d2a3_1207bbf8 , 
    R_1c0_1203c0b8 , 
    R_14f_12b25778 , 
    R_8472_126654e8 , 
    R_1483d_11ce0d48 , 
    R_12b67_11cdf3a8 , 
    R_11346_12655448 , 
    R_13893_12084d98 , 
    R_103f0_1207ecb8 , 
    R_1308d_1379eea8 , 
    R_f8ce_102f10c8 , 
    R_13f82_11543978 , 
    R_12359_133022e8 , 
    R_12cd3_13a1f728 , 
    R_13546_1153efb8 , 
    R_143b6_115408b8 , 
    R_148e5_10568518 , 
    R_10a79_11545278 , 
    R_1368d_102f3be8 , 
    R_14002_12047518 , 
    R_febc_1207caf8 , 
    R_14987_10571d98 , 
    R_14894_126569e8 , 
    R_13e23_102f1708 , 
    R_12304_10569e18 , 
    R_12daa_f8cc218 , 
    R_1289e_13316128 , 
    R_146ea_132fd6a8 , 
    R_104_12b414d8 , 
    R_e9_12055a78 , 
    R_226_12652568 , 
    R_20b_12656bc8 , 
    R_1484c_1056c078 , 
    R_149fc_12077a58 , 
    R_143f0_120442b8 , 
    R_107_1203f538 , 
    R_208_12b260d8 , 
    R_1d2_1203ce78 , 
    R_1442a_102f6668 , 
    R_13d_1379c568 , 
    R_134be_13a19148 , 
    R_145cf_13304328 , 
    R_12fa4_1153e0b8 , 
    R_1053d_12079858 , 
    R_ee_f8c86b8 , 
    R_221_12652888 , 
    R_13eb5_132f7ac8 , 
    R_190_133178e8 , 
    R_17f_115396f8 , 
    R_137af_11ce6e28 , 
    R_1455a_102ed748 , 
    R_10db8_102f74c8 , 
    R_ab_1264cde8 , 
    R_1187e_12077698 , 
    R_5a_126653a8 , 
    R_7e57_13a1a188 , 
    R_146ed_1153a238 , 
    R_1b0_12b29918 , 
    R_15f_1265f188 , 
    R_138b8_1264a368 , 
    R_13bd6_102f9188 , 
    R_14a17_102f0ee8 , 
    R_143a6_133121a8 , 
    R_11f57_12649328 , 
    R_14972_13302608 , 
    R_10701_1207f1b8 , 
    R_14503_1203e3b8 , 
    R_a4_12b36e98 , 
    R_6a_12b40178 , 
    R_aeba_105624d8 , 
    R_1379b_11ce6ec8 , 
    R_134e2_13a1e3c8 , 
    R_10973_12663008 , 
    R_11c66_102f7ba8 , 
    R_1325f_126468a8 , 
    R_1327d_10570d58 , 
    R_13417_102f3968 , 
    R_101_1264f048 , 
    R_95_133017a8 , 
    R_20e_1265e788 , 
    R_13c59_105b5638 , 
    R_13ca1_12652f68 , 
    R_1481c_11cdb988 , 
    R_14611_11545458 , 
    R_12fae_102f7388 , 
    R_1469f_1207d138 , 
    R_142dd_13314828 , 
    R_1279d_12079fd8 , 
    R_12646_1056b2b8 , 
    R_11486_102ee788 , 
    R_13389_1207fb18 , 
    R_1492d_11ce64c8 , 
    R_12d46_12648928 , 
    R_145b7_12b3d5b8 , 
    R_b211_12048c38 , 
    R_143aa_13795c68 , 
    R_1110c_11cdc928 , 
    R_1a5_12b3c618 , 
    R_16a_137a1248 , 
    R_df67_1207b8d8 , 
    R_124f6_1264f2c8 , 
    R_12b54_102f2248 , 
    R_d7dc_13a17de8 , 
    R_1247b_11ce4808 , 
    R_149ea_11540598 , 
    R_10a_12b30678 , 
    R_13c77_13a1cc08 , 
    R_205_12653dc8 , 
    R_14753_1264efa8 , 
    R_191_12043d18 , 
    R_17e_132f8568 , 
    R_11c4b_13a15c28 , 
    R_13208_11542758 , 
    R_e0ad_133021a8 , 
    R_11a3f_12b3e9b8 , 
    R_1230e_f8cb598 , 
    R_eee_1056adb8 , 
    R_14444_12648108 , 
    R_1dc_11538d98 , 
    R_12b7a_1264f188 , 
    R_133_13313888 , 
    R_147b1_105b5a98 , 
    R_f116_11ce1068 , 
    R_13a5c_1379a268 , 
    R_14340_12078458 , 
    R_e522_1330ed28 , 
    R_146f0_1153da78 , 
    R_136f4_12649148 , 
    R_119e8_1153e798 , 
    R_1391b_12b277f8 , 
    R_fd37_120394f8 , 
    R_1461d_11539dd8 , 
    R_ee50_102eb9e8 , 
    R_dd_132f61c8 , 
    R_232_105afa58 , 
    R_4c_12652b08 , 
    R_135a0_1153f0f8 , 
    R_125d0_12b3f6d8 , 
    R_b4_13302988 , 
    R_51_13309648 , 
    R_f925_12048b98 , 
    R_14034_f8cf198 , 
    R_123e9_f8c0eb8 , 
    R_14726_1203bc58 , 
    R_10894_1153ad78 , 
    R_1b9_1379b7a8 , 
    R_156_137927e8 , 
    R_1471a_1379da08 , 
    R_13d4e_11544f58 , 
    R_112ae_115429d8 , 
    R_dcb0_10564e18 , 
    R_13ae3_12083498 , 
    R_11a90_13a1ba88 , 
    R_13f1a_10566998 , 
    R_fdd5_1264d068 , 
    R_13acb_13a17988 , 
    R_ef1_13a16ee8 , 
    R_145e1_12b40d58 , 
    R_14915_102f7748 , 
    R_ed3c_120760b8 , 
    R_13cdc_11542398 , 
    R_f544_102f5d08 , 
    R_147e7_13793fa8 , 
    R_e4_133095a8 , 
    R_8d_1153d078 , 
    R_78_12044178 , 
    R_22b_12b3b538 , 
    R_128ff_105b6178 , 
    R_148ac_102f0f88 , 
    R_1e9_133208a8 , 
    R_192_12b44a98 , 
    R_17d_12661f28 , 
    R_12b83_13305e08 , 
    R_fbb3_10567078 , 
    R_126_12660588 , 
    R_cfc6_1264a868 , 
    R_1492a_13a1e1e8 , 
    R_116bb_1207d6d8 , 
    R_144d8_1330d9c8 , 
    R_e6f2_102ecc08 , 
    R_14a14_1207bdd8 , 
    R_10f70_11544a58 , 
    R_119fa_1207f2f8 , 
    R_cef5_1265b6c8 , 
    R_115b3_12082458 , 
    R_211_1265c028 , 
    R_146cc_11542618 , 
    R_fe_120448f8 , 
    R_119df_1056bad8 , 
    R_13787_11ce21e8 , 
    R_147dd_11ce6068 , 
    R_14695_11cdf8a8 , 
    R_149b1_102fa128 , 
    R_110af_1379aee8 , 
    R_14560_1330b3a8 , 
    R_143ff_11cdca68 , 
    R_d4_12654a48 , 
    R_23b_13799408 , 
    R_1c7_132fc0c8 , 
    R_148_105aacd8 , 
    R_13d6d_13a17668 , 
    R_ce64_1056f9f8 , 
    R_14474_13307a28 , 
    R_12bde_102f62a8 , 
    R_1436a_102eefa8 , 
    R_14957_11540db8 , 
    R_b634_11cdc068 , 
    R_1460e_11ce2dc8 , 
    R_f24f_11ce2fa8 , 
    R_13763_105679d8 , 
    R_f0b2_102f7f68 , 
    R_14620_11ce6108 , 
    R_131f5_12084618 , 
    R_1490f_12651e88 , 
    R_136cc_1264fcc8 , 
    R_f227_1207a398 , 
    R_13959_1153f918 , 
    R_142cf_12659aa8 , 
    R_f6b2_11cdfb28 , 
    R_1ed_1203f5d8 , 
    R_a2f6_11cdb3e8 , 
    R_fc5e_13a18888 , 
    R_122_12663d28 , 
    R_13f67_12083b78 , 
    R_13740_11cdb348 , 
    R_146c9_1153fd78 , 
    R_145db_13a12b68 , 
    R_101ae_13a1fae8 , 
    R_bb03_12b29ff8 , 
    R_1101b_12045f38 , 
    R_12bfd_10564b98 , 
    R_121a5_1056a138 , 
    R_127df_1330a728 , 
    R_11617_105656d8 , 
    R_13f90_12080518 , 
    R_13be9_12662388 , 
    R_12760_1331ab88 , 
    R_126bb_10563b58 , 
    R_147c6_12081cd8 , 
    R_21c_12b41398 , 
    R_13b33_102f0588 , 
    R_1f8_132f5fe8 , 
    R_11d2f_105665d8 , 
    R_1227d_1265f2c8 , 
    R_11a35_102f44a8 , 
    R_1479c_1056c758 , 
    R_116e4_12659828 , 
    R_14662_1207ceb8 , 
    R_14515_12079ad8 , 
    R_117_12650c68 , 
    R_115ca_11ce5fc8 , 
    R_f3_1379bde8 , 
    R_e229_102ecca8 , 
    R_202_12b3f098 , 
    R_1e5_1203a218 , 
    R_12a_1331fea8 , 
    R_10d_1330bda8 , 
    R_135d6_1056fef8 , 
    R_14918_13a1d888 , 
    R_1452a_10564378 , 
    R_14984_1056bc18 , 
    R_1cd_1265c8e8 , 
    R_eb34_11cda628 , 
    R_125ac_11ce4308 , 
    R_193_f8c7cb8 , 
    R_1216d_1264d7e8 , 
    R_17c_132fe648 , 
    R_142_13792ce8 , 
    R_cdb8_102f4f48 , 
    R_144bd_11cdeb88 , 
    R_131ae_1056bd58 , 
    R_14909_1379f768 , 
    R_14924_12b3adb8 , 
    R_102a2_12b41e38 , 
    R_13aa8_120525f8 , 
    R_d3ca_102ef7c8 , 
    R_1459f_120792b8 , 
    R_120b3_12b407b8 , 
    R_127a7_105683d8 , 
    R_14545_1056b218 , 
    R_12056_1204f178 , 
    R_11f2a_10563ab8 , 
    R_e021_12b26718 , 
    R_f377_1056d1f8 , 
    R_127ca_13a16da8 , 
    R_14689_120838f8 , 
    R_11be7_1207a6b8 , 
    R_139a1_1264c668 , 
    R_14536_12b42978 , 
    R_13c2d_11cdd828 , 
    R_14906_11544ff8 , 
    R_11a5d_132f52c8 , 
    R_ca63_1331c8e8 , 
    R_14714_102f77e8 , 
    R_14799_137933c8 , 
    R_1390f_13a14828 , 
    R_1234f_12083858 , 
    R_142c6_12081738 , 
    R_127ae_12b3ccf8 , 
    R_13590_12079a38 , 
    R_148b8_102eaa48 , 
    R_5735_137a0988 , 
    R_1a6_12038698 , 
    R_169_1203e458 , 
    R_127c1_12082638 , 
    R_1288a_137a1ec8 , 
    R_1488e_102f6708 , 
    R_113b9_1264ea08 , 
    R_1430f_11cd8fa8 , 
    R_f97f_13304dc8 , 
    R_104fa_120761f8 , 
    R_119ae_11cdfa88 , 
    R_12c78_1207ca58 , 
    R_d606_11ce46c8 , 
    R_146a5_102f90e8 , 
    R_14900_120781d8 , 
    R_1374f_13a16808 , 
    R_ff3c_11ce1f68 , 
    R_e834_10564238 , 
    R_14a5e_105aa4b8 , 
    R_13465_13316bc8 , 
    R_13d25_11540b38 , 
    R_56_13308248 , 
    R_ef7_1153e838 , 
    R_13193_102ec7a8 , 
    R_132f1_13a145a8 , 
    R_1291e_1056ee18 , 
    R_14921_105640f8 , 
    R_1371a_12083fd8 , 
    R_14837_132f32e8 , 
    R_13a37_12b3d338 , 
    R_dad2_1379c6a8 , 
    R_1495d_12b43878 , 
    R_149f3_12b27c58 , 
    R_107c6_1203f998 , 
    R_1456c_12b437d8 , 
    R_11888_13794868 , 
    R_13b62_13a13428 , 
    R_1360f_10563158 , 
    R_1b1_12657ac8 , 
    R_10844_1153e1f8 , 
    R_194_1331d4c8 , 
    R_17b_1265ea08 , 
    R_15e_126544a8 , 
    R_be25_102ec028 , 
    R_148fd_102eb768 , 
    R_14683_13a1d9c8 , 
    R_a069_12080298 , 
    R_1233a_13a143c8 , 
    R_6e_13304b48 , 
    R_1334f_1204e598 , 
    R_121e7_1207ff78 , 
    R_12bb7_102f3e68 , 
    R_12bcc_12652608 , 
    R_f783_13797b08 , 
    R_14680_12076fb8 , 
    R_13d2b_12085338 , 
    R_11bbe_1153de38 , 
    R_148e8_1264bda8 , 
    R_148fa_102f5948 , 
    R_149d8_132fc168 , 
    R_148ee_120808d8 , 
    R_148f4_11cd8468 , 
    R_ff98_12b41618 , 
    R_13bc3_102f8d28 , 
    R_12b1f_120564d8 , 
    R_c961_12080f18 , 
    R_214_12655588 , 
    R_dff5_102ed9c8 , 
    R_13d49_13a16bc8 , 
    R_fb_1379f808 , 
    R_12958_102f1848 , 
    R_12220_1379e908 , 
    R_144de_12076798 , 
    R_c6d1_10566178 , 
    R_11547_1264cc08 , 
    R_138ac_102eb128 , 
    R_12853_105b58b8 , 
    R_1f1_12655268 , 
    R_11e_12b29b98 , 
    R_13d30_1207b658 , 
    R_b2_105aa0f8 , 
    R_d5a1_105690f8 , 
    R_c700_13304788 , 
    R_a359_12662888 , 
    R_1449f_12055898 , 
    R_14587_10565ef8 , 
    R_14759_1056e378 , 
    R_1385d_1056ab38 , 
    R_1401f_132fb588 , 
    R_1245b_12658f68 , 
    R_fe3a_11cdb168 , 
    R_a47d_13a18f68 , 
    R_145ea_1056c438 , 
    R_99a4_102f5bc8 , 
    R_1491e_12661528 , 
    R_1c1_126618e8 , 
    R_b180_12039a98 , 
    R_14e_12b29e18 , 
    R_13b1f_12052c38 , 
    R_146e4_f8cb638 , 
    R_14581_10571b18 , 
    R_1354d_12040078 , 
    R_13508_120842f8 , 
    R_148d9_13a14d28 , 
    R_149c0_102ed068 , 
    R_1477e_10568fb8 , 
    R_14735_105680b8 , 
    R_13d35_11ce1108 , 
    R_4d49_102f8dc8 , 
    R_133aa_11545b38 , 
    R_14518_102f67a8 , 
    R_bf1d_1153d618 , 
    R_a9_1204d4b8 , 
    R_14702_12b3d0b8 , 
    R_1431c_11cde188 , 
    R_9323_1331d068 , 
    R_14a2f_12075ed8 , 
    R_1e1_13321ca8 , 
    R_12e_105af9b8 , 
    R_9d_1379c9c8 , 
    R_12caa_126508a8 , 
    R_115df_10566c18 , 
    R_144fd_102f1b68 , 
    R_127f1_12b2a098 , 
    R_137eb_12082138 , 
    R_11b9a_12b3f278 , 
    R_1483a_12081f58 , 
    R_7d2b_11ce4948 , 
    R_13a49_102f8e68 , 
    R_1493c_11cdc568 , 
    R_14a3e_102ed428 , 
    R_195_12045cb8 , 
    R_14489_12b3fe58 , 
    R_17a_1330dc48 , 
    R_1066b_1264a228 , 
    R_139b5_11536318 , 
    R_12775_126513e8 , 
    R_13d43_13a1c168 , 
    R_13e78_1056a598 , 
    R_90_f8cccb8 , 
    R_75_12b443b8 , 
    R_14816_10565db8 , 
    R_e4c7_10571398 , 
    R_14354_13317348 , 
    R_146c3_12b3bfd8 , 
    R_db95_12b2ff98 , 
    R_b45b_11ce7508 , 
    R_145de_1056b5d8 , 
    R_13c7d_1056d798 , 
    R_c7c0_102ed4c8 , 
    R_1ff_13315c28 , 
    R_1361a_102f01c8 , 
    R_110_1204b938 , 
    R_10c17_13a13888 , 
    R_d6_1264b1c8 , 
    R_239_12b2a958 , 
    R_144a8_115369f8 , 
    R_12516_13305188 , 
    R_14699_10567e38 , 
    R_12de4_12045b18 , 
    R_10fd9_11ce1928 , 
    R_145c6_13a1cb68 , 
    R_147c3_13a177a8 , 
    R_1313e_1207a1b8 , 
    R_e9a6_1153dcf8 , 
    R_123a6_12077418 , 
    R_e669_1056eb98 , 
    R_eea5_13793c88 , 
    R_8e12_f8c7538 , 
    R_11a2c_12b3f1d8 , 
    R_bc89_12664548 , 
    R_b132_13300a88 , 
    R_14626_102f4ae8 , 
    R_125c9_11ce5c08 , 
    R_14891_1265e0a8 , 
    R_13ba9_1056f4f8 , 
    R_11299_1056a4f8 , 
    R_1395f_1207ba18 , 
    R_1085f_13312a28 , 
    R_c642_12b41b18 , 
    R_1445c_f8ce478 , 
    R_14981_12b3f598 , 
    R_148e2_12650b28 , 
    R_988f_13a1e968 , 
    R_962b_105647d8 , 
    R_124a7_12079498 , 
    R_fe64_1153f378 , 
    R_11f16_102eb088 , 
    R_13e03_1379bf28 , 
    R_14927_11cdf808 , 
    R_1ba_1330eb48 , 
    R_14471_13793be8 , 
    R_121fd_11ce3048 , 
    R_14499_1207a9d8 , 
    R_155_12b43f58 , 
    R_98_12048af8 , 
    R_e916_105699b8 , 
    R_e1ea_1056b998 , 
    R_11af3_13793788 , 
    R_13bcf_12650948 , 
    R_10070_12077e18 , 
    R_f2f6_126613e8 , 
    R_104a3_11542d98 , 
    R_149ae_10565138 , 
    R_1430b_1204c8d8 , 
    R_ede8_1056dfb8 , 
    R_13495_13a1e008 , 
    R_df_132f6808 , 
    R_230_12664a48 , 
    R_136ac_102eacc8 , 
    R_dd20_137974c8 , 
    R_14741_132f2c08 , 
    R_137c1_11543dd8 , 
    R_14364_11ce6568 , 
    R_11d60_132fc8e8 , 
    R_14a44_105b60d8 , 
    R_13749_11543518 , 
    R_854a_1207fed8 , 
    R_14a11_12045a78 , 
    R_1a7_12659b48 , 
    R_168_105b3158 , 
    R_f03_13a17208 , 
    R_1274c_12653fa8 , 
    R_147b7_12079df8 , 
    R_a2_1379e228 , 
    R_63_f8c7b78 , 
    R_13c49_102ecac8 , 
    R_d68f_12078a98 , 
    R_148f1_11cde688 , 
    R_196_11536778 , 
    R_179_13301c08 , 
    R_11c1b_120757f8 , 
    R_1181a_10565098 , 
    R_14912_13300628 , 
    R_10c93_13310768 , 
    R_147f2_10571618 , 
    R_c832_12075f78 , 
    R_14530_11540778 , 
    R_e8ba_11ce3b88 , 
    R_14903_11ce50c8 , 
    R_14629_115412b8 , 
    R_11966_10562118 , 
    R_f8fa_105b4d78 , 
    R_1d8_1331f5e8 , 
    R_1281b_1207f6b8 , 
    R_137_1331a7c8 , 
    R_5f_12b428d8 , 
    R_12288_126495a8 , 
    R_a469_13a14648 , 
    R_130cc_13a17348 , 
    R_136e6_11cdcb08 , 
    R_d806_102f5a88 , 
    R_fd98_12052d78 , 
    R_144b4_1153eab8 , 
    R_1482b_12b3b3f8 , 
    R_13858_12081e18 , 
    R_1d3_1265ae08 , 
    R_13c_1265b1c8 , 
    R_14596_12048558 , 
    R_eb_1153bf98 , 
    R_224_12b29698 , 
    R_13d3c_132f70c8 , 
    R_c353_102f31e8 , 
    R_1092e_13a140a8 , 
    R_1018e_10563478 , 
    R_12875_1153eb58 , 
    R_13693_13795448 , 
    R_123bb_11ce7008 , 
    R_dfc9_12647208 , 
    R_da6d_12082098 , 
    R_1198e_1153d758 , 
    R_149ff_1264c848 , 
    R_1180e_12648248 , 
    R_12535_126604e8 , 
    R_12780_10568b58 , 
    R_9dc0_102f6f28 , 
    R_c4a7_1330a908 , 
    R_11bfb_12649968 , 
    R_13fe4_105622f8 , 
    R_12e0c_13797388 , 
    R_1454e_11ce1c48 , 
    R_14069_1153db18 , 
    R_10c0e_120464d8 , 
    R_13c1f_f8c8938 , 
    R_d910_1056e418 , 
    R_cfae_13a15368 , 
    R_10806_1264d608 , 
    R_13706_13319b48 , 
    R_12e21_1330cb68 , 
    R_f8_12665808 , 
    R_67_105aac38 , 
    R_217_105b3fb8 , 
    R_12a8e_1264ef08 , 
    R_e5ea_115436f8 , 
    R_14858_10571c58 , 
    R_111b8_102ebbc8 , 
    R_12ba4_12b28ab8 , 
    R_108f1_102f35a8 , 
    R_138a5_1264e468 , 
    R_131ff_13a1eaa8 , 
    R_11448_11ce41c8 , 
    R_11534_13a13ce8 , 
    R_12d1d_1207c238 , 
    R_134e8_13a1e8c8 , 
    R_b82e_1153c2b8 , 
    R_11572_11ce43a8 , 
    R_14897_1265c988 , 
    R_125fa_1265b128 , 
    R_b95d_102f8008 , 
    R_14436_10570718 , 
    R_f951_132fcde8 , 
    R_10246_1056ae58 , 
    R_12041_11ce0ac8 , 
    R_138cd_1153e018 , 
    R_1b2_12660f88 , 
    R_197_1379a768 , 
    R_121dd_12659328 , 
    R_178_12658d88 , 
    R_15d_133195a8 , 
    R_13f24_13318428 , 
    R_146f6_132fbc68 , 
    R_b880_12083d58 , 
    R_12ab4_132f57c8 , 
    R_ed14_133110c8 , 
    R_144f0_132ff0e8 , 
    R_10aa5_12053f98 , 
    R_1290a_11ce1388 , 
    R_9d4e_11cddbe8 , 
    R_e6_12b344f8 , 
    R_b0_12b3f458 , 
    R_229_126659e8 , 
    R_12b3f_105b6538 , 
    R_1f5_1203e958 , 
    R_f624_1265b808 , 
    R_14711_11ce2828 , 
    R_fe05_102f9548 , 
    R_1118b_11cdb8e8 , 
    R_1c8_f8c6b38 , 
    R_147_12b38c98 , 
    R_11a_1204b438 , 
    R_14778_13a1f688 , 
    R_137fd_11544418 , 
    R_f0_13795d08 , 
    R_c3_132ff188 , 
    R_21f_1265a2c8 , 
    R_12e60_132f3a68 , 
    R_4a02_12646e48 , 
    R_c5_12657e88 , 
    R_132ae_1056ef58 , 
    R_d400_133126a8 , 
    R_128a8_f8c9978 , 
    R_ecbd_12040a78 , 
    R_146ba_11cd8c88 , 
    R_ea59_102f5088 , 
    R_1183a_1204a498 , 
    R_13d1f_1207ddb8 , 
    R_136e0_11ce7148 , 
    R_ddb7_12078b38 , 
    R_14575_13307c08 , 
    R_14864_13a1b768 , 
    R_1471d_12040bb8 , 
    R_11237_1056f958 , 
    R_13fee_12663288 , 
    R_c1_1204fd58 , 
    R_14632_11cd85a8 , 
    R_4d_12662d88 , 
    R_b895_1264a4a8 , 
    R_11b87_12648b08 , 
    R_111c4_12076658 , 
    R_a534_12b3d018 , 
    R_11805_12b41578 , 
    R_c901_126603a8 , 
    R_13bde_13a1bbc8 , 
    R_149b4_10564d78 , 
    R_c7_126589c8 , 
    R_248_1331ef08 , 
    R_5b_12655088 , 
    R_13720_102f3f08 , 
    R_b9b1_1056c9d8 , 
    R_f1cc_10567ed8 , 
    R_cd0b_11542f78 , 
    R_1497b_11cdfda8 , 
    R_12d6f_13799b88 , 
    R_14305_120844d8 , 
    R_145ae_102efe08 , 
    R_147d6_12b27b18 , 
    R_13dc3_11cdbf28 , 
    R_dc22_1153d438 , 
    R_5970_11cdbe88 , 
    R_113_1265c528 , 
    R_82_f8cbc78 , 
    R_1fc_12050078 , 
    R_b00a_1153e658 , 
    R_1346e_10567bb8 , 
    R_1dd_12b395f8 , 
    R_10390_1207ed58 , 
    R_12cf4_13310ee8 , 
    R_10675_1203cab8 , 
    R_1399b_1264c3e8 , 
    R_132_120518d8 , 
    R_d8_12b3c938 , 
    R_237_105a9fb8 , 
    R_d4b2_1265bda8 , 
    R_14453_12649d28 , 
    R_10e2c_102ecde8 , 
    R_52_13799868 , 
    R_143dc_120824f8 , 
    R_13ebe_11ce4128 , 
    R_14053_102f21a8 , 
    R_10960_133050e8 , 
    R_1037b_1264a048 , 
    R_7fe6_12b3f638 , 
    R_12685_11cdf088 , 
    R_135e9_11ce0de8 , 
    R_bf_1379fa88 , 
    R_85_12b41898 , 
    R_149d5_11541358 , 
    R_13f4d_10561fd8 , 
    R_d0f1_1056a1d8 , 
    R_a3f3_12646da8 , 
    R_1311d_13a131a8 , 
    R_1026e_11541ad8 , 
    R_139de_13310588 , 
    R_144cc_11ce23c8 , 
    R_1403a_1331cc08 , 
    R_1ce_12656628 , 
    R_198_12b3fdb8 , 
    R_d37f_1379a1c8 , 
    R_177_1330de28 , 
    R_141_12b3cf78 , 
    R_14500_102f92c8 , 
    R_c9_12b28fb8 , 
    R_246_1203df58 , 
    R_93_12659be8 , 
    R_72_132fe788 , 
    R_125bf_105685b8 , 
    R_1a8_137a0d48 , 
    R_147a5_1264a728 , 
    R_167_1204f678 , 
    R_7f_105ac998 , 
    R_149f0_13a1fea8 , 
    R_12210_13793aa8 , 
    R_13db7_11ce11a8 , 
    R_100e9_132f3ec8 , 
    R_5362_13a18108 , 
    R_124d7_13a18e28 , 
    R_14a55_133001c8 , 
    R_12419_1153d398 , 
    R_108b6_1264e0a8 , 
    R_10d4d_11cded68 , 
    R_1464a_13a15b88 , 
    R_c7f2_11cdc748 , 
    R_13c83_11544698 , 
    R_1489a_f8c6c78 , 
    R_125b6_12040b18 , 
    R_c00b_12079718 , 
    R_eeb_13a13608 , 
    R_f088_1330ba88 , 
    R_1365e_1207b838 , 
    R_fa81_12052198 , 
    R_145f3_13a14788 , 
    R_10995_102f3148 , 
    R_123f8_13a13388 , 
    R_6358_1204fe98 , 
    R_14763_11ce4c68 , 
    R_1433c_12077c38 , 
    R_dde7_13a141e8 , 
    R_13ef9_1204a858 , 
    R_14810_1056db58 , 
    R_13fdc_102f15c8 , 
    R_d995_11ce0fc8 , 
    R_117fc_12056078 , 
    R_8d57_11ce53e8 , 
    R_11bb4_12b39cd8 , 
    R_13b97_1207a438 , 
    R_14068_11cdc108 , 
    R_1335a_105b5ef8 , 
    R_1043d_13a1c5c8 , 
    R_128cf_11cdabc8 , 
    R_1219b_1207a938 , 
    R_10dce_105631f8 , 
    R_bbfa_10564418 , 
    R_11864_12b44318 , 
    R_12435_11ce4088 , 
    R_a7_1265a5e8 , 
    R_111f4_11cdf6c8 , 
    R_135cf_1207eb78 , 
    R_102ef_1153c218 , 
    R_12ca0_11ce0668 , 
    R_1c2_1330f228 , 
    R_c6f4_12056438 , 
    R_1404f_12b3e738 , 
    R_ee7b_1379a628 , 
    R_127e9_f8c8078 , 
    R_14d_1203cbf8 , 
    R_bd_1203f3f8 , 
    R_48_13301848 , 
    R_10afa_13a15d68 , 
    R_ed66_11ce3368 , 
    R_13a92_102f0bc8 , 
    R_e9fb_12646268 , 
    R_10d30_12084078 , 
    R_149ab_1153d7f8 , 
    R_88_13300d08 , 
    R_6b_105aaff8 , 
    R_11c31_115418f8 , 
    R_13677_102f9868 , 
    R_133f2_1379f088 , 
    R_13edf_120837b8 , 
    R_d399_137980a8 , 
    R_1446e_1207d958 , 
    R_1382d_1207d9f8 , 
    R_cb_1331fa48 , 
    R_244_1264c708 , 
    R_12dc8_13a1f548 , 
    R_12299_1265d1a8 , 
    R_1474a_12076dd8 , 
    R_13844_12663aa8 , 
    R_13c11_1153d578 , 
    R_14650_1056f278 , 
    R_146fc_12647848 , 
    R_10f84_1207bab8 , 
    R_131cc_12b272f8 , 
    R_1451b_10567cf8 , 
    R_14390_10567c58 , 
    R_13754_12082318 , 
    R_1bb_12664868 , 
    R_154_1204e1d8 , 
    R_14831_1264f408 , 
    R_7c_105b1cb8 , 
    R_f1a0_12075938 , 
    R_e9d0_1153f558 , 
    R_f0eb_102f7568 , 
    R_fb0c_1331a368 , 
    R_1397b_1331b268 , 
    R_e589_1379bb68 , 
    R_1381a_120547b8 , 
    R_1463e_105703f8 , 
    R_12e76_11cd9908 , 
    R_199_132fb3a8 , 
    R_176_12b265d8 , 
    R_125_13798008 , 
    R_11ad2_102ed108 , 
    R_1ea_1265a868 , 
    R_10764_11cd9548 , 
    R_14563_1264d6a8 , 
    R_12c1a_102f0268 , 
    R_146d2_1203a998 , 
    R_147bd_102f9048 , 
    R_fa57_1207f398 , 
    R_c5a3_120849d8 , 
    R_11dc9_f8c9b58 , 
    R_11d95_1153f198 , 
    R_1329b_11cd95e8 , 
    R_14861_f8c41f8 , 
    R_1064a_10561f38 , 
    R_ce07_f8c8f78 , 
    R_14720_11ce07a8 , 
    R_13ca7_12078098 , 
    R_147f5_1207a078 , 
    R_142d3_12036758 , 
    R_13dee_12083a38 , 
    R_ec91_126490a8 , 
    R_13421_11544c38 , 
    R_cf92_11cdfee8 , 
    R_4c49_13a1d748 , 
    R_114d1_13307de8 , 
    R_cff7_12076bf8 , 
    R_142ff_11ce1b08 , 
    R_139c0_13a1e5a8 , 
    R_143cc_1056e738 , 
    R_ba4e_13a1d388 , 
    R_12485_105b6358 , 
    R_11f0c_13a1aea8 , 
    R_14867_12054b78 , 
    R_137b5_10569cd8 , 
    R_11d1b_12649288 , 
    R_13d7b_102f56c8 , 
    R_14a2c_102f12a8 , 
    R_14608_13a155e8 , 
    R_144c9_10571578 , 
    R_fc0a_11541858 , 
    R_144fa_120775f8 , 
    R_129_1331c988 , 
    R_13561_1330d068 , 
    R_e1_12661708 , 
    R_1299a_1207b158 , 
    R_1489d_105686f8 , 
    R_22e_132f2ac8 , 
    R_6d01_102f72e8 , 
    R_ffc3_12656e48 , 
    R_1496f_102f9908 , 
    R_1e6_13792a68 , 
    R_14760_11ce3868 , 
    R_d2d1_13793468 , 
    R_12145_1207b978 , 
    R_f5_11537038 , 
    R_bb_13799cc8 , 
    R_21a_1265b088 , 
    R_14975_11541998 , 
    R_147c0_11ce20a8 , 
    R_13b7f_1153a198 , 
    R_13615_12084c58 , 
    R_14a29_10571438 , 
    R_13526_102f49a8 , 
    R_11215_12075b18 , 
    R_10e4c_13a169e8 , 
    R_13d97_105651d8 , 
    R_1b3_1379b348 , 
    R_13fab_11538758 , 
    R_10ff9_105aad78 , 
    R_145c0_11cd7f68 , 
    R_145fc_120476f8 , 
    R_15c_137992c8 , 
    R_67bc_13311028 , 
    R_efc2_11cdefe8 , 
    R_145cc_132f8388 , 
    R_ae_1379c1a8 , 
    R_1263c_11cdf768 , 
    R_57_126522e8 , 
    R_14659_1264e1e8 , 
    R_13899_133075c8 , 
    R_125e5_13311348 , 
    R_113fb_11ce7288 , 
    R_11e0e_102f4908 , 
    R_11270_12b29a58 , 
    R_f61a_13305cc8 , 
    R_1499f_133198c8 , 
    R_121_13795808 , 
    R_106_12b25a98 , 
    R_1458a_102eb268 , 
    R_126cf_13a19788 , 
    R_209_1379cb08 , 
    R_1ee_12656268 , 
    R_12c5a_102ef688 , 
    R_1270e_11cdb708 , 
    R_e437_102f2c48 , 
    R_147cf_11ce5168 , 
    R_e233_1056d338 , 
    R_13bbe_11ce55c8 , 
    R_11e6b_1207d458 , 
    R_13f0b_12b42f18 , 
    R_103_12b41c58 , 
    R_cd_12b39a58 , 
    R_242_12654688 , 
    R_20c_12b43c38 , 
    R_11ce5_1379e048 , 
    R_ef4_1056dc98 , 
    R_11823_13a15fe8 , 
    R_130b8_13a12988 , 
    R_12baf_12648ba8 , 
    R_119a4_102f3288 , 
    R_f4e5_1264b308 , 
    R_12c6f_11cdea48 , 
    R_1473b_102fa308 , 
    R_8b_132f8608 , 
    R_11467_105659f8 , 
    R_11b4a_11ce1568 , 
    R_137f7_12077878 , 
    R_e5b5_1153d938 , 
    R_14775_13a1bda8 , 
    R_14671_1264ab88 , 
    R_14066_12084258 , 
    R_13954_12076518 , 
    R_de4d_12b26538 , 
    R_149f6_11cda308 , 
    R_aff6_102f4a48 , 
    R_d75d_1207c0f8 , 
    R_10f46_12081ff8 , 
    R_c50b_11cdd3c8 , 
    R_136ed_12082ef8 , 
    R_101d1_1056e198 , 
    R_1a9_12037658 , 
    R_166_120507f8 , 
    R_9b_12b3b178 , 
    R_bb16_12650268 , 
    R_1265a_105635b8 , 
    R_b802_1265dba8 , 
    R_131ea_102f4cc8 , 
    R_14a0e_10570e98 , 
    R_19a_12662068 , 
    R_175_12b3fc78 , 
    R_109_12b2c7f8 , 
    R_206_105b5b38 , 
    R_146b4_1153fcd8 , 
    R_11e21_11cd9e08 , 
    R_104ba_f8c7218 , 
    R_13fbc_11541218 , 
    R_144ba_102f8c88 , 
    R_11622_102ed388 , 
    R_13c02_12b29198 , 
    R_13ba3_105626b8 , 
    R_ff0f_12081918 , 
    R_123d6_11541e98 , 
    R_fd64_102f3328 , 
    R_14486_102ef728 , 
    R_13776_1379fd08 , 
    R_14665_132f5ae8 , 
    R_10098_13793968 , 
    R_11072_13a1ed28 , 
    R_14554_10565778 , 
    R_137a8_1056b678 , 
    R_11b55_12649a08 , 
    R_14411_12663508 , 
    R_84a7_12b40fd8 , 
    R_133fc_1153ee78 , 
    R_da_1331b088 , 
    R_a0_1379b2a8 , 
    R_235_1264d4c8 , 
    R_1333b_11542c58 , 
    R_132e7_11ce28c8 , 
    R_1357d_1153feb8 , 
    R_14644_1056d978 , 
    R_100_1265f0e8 , 
    R_79_137a1388 , 
    R_e0d7_126556c8 , 
    R_11b42_1264b6c8 , 
    R_20f_12b28018 , 
    R_f4db_1207bfb8 , 
    R_1193e_13a19968 , 
    R_138d5_1379b848 , 
    R_13e4c_1207f118 , 
    R_13a7e_102f6ac8 , 
    R_12d79_102ee468 , 
    R_116a8_12084398 , 
    R_116_1265f868 , 
    R_148a3_11cdecc8 , 
    R_13273_13a1a688 , 
    R_1f9_1379ddc8 , 
    R_1025b_1330bee8 , 
    R_122e8_12b39878 , 
    R_11ba2_11544738 , 
    R_12521_1056c258 , 
    R_e8e6_f8cf4b8 , 
    R_8cd2_1264ac28 , 
    R_11a11_126477a8 , 
    R_143c6_120850b8 , 
    R_13e99_12039e58 , 
    R_1466b_13306808 , 
    R_14465_1207a758 , 
    R_134b3_102f3468 , 
    R_11fe7_1330c3e8 , 
    R_1258d_13a14dc8 , 
    R_14677_105712f8 , 
    R_1367d_102eb628 , 
    R_1e2_12663c88 , 
    R_b9_12661848 , 
    R_12d_12660268 , 
    R_f47c_1153ded8 , 
    R_1468c_13a1aae8 , 
    R_145ba_120815f8 , 
    R_14790_11cd9cc8 , 
    R_14419_12048f58 , 
    R_13bb3_1207b6f8 , 
    R_1046b_105688d8 , 
    R_1232e_13314008 , 
    R_1170d_1264c528 , 
    R_14a41_1056fa98 , 
    R_14459_11cd92c8 , 
    R_14480_11cdcf68 , 
    R_13a88_11ce3f48 , 
    R_c8f0_102f0d08 , 
    R_134ff_1056bf38 , 
    R_aac5_13a18748 , 
    R_14509_13a1e148 , 
    R_cebc_12039d18 , 
    R_135bd_12081058 , 
    R_147ba_12078ef8 , 
    R_f4a6_105654f8 , 
    R_1182e_13a19aa8 , 
    R_142eb_11cdec28 , 
    R_13bf5_10568ab8 , 
    R_12093_12077058 , 
    R_13dac_13a15688 , 
    R_dc51_13304f08 , 
    R_13e8f_1264a0e8 , 
    R_13c89_12b39f58 , 
    R_f0be_102f1de8 , 
    R_9373_10563e78 , 
    R_11a48_13a195a8 , 
    R_f3f9_1153f9b8 , 
    R_1d4_12b42fb8 , 
    R_e3f1_12b25bd8 , 
    R_13c27_13309b48 , 
    R_240_105ab4f8 , 
    R_cf_13311a28 , 
    R_13c38_1204a3f8 , 
    R_13b_13300f88 , 
    R_11ef6_11cd7888 , 
    R_135c9_11ce6888 , 
    R_116d1_1153d898 , 
    R_149d2_12080158 , 
    R_ba5b_12b403f8 , 
    R_ea84_1330ca28 , 
    R_f59a_11ce3908 , 
    R_1496c_1331e968 , 
    R_12bd5_11ce3fe8 , 
    R_1253e_105b6678 , 
    R_14873_11cd79c8 , 
    R_149a5_132ff868 , 
    R_14512_11540bd8 , 
    R_14756_10565318 , 
    R_1c9_13313a68 , 
    R_d09b_12660948 , 
    R_203_12050cf8 , 
    R_10c_12038058 , 
    R_146_12b42298 , 
    R_136c1_12b276b8 , 
    R_1480a_12649e68 , 
    R_1d9_1379e7c8 , 
    R_13e84_1056ad18 , 
    R_1021c_1056fc78 , 
    R_136_132fe6e8 , 
    R_145ff_102ef2c8 , 
    R_19b_12b28dd8 , 
    R_1031a_11540e58 , 
    R_1f2_11538438 , 
    R_13114_102f3648 , 
    R_ec36_12042af8 , 
    R_222_133189c8 , 
    R_6f_12b3a458 , 
    R_96_1203c838 , 
    R_ed_1203deb8 , 
    R_11d_1204c838 , 
    R_174_13318928 , 
    R_119f1_13316588 , 
    R_1486a_13a1d428 , 
    R_11717_1207d778 , 
    R_14781_115447d8 , 
    R_13995_12038738 , 
    R_e4f5_12049598 , 
    R_74a9_12645d68 , 
    R_10208_12038558 , 
    R_145ab_12b3f9f8 , 
    R_227_1331e508 , 
    R_e8_133028e8 , 
    R_13809_1153faf8 , 
    R_f732_12649008 , 
    R_14524_137968e8 , 
    R_146d8_11cd94a8 , 
    R_14064_1264d2e8 , 
    R_12dfa_11cd88c8 , 
    R_135ef_102f0a88 , 
    R_10ee5_12047798 , 
    R_14548_120493b8 , 
    R_11030_11cdbca8 , 
    R_1400f_13a1a368 , 
    R_f051_1264e6e8 , 
    R_de7c_102eafe8 , 
    R_13538_120754d8 , 
    R_13e56_12b297d8 , 
    R_84eb_1331c2a8 , 
    R_1498a_1207e3f8 , 
    R_148a6_115459f8 , 
    R_212_1330bd08 , 
    R_fd_13307d48 , 
    R_144a5_13a1c028 , 
    R_10110_120369d8 , 
    R_12b5e_12651208 , 
    R_149ed_13303428 , 
    R_144db_12078598 , 
    R_bf9f_11cd9b88 , 
    R_14017_f8c20d8 , 
    R_13a3d_f8ca918 , 
    R_13b2d_120830d8 , 
    R_8e_132f37e8 , 
    R_12aeb_120810f8 , 
    R_a23e_11ce5ca8 , 
    R_12ce9_12081c38 , 
    R_f00_1207c058 , 
    R_c1fe_1264be48 , 
    R_f2d2_11cdf948 , 
    R_14385_12044c18 , 
    R_143c0_1265fb88 , 
    R_14496_13a1c668 , 
    R_14738_12b28bf8 , 
    R_cab9_102f99a8 , 
    R_1255c_f8c61d8 , 
    R_143ba_11cde868 , 
    R_147c9_13a18ce8 , 
    R_13311_13a198c8 , 
    R_147a2_102f2ce8 , 
    R_fbe0_13a1b628 , 
    R_dcc6_12664ae8 , 
    R_103cf_12085158 , 
    R_13909_1204f5d8 , 
    R_1197b_115433d8 , 
    R_144e1_13a1f4a8 , 
    R_145a2_11cd7ce8 , 
    R_12d50_120851f8 , 
    R_12380_10563338 , 
    R_107a7_1379f9e8 , 
    R_10e8a_102ea688 , 
    R_122fb_13a17708 , 
    R_12aa7_12037798 , 
    R_12107_1264d428 , 
    R_14533_1330c8e8 , 
    R_14542_120759d8 , 
    R_4276_102effe8 , 
    R_1478d_115453b8 , 
    R_130c1_11542258 , 
    R_13ff8_102f9fe8 , 
    R_1aa_13795268 , 
    R_116b1_13a159a8 , 
    R_1bc_126536e8 , 
    R_b76e_1153c8f8 , 
    R_4e_13792e28 , 
    R_60_12b44bd8 , 
    R_a5_13311668 , 
    R_b7_1379f948 , 
    R_153_13793288 , 
    R_165_13306948 , 
    R_f9fe_102f9408 , 
    R_14431_12080478 , 
    R_1c3_12047158 , 
    R_64_f8c1bd8 , 
    R_14c_120387d8 , 
    R_12471_102f7068 , 
    R_148c1_13316f88 , 
    R_11433_1265f048 , 
    R_13ce2_1264aa48 , 
    R_121bd_115449b8 , 
    R_14813_10566d58 , 
    R_147fb_102f83c8 , 
    R_146ab_12051658 , 
    R_12c65_1264cb68 , 
    R_e2b4_f8c0f58 , 
    R_10c61_120805b8 , 
    R_10f1d_10566df8 , 
    R_10de4_1379b5c8 , 
    R_ae51_105ab098 , 
    R_146f3_12659d28 , 
    R_d03f_126484c8 , 
    R_9fe2_11543fb8 , 
    R_10b79_12657028 , 
    R_64c2_12662748 , 
    R_139d0_102f1fc8 , 
    R_13639_1207f578 , 
    R_1b4_12654728 , 
    R_1cf_133184c8 , 
    R_e214_1207ae38 , 
    R_140_12665448 , 
    R_15b_f8c0378 , 
    R_1435c_13304d28 , 
    R_10745_12056898 , 
    R_1044f_120557f8 , 
    R_10824_11ce3188 , 
    R_13820_12b41438 , 
    R_69b8_11cdc888 , 
    R_124b9_1056d658 , 
    R_143f4_102edd88 , 
    R_142f5_1264a908 , 
    R_76_f8ca198 , 
    R_ac_12660a88 , 
    R_1269b_11cd9368 , 
    R_147b4_120766f8 , 
    R_14834_13a16a88 , 
    R_12e88_102f8a08 , 
    R_f021_102ec168 , 
    R_f6dd_13a163a8 , 
    R_145e4_126463a8 , 
    R_14723_1264db08 , 
    R_173_f8c3438 , 
    R_19c_12b40218 , 
    R_11142_10562f78 , 
    R_23e_1265bc68 , 
    R_d1_13311f28 , 
    R_13512_12080dd8 , 
    R_7859_11cdaee8 , 
    R_14593_115458b8 , 
    R_148a9_12647ac8 , 
    R_10577_11545318 , 
    R_133ca_1203e098 , 
    R_13b92_13a14be8 , 
    R_10efd_102ec3e8 , 
    R_f0b_1153f4b8 , 
    R_12e15_10568018 , 
    R_200_12b29eb8 , 
    R_21d_137a03e8 , 
    R_f2_12652ec8 , 
    R_10f_12b3e5f8 , 
    R_ca13_11ce4628 , 
    R_14966_11546218 , 
    R_13ad8_1203a358 , 
    R_12d8d_105b5db8 , 
    R_10165_1264cac8 , 
    R_1337f_13a12c08 , 
    R_53_f8c2a38 , 
    R_149c9_132f4fa8 , 
    R_10aae_1207c558 , 
    R_13aad_11541a38 , 
    R_12362_10563dd8 , 
    R_5c4e_1056ced8 , 
    R_130f5_1056a098 , 
    R_12a7c_11cdde68 , 
    R_14415_12b2a318 , 
    R_1488b_13a189c8 , 
    R_14062_1204cf18 , 
    R_14784_11cd8508 , 
    R_1032f_10570f38 , 
    R_9bdf_102ee5a8 , 
    R_13bf0_1331c528 , 
    R_11b90_11ce0208 , 
    R_149cf_13a17b68 , 
    R_12021_11ce25a8 , 
    R_1de_12056d98 , 
    R_49_1331f4a8 , 
    R_131_105ab3b8 , 
    R_1462f_13794688 , 
    R_10628_1203d2d8 , 
    R_122bf_10570038 , 
    R_11387_11540d18 , 
    R_11fa6_13306308 , 
    R_85b5_120819b8 , 
    R_142ef_102eec88 , 
    R_1434c_102f13e8 , 
    R_22c_1379b708 , 
    R_5c_137944a8 , 
    R_e3_1203e778 , 
    R_b948_1153a5f8 , 
    R_e169_11cd7a68 , 
    R_d051_11536ef8 , 
    R_10e01_120551b8 , 
    R_233_12b392d8 , 
    R_68_12b283d8 , 
    R_dc_13300768 , 
    R_13bfb_13316a88 , 
    R_10ad6_10565598 , 
    R_14870_10570538 , 
    R_12260_13a1b268 , 
    R_d661_1265cfc8 , 
    R_14572_11cd9d68 , 
    R_130ff_12078318 , 
    R_a98a_11cdaf88 , 
    R_14978_12b321f8 , 
    R_14a1a_115445f8 , 
    R_14a26_13792568 , 
    R_b327_12648568 , 
    R_108fb_105b5e58 , 
    R_1440d_11544238 , 
    R_10cff_13a1dc48 , 
    R_139ae_11cd8b48 , 
    R_14338_11cda808 , 
    R_106b3_13a16088 , 
    R_c4f8_11ce12e8 , 
    R_215_1265b948 , 
    R_fa_133070c8 , 
    R_11b68_1264ec88 , 
    R_129b1_1056f098 , 
    R_13670_10564558 , 
    R_1439c_11cdd148 , 
    R_107e6_11cdbc08 , 
    R_f279_13a1acc8 , 
    R_12ed9_102edf68 , 
    R_12bc1_13a1f048 , 
    R_13b19_12b2ba38 , 
    R_e361_120812d8 , 
    R_bef9_11ce0528 , 
    R_13ce8_120793f8 , 
    R_a235_12084a78 , 
    R_14521_1264f228 , 
    R_13cad_13a1edc8 , 
    R_148af_11540098 , 
    R_10968_13304968 , 
    R_13fcb_102f0c68 , 
    R_11645_13304e68 , 
    R_bf09_1056b498 , 
    R_12553_13310308 , 
    R_145d5_132fa228 , 
    R_146a2_1207bf18 , 
    R_136fc_12076018 , 
    R_149a2_1264d1a8 , 
    R_12b9a_13a14968 , 
    R_137cc_10569af8 , 
    R_c5ef_12081238 , 
    R_1184d_11cd9188 , 
    R_13c8f_102ed568 , 
    R_109bf_1379c248 , 
    R_14326_13301528 , 
    R_11123_12045258 , 
    R_e197_11ce3228 , 
    R_172_126656c8 , 
    R_19d_132ffb88 , 
    R_c306_f8c5418 , 
    R_b5_133157c8 , 
    R_13902_13799ae8 , 
    R_14348_1056c398 , 
    R_1457b_102f5628 , 
    R_14766_105674d8 , 
    R_d2c1_12036e38 , 
    R_1f6_1330dce8 , 
    R_10c28_12080e78 , 
    R_119_133166c8 , 
    R_1300e_12646bc8 , 
    R_13129_10567b18 , 
    R_1394d_1056f318 , 
    R_14846_13798b48 , 
    R_146cf_1379e868 , 
    R_10019_11542118 , 
    R_fb35_132fb4e8 , 
    R_11a23_126506c8 , 
    R_9aae_1056dbf8 , 
    R_14468_1264aea8 , 
    R_7aaf_f8c22b8 , 
    R_b5af_1264e508 , 
    R_13f11_11cd7b08 , 
    R_e6c6_12075cf8 , 
    R_14374_102f0768 , 
    R_14605_13a182e8 , 
    R_13de4_102f94a8 , 
    R_102c2_1264ed28 , 
    R_91_13799548 , 
    R_135f5_11cda4e8 , 
    R_14807_1331e288 , 
    R_14a08_11cdc388 , 
    R_cb44_12b3ee18 , 
    R_13a63_11544198 , 
    R_109ca_1264cd48 , 
    R_12e41_10569198 , 
    R_e46a_13a181a8 , 
    R_12963_13a1afe8 , 
    R_14a5a_12b42158 , 
    R_13e38_1207efd8 , 
    R_144ea_1264f5e8 , 
    R_11668_137a1d88 , 
    R_13ec7_11540318 , 
    R_ff67_13799688 , 
    R_13b27_102eb588 , 
    R_fa2a_1056e0f8 , 
    R_145a5_132f4dc8 , 
    R_14060_13a15ae8 , 
    R_164_12b27118 , 
    R_104d9_120779b8 , 
    R_1ab_f8c2998 , 
    R_23c_13319328 , 
    R_bbdf_133063a8 , 
    R_d3_12659968 , 
    R_cc7b_13a1b128 , 
    R_12ffe_1331cd48 , 
    R_1323e_126561c8 , 
    R_1207f_133190a8 , 
    R_10f99_126549a8 , 
    R_913d_12646b28 , 
    R_c3ee_102f6848 , 
    R_13b12_13a1a728 , 
    R_10a0c_11cdf1c8 , 
    R_13974_13a19008 , 
    R_13602_126635a8 , 
    R_124e1_11cdb668 , 
    R_142d7_12b30d58 , 
    R_14960_105b5598 , 
    R_f86d_120385f8 , 
    R_148a0_12b38ab8 , 
    R_e63f_f8cb9f8 , 
    R_12741_105642d8 , 
    R_684e_1056aa98 , 
    R_13b04_12081558 , 
    R_1453f_11ce2328 , 
    R_148b5_1207f898 , 
    R_1499c_12080658 , 
    R_128e2_12647668 , 
    R_13345_11ce0988 , 
    R_cd4f_102f2f68 , 
    R_13dd3_1204cd38 , 
    R_13ea4_11ce0708 , 
    R_f16b_11cda448 , 
    R_139fe_1153e5b8 , 
    R_12eed_102ee1e8 , 
    R_13479_13306b28 , 
    R_1135b_1056d158 , 
    R_131a5_1153dc58 , 
    R_14744_1264b3a8 , 
    R_144c6_1056d5b8 , 
    R_13109_f8c4798 , 
    R_137bb_10564058 , 
    R_146db_1056a818 , 
    R_119c2_13a1a548 , 
    R_eb5e_1056d018 , 
    R_b0d7_1153e3d8 , 
    R_13b9e_12083038 , 
    R_1116a_13a15868 , 
    R_12a65_10564c38 , 
    R_14969_11cdb2a8 , 
    R_1464d_12075618 , 
    R_e3c5_12080a18 , 
    R_1469c_120511f8 , 
    R_d50f_12663828 , 
    R_137f0_12079358 , 
    R_11593_1207a258 , 
    R_14350_1207d8b8 , 
    R_cbe2_11536a98 , 
    R_110ed_10563d38 , 
    R_1125d_102f86e8 , 
    R_13c09_11ce4268 , 
    R_135fc_13795948 , 
    R_14557_11cdcec8 , 
    R_112_13312248 , 
    R_1fd_133221a8 , 
    R_9e_11539838 , 
    R_143b2_11cddd28 , 
    R_12fec_102efea8 , 
    R_c4d7_13a1f408 , 
    R_1398e_13320bc8 , 
    R_12894_11ce1428 , 
    R_b6f4_102f9ea8 , 
    R_fcb3_12649be8 , 
    R_12375_1207edf8 , 
    R_146b1_102ed248 , 
    R_11b11_11545818 , 
    R_58_13317a28 , 
    R_73_12b3e0f8 , 
    R_bd7c_11ce2be8 , 
    R_12fd8_10565278 , 
    R_14876_12054678 , 
    R_138da_1153dbb8 , 
    R_14825_12647168 , 
    R_14a4d_12646ee8 , 
    R_124_1203edb8 , 
    R_15a_f8c6958 , 
    R_1b5_1331afe8 , 
    R_1eb_12038d78 , 
    R_1475d_11546038 , 
    R_171_105aa5f8 , 
    R_106ea_102f6528 , 
    R_19e_1331e788 , 
    R_11a86_1204ffd8 , 
    R_fad7_102f5ee8 , 
    R_e21e_1056b7b8 , 
    R_12933_11cd7c48 , 
    R_6c_12040938 , 
    R_99_12b27618 , 
    R_1353d_1153d9d8 , 
    R_b283_1330acc8 , 
    R_143ae_13a1cca8 , 
    R_14801_11540c78 , 
    R_149e7_10568298 , 
    R_14708_1203c018 , 
    R_14450_13a17028 , 
    R_128_12b43b98 , 
    R_145_1265aa48 , 
    R_1ca_1265ff48 , 
    R_1e7_12b3d798 , 
    R_7741_13a16128 , 
    R_da39_12b40718 , 
    R_e38d_12651168 , 
    R_12fc4_11544878 , 
    R_145e7_11544058 , 
    R_1465f_105676b8 , 
    R_10fc1_12078638 , 
    R_704f_11ce4da8 , 
    R_13a8d_13318108 , 
    R_145c3_1264da68 , 
    R_faad_13a1fd68 , 
    R_12738_10570678 , 
    R_11935_13a1ff48 , 
    R_11720_1330eaa8 , 
    R_d16a_11ce5de8 , 
    R_13e0d_13a1b4e8 , 
    R_1447d_11ce3a48 , 
    R_152_12b3c4d8 , 
    R_105ba_13306bc8 , 
    R_b1aa_12649468 , 
    R_1bd_12653be8 , 
    R_14a50_13a161c8 , 
    R_13a83_10567a78 , 
    R_123c2_13797108 , 
    R_144b7_13305d68 , 
    R_13814_137926a8 , 
    R_12cbd_13a14328 , 
    R_11bab_120768d8 , 
    R_c07e_13a18b08 , 
    R_142f9_11545e58 , 
    R_1478a_12652928 , 
    R_14a3b_11ce2d28 , 
    R_c3a2_13a19508 , 
    R_aa_126535a8 , 
    R_146e7_10566538 , 
    R_138fb_12082778 , 
    R_13988_133186a8 , 
    R_13c43_1264cca8 , 
    R_14590_132f3b08 , 
    R_110cf_137940e8 , 
    R_13326_12648d88 , 
    R_13153_10567118 , 
    R_1405e_f8c95b8 , 
    R_1051f_13793b48 , 
    R_f518_12075bb8 , 
    R_143a2_12079038 , 
    R_147a8_12657de8 , 
    R_13cb3_102f6fc8 , 
    R_10c3d_f8c5b98 , 
    R_e7ab_1264f7c8 , 
    R_13449_12077378 , 
    R_14403_12b29418 , 
    R_148b2_132fc708 , 
    R_1468f_10562cf8 , 
    R_f7_13309828 , 
    R_13f54_102f4e08 , 
    R_218_12050258 , 
    R_83_1379cd88 , 
    R_12f16_137a0b68 , 
    R_10598_102ead68 , 
    R_10365_12051478 , 
    R_13ab4_13a12ca8 , 
    R_13393_10568a18 , 
    R_13683_1207cf58 , 
    R_13a_105ac2b8 , 
    R_127d5_11cdf268 , 
    R_11917_11ce1248 , 
    R_1d5_1265e468 , 
    R_12e98_1204e778 , 
    R_b3_12655ea8 , 
    R_149cc_10564cd8 , 
    R_134d9_10565f98 , 
    R_fd0b_102ec488 , 
    R_af25_133136a8 , 
    R_11948_12b288d8 , 
    R_149c6_1207b018 , 
    R_14b_12b28a18 , 
    R_1c4_12652e28 , 
    R_10199_13a1f368 , 
    R_80_12055438 , 
    R_10b70_f8cd438 , 
    R_10cdf_115401d8 , 
    R_11a66_1207dc78 , 
    R_132fc_13307708 , 
    R_8c7b_12076b58 , 
    R_1495a_1207a2f8 , 
    R_1201a_10570218 , 
    R_132d6_11ce0348 , 
    R_14963_13304be8 , 
    R_1285e_11545c78 , 
    R_130de_102f58a8 , 
    R_fb5f_13a1e288 , 
    R_13ecf_1207c5f8 , 
    R_1456f_13a1f5e8 , 
    R_ea_1331a9a8 , 
    R_120_12b400d8 , 
    R_13eac_11ce2a08 , 
    R_12568_1056b0d8 , 
    R_e3ba_1207df98 , 
    R_dcf2_12085298 , 
    R_1ef_f8c2cb8 , 
    R_225_12b3a318 , 
    R_f7da_1204e9f8 , 
    R_f857_13a13748 , 
    R_1461a_13301988 , 
    R_146b7_13a15228 , 
    R_1384a_126503a8 , 
    R_c8e7_105b6498 , 
    R_86_137a1a68 , 
    R_a3_126621a8 , 
    R_f862_13a1a908 , 
    R_10ab7_102f7b08 , 
    R_11890_102eb308 , 
    R_df3c_120774b8 , 
    R_1369b_1330c2a8 , 
    R_12e03_132ff368 , 
    R_1356b_102f5da8 , 
    R_10e42_1207e718 , 
    R_10f59_f8c2c18 , 
    R_127b6_12b412f8 , 
    R_120e7_12b44818 , 
    R_12492_1265b9e8 , 
    R_10d12_13792b08 , 
    R_130ae_12044b78 , 
    R_13652_11ce1ce8 , 
    R_117a7_12080fb8 , 
    R_14674_13a13ba8 , 
    R_11306_11540638 , 
    R_d5_126617a8 , 
    R_de_1265ce88 , 
    R_12c_1379b488 , 
    R_135_f8c6f98 , 
    R_1da_12664b88 , 
    R_1e3_1153c498 , 
    R_122dd_13a1b6c8 , 
    R_231_1379a6c8 , 
    R_23a_12660b28 , 
    R_1240e_13a150e8 , 
    R_14686_13a137e8 , 
    R_146c6_f8cf918 , 
    R_13f5b_1207c738 , 
    R_ebb7_102efd68 , 
    R_1447a_105697d8 , 
    R_13c95_12650ee8 , 
    R_11de0_12083cb8 , 
    R_11552_12648c48 , 
    R_11cb2_1207ab18 , 
    R_14849_11ce0028 , 
    R_13f45_13a134c8 , 
    R_13726_12084f78 , 
    R_121f2_102f30a8 , 
    R_ef_1379b0c8 , 
    R_163_12b38a18 , 
    R_1ac_12b29558 , 
    R_220_12b25638 , 
    R_14623_13a12a28 , 
    R_1393a_11ce3408 , 
    R_139ea_11cd8828 , 
    R_cf49_11541718 , 
    R_b889_1056a458 , 
    R_1349f_1204fdf8 , 
    R_170_120440d8 , 
    R_19f_133087e8 , 
    R_a9d8_102f22e8 , 
    R_7d_12660308 , 
    R_1460b_10569a58 , 
    R_11983_13318568 , 
    R_a6e4_13314648 , 
    R_144b1_1207b478 , 
    R_14614_12664f48 , 
    R_139d7_132fda68 , 
    R_ec64_11ce6248 , 
    R_12d32_115454f8 , 
    R_82bb_1204a678 , 
    R_1472c_13a139c8 , 
    R_144f7_10565e58 , 
    R_10dad_12082f98 , 
    R_b05c_1330b4e8 , 
    R_13ef1_105714d8 , 
    R_14635_12b3b038 , 
    R_117b5_1056fdb8 , 
    R_14692_11cdf128 , 
    R_13f_1203dd78 , 
    R_1055c_105672f8 , 
    R_1d0_12040258 , 
    R_13aba_1265cde8 , 
    R_131e1_102f2ec8 , 
    R_eb07_1153ef18 , 
    R_9c9a_1056c578 , 
    R_10605_11545d18 , 
    R_13a97_12079218 , 
    R_1331b_102efc28 , 
    R_14879_11ce58e8 , 
    R_14996_102eb3a8 , 
    R_1405c_11ce34a8 , 
    R_14945_1056e238 , 
    R_b65f_11cdba28 , 
    R_13f3e_13a1e508 , 
    R_dbc0_132fb9e8 , 
    R_1351c_13797068 , 
    R_14804_120788b8 , 
    R_14a0b_133206c8 , 
    R_89_126595a8 , 
    R_13c33_11ce3688 , 
    R_4f_12b44d18 , 
    R_cb5a_12b256d8 , 
    R_13b85_10571258 , 
    R_138f4_1330a9a8 , 
    R_ee1a_1264fae8 , 
    R_10411_102f8828 , 
    R_14331_1056be98 , 
    R_14717_1153a378 , 
    R_94_1330ee68 , 
    R_e5_1153cfd8 , 
    R_22a_12b43698 , 
    R_cba1_13a16e48 , 
    R_129d1_12047978 , 
    R_143d8_11cdc2e8 , 
    R_13070_1264b268 , 
    R_12915_1056d518 , 
    R_12942_11cdd0a8 , 
    R_145a8_12662608 , 
    R_fda2_1264e328 , 
    R_ee25_13a16588 , 
    R_13a1f_11cde2c8 , 
    R_1432d_11cdddc8 , 
    R_13be3_12036bb8 , 
    R_fe10_13a14468 , 
    R_12610_1204bcf8 , 
    R_13701_11cdc608 , 
    R_12597_105711b8 , 
    R_1441d_12035d58 , 
    R_1443c_137979c8 , 
    R_139a7_11ce70a8 , 
    R_13ad3_1056bdf8 , 
    R_143e0_102efcc8 , 
    R_147cc_13315ae8 , 
    R_1444b_11cdad08 , 
    R_12631_12036c58 , 
    R_13dda_102f4fe8 , 
    R_efd_13a14fa8 , 
    R_14954_12054358 , 
    R_1287f_115422f8 , 
    R_1169f_102f8968 , 
    R_13a2b_1264b628 , 
    R_11285_102f9e08 , 
    R_12548_1056ce38 , 
    R_1173e_12649fa8 , 
    R_10b51_13a18a68 , 
    R_148ca_13a18c48 , 
    R_12c82_102f0448 , 
    R_13b79_11543d38 , 
    R_14057_f8cd618 , 
    R_a2e4_1056c618 , 
    R_101e6_1330c7a8 , 
    R_13a56_f8c0a58 , 
    R_d6bc_13a1ca28 , 
    R_4a_1265e648 , 
    R_115_13316c68 , 
    R_1224c_12b3d478 , 
    R_1fa_1265d388 , 
    R_eeda_11cd81e8 , 
    R_1455d_11cd9fe8 , 
    R_1402e_1264dc48 , 
    R_c753_12039098 , 
    R_1283c_13a1da68 , 
    R_aeda_13a1d6a8 , 
    R_14939_1379f448 , 
    R_14a20_13a13e28 , 
    R_13a9d_12081698 , 
    R_117c0_11ce3e08 , 
    R_114e1_132f28e8 , 
    R_1476f_132fb768;
wire 
    n10016 , 
    n10017 , 
    n10018 , 
    n10019 , 
    n10020 , 
    n10021 , 
    n10022 , 
    n10023 , 
    n10024 , 
    n10025 , 
    n10026 , 
    n10027 , 
    n10028 , 
    n10029 , 
    n10030 , 
    n10031 , 
    n10032 , 
    n10033 , 
    n10034 , 
    n10035 , 
    n10036 , 
    n10037 , 
    n10038 , 
    n10039 , 
    n10040 , 
    n10041 , 
    n10042 , 
    n10043 , 
    n10044 , 
    n10045 , 
    n10046 , 
    n10047 , 
    n10048 , 
    n10049 , 
    n10050 , 
    n10051 , 
    n10052 , 
    n10053 , 
    n10054 , 
    n10055 , 
    n10056 , 
    n10057 , 
    n10058 , 
    n10059 , 
    n10060 , 
    n10061 , 
    n10062 , 
    n10063 , 
    n10064 , 
    n10065 , 
    n10066 , 
    n10067 , 
    n10068 , 
    n10069 , 
    n10070 , 
    n10071 , 
    n10072 , 
    n10073 , 
    n10074 , 
    n10075 , 
    n10076 , 
    n10077 , 
    n10078 , 
    n10079 , 
    n10080 , 
    n10081 , 
    n10082 , 
    n10083 , 
    n10084 , 
    n10085 , 
    n10086 , 
    n10087 , 
    n10088 , 
    n10089 , 
    n10090 , 
    n10091 , 
    n10092 , 
    n10093 , 
    n10094 , 
    n10095 , 
    n10096 , 
    n10097 , 
    n10098 , 
    n10099 , 
    n10100 , 
    n10101 , 
    n10102 , 
    n10103 , 
    n10104 , 
    n10105 , 
    n10106 , 
    n10107 , 
    n10108 , 
    n10109 , 
    n10110 , 
    n10111 , 
    n10112 , 
    n10113 , 
    n10114 , 
    n10115 , 
    n10116 , 
    n10117 , 
    n10118 , 
    n10119 , 
    n10120 , 
    n10121 , 
    n10122 , 
    n10123 , 
    n10124 , 
    n10125 , 
    n10126 , 
    n10127 , 
    n10128 , 
    n10129 , 
    n10130 , 
    n10131 , 
    n10132 , 
    n10133 , 
    n10134 , 
    n10135 , 
    n10136 , 
    n10137 , 
    n10138 , 
    n10139 , 
    n10140 , 
    n10141 , 
    n10142 , 
    n10143 , 
    n10144 , 
    n10145 , 
    n10146 , 
    n10147 , 
    n10148 , 
    n10149 , 
    n10150 , 
    n10151 , 
    n10152 , 
    n10153 , 
    n10154 , 
    n10155 , 
    n10156 , 
    n10157 , 
    n10158 , 
    n10159 , 
    n10160 , 
    n10161 , 
    n10162 , 
    n10163 , 
    n10164 , 
    n10165 , 
    n10166 , 
    n10167 , 
    n10168 , 
    n10169 , 
    n10170 , 
    n10171 , 
    n10172 , 
    n10173 , 
    n10174 , 
    n10175 , 
    n10176 , 
    n10177 , 
    n10178 , 
    n10179 , 
    n10180 , 
    n10181 , 
    n10182 , 
    n10183 , 
    n10184 , 
    n10185 , 
    n10186 , 
    n10187 , 
    n10188 , 
    n10189 , 
    n10190 , 
    n10191 , 
    n10192 , 
    n10193 , 
    n10194 , 
    n10195 , 
    n10196 , 
    n10197 , 
    n10198 , 
    n10199 , 
    n10200 , 
    n10201 , 
    n10202 , 
    n10203 , 
    n10204 , 
    n10205 , 
    n10206 , 
    n10207 , 
    n10208 , 
    n10209 , 
    n10210 , 
    n10211 , 
    n10212 , 
    n10213 , 
    n10214 , 
    n10215 , 
    n10216 , 
    n10217 , 
    n10218 , 
    n10219 , 
    n10220 , 
    n10221 , 
    n10222 , 
    n10223 , 
    n10224 , 
    n10225 , 
    n10226 , 
    n10227 , 
    n10228 , 
    n10229 , 
    n10230 , 
    n10231 , 
    n10232 , 
    n10233 , 
    n10234 , 
    n10235 , 
    n10236 , 
    n10237 , 
    n10238 , 
    n10239 , 
    n10240 , 
    n10241 , 
    n10242 , 
    n10243 , 
    n10244 , 
    n10245 , 
    n10246 , 
    n10247 , 
    n10248 , 
    n10249 , 
    n10250 , 
    n10251 , 
    n10252 , 
    n10253 , 
    n10254 , 
    n10255 , 
    n10256 , 
    n10257 , 
    n10258 , 
    n10259 , 
    n10260 , 
    n10261 , 
    n10262 , 
    n10263 , 
    n10264 , 
    n10265 , 
    n10266 , 
    n10267 , 
    n10268 , 
    n10269 , 
    n10270 , 
    n10271 , 
    n10272 , 
    n10273 , 
    n10274 , 
    n10275 , 
    n10276 , 
    n10277 , 
    n10278 , 
    n10279 , 
    n10280 , 
    n10281 , 
    n10282 , 
    n10283 , 
    n10284 , 
    n10285 , 
    n10286 , 
    n10287 , 
    n10288 , 
    n10289 , 
    n10290 , 
    n10291 , 
    n10292 , 
    n10293 , 
    n10294 , 
    n10295 , 
    n10296 , 
    n10297 , 
    n10298 , 
    n10299 , 
    n10300 , 
    n10301 , 
    n10302 , 
    n10303 , 
    n10304 , 
    n10305 , 
    n10306 , 
    n10307 , 
    n10308 , 
    n10309 , 
    n10310 , 
    n10311 , 
    n10312 , 
    n10313 , 
    n10314 , 
    n10315 , 
    n10316 , 
    n10317 , 
    n10318 , 
    n10319 , 
    n10320 , 
    n10321 , 
    n10322 , 
    n10323 , 
    n10324 , 
    n10325 , 
    n10326 , 
    n10327 , 
    n10328 , 
    n10329 , 
    n10330 , 
    n10331 , 
    n10332 , 
    n10333 , 
    n10334 , 
    n10335 , 
    n10336 , 
    n10337 , 
    n10338 , 
    n10339 , 
    n10340 , 
    n10341 , 
    n10342 , 
    n10343 , 
    n10344 , 
    n10345 , 
    n10346 , 
    n10347 , 
    n10348 , 
    n10349 , 
    n10350 , 
    n10351 , 
    n10352 , 
    n10353 , 
    n10354 , 
    n10355 , 
    n10356 , 
    n10357 , 
    n10358 , 
    n10359 , 
    n10360 , 
    n10361 , 
    n10362 , 
    n10363 , 
    n10364 , 
    n10365 , 
    n10366 , 
    n10367 , 
    n10368 , 
    n10369 , 
    n10370 , 
    n10371 , 
    n10372 , 
    n10373 , 
    n10374 , 
    n10375 , 
    n10376 , 
    n10377 , 
    n10378 , 
    n10379 , 
    n10380 , 
    n10381 , 
    n10382 , 
    n10383 , 
    n10384 , 
    n10385 , 
    n10386 , 
    n10387 , 
    n10388 , 
    n10389 , 
    n10390 , 
    n10391 , 
    n10392 , 
    n10393 , 
    n10394 , 
    n10395 , 
    n10396 , 
    n10397 , 
    n10398 , 
    n10399 , 
    n10400 , 
    n10401 , 
    n10402 , 
    n10403 , 
    n10404 , 
    n10405 , 
    n10406 , 
    n10407 , 
    n10408 , 
    n10409 , 
    n10410 , 
    n10411 , 
    n10412 , 
    n10413 , 
    n10414 , 
    n10415 , 
    n10416 , 
    n10417 , 
    n10418 , 
    n10419 , 
    n10420 , 
    n10421 , 
    n10422 , 
    n10423 , 
    n10424 , 
    n10425 , 
    n10426 , 
    n10427 , 
    n10428 , 
    n10429 , 
    n10430 , 
    n10431 , 
    n10432 , 
    n10433 , 
    n10434 , 
    n10435 , 
    n10436 , 
    n10437 , 
    n10438 , 
    n10439 , 
    n10440 , 
    n10441 , 
    n10442 , 
    n10443 , 
    n10444 , 
    n10445 , 
    n10446 , 
    n10447 , 
    n10448 , 
    n10449 , 
    n10450 , 
    n10451 , 
    n10452 , 
    n10453 , 
    n10454 , 
    n10455 , 
    n10456 , 
    n10457 , 
    n10458 , 
    n10459 , 
    n10460 , 
    n10461 , 
    n10462 , 
    n10463 , 
    n10464 , 
    n10465 , 
    n10466 , 
    n10467 , 
    n10468 , 
    n10469 , 
    n10470 , 
    n10471 , 
    n10472 , 
    n10473 , 
    n10474 , 
    n10475 , 
    n10476 , 
    n10477 , 
    n10478 , 
    n10479 , 
    n10480 , 
    n10481 , 
    n10482 , 
    n10483 , 
    n10484 , 
    n10485 , 
    n10486 , 
    n10487 , 
    n10488 , 
    n10489 , 
    n10490 , 
    n10491 , 
    n10492 , 
    n10493 , 
    n10494 , 
    n10495 , 
    n10496 , 
    n10497 , 
    n10498 , 
    n10499 , 
    n10500 , 
    n10501 , 
    n10502 , 
    n10503 , 
    n10504 , 
    n10505 , 
    n10506 , 
    n10507 , 
    n10508 , 
    n10509 , 
    n10510 , 
    n10511 , 
    n10512 , 
    n10513 , 
    n10514 , 
    n10515 , 
    n10516 , 
    n10517 , 
    n10518 , 
    n10519 , 
    n10520 , 
    n10521 , 
    n10522 , 
    n10523 , 
    n10524 , 
    n10525 , 
    n10526 , 
    n10527 , 
    n10528 , 
    n10529 , 
    n10530 , 
    n10531 , 
    n10532 , 
    n10533 , 
    n10534 , 
    n10535 , 
    n10536 , 
    n10537 , 
    n10538 , 
    n10539 , 
    n10540 , 
    n10541 , 
    n10542 , 
    n10543 , 
    n10544 , 
    n10545 , 
    n10546 , 
    n10547 , 
    n10548 , 
    n10549 , 
    n10550 , 
    n10551 , 
    n10552 , 
    n10553 , 
    n10554 , 
    n10555 , 
    n10556 , 
    n10557 , 
    n10558 , 
    n10559 , 
    n10560 , 
    n10561 , 
    n10562 , 
    n10563 , 
    n10564 , 
    n10565 , 
    n10566 , 
    n10567 , 
    n10568 , 
    n10569 , 
    n10570 , 
    n10571 , 
    n10572 , 
    n10573 , 
    n10574 , 
    n10575 , 
    n10576 , 
    n10577 , 
    n10578 , 
    n10579 , 
    n10580 , 
    n10581 , 
    n10582 , 
    n10583 , 
    n10584 , 
    n10585 , 
    n10586 , 
    n10587 , 
    n10588 , 
    n10589 , 
    n10590 , 
    n10591 , 
    n10592 , 
    n10593 , 
    n10594 , 
    n10595 , 
    n10596 , 
    n10597 , 
    n10598 , 
    n10599 , 
    n10600 , 
    n10601 , 
    n10602 , 
    n10603 , 
    n10604 , 
    n10605 , 
    n10606 , 
    n10607 , 
    n10608 , 
    n10609 , 
    n10610 , 
    n10611 , 
    n10612 , 
    n10613 , 
    n10614 , 
    n10615 , 
    n10616 , 
    n10617 , 
    n10618 , 
    n10619 , 
    n10620 , 
    n10621 , 
    n10622 , 
    n10623 , 
    n10624 , 
    n10625 , 
    n10626 , 
    n10627 , 
    n10628 , 
    n10629 , 
    n10630 , 
    n10631 , 
    n10632 , 
    n10633 , 
    n10634 , 
    n10635 , 
    n10636 , 
    n10637 , 
    n10638 , 
    n10639 , 
    n10640 , 
    n10641 , 
    n10642 , 
    n10643 , 
    n10644 , 
    n10645 , 
    n10646 , 
    n10647 , 
    n10648 , 
    n10649 , 
    n10650 , 
    n10651 , 
    n10652 , 
    n10653 , 
    n10654 , 
    n10655 , 
    n10656 , 
    n10657 , 
    n10658 , 
    n10659 , 
    n10660 , 
    n10661 , 
    n10662 , 
    n10663 , 
    n10664 , 
    n10665 , 
    n10666 , 
    n10667 , 
    n10668 , 
    n10669 , 
    n10670 , 
    n10671 , 
    n10672 , 
    n10673 , 
    n10674 , 
    n10675 , 
    n10676 , 
    n10677 , 
    n10678 , 
    n10679 , 
    n10680 , 
    n10681 , 
    n10682 , 
    n10683 , 
    n10684 , 
    n10685 , 
    n10686 , 
    n10687 , 
    n10688 , 
    n10689 , 
    n10690 , 
    n10691 , 
    n10692 , 
    n10693 , 
    n10694 , 
    n10695 , 
    n10696 , 
    n10697 , 
    n10698 , 
    n10699 , 
    n10700 , 
    n10701 , 
    n10702 , 
    n10703 , 
    n10704 , 
    n10705 , 
    n10706 , 
    n10707 , 
    n10708 , 
    n10709 , 
    n10710 , 
    n10711 , 
    n10712 , 
    n10713 , 
    n10714 , 
    n10715 , 
    n10716 , 
    n10717 , 
    n10718 , 
    n10719 , 
    n10720 , 
    n10721 , 
    n10722 , 
    n10723 , 
    n10724 , 
    n10725 , 
    n10726 , 
    n10727 , 
    n10728 , 
    n10729 , 
    n10730 , 
    n10731 , 
    n10732 , 
    n10733 , 
    n10734 , 
    n10735 , 
    n10736 , 
    n10737 , 
    n10738 , 
    n10739 , 
    n10740 , 
    n10741 , 
    n10742 , 
    n10743 , 
    n10744 , 
    n10745 , 
    n10746 , 
    n10747 , 
    n10748 , 
    n10749 , 
    n10750 , 
    n10751 , 
    n10752 , 
    n10753 , 
    n10754 , 
    n10755 , 
    n10756 , 
    n10757 , 
    n10758 , 
    n10759 , 
    n10760 , 
    n10761 , 
    n10762 , 
    n10763 , 
    n10764 , 
    n10765 , 
    n10766 , 
    n10767 , 
    n10768 , 
    n10769 , 
    n10770 , 
    n10771 , 
    n10772 , 
    n10773 , 
    n10774 , 
    n10775 , 
    n10776 , 
    n10777 , 
    n10778 , 
    n10779 , 
    n10780 , 
    n10781 , 
    n10782 , 
    n10783 , 
    n10784 , 
    n10785 , 
    n10786 , 
    n10787 , 
    n10788 , 
    n10789 , 
    n10790 , 
    n10791 , 
    n10792 , 
    n10793 , 
    n10794 , 
    n10795 , 
    n10796 , 
    n10797 , 
    n10798 , 
    n10799 , 
    n10800 , 
    n10801 , 
    n10802 , 
    n10803 , 
    n10804 , 
    n10805 , 
    n10806 , 
    n10807 , 
    n10808 , 
    n10809 , 
    n10810 , 
    n10811 , 
    n10812 , 
    n10813 , 
    n10814 , 
    n10815 , 
    n10816 , 
    n10817 , 
    n10818 , 
    n10819 , 
    n10820 , 
    n10821 , 
    n10822 , 
    n10823 , 
    n10824 , 
    n10825 , 
    n10826 , 
    n10827 , 
    n10828 , 
    n10829 , 
    n10830 , 
    n10831 , 
    n10832 , 
    n10833 , 
    n10834 , 
    n10835 , 
    n10836 , 
    n10837 , 
    n10838 , 
    n10839 , 
    n10840 , 
    n10841 , 
    n10842 , 
    n10843 , 
    n10844 , 
    n10845 , 
    n10846 , 
    n10847 , 
    n10848 , 
    n10849 , 
    n10850 , 
    n10851 , 
    n10852 , 
    n10853 , 
    n10854 , 
    n10855 , 
    n10856 , 
    n10857 , 
    n10858 , 
    n10859 , 
    n10860 , 
    n10861 , 
    n10862 , 
    n10863 , 
    n10864 , 
    n10865 , 
    n10866 , 
    n10867 , 
    n10868 , 
    n10869 , 
    n10870 , 
    n10871 , 
    n10872 , 
    n10873 , 
    n10874 , 
    n10875 , 
    n10876 , 
    n10877 , 
    n10878 , 
    n10879 , 
    n10880 , 
    n10881 , 
    n10882 , 
    n10883 , 
    n10884 , 
    n10885 , 
    n10886 , 
    n10887 , 
    n10888 , 
    n10889 , 
    n10890 , 
    n10891 , 
    n10892 , 
    n10893 , 
    n10894 , 
    n10895 , 
    n10896 , 
    n10897 , 
    n10898 , 
    n10899 , 
    n10900 , 
    n10901 , 
    n10902 , 
    n10903 , 
    n10904 , 
    n10905 , 
    n10906 , 
    n10907 , 
    n10908 , 
    n10909 , 
    n10910 , 
    n10911 , 
    n10912 , 
    n10913 , 
    n10914 , 
    n10915 , 
    n10916 , 
    n10917 , 
    n10918 , 
    n10919 , 
    n10920 , 
    n10921 , 
    n10922 , 
    n10923 , 
    n10924 , 
    n10925 , 
    n10926 , 
    n10927 , 
    n10928 , 
    n10929 , 
    n10930 , 
    n10931 , 
    n10932 , 
    n10933 , 
    n10934 , 
    n10935 , 
    n10936 , 
    n10937 , 
    n10938 , 
    n10939 , 
    n10940 , 
    n10941 , 
    n10942 , 
    n10943 , 
    n10944 , 
    n10945 , 
    n10946 , 
    n10947 , 
    n10948 , 
    n10949 , 
    n10950 , 
    n10951 , 
    n10952 , 
    n10953 , 
    n10954 , 
    n10955 , 
    n10956 , 
    n10957 , 
    n10958 , 
    n10959 , 
    n10960 , 
    n10961 , 
    n10962 , 
    n10963 , 
    n10964 , 
    n10965 , 
    n10966 , 
    n10967 , 
    n10968 , 
    n10969 , 
    n10970 , 
    n10971 , 
    n10972 , 
    n10973 , 
    n10974 , 
    n10975 , 
    n10976 , 
    n10977 , 
    n10978 , 
    n10979 , 
    n10980 , 
    n10981 , 
    n10982 , 
    n10983 , 
    n10984 , 
    n10985 , 
    n10986 , 
    n10987 , 
    n10988 , 
    n10989 , 
    n10990 , 
    n10991 , 
    n10992 , 
    n10993 , 
    n10994 , 
    n10995 , 
    n10996 , 
    n10997 , 
    n10998 , 
    n10999 , 
    n11000 , 
    n11001 , 
    n11002 , 
    n11003 , 
    n11004 , 
    n11005 , 
    n11006 , 
    n11007 , 
    n11008 , 
    n11009 , 
    n11010 , 
    n11011 , 
    n11012 , 
    n11013 , 
    n11014 , 
    n11015 , 
    n11016 , 
    n11017 , 
    n11018 , 
    n11019 , 
    n11020 , 
    n11021 , 
    n11022 , 
    n11023 , 
    n11024 , 
    n11025 , 
    n11026 , 
    n11027 , 
    n11028 , 
    n11029 , 
    n11030 , 
    n11031 , 
    n11032 , 
    n11033 , 
    n11034 , 
    n11035 , 
    n11036 , 
    n11037 , 
    n11038 , 
    n11039 , 
    n11040 , 
    n11041 , 
    n11042 , 
    n11043 , 
    n11044 , 
    n11045 , 
    n11046 , 
    n11047 , 
    n11048 , 
    n11049 , 
    n11050 , 
    n11051 , 
    n11052 , 
    n11053 , 
    n11054 , 
    n11055 , 
    n11056 , 
    n11057 , 
    n11058 , 
    n11059 , 
    n11060 , 
    n11061 , 
    n11062 , 
    n11063 , 
    n11064 , 
    n11065 , 
    n11066 , 
    n11067 , 
    n11068 , 
    n11069 , 
    n11070 , 
    n11071 , 
    n11072 , 
    n11073 , 
    n11074 , 
    n11075 , 
    n11076 , 
    n11077 , 
    n11078 , 
    n11079 , 
    n11080 , 
    n11081 , 
    n11082 , 
    n11083 , 
    n11084 , 
    n11085 , 
    n11086 , 
    n11087 , 
    n11088 , 
    n11089 , 
    n11090 , 
    n11091 , 
    n11092 , 
    n11093 , 
    n11094 , 
    n11095 , 
    n11096 , 
    n11097 , 
    n11098 , 
    n11099 , 
    n11100 , 
    n11101 , 
    n11102 , 
    n11103 , 
    n11104 , 
    n11105 , 
    n11106 , 
    n11107 , 
    n11108 , 
    n11109 , 
    n11110 , 
    n11111 , 
    n11112 , 
    n11113 , 
    n11114 , 
    n11115 , 
    n11116 , 
    n11117 , 
    n11118 , 
    n11119 , 
    n11120 , 
    n11121 , 
    n11122 , 
    n11123 , 
    n11124 , 
    n11125 , 
    n11126 , 
    n11127 , 
    n11128 , 
    n11129 , 
    n11130 , 
    n11131 , 
    n11132 , 
    n11133 , 
    n11134 , 
    n11135 , 
    n11136 , 
    n11137 , 
    n11138 , 
    n11139 , 
    n11140 , 
    n11141 , 
    n11142 , 
    n11143 , 
    n11144 , 
    n11145 , 
    n11146 , 
    n11147 , 
    n11148 , 
    n11149 , 
    n11150 , 
    n11151 , 
    n11152 , 
    n11153 , 
    n11154 , 
    n11155 , 
    n11156 , 
    n11157 , 
    n11158 , 
    n11159 , 
    n11160 , 
    n11161 , 
    n11162 , 
    n11163 , 
    n11164 , 
    n11165 , 
    n11166 , 
    n11167 , 
    n11168 , 
    n11169 , 
    n11170 , 
    n11171 , 
    n11172 , 
    n11173 , 
    n11174 , 
    n11175 , 
    n11176 , 
    n11177 , 
    n11178 , 
    n11179 , 
    n11180 , 
    n11181 , 
    n11182 , 
    n11183 , 
    n11184 , 
    n11185 , 
    n11186 , 
    n11187 , 
    n11188 , 
    n11189 , 
    n11190 , 
    n11191 , 
    n11192 , 
    n11193 , 
    n11194 , 
    n11195 , 
    n11196 , 
    n11197 , 
    n11198 , 
    n11199 , 
    n11200 , 
    n11201 , 
    n11202 , 
    n11203 , 
    n11204 , 
    n11205 , 
    n11206 , 
    n11207 , 
    n11208 , 
    n11209 , 
    n11210 , 
    n11211 , 
    n11212 , 
    n11213 , 
    n11214 , 
    n11215 , 
    n11216 , 
    n11217 , 
    n11218 , 
    n11219 , 
    n11220 , 
    n11221 , 
    n11222 , 
    n11223 , 
    n11224 , 
    n11225 , 
    n11226 , 
    n11227 , 
    n11228 , 
    n11229 , 
    n11230 , 
    n11231 , 
    n11232 , 
    n11233 , 
    n11234 , 
    n11235 , 
    n11236 , 
    n11237 , 
    n11238 , 
    n11239 , 
    n11240 , 
    n11241 , 
    n11242 , 
    n11243 , 
    n11244 , 
    n11245 , 
    n11246 , 
    n11247 , 
    n11248 , 
    n11249 , 
    n11250 , 
    n11251 , 
    n11252 , 
    n11253 , 
    n11254 , 
    n11255 , 
    n11256 , 
    n11257 , 
    n11258 , 
    n11259 , 
    n11260 , 
    n11261 , 
    n11262 , 
    n11263 , 
    n11264 , 
    n11265 , 
    n11266 , 
    n11267 , 
    n11268 , 
    n11269 , 
    n11270 , 
    n11271 , 
    n11272 , 
    n11273 , 
    n11274 , 
    n11275 , 
    n11276 , 
    n11277 , 
    n11278 , 
    n11279 , 
    n11280 , 
    n11281 , 
    n11282 , 
    n11283 , 
    n11284 , 
    n11285 , 
    n11286 , 
    n11287 , 
    n11288 , 
    n11289 , 
    n11290 , 
    n11291 , 
    n11292 , 
    n11293 , 
    n11294 , 
    n11295 , 
    n11296 , 
    n11297 , 
    n11298 , 
    n11299 , 
    n11300 , 
    n11301 , 
    n11302 , 
    n11303 , 
    n11304 , 
    n11305 , 
    n11306 , 
    n11307 , 
    n11308 , 
    n11309 , 
    n11310 , 
    n11311 , 
    n11312 , 
    n11313 , 
    n11314 , 
    n11315 , 
    n11316 , 
    n11317 , 
    n11318 , 
    n11319 , 
    n11320 , 
    n11321 , 
    n11322 , 
    n11323 , 
    n11324 , 
    n11325 , 
    n11326 , 
    n11327 , 
    n11328 , 
    n11329 , 
    n11330 , 
    n11331 , 
    n11332 , 
    n11333 , 
    n11334 , 
    n11335 , 
    n11336 , 
    n11337 , 
    n11338 , 
    n11339 , 
    n11340 , 
    n11341 , 
    n11342 , 
    n11343 , 
    n11344 , 
    n11345 , 
    n11346 , 
    n11347 , 
    n11348 , 
    n11349 , 
    n11350 , 
    n11351 , 
    n11352 , 
    n11353 , 
    n11354 , 
    n11355 , 
    n11356 , 
    n11357 , 
    n11358 , 
    n11359 , 
    n11360 , 
    n11361 , 
    n11362 , 
    n11363 , 
    n11364 , 
    n11365 , 
    n11366 , 
    n11367 , 
    n11368 , 
    n11369 , 
    n11370 , 
    n11371 , 
    n11372 , 
    n11373 , 
    n11374 , 
    n11375 , 
    n11376 , 
    n11377 , 
    n11378 , 
    n11379 , 
    n11380 , 
    n11381 , 
    n11382 , 
    n11383 , 
    n11384 , 
    n11385 , 
    n11386 , 
    n11387 , 
    n11388 , 
    n11389 , 
    n11390 , 
    n11391 , 
    n11392 , 
    n11393 , 
    n11394 , 
    n11395 , 
    n11396 , 
    n11397 , 
    n11398 , 
    n11399 , 
    n11400 , 
    n11401 , 
    n11402 , 
    n11403 , 
    n11404 , 
    n11405 , 
    n11406 , 
    n11407 , 
    n11408 , 
    n11409 , 
    n11410 , 
    n11411 , 
    n11412 , 
    n11413 , 
    n11414 , 
    n11415 , 
    n11416 , 
    n11417 , 
    n11418 , 
    n11419 , 
    n11420 , 
    n11421 , 
    n11422 , 
    n11423 , 
    n11424 , 
    n11425 , 
    n11426 , 
    n11427 , 
    n11428 , 
    n11429 , 
    n11430 , 
    n11431 , 
    n11432 , 
    n11433 , 
    n11434 , 
    n11435 , 
    n11436 , 
    n11437 , 
    n11438 , 
    n11439 , 
    n11440 , 
    n11441 , 
    n11442 , 
    n11443 , 
    n11444 , 
    n11445 , 
    n11446 , 
    n11447 , 
    n11448 , 
    n11449 , 
    n11450 , 
    n11451 , 
    n11452 , 
    n11453 , 
    n11454 , 
    n11455 , 
    n11456 , 
    n11457 , 
    n11458 , 
    n11459 , 
    n11460 , 
    n11461 , 
    n11462 , 
    n11463 , 
    n11464 , 
    n11465 , 
    n11466 , 
    n11467 , 
    n11468 , 
    n11469 , 
    n11470 , 
    n11471 , 
    n11472 , 
    n11473 , 
    n11474 , 
    n11475 , 
    n11476 , 
    n11477 , 
    n11478 , 
    n11479 , 
    n11480 , 
    n11481 , 
    n11482 , 
    n11483 , 
    n11484 , 
    n11485 , 
    n11486 , 
    n11487 , 
    n11488 , 
    n11489 , 
    n11490 , 
    n11491 , 
    n11492 , 
    n11493 , 
    n11494 , 
    n11495 , 
    n11496 , 
    n11497 , 
    n11498 , 
    n11499 , 
    n11500 , 
    n11501 , 
    n11502 , 
    n11503 , 
    n11504 , 
    n11505 , 
    n11506 , 
    n11507 , 
    n11508 , 
    n11509 , 
    n11510 , 
    n11511 , 
    n11512 , 
    n11513 , 
    n11514 , 
    n11515 , 
    n11516 , 
    n11517 , 
    n11518 , 
    n11519 , 
    n11520 , 
    n11521 , 
    n11522 , 
    n11523 , 
    n11524 , 
    n11525 , 
    n11526 , 
    n11527 , 
    n11528 , 
    n11529 , 
    n11530 , 
    n11531 , 
    n11532 , 
    n11533 , 
    n11534 , 
    n11535 , 
    n11536 , 
    n11537 , 
    n11538 , 
    n11539 , 
    n11540 , 
    n11541 , 
    n11542 , 
    n11543 , 
    n11544 , 
    n11545 , 
    n11546 , 
    n11547 , 
    n11548 , 
    n11549 , 
    n11550 , 
    n11551 , 
    n11552 , 
    n11553 , 
    n11554 , 
    n11555 , 
    n11556 , 
    n11557 , 
    n11558 , 
    n11559 , 
    n11560 , 
    n11561 , 
    n11562 , 
    n11563 , 
    n11564 , 
    n11565 , 
    n11566 , 
    n11567 , 
    n11568 , 
    n11569 , 
    n11570 , 
    n11571 , 
    n11572 , 
    n11573 , 
    n11574 , 
    n11575 , 
    n11576 , 
    n11577 , 
    n11578 , 
    n11579 , 
    n11580 , 
    n11581 , 
    n11582 , 
    n11583 , 
    n11584 , 
    n11585 , 
    n11586 , 
    n11587 , 
    n11588 , 
    n11589 , 
    n11590 , 
    n11591 , 
    n11592 , 
    n11593 , 
    n11594 , 
    n11595 , 
    n11596 , 
    n11597 , 
    n11598 , 
    n11599 , 
    n11600 , 
    n11601 , 
    n11602 , 
    n11603 , 
    n11604 , 
    n11605 , 
    n11606 , 
    n11607 , 
    n11608 , 
    n11609 , 
    n11610 , 
    n11611 , 
    n11612 , 
    n11613 , 
    n11614 , 
    n11615 , 
    n11616 , 
    n11617 , 
    n11618 , 
    n11619 , 
    n11620 , 
    n11621 , 
    n11622 , 
    n11623 , 
    n11624 , 
    n11625 , 
    n11626 , 
    n11627 , 
    n11628 , 
    n11629 , 
    n11630 , 
    n11631 , 
    n11632 , 
    n11633 , 
    n11634 , 
    n11635 , 
    n11636 , 
    n11637 , 
    n11638 , 
    n11639 , 
    n11640 , 
    n11641 , 
    n11642 , 
    n11643 , 
    n11644 , 
    n11645 , 
    n11646 , 
    n11647 , 
    n11648 , 
    n11649 , 
    n11650 , 
    n11651 , 
    n11652 , 
    n11653 , 
    n11654 , 
    n11655 , 
    n11656 , 
    n11657 , 
    n11658 , 
    n11659 , 
    n11660 , 
    n11661 , 
    n11662 , 
    n11663 , 
    n11664 , 
    n11665 , 
    n11666 , 
    n11667 , 
    n11668 , 
    n11669 , 
    n11670 , 
    n11671 , 
    n11672 , 
    n11673 , 
    n11674 , 
    n11675 , 
    n11676 , 
    n11677 , 
    n11678 , 
    n11679 , 
    n11680 , 
    n11681 , 
    n11682 , 
    n11683 , 
    n11684 , 
    n11685 , 
    n11686 , 
    n11687 , 
    n11688 , 
    n11689 , 
    n11690 , 
    n11691 , 
    n11692 , 
    n11693 , 
    n11694 , 
    n11695 , 
    n11696 , 
    n11697 , 
    n11698 , 
    n11699 , 
    n11700 , 
    n11701 , 
    n11702 , 
    n11703 , 
    n11704 , 
    n11705 , 
    n11706 , 
    n11707 , 
    n11708 , 
    n11709 , 
    n11710 , 
    n11711 , 
    n11712 , 
    n11713 , 
    n11714 , 
    n11715 , 
    n11716 , 
    n11717 , 
    n11718 , 
    n11719 , 
    n11720 , 
    n11721 , 
    n11722 , 
    n11723 , 
    n11724 , 
    n11725 , 
    n11726 , 
    n11727 , 
    n11728 , 
    n11729 , 
    n11730 , 
    n11731 , 
    n11732 , 
    n11733 , 
    n11734 , 
    n11735 , 
    n11736 , 
    n11737 , 
    n11738 , 
    n11739 , 
    n11740 , 
    n11741 , 
    n11742 , 
    n11743 , 
    n11744 , 
    n11745 , 
    n11746 , 
    n11747 , 
    n11748 , 
    n11749 , 
    n11750 , 
    n11751 , 
    n11752 , 
    n11753 , 
    n11754 , 
    n11755 , 
    n11756 , 
    n11757 , 
    n11758 , 
    n11759 , 
    n11760 , 
    n11761 , 
    n11762 , 
    n11763 , 
    n11764 , 
    n11765 , 
    n11766 , 
    n11767 , 
    n11768 , 
    n11769 , 
    n11770 , 
    n11771 , 
    n11772 , 
    n11773 , 
    n11774 , 
    n11775 , 
    n11776 , 
    n11777 , 
    n11778 , 
    n11779 , 
    n11780 , 
    n11781 , 
    n11782 , 
    n11783 , 
    n11784 , 
    n11785 , 
    n11786 , 
    n11787 , 
    n11788 , 
    n11789 , 
    n11790 , 
    n11791 , 
    n11792 , 
    n11793 , 
    n11794 , 
    n11795 , 
    n11796 , 
    n11797 , 
    n11798 , 
    n11799 , 
    n11800 , 
    n11801 , 
    n11802 , 
    n11803 , 
    n11804 , 
    n11805 , 
    n11806 , 
    n11807 , 
    n11808 , 
    n11809 , 
    n11810 , 
    n11811 , 
    n11812 , 
    n11813 , 
    n11814 , 
    n11815 , 
    n11816 , 
    n11817 , 
    n11818 , 
    n11819 , 
    n11820 , 
    n11821 , 
    n11822 , 
    n11823 , 
    n11824 , 
    n11825 , 
    n11826 , 
    n11827 , 
    n11828 , 
    n11829 , 
    n11830 , 
    n11831 , 
    n11832 , 
    n11833 , 
    n11834 , 
    n11835 , 
    n11836 , 
    n11837 , 
    n11838 , 
    n11839 , 
    n11840 , 
    n11841 , 
    n11842 , 
    n11843 , 
    n11844 , 
    n11845 , 
    n11846 , 
    n11847 , 
    n11848 , 
    n11849 , 
    n11850 , 
    n11851 , 
    n11852 , 
    n11853 , 
    n11854 , 
    n11855 , 
    n11856 , 
    n11857 , 
    n11858 , 
    n11859 , 
    n11860 , 
    n11861 , 
    n11862 , 
    n11863 , 
    n11864 , 
    n11865 , 
    n11866 , 
    n11867 , 
    n11868 , 
    n11869 , 
    n11870 , 
    n11871 , 
    n11872 , 
    n11873 , 
    n11874 , 
    n11875 , 
    n11876 , 
    n11877 , 
    n11878 , 
    n11879 , 
    n11880 , 
    n11881 , 
    n11882 , 
    n11883 , 
    n11884 , 
    n11885 , 
    n11886 , 
    n11887 , 
    n11888 , 
    n11889 , 
    n11890 , 
    n11891 , 
    n11892 , 
    n11893 , 
    n11894 , 
    n11895 , 
    n11896 , 
    n11897 , 
    n11898 , 
    n11899 , 
    n11900 , 
    n11901 , 
    n11902 , 
    n11903 , 
    n11904 , 
    n11905 , 
    n11906 , 
    n11907 , 
    n11908 , 
    n11909 , 
    n11910 , 
    n11911 , 
    n11912 , 
    n11913 , 
    n11914 , 
    n11915 , 
    n11916 , 
    n11917 , 
    n11918 , 
    n11919 , 
    n11920 , 
    n11921 , 
    n11922 , 
    n11923 , 
    n11924 , 
    n11925 , 
    n11926 , 
    n11927 , 
    n11928 , 
    n11929 , 
    n11930 , 
    n11931 , 
    n11932 , 
    n11933 , 
    n11934 , 
    n11935 , 
    n11936 , 
    n11937 , 
    n11938 , 
    n11939 , 
    n11940 , 
    n11941 , 
    n11942 , 
    n11943 , 
    n11944 , 
    n11945 , 
    n11946 , 
    n11947 , 
    n11948 , 
    n11949 , 
    n11950 , 
    n11951 , 
    n11952 , 
    n11953 , 
    n11954 , 
    n11955 , 
    n11956 , 
    n11957 , 
    n11958 , 
    n11959 , 
    n11960 , 
    n11961 , 
    n11962 , 
    n11963 , 
    n11964 , 
    n11965 , 
    n11966 , 
    n11967 , 
    n11968 , 
    n11969 , 
    n11970 , 
    n11971 , 
    n11972 , 
    n11973 , 
    n11974 , 
    n11975 , 
    n11976 , 
    n11977 , 
    n11978 , 
    n11979 , 
    n11980 , 
    n11981 , 
    n11982 , 
    n11983 , 
    n11984 , 
    n11985 , 
    n11986 , 
    n11987 , 
    n11988 , 
    n11989 , 
    n11990 , 
    n11991 , 
    n11992 , 
    n11993 , 
    n11994 , 
    n11995 , 
    n11996 , 
    n11997 , 
    n11998 , 
    n11999 , 
    n12000 , 
    n12001 , 
    n12002 , 
    n12003 , 
    n12004 , 
    n12005 , 
    n12006 , 
    n12007 , 
    n12008 , 
    n12009 , 
    n12010 , 
    n12011 , 
    n12012 , 
    n12013 , 
    n12014 , 
    n12015 , 
    n12016 , 
    n12017 , 
    n12018 , 
    n12019 , 
    n12020 , 
    n12021 , 
    n12022 , 
    n12023 , 
    n12024 , 
    n12025 , 
    n12026 , 
    n12027 , 
    n12028 , 
    n12029 , 
    n12030 , 
    n12031 , 
    n12032 , 
    n12033 , 
    n12034 , 
    n12035 , 
    n12036 , 
    n12037 , 
    n12038 , 
    n12039 , 
    n12040 , 
    n12041 , 
    n12042 , 
    n12043 , 
    n12044 , 
    n12045 , 
    n12046 , 
    n12047 , 
    n12048 , 
    n12049 , 
    n12050 , 
    n12051 , 
    n12052 , 
    n12053 , 
    n12054 , 
    n12055 , 
    n12056 , 
    n12057 , 
    n12058 , 
    n12059 , 
    n12060 , 
    n12061 , 
    n12062 , 
    n12063 , 
    n12064 , 
    n12065 , 
    n12066 , 
    n12067 , 
    n12068 , 
    n12069 , 
    n12070 , 
    n12071 , 
    n12072 , 
    n12073 , 
    n12074 , 
    n12075 , 
    n12076 , 
    n12077 , 
    n12078 , 
    n12079 , 
    n12080 , 
    n12081 , 
    n12082 , 
    n12083 , 
    n12084 , 
    n12085 , 
    n12086 , 
    n12087 , 
    n12088 , 
    n12089 , 
    n12090 , 
    n12091 , 
    n12092 , 
    n12093 , 
    n12094 , 
    n12095 , 
    n12096 , 
    n12097 , 
    n12098 , 
    n12099 , 
    n12100 , 
    n12101 , 
    n12102 , 
    n12103 , 
    n12104 , 
    n12105 , 
    n12106 , 
    n12107 , 
    n12108 , 
    n12109 , 
    n12110 , 
    n12111 , 
    n12112 , 
    n12113 , 
    n12114 , 
    n12115 , 
    n12116 , 
    n12117 , 
    n12118 , 
    n12119 , 
    n12120 , 
    n12121 , 
    n12122 , 
    n12123 , 
    n12124 , 
    n12125 , 
    n12126 , 
    n12127 , 
    n12128 , 
    n12129 , 
    n12130 , 
    n12131 , 
    n12132 , 
    n12133 , 
    n12134 , 
    n12135 , 
    n12136 , 
    n12137 , 
    n12138 , 
    n12139 , 
    n12140 , 
    n12141 , 
    n12142 , 
    n12143 , 
    n12144 , 
    n12145 , 
    n12146 , 
    n12147 , 
    n12148 , 
    n12149 , 
    n12150 , 
    n12151 , 
    n12152 , 
    n12153 , 
    n12154 , 
    n12155 , 
    n12156 , 
    n12157 , 
    n12158 , 
    n12159 , 
    n12160 , 
    n12161 , 
    n12162 , 
    n12163 , 
    n12164 , 
    n12165 , 
    n12166 , 
    n12167 , 
    n12168 , 
    n12169 , 
    n12170 , 
    n12171 , 
    n12172 , 
    n12173 , 
    n12174 , 
    n12175 , 
    n12176 , 
    n12177 , 
    n12178 , 
    n12179 , 
    n12180 , 
    n12181 , 
    n12182 , 
    n12183 , 
    n12184 , 
    n12185 , 
    n12186 , 
    n12187 , 
    n12188 , 
    n12189 , 
    n12190 , 
    n12191 , 
    n12192 , 
    n12193 , 
    n12194 , 
    n12195 , 
    n12196 , 
    n12197 , 
    n12198 , 
    n12199 , 
    n12200 , 
    n12201 , 
    n12202 , 
    n12203 , 
    n12204 , 
    n12205 , 
    n12206 , 
    n12207 , 
    n12208 , 
    n12209 , 
    n12210 , 
    n12211 , 
    n12212 , 
    n12213 , 
    n12214 , 
    n12215 , 
    n12216 , 
    n12217 , 
    n12218 , 
    n12219 , 
    n12220 , 
    n12221 , 
    n12222 , 
    n12223 , 
    n12224 , 
    n12225 , 
    n12226 , 
    n12227 , 
    n12228 , 
    n12229 , 
    n12230 , 
    n12231 , 
    n12232 , 
    n12233 , 
    n12234 , 
    n12235 , 
    n12236 , 
    n12237 , 
    n12238 , 
    n12239 , 
    n12240 , 
    n12241 , 
    n12242 , 
    n12243 , 
    n12244 , 
    n12245 , 
    n12246 , 
    n12247 , 
    n12248 , 
    n12249 , 
    n12250 , 
    n12251 , 
    n12252 , 
    n12253 , 
    n12254 , 
    n12255 , 
    n12256 , 
    n12257 , 
    n12258 , 
    n12259 , 
    n12260 , 
    n12261 , 
    n12262 , 
    n12263 , 
    n12264 , 
    n12265 , 
    n12266 , 
    n12267 , 
    n12268 , 
    n12269 , 
    n12270 , 
    n12271 , 
    n12272 , 
    n12273 , 
    n12274 , 
    n12275 , 
    n12276 , 
    n12277 , 
    n12278 , 
    n12279 , 
    n12280 , 
    n12281 , 
    n12282 , 
    n12283 , 
    n12284 , 
    n12285 , 
    n12286 , 
    n12287 , 
    n12288 , 
    n12289 , 
    n12290 , 
    n12291 , 
    n12292 , 
    n12293 , 
    n12294 , 
    n12295 , 
    n12296 , 
    n12297 , 
    n12298 , 
    n12299 , 
    n12300 , 
    n12301 , 
    n12302 , 
    n12303 , 
    n12304 , 
    n12305 , 
    n12306 , 
    n12307 , 
    n12308 , 
    n12309 , 
    n12310 , 
    n12311 , 
    n12312 , 
    n12313 , 
    n12314 , 
    n12315 , 
    n12316 , 
    n12317 , 
    n12318 , 
    n12319 , 
    n12320 , 
    n12321 , 
    n12322 , 
    n12323 , 
    n12324 , 
    n12325 , 
    n12326 , 
    n12327 , 
    n12328 , 
    n12329 , 
    n12330 , 
    n12331 , 
    n12332 , 
    n12333 , 
    n12334 , 
    n12335 , 
    n12336 , 
    n12337 , 
    n12338 , 
    n12339 , 
    n12340 , 
    n12341 , 
    n12342 , 
    n12343 , 
    n12344 , 
    n12345 , 
    n12346 , 
    n12347 , 
    n12348 , 
    n12349 , 
    n12350 , 
    n12351 , 
    n12352 , 
    n12353 , 
    n12354 , 
    n12355 , 
    n12356 , 
    n12357 , 
    n12358 , 
    n12359 , 
    n12360 , 
    n12361 , 
    n12362 , 
    n12363 , 
    n12364 , 
    n12365 , 
    n12366 , 
    n12367 , 
    n12368 , 
    n12369 , 
    n12370 , 
    n12371 , 
    n12372 , 
    n12373 , 
    n12374 , 
    n12375 , 
    n12376 , 
    n12377 , 
    n12378 , 
    n12379 , 
    n12380 , 
    n12381 , 
    n12382 , 
    n12383 , 
    n12384 , 
    n12385 , 
    n12386 , 
    n12387 , 
    n12388 , 
    n12389 , 
    n12390 , 
    n12391 , 
    n12392 , 
    n12393 , 
    n12394 , 
    n12395 , 
    n12396 , 
    n12397 , 
    n12398 , 
    n12399 , 
    n12400 , 
    n12401 , 
    n12402 , 
    n12403 , 
    n12404 , 
    n12405 , 
    n12406 , 
    n12407 , 
    n12408 , 
    n12409 , 
    n12410 , 
    n12411 , 
    n12412 , 
    n12413 , 
    n12414 , 
    n12415 , 
    n12416 , 
    n12417 , 
    n12418 , 
    n12419 , 
    n12420 , 
    n12421 , 
    n12422 , 
    n12423 , 
    n12424 , 
    n12425 , 
    n12426 , 
    n12427 , 
    n12428 , 
    n12429 , 
    n12430 , 
    n12431 , 
    n12432 , 
    n12433 , 
    n12434 , 
    n12435 , 
    n12436 , 
    n12437 , 
    n12438 , 
    n12439 , 
    n12440 , 
    n12441 , 
    n12442 , 
    n12443 , 
    n12444 , 
    n12445 , 
    n12446 , 
    n12447 , 
    n12448 , 
    n12449 , 
    n12450 , 
    n12451 , 
    n12452 , 
    n12453 , 
    n12454 , 
    n12455 , 
    n12456 , 
    n12457 , 
    n12458 , 
    n12459 , 
    n12460 , 
    n12461 , 
    n12462 , 
    n12463 , 
    n12464 , 
    n12465 , 
    n12466 , 
    n12467 , 
    n12468 , 
    n12469 , 
    n12470 , 
    n12471 , 
    n12472 , 
    n12473 , 
    n12474 , 
    n12475 , 
    n12476 , 
    n12477 , 
    n12478 , 
    n12479 , 
    n12480 , 
    n12481 , 
    n12482 , 
    n12483 , 
    n12484 , 
    n12485 , 
    n12486 , 
    n12487 , 
    n12488 , 
    n12489 , 
    n12490 , 
    n12491 , 
    n12492 , 
    n12493 , 
    n12494 , 
    n12495 , 
    n12496 , 
    n12497 , 
    n12498 , 
    n12499 , 
    n12500 , 
    n12501 , 
    n12502 , 
    n12503 , 
    n12504 , 
    n12505 , 
    n12506 , 
    n12507 , 
    n12508 , 
    n12509 , 
    n12510 , 
    n12511 , 
    n12512 , 
    n12513 , 
    n12514 , 
    n12515 , 
    n12516 , 
    n12517 , 
    n12518 , 
    n12519 , 
    n12520 , 
    n12521 , 
    n12522 , 
    n12523 , 
    n12524 , 
    n12525 , 
    n12526 , 
    n12527 , 
    n12528 , 
    n12529 , 
    n12530 , 
    n12531 , 
    n12532 , 
    n12533 , 
    n12534 , 
    n12535 , 
    n12536 , 
    n12537 , 
    n12538 , 
    n12539 , 
    n12540 , 
    n12541 , 
    n12542 , 
    n12543 , 
    n12544 , 
    n12545 , 
    n12546 , 
    n12547 , 
    n12548 , 
    n12549 , 
    n12550 , 
    n12551 , 
    n12552 , 
    n12553 , 
    n12554 , 
    n12555 , 
    n12556 , 
    n12557 , 
    n12558 , 
    n12559 , 
    n12560 , 
    n12561 , 
    n12562 , 
    n12563 , 
    n12564 , 
    n12565 , 
    n12566 , 
    n12567 , 
    n12568 , 
    n12569 , 
    n12570 , 
    n12571 , 
    n12572 , 
    n12573 , 
    n12574 , 
    n12575 , 
    n12576 , 
    n12577 , 
    n12578 , 
    n12579 , 
    n12580 , 
    n12581 , 
    n12582 , 
    n12583 , 
    n12584 , 
    n12585 , 
    n12586 , 
    n12587 , 
    n12588 , 
    n12589 , 
    n12590 , 
    n12591 , 
    n12592 , 
    n12593 , 
    n12594 , 
    n12595 , 
    n12596 , 
    n12597 , 
    n12598 , 
    n12599 , 
    n12600 , 
    n12601 , 
    n12602 , 
    n12603 , 
    n12604 , 
    n12605 , 
    n12606 , 
    n12607 , 
    n12608 , 
    n12609 , 
    n12610 , 
    n12611 , 
    n12612 , 
    n12613 , 
    n12614 , 
    n12615 , 
    n12616 , 
    n12617 , 
    n12618 , 
    n12619 , 
    n12620 , 
    n12621 , 
    n12622 , 
    n12623 , 
    n12624 , 
    n12625 , 
    n12626 , 
    n12627 , 
    n12628 , 
    n12629 , 
    n12630 , 
    n12631 , 
    n12632 , 
    n12633 , 
    n12634 , 
    n12635 , 
    n12636 , 
    n12637 , 
    n12638 , 
    n12639 , 
    n12640 , 
    n12641 , 
    n12642 , 
    n12643 , 
    n12644 , 
    n12645 , 
    n12646 , 
    n12647 , 
    n12648 , 
    n12649 , 
    n12650 , 
    n12651 , 
    n12652 , 
    n12653 , 
    n12654 , 
    n12655 , 
    n12656 , 
    n12657 , 
    n12658 , 
    n12659 , 
    n12660 , 
    n12661 , 
    n12662 , 
    n12663 , 
    n12664 , 
    n12665 , 
    n12666 , 
    n12667 , 
    n12668 , 
    n12669 , 
    n12670 , 
    n12671 , 
    n12672 , 
    n12673 , 
    n12674 , 
    n12675 , 
    n12676 , 
    n12677 , 
    n12678 , 
    n12679 , 
    n12680 , 
    n12681 , 
    n12682 , 
    n12683 , 
    n12684 , 
    n12685 , 
    n12686 , 
    n12687 , 
    n12688 , 
    n12689 , 
    n12690 , 
    n12691 , 
    n12692 , 
    n12693 , 
    n12694 , 
    n12695 , 
    n12696 , 
    n12697 , 
    n12698 , 
    n12699 , 
    n12700 , 
    n12701 , 
    n12702 , 
    n12703 , 
    n12704 , 
    n12705 , 
    n12706 , 
    n12707 , 
    n12708 , 
    n12709 , 
    n12710 , 
    n12711 , 
    n12712 , 
    n12713 , 
    n12714 , 
    n12715 , 
    n12716 , 
    n12717 , 
    n12718 , 
    n12719 , 
    n12720 , 
    n12721 , 
    n12722 , 
    n12723 , 
    n12724 , 
    n12725 , 
    n12726 , 
    n12727 , 
    n12728 , 
    n12729 , 
    n12730 , 
    n12731 , 
    n12732 , 
    n12733 , 
    n12734 , 
    n12735 , 
    n12736 , 
    n12737 , 
    n12738 , 
    n12739 , 
    n12740 , 
    n12741 , 
    n12742 , 
    n12743 , 
    n12744 , 
    n12745 , 
    n12746 , 
    n12747 , 
    n12748 , 
    n12749 , 
    n12750 , 
    n12751 , 
    n12752 , 
    n12753 , 
    n12754 , 
    n12755 , 
    n12756 , 
    n12757 , 
    n12758 , 
    n12759 , 
    n12760 , 
    n12761 , 
    n12762 , 
    n12763 , 
    n12764 , 
    n12765 , 
    n12766 , 
    n12767 , 
    n12768 , 
    n12769 , 
    n12770 , 
    n12771 , 
    n12772 , 
    n12773 , 
    n12774 , 
    n12775 , 
    n12776 , 
    n12777 , 
    n12778 , 
    n12779 , 
    n12780 , 
    n12781 , 
    n12782 , 
    n12783 , 
    n12784 , 
    n12785 , 
    n12786 , 
    n12787 , 
    n12788 , 
    n12789 , 
    n12790 , 
    n12791 , 
    n12792 , 
    n12793 , 
    n12794 , 
    n12795 , 
    n12796 , 
    n12797 , 
    n12798 , 
    n12799 , 
    n12800 , 
    n12801 , 
    n12802 , 
    n12803 , 
    n12804 , 
    n12805 , 
    n12806 , 
    n12807 , 
    n12808 , 
    n12809 , 
    n12810 , 
    n12811 , 
    n12812 , 
    n12813 , 
    n12814 , 
    n12815 , 
    n12816 , 
    n12817 , 
    n12818 , 
    n12819 , 
    n12820 , 
    n12821 , 
    n12822 , 
    n12823 , 
    n12824 , 
    n12825 , 
    n12826 , 
    n12827 , 
    n12828 , 
    n12829 , 
    n12830 , 
    n12831 , 
    n12832 , 
    n12833 , 
    n12834 , 
    n12835 , 
    n12836 , 
    n12837 , 
    n12838 , 
    n12839 , 
    n12840 , 
    n12841 , 
    n12842 , 
    n12843 , 
    n12844 , 
    n12845 , 
    n12846 , 
    n12847 , 
    n12848 , 
    n12849 , 
    n12850 , 
    n12851 , 
    n12852 , 
    n12853 , 
    n12854 , 
    n12855 , 
    n12856 , 
    n12857 , 
    n12858 , 
    n12859 , 
    n12860 , 
    n12861 , 
    n12862 , 
    n12863 , 
    n12864 , 
    n12865 , 
    n12866 , 
    n12867 , 
    n12868 , 
    n12869 , 
    n12870 , 
    n12871 , 
    n12872 , 
    n12873 , 
    n12874 , 
    n12875 , 
    n12876 , 
    n12877 , 
    n12878 , 
    n12879 , 
    n12880 , 
    n12881 , 
    n12882 , 
    n12883 , 
    n12884 , 
    n12885 , 
    n12886 , 
    n12887 , 
    n12888 , 
    n12889 , 
    n12890 , 
    n12891 , 
    n12892 , 
    n12893 , 
    n12894 , 
    n12895 , 
    n12896 , 
    n12897 , 
    n12898 , 
    n12899 , 
    n12900 , 
    n12901 , 
    n12902 , 
    n12903 , 
    n12904 , 
    n12905 , 
    n12906 , 
    n12907 , 
    n12908 , 
    n12909 , 
    n12910 , 
    n12911 , 
    n12912 , 
    n12913 , 
    n12914 , 
    n12915 , 
    n12916 , 
    n12917 , 
    n12918 , 
    n12919 , 
    n12920 , 
    n12921 , 
    n12922 , 
    n12923 , 
    n12924 , 
    n12925 , 
    n12926 , 
    n12927 , 
    n12928 , 
    n12929 , 
    n12930 , 
    n12931 , 
    n12932 , 
    n12933 , 
    n12934 , 
    n12935 , 
    n12936 , 
    n12937 , 
    n12938 , 
    n12939 , 
    n12940 , 
    n12941 , 
    n12942 , 
    n12943 , 
    n12944 , 
    n12945 , 
    n12946 , 
    n12947 , 
    n12948 , 
    n12949 , 
    n12950 , 
    n12951 , 
    n12952 , 
    n12953 , 
    n12954 , 
    n12955 , 
    n12956 , 
    n12957 , 
    n12958 , 
    n12959 , 
    n12960 , 
    n12961 , 
    n12962 , 
    n12963 , 
    n12964 , 
    n12965 , 
    n12966 , 
    n12967 , 
    n12968 , 
    n12969 , 
    n12970 , 
    n12971 , 
    n12972 , 
    n12973 , 
    n12974 , 
    n12975 , 
    n12976 , 
    n12977 , 
    n12978 , 
    n12979 , 
    n12980 , 
    n12981 , 
    n12982 , 
    n12983 , 
    n12984 , 
    n12985 , 
    n12986 , 
    n12987 , 
    n12988 , 
    n12989 , 
    n12990 , 
    n12991 , 
    n12992 , 
    n12993 , 
    n12994 , 
    n12995 , 
    n12996 , 
    n12997 , 
    n12998 , 
    n12999 , 
    n13000 , 
    n13001 , 
    n13002 , 
    n13003 , 
    n13004 , 
    n13005 , 
    n13006 , 
    n13007 , 
    n13008 , 
    n13009 , 
    n13010 , 
    n13011 , 
    n13012 , 
    n13013 , 
    n13014 , 
    n13015 , 
    n13016 , 
    n13017 , 
    n13018 , 
    n13019 , 
    n13020 , 
    n13021 , 
    n13022 , 
    n13023 , 
    n13024 , 
    n13025 , 
    n13026 , 
    n13027 , 
    n13028 , 
    n13029 , 
    n13030 , 
    n13031 , 
    n13032 , 
    n13033 , 
    n13034 , 
    n13035 , 
    n13036 , 
    n13037 , 
    n13038 , 
    n13039 , 
    n13040 , 
    n13041 , 
    n13042 , 
    n13043 , 
    n13044 , 
    n13045 , 
    n13046 , 
    n13047 , 
    n13048 , 
    n13049 , 
    n13050 , 
    n13051 , 
    n13052 , 
    n13053 , 
    n13054 , 
    n13055 , 
    n13056 , 
    n13057 , 
    n13058 , 
    n13059 , 
    n13060 , 
    n13061 , 
    n13062 , 
    n13063 , 
    n13064 , 
    n13065 , 
    n13066 , 
    n13067 , 
    n13068 , 
    n13069 , 
    n13070 , 
    n13071 , 
    n13072 , 
    n13073 , 
    n13074 , 
    n13075 , 
    n13076 , 
    n13077 , 
    n13078 , 
    n13079 , 
    n13080 , 
    n13081 , 
    n13082 , 
    n13083 , 
    n13084 , 
    n13085 , 
    n13086 , 
    n13087 , 
    n13088 , 
    n13089 , 
    n13090 , 
    n13091 , 
    n13092 , 
    n13093 , 
    n13094 , 
    n13095 , 
    n13096 , 
    n13097 , 
    n13098 , 
    n13099 , 
    n13100 , 
    n13101 , 
    n13102 , 
    n13103 , 
    n13104 , 
    n13105 , 
    n13106 , 
    n13107 , 
    n13108 , 
    n13109 , 
    n13110 , 
    n13111 , 
    n13112 , 
    n13113 , 
    n13114 , 
    n13115 , 
    n13116 , 
    n13117 , 
    n13118 , 
    n13119 , 
    n13120 , 
    n13121 , 
    n13122 , 
    n13123 , 
    n13124 , 
    n13125 , 
    n13126 , 
    n13127 , 
    n13128 , 
    n13129 , 
    n13130 , 
    n13131 , 
    n13132 , 
    n13133 , 
    n13134 , 
    n13135 , 
    n13136 , 
    n13137 , 
    n13138 , 
    n13139 , 
    n13140 , 
    n13141 , 
    n13142 , 
    n13143 , 
    n13144 , 
    n13145 , 
    n13146 , 
    n13147 , 
    n13148 , 
    n13149 , 
    n13150 , 
    n13151 , 
    n13152 , 
    n13153 , 
    n13154 , 
    n13155 , 
    n13156 , 
    n13157 , 
    n13158 , 
    n13159 , 
    n13160 , 
    n13161 , 
    n13162 , 
    n13163 , 
    n13164 , 
    n13165 , 
    n13166 , 
    n13167 , 
    n13168 , 
    n13169 , 
    n13170 , 
    n13171 , 
    n13172 , 
    n13173 , 
    n13174 , 
    n13175 , 
    n13176 , 
    n13177 , 
    n13178 , 
    n13179 , 
    n13180 , 
    n13181 , 
    n13182 , 
    n13183 , 
    n13184 , 
    n13185 , 
    n13186 , 
    n13187 , 
    n13188 , 
    n13189 , 
    n13190 , 
    n13191 , 
    n13192 , 
    n13193 , 
    n13194 , 
    n13195 , 
    n13196 , 
    n13197 , 
    n13198 , 
    n13199 , 
    n13200 , 
    n13201 , 
    n13202 , 
    n13203 , 
    n13204 , 
    n13205 , 
    n13206 , 
    n13207 , 
    n13208 , 
    n13209 , 
    n13210 , 
    n13211 , 
    n13212 , 
    n13213 , 
    n13214 , 
    n13215 , 
    n13216 , 
    n13217 , 
    n13218 , 
    n13219 , 
    n13220 , 
    n13221 , 
    n13222 , 
    n13223 , 
    n13224 , 
    n13225 , 
    n13226 , 
    n13227 , 
    n13228 , 
    n13229 , 
    n13230 , 
    n13231 , 
    n13232 , 
    n13233 , 
    n13234 , 
    n13235 , 
    n13236 , 
    n13237 , 
    n13238 , 
    n13239 , 
    n13240 , 
    n13241 , 
    n13242 , 
    n13243 , 
    n13244 , 
    n13245 , 
    n13246 , 
    n13247 , 
    n13248 , 
    n13249 , 
    n13250 , 
    n13251 , 
    n13252 , 
    n13253 , 
    n13254 , 
    n13255 , 
    n13256 , 
    n13257 , 
    n13258 , 
    n13259 , 
    n13260 , 
    n13261 , 
    n13262 , 
    n13263 , 
    n13264 , 
    n13265 , 
    n13266 , 
    n13267 , 
    n13268 , 
    n13269 , 
    n13270 , 
    n13271 , 
    n13272 , 
    n13273 , 
    n13274 , 
    n13275 , 
    n13276 , 
    n13277 , 
    n13278 , 
    n13279 , 
    n13280 , 
    n13281 , 
    n13282 , 
    n13283 , 
    n13284 , 
    n13285 , 
    n13286 , 
    n13287 , 
    n13288 , 
    n13289 , 
    n13290 , 
    n13291 , 
    n13292 , 
    n13293 , 
    n13294 , 
    n13295 , 
    n13296 , 
    n13297 , 
    n13298 , 
    n13299 , 
    n13300 , 
    n13301 , 
    n13302 , 
    n13303 , 
    n13304 , 
    n13305 , 
    n13306 , 
    n13307 , 
    n13308 , 
    n13309 , 
    n13310 , 
    n13311 , 
    n13312 , 
    n13313 , 
    n13314 , 
    n13315 , 
    n13316 , 
    n13317 , 
    n13318 , 
    n13319 , 
    n13320 , 
    n13321 , 
    n13322 , 
    n13323 , 
    n13324 , 
    n13325 , 
    n13326 , 
    n13327 , 
    n13328 , 
    n13329 , 
    n13330 , 
    n13331 , 
    n13332 , 
    n13333 , 
    n13334 , 
    n13335 , 
    n13336 , 
    n13337 , 
    n13338 , 
    n13339 , 
    n13340 , 
    n13341 , 
    n13342 , 
    n13343 , 
    n13344 , 
    n13345 , 
    n13346 , 
    n13347 , 
    n13348 , 
    n13349 , 
    n13350 , 
    n13351 , 
    n13352 , 
    n13353 , 
    n13354 , 
    n13355 , 
    n13356 , 
    n13357 , 
    n13358 , 
    n13359 , 
    n13360 , 
    n13361 , 
    n13362 , 
    n13363 , 
    n13364 , 
    n13365 , 
    n13366 , 
    n13367 , 
    n13368 , 
    n13369 , 
    n13370 , 
    n13371 , 
    n13372 , 
    n13373 , 
    n13374 , 
    n13375 , 
    n13376 , 
    n13377 , 
    n13378 , 
    n13379 , 
    n13380 , 
    n13381 , 
    n13382 , 
    n13383 , 
    n13384 , 
    n13385 , 
    n13386 , 
    n13387 , 
    n13388 , 
    n13389 , 
    n13390 , 
    n13391 , 
    n13392 , 
    n13393 , 
    n13394 , 
    n13395 , 
    n13396 , 
    n13397 , 
    n13398 , 
    n13399 , 
    n13400 , 
    n13401 , 
    n13402 , 
    n13403 , 
    n13404 , 
    n13405 , 
    n13406 , 
    n13407 , 
    n13408 , 
    n13409 , 
    n13410 , 
    n13411 , 
    n13412 , 
    n13413 , 
    n13414 , 
    n13415 , 
    n13416 , 
    n13417 , 
    n13418 , 
    n13419 , 
    n13420 , 
    n13421 , 
    n13422 , 
    n13423 , 
    n13424 , 
    n13425 , 
    n13426 , 
    n13427 , 
    n13428 , 
    n13429 , 
    n13430 , 
    n13431 , 
    n13432 , 
    n13433 , 
    n13434 , 
    n13435 , 
    n13436 , 
    n13437 , 
    n13438 , 
    n13439 , 
    n13440 , 
    n13441 , 
    n13442 , 
    n13443 , 
    n13444 , 
    n13445 , 
    n13446 , 
    n13447 , 
    n13448 , 
    n13449 , 
    n13450 , 
    n13451 , 
    n13452 , 
    n13453 , 
    n13454 , 
    n13455 , 
    n13456 , 
    n13457 , 
    n13458 , 
    n13459 , 
    n13460 , 
    n13461 , 
    n13462 , 
    n13463 , 
    n13464 , 
    n13465 , 
    n13466 , 
    n13467 , 
    n13468 , 
    n13469 , 
    n13470 , 
    n13471 , 
    n13472 , 
    n13473 , 
    n13474 , 
    n13475 , 
    n13476 , 
    n13477 , 
    n13478 , 
    n13479 , 
    n13480 , 
    n13481 , 
    n13482 , 
    n13483 , 
    n13484 , 
    n13485 , 
    n13486 , 
    n13487 , 
    n13488 , 
    n13489 , 
    n13490 , 
    n13491 , 
    n13492 , 
    n13493 , 
    n13494 , 
    n13495 , 
    n13496 , 
    n13497 , 
    n13498 , 
    n13499 , 
    n13500 , 
    n13501 , 
    n13502 , 
    n13503 , 
    n13504 , 
    n13505 , 
    n13506 , 
    n13507 , 
    n13508 , 
    n13509 , 
    n13510 , 
    n13511 , 
    n13512 , 
    n13513 , 
    n13514 , 
    n13515 , 
    n13516 , 
    n13517 , 
    n13518 , 
    n13519 , 
    n13520 , 
    n13521 , 
    n13522 , 
    n13523 , 
    n13524 , 
    n13525 , 
    n13526 , 
    n13527 , 
    n13528 , 
    n13529 , 
    n13530 , 
    n13531 , 
    n13532 , 
    n13533 , 
    n13534 , 
    n13535 , 
    n13536 , 
    n13537 , 
    n13538 , 
    n13539 , 
    n13540 , 
    n13541 , 
    n13542 , 
    n13543 , 
    n13544 , 
    n13545 , 
    n13546 , 
    n13547 , 
    n13548 , 
    n13549 , 
    n13550 , 
    n13551 , 
    n13552 , 
    n13553 , 
    n13554 , 
    n13555 , 
    n13556 , 
    n13557 , 
    n13558 , 
    n13559 , 
    n13560 , 
    n13561 , 
    n13562 , 
    n13563 , 
    n13564 , 
    n13565 , 
    n13566 , 
    n13567 , 
    n13568 , 
    n13569 , 
    n13570 , 
    n13571 , 
    n13572 , 
    n13573 , 
    n13574 , 
    n13575 , 
    n13576 , 
    n13577 , 
    n13578 , 
    n13579 , 
    n13580 , 
    n13581 , 
    n13582 , 
    n13583 , 
    n13584 , 
    n13585 , 
    n13586 , 
    n13587 , 
    n13588 , 
    n13589 , 
    n13590 , 
    n13591 , 
    n13592 , 
    n13593 , 
    n13594 , 
    n13595 , 
    n13596 , 
    n13597 , 
    n13598 , 
    n13599 , 
    n13600 , 
    n13601 , 
    n13602 , 
    n13603 , 
    n13604 , 
    n13605 , 
    n13606 , 
    n13607 , 
    n13608 , 
    n13609 , 
    n13610 , 
    n13611 , 
    n13612 , 
    n13613 , 
    n13614 , 
    n13615 , 
    n13616 , 
    n13617 , 
    n13618 , 
    n13619 , 
    n13620 , 
    n13621 , 
    n13622 , 
    n13623 , 
    n13624 , 
    n13625 , 
    n13626 , 
    n13627 , 
    n13628 , 
    n13629 , 
    n13630 , 
    n13631 , 
    n13632 , 
    n13633 , 
    n13634 , 
    n13635 , 
    n13636 , 
    n13637 , 
    n13638 , 
    n13639 , 
    n13640 , 
    n13641 , 
    n13642 , 
    n13643 , 
    n13644 , 
    n13645 , 
    n13646 , 
    n13647 , 
    n13648 , 
    n13649 , 
    n13650 , 
    n13651 , 
    n13652 , 
    n13653 , 
    n13654 , 
    n13655 , 
    n13656 , 
    n13657 , 
    n13658 , 
    n13659 , 
    n13660 , 
    n13661 , 
    n13662 , 
    n13663 , 
    n13664 , 
    n13665 , 
    n13666 , 
    n13667 , 
    n13668 , 
    n13669 , 
    n13670 , 
    n13671 , 
    n13672 , 
    n13673 , 
    n13674 , 
    n13675 , 
    n13676 , 
    n13677 , 
    n13678 , 
    n13679 , 
    n13680 , 
    n13681 , 
    n13682 , 
    n13683 , 
    n13684 , 
    n13685 , 
    n13686 , 
    n13687 , 
    n13688 , 
    n13689 , 
    n13690 , 
    n13691 , 
    n13692 , 
    n13693 , 
    n13694 , 
    n13695 , 
    n13696 , 
    n13697 , 
    n13698 , 
    n13699 , 
    n13700 , 
    n13701 , 
    n13702 , 
    n13703 , 
    n13704 , 
    n13705 , 
    n13706 , 
    n13707 , 
    n13708 , 
    n13709 , 
    n13710 , 
    n13711 , 
    n13712 , 
    n13713 , 
    n13714 , 
    n13715 , 
    n13716 , 
    n13717 , 
    n13718 , 
    n13719 , 
    n13720 , 
    n13721 , 
    n13722 , 
    n13723 , 
    n13724 , 
    n13725 , 
    n13726 , 
    n13727 , 
    n13728 , 
    n13729 , 
    n13730 , 
    n13731 , 
    n13732 , 
    n13733 , 
    n13734 , 
    n13735 , 
    n13736 , 
    n13737 , 
    n13738 , 
    n13739 , 
    n13740 , 
    n13741 , 
    n13742 , 
    n13743 , 
    n13744 , 
    n13745 , 
    n13746 , 
    n13747 , 
    n13748 , 
    n13749 , 
    n13750 , 
    n13751 , 
    n13752 , 
    n13753 , 
    n13754 , 
    n13755 , 
    n13756 , 
    n13757 , 
    n13758 , 
    n13759 , 
    n13760 , 
    n13761 , 
    n13762 , 
    n13763 , 
    n13764 , 
    n13765 , 
    n13766 , 
    n13767 , 
    n13768 , 
    n13769 , 
    n13770 , 
    n13771 , 
    n13772 , 
    n13773 , 
    n13774 , 
    n13775 , 
    n13776 , 
    n13777 , 
    n13778 , 
    n13779 , 
    n13780 , 
    n13781 , 
    n13782 , 
    n13783 , 
    n13784 , 
    n13785 , 
    n13786 , 
    n13787 , 
    n13788 , 
    n13789 , 
    n13790 , 
    n13791 , 
    n13792 , 
    n13793 , 
    n13794 , 
    n13795 , 
    n13796 , 
    n13797 , 
    n13798 , 
    n13799 , 
    n13800 , 
    n13801 , 
    n13802 , 
    n13803 , 
    n13804 , 
    n13805 , 
    n13806 , 
    n13807 , 
    n13808 , 
    n13809 , 
    n13810 , 
    n13811 , 
    n13812 , 
    n13813 , 
    n13814 , 
    n13815 , 
    n13816 , 
    n13817 , 
    n13818 , 
    n13819 , 
    n13820 , 
    n13821 , 
    n13822 , 
    n13823 , 
    n13824 , 
    n13825 , 
    n13826 , 
    n13827 , 
    n13828 , 
    n13829 , 
    n13830 , 
    n13831 , 
    n13832 , 
    n13833 , 
    n13834 , 
    n13835 , 
    n13836 , 
    n13837 , 
    n13838 , 
    n13839 , 
    n13840 , 
    n13841 , 
    n13842 , 
    n13843 , 
    n13844 , 
    n13845 , 
    n13846 , 
    n13847 , 
    n13848 , 
    n13849 , 
    n13850 , 
    n13851 , 
    n13852 , 
    n13853 , 
    n13854 , 
    n13855 , 
    n13856 , 
    n13857 , 
    n13858 , 
    n13859 , 
    n13860 , 
    n13861 , 
    n13862 , 
    n13863 , 
    n13864 , 
    n13865 , 
    n13866 , 
    n13867 , 
    n13868 , 
    n13869 , 
    n13870 , 
    n13871 , 
    n13872 , 
    n13873 , 
    n13874 , 
    n13875 , 
    n13876 , 
    n13877 , 
    n13878 , 
    n13879 , 
    n13880 , 
    n13881 , 
    n13882 , 
    n13883 , 
    n13884 , 
    n13885 , 
    n13886 , 
    n13887 , 
    n13888 , 
    n13889 , 
    n13890 , 
    n13891 , 
    n13892 , 
    n13893 , 
    n13894 , 
    n13895 , 
    n13896 , 
    n13897 , 
    n13898 , 
    n13899 , 
    n13900 , 
    n13901 , 
    n13902 , 
    n13903 , 
    n13904 , 
    n13905 , 
    n13906 , 
    n13907 , 
    n13908 , 
    n13909 , 
    n13910 , 
    n13911 , 
    n13912 , 
    n13913 , 
    n13914 , 
    n13915 , 
    n13916 , 
    n13917 , 
    n13918 , 
    n13919 , 
    n13920 , 
    n13921 , 
    n13922 , 
    n13923 , 
    n13924 , 
    n13925 , 
    n13926 , 
    n13927 , 
    n13928 , 
    n13929 , 
    n13930 , 
    n13931 , 
    n13932 , 
    n13933 , 
    n13934 , 
    n13935 , 
    n13936 , 
    n13937 , 
    n13938 , 
    n13939 , 
    n13940 , 
    n13941 , 
    n13942 , 
    n13943 , 
    n13944 , 
    n13945 , 
    n13946 , 
    n13947 , 
    n13948 , 
    n13949 , 
    n13950 , 
    n13951 , 
    n13952 , 
    n13953 , 
    n13954 , 
    n13955 , 
    n13956 , 
    n13957 , 
    n13958 , 
    n13959 , 
    n13960 , 
    n13961 , 
    n13962 , 
    n13963 , 
    n13964 , 
    n13965 , 
    n13966 , 
    n13967 , 
    n13968 , 
    n13969 , 
    n13970 , 
    n13971 , 
    n13972 , 
    n13973 , 
    n13974 , 
    n13975 , 
    n13976 , 
    n13977 , 
    n13978 , 
    n13979 , 
    n13980 , 
    n13981 , 
    n13982 , 
    n13983 , 
    n13984 , 
    n13985 , 
    n13986 , 
    n13987 , 
    n13988 , 
    n13989 , 
    n13990 , 
    n13991 , 
    n13992 , 
    n13993 , 
    n13994 , 
    n13995 , 
    n13996 , 
    n13997 , 
    n13998 , 
    n13999 , 
    n14000 , 
    n14001 , 
    n14002 , 
    n14003 , 
    n14004 , 
    n14005 , 
    n14006 , 
    n14007 , 
    n14008 , 
    n14009 , 
    n14010 , 
    n14011 , 
    n14012 , 
    n14013 , 
    n14014 , 
    n14015 , 
    n14016 , 
    n14017 , 
    n14018 , 
    n14019 , 
    n14020 , 
    n14021 , 
    n14022 , 
    n14023 , 
    n14024 , 
    n14025 , 
    n14026 , 
    n14027 , 
    n14028 , 
    n14029 , 
    n14030 , 
    n14031 , 
    n14032 , 
    n14033 , 
    n14034 , 
    n14035 , 
    n14036 , 
    n14037 , 
    n14038 , 
    n14039 , 
    n14040 , 
    n14041 , 
    n14042 , 
    n14043 , 
    n14044 , 
    n14045 , 
    n14046 , 
    n14047 , 
    n14048 , 
    n14049 , 
    n14050 , 
    n14051 , 
    n14052 , 
    n14053 , 
    n14054 , 
    n14055 , 
    n14056 , 
    n14057 , 
    n14058 , 
    n14059 , 
    n14060 , 
    n14061 , 
    n14062 , 
    n14063 , 
    n14064 , 
    n14065 , 
    n14066 , 
    n14067 , 
    n14068 , 
    n14069 , 
    n14070 , 
    n14071 , 
    n14072 , 
    n14073 , 
    n14074 , 
    n14075 , 
    n14076 , 
    n14077 , 
    n14078 , 
    n14079 , 
    n14080 , 
    n14081 , 
    n14082 , 
    n14083 , 
    n14084 , 
    n14085 , 
    n14086 , 
    n14087 , 
    n14088 , 
    n14089 , 
    n14090 , 
    n14091 , 
    n14092 , 
    n14093 , 
    n14094 , 
    n14095 , 
    n14096 , 
    n14097 , 
    n14098 , 
    n14099 , 
    n14100 , 
    n14101 , 
    n14102 , 
    n14103 , 
    n14104 , 
    n14105 , 
    n14106 , 
    n14107 , 
    n14108 , 
    n14109 , 
    n14110 , 
    n14111 , 
    n14112 , 
    n14113 , 
    n14114 , 
    n14115 , 
    n14116 , 
    n14117 , 
    n14118 , 
    n14119 , 
    n14120 , 
    n14121 , 
    n14122 , 
    n14123 , 
    n14124 , 
    n14125 , 
    n14126 , 
    n14127 , 
    n14128 , 
    n14129 , 
    n14130 , 
    n14131 , 
    n14132 , 
    n14133 , 
    n14134 , 
    n14135 , 
    n14136 , 
    n14137 , 
    n14138 , 
    n14139 , 
    n14140 , 
    n14141 , 
    n14142 , 
    n14143 , 
    n14144 , 
    n14145 , 
    n14146 , 
    n14147 , 
    n14148 , 
    n14149 , 
    n14150 , 
    n14151 , 
    n14152 , 
    n14153 , 
    n14154 , 
    n14155 , 
    n14156 , 
    n14157 , 
    n14158 , 
    n14159 , 
    n14160 , 
    n14161 , 
    n14162 , 
    n14163 , 
    n14164 , 
    n14165 , 
    n14166 , 
    n14167 , 
    n14168 , 
    n14169 , 
    n14170 , 
    n14171 , 
    n14172 , 
    n14173 , 
    n14174 , 
    n14175 , 
    n14176 , 
    n14177 , 
    n14178 , 
    n14179 , 
    n14180 , 
    n14181 , 
    n14182 , 
    n14183 , 
    n14184 , 
    n14185 , 
    n14186 , 
    n14187 , 
    n14188 , 
    n14189 , 
    n14190 , 
    n14191 , 
    n14192 , 
    n14193 , 
    n14194 , 
    n14195 , 
    n14196 , 
    n14197 , 
    n14198 , 
    n14199 , 
    n14200 , 
    n14201 , 
    n14202 , 
    n14203 , 
    n14204 , 
    n14205 , 
    n14206 , 
    n14207 , 
    n14208 , 
    n14209 , 
    n14210 , 
    n14211 , 
    n14212 , 
    n14213 , 
    n14214 , 
    n14215 , 
    n14216 , 
    n14217 , 
    n14218 , 
    n14219 , 
    n14220 , 
    n14221 , 
    n14222 , 
    n14223 , 
    n14224 , 
    n14225 , 
    n14226 , 
    n14227 , 
    n14228 , 
    n14229 , 
    n14230 , 
    n14231 , 
    n14232 , 
    n14233 , 
    n14234 , 
    n14235 , 
    n14236 , 
    n14237 , 
    n14238 , 
    n14239 , 
    n14240 , 
    n14241 , 
    n14242 , 
    n14243 , 
    n14244 , 
    n14245 , 
    n14246 , 
    n14247 , 
    n14248 , 
    n14249 , 
    n14250 , 
    n14251 , 
    n14252 , 
    n14253 , 
    n14254 , 
    n14255 , 
    n14256 , 
    n14257 , 
    n14258 , 
    n14259 , 
    n14260 , 
    n14261 , 
    n14262 , 
    n14263 , 
    n14264 , 
    n14265 , 
    n14266 , 
    n14267 , 
    n14268 , 
    n14269 , 
    n14270 , 
    n14271 , 
    n14272 , 
    n14273 , 
    n14274 , 
    n14275 , 
    n14276 , 
    n14277 , 
    n14278 , 
    n14279 , 
    n14280 , 
    n14281 , 
    n14282 , 
    n14283 , 
    n14284 , 
    n14285 , 
    n14286 , 
    n14287 , 
    n14288 , 
    n14289 , 
    n14290 , 
    n14291 , 
    n14292 , 
    n14293 , 
    n14294 , 
    n14295 , 
    n14296 , 
    n14297 , 
    n14298 , 
    n14299 , 
    n14300 , 
    n14301 , 
    n14302 , 
    n14303 , 
    n14304 , 
    n14305 , 
    n14306 , 
    n14307 , 
    n14308 , 
    n14309 , 
    n14310 , 
    n14311 , 
    n14312 , 
    n14313 , 
    n14314 , 
    n14315 , 
    n14316 , 
    n14317 , 
    n14318 , 
    n14319 , 
    n14320 , 
    n14321 , 
    n14322 , 
    n14323 , 
    n14324 , 
    n14325 , 
    n14326 , 
    n14327 , 
    n14328 , 
    n14329 , 
    n14330 , 
    n14331 , 
    n14332 , 
    n14333 , 
    n14334 , 
    n14335 , 
    n14336 , 
    n14337 , 
    n14338 , 
    n14339 , 
    n14340 , 
    n14341 , 
    n14342 , 
    n14343 , 
    n14344 , 
    n14345 , 
    n14346 , 
    n14347 , 
    n14348 , 
    n14349 , 
    n14350 , 
    n14351 , 
    n14352 , 
    n14353 , 
    n14354 , 
    n14355 , 
    n14356 , 
    n14357 , 
    n14358 , 
    n14359 , 
    n14360 , 
    n14361 , 
    n14362 , 
    n14363 , 
    n14364 , 
    n14365 , 
    n14366 , 
    n14367 , 
    n14368 , 
    n14369 , 
    n14370 , 
    n14371 , 
    n14372 , 
    n14373 , 
    n14374 , 
    n14375 , 
    n14376 , 
    n14377 , 
    n14378 , 
    n14379 , 
    n14380 , 
    n14381 , 
    n14382 , 
    n14383 , 
    n14384 , 
    n14385 , 
    n14386 , 
    n14387 , 
    n14388 , 
    n14389 , 
    n14390 , 
    n14391 , 
    n14392 , 
    n14393 , 
    n14394 , 
    n14395 , 
    n14396 , 
    n14397 , 
    n14398 , 
    n14399 , 
    n14400 , 
    n14401 , 
    n14402 , 
    n14403 , 
    n14404 , 
    n14405 , 
    n14406 , 
    n14407 , 
    n14408 , 
    n14409 , 
    n14410 , 
    n14411 , 
    n14412 , 
    n14413 , 
    n14414 , 
    n14415 , 
    n14416 , 
    n14417 , 
    n14418 , 
    n14419 , 
    n14420 , 
    n14421 , 
    n14422 , 
    n14423 , 
    n14424 , 
    n14425 , 
    n14426 , 
    n14427 , 
    n14428 , 
    n14429 , 
    n14430 , 
    n14431 , 
    n14432 , 
    n14433 , 
    n14434 , 
    n14435 , 
    n14436 , 
    n14437 , 
    n14438 , 
    n14439 , 
    n14440 , 
    n14441 , 
    n14442 , 
    n14443 , 
    n14444 , 
    n14445 , 
    n14446 , 
    n14447 , 
    n14448 , 
    n14449 , 
    n14450 , 
    n14451 , 
    n14452 , 
    n14453 , 
    n14454 , 
    n14455 , 
    n14456 , 
    n14457 , 
    n14458 , 
    n14459 , 
    n14460 , 
    n14461 , 
    n14462 , 
    n14463 , 
    n14464 , 
    n14465 , 
    n14466 , 
    n14467 , 
    n14468 , 
    n14469 , 
    n14470 , 
    n14471 , 
    n14472 , 
    n14473 , 
    n14474 , 
    n14475 , 
    n14476 , 
    n14477 , 
    n14478 , 
    n14479 , 
    n14480 , 
    n14481 , 
    n14482 , 
    n14483 , 
    n14484 , 
    n14485 , 
    n14486 , 
    n14487 , 
    n14488 , 
    n14489 , 
    n14490 , 
    n14491 , 
    n14492 , 
    n14493 , 
    n14494 , 
    n14495 , 
    n14496 , 
    n14497 , 
    n14498 , 
    n14499 , 
    n14500 , 
    n14501 , 
    n14502 , 
    n14503 , 
    n14504 , 
    n14505 , 
    n14506 , 
    n14507 , 
    n14508 , 
    n14509 , 
    n14510 , 
    n14511 , 
    n14512 , 
    n14513 , 
    n14514 , 
    n14515 , 
    n14516 , 
    n14517 , 
    n14518 , 
    n14519 , 
    n14520 , 
    n14521 , 
    n14522 , 
    n14523 , 
    n14524 , 
    n14525 , 
    n14526 , 
    n14527 , 
    n14528 , 
    n14529 , 
    n14530 , 
    n14531 , 
    n14532 , 
    n14533 , 
    n14534 , 
    n14535 , 
    n14536 , 
    n14537 , 
    n14538 , 
    n14539 , 
    n14540 , 
    n14541 , 
    n14542 , 
    n14543 , 
    n14544 , 
    n14545 , 
    n14546 , 
    n14547 , 
    n14548 , 
    n14549 , 
    n14550 , 
    n14551 , 
    n14552 , 
    n14553 , 
    n14554 , 
    n14555 , 
    n14556 , 
    n14557 , 
    n14558 , 
    n14559 , 
    n14560 , 
    n14561 , 
    n14562 , 
    n14563 , 
    n14564 , 
    n14565 , 
    n14566 , 
    n14567 , 
    n14568 , 
    n14569 , 
    n14570 , 
    n14571 , 
    n14572 , 
    n14573 , 
    n14574 , 
    n14575 , 
    n14576 , 
    n14577 , 
    n14578 , 
    n14579 , 
    n14580 , 
    n14581 , 
    n14582 , 
    n14583 , 
    n14584 , 
    n14585 , 
    n14586 , 
    n14587 , 
    n14588 , 
    n14589 , 
    n14590 , 
    n14591 , 
    n14592 , 
    n14593 , 
    n14594 , 
    n14595 , 
    n14596 , 
    n14597 , 
    n14598 , 
    n14599 , 
    n14600 , 
    n14601 , 
    n14602 , 
    n14603 , 
    n14604 , 
    n14605 , 
    n14606 , 
    n14607 , 
    n14608 , 
    n14609 , 
    n14610 , 
    n14611 , 
    n14612 , 
    n14613 , 
    n14614 , 
    n14615 , 
    n14616 , 
    n14617 , 
    n14618 , 
    n14619 , 
    n14620 , 
    n14621 , 
    n14622 , 
    n14623 , 
    n14624 , 
    n14625 , 
    n14626 , 
    n14627 , 
    n14628 , 
    n14629 , 
    n14630 , 
    n14631 , 
    n14632 , 
    n14633 , 
    n14634 , 
    n14635 , 
    n14636 , 
    n14637 , 
    n14638 , 
    n14639 , 
    n14640 , 
    n14641 , 
    n14642 , 
    n14643 , 
    n14644 , 
    n14645 , 
    n14646 , 
    n14647 , 
    n14648 , 
    n14649 , 
    n14650 , 
    n14651 , 
    n14652 , 
    n14653 , 
    n14654 , 
    n14655 , 
    n14656 , 
    n14657 , 
    n14658 , 
    n14659 , 
    n14660 , 
    n14661 , 
    n14662 , 
    n14663 , 
    n14664 , 
    n14665 , 
    n14666 , 
    n14667 , 
    n14668 , 
    n14669 , 
    n14670 , 
    n14671 , 
    n14672 , 
    n14673 , 
    n14674 , 
    n14675 , 
    n14676 , 
    n14677 , 
    n14678 , 
    n14679 , 
    n14680 , 
    n14681 , 
    n14682 , 
    n14683 , 
    n14684 , 
    n14685 , 
    n14686 , 
    n14687 , 
    n14688 , 
    n14689 , 
    n14690 , 
    n14691 , 
    n14692 , 
    n14693 , 
    n14694 , 
    n14695 , 
    n14696 , 
    n14697 , 
    n14698 , 
    n14699 , 
    n14700 , 
    n14701 , 
    n14702 , 
    n14703 , 
    n14704 , 
    n14705 , 
    n14706 , 
    n14707 , 
    n14708 , 
    n14709 , 
    n14710 , 
    n14711 , 
    n14712 , 
    n14713 , 
    n14714 , 
    n14715 , 
    n14716 , 
    n14717 , 
    n14718 , 
    n14719 , 
    n14720 , 
    n14721 , 
    n14722 , 
    n14723 , 
    n14724 , 
    n14725 , 
    n14726 , 
    n14727 , 
    n14728 , 
    n14729 , 
    n14730 , 
    n14731 , 
    n14732 , 
    n14733 , 
    n14734 , 
    n14735 , 
    n14736 , 
    n14737 , 
    n14738 , 
    n14739 , 
    n14740 , 
    n14741 , 
    n14742 , 
    n14743 , 
    n14744 , 
    n14745 , 
    n14746 , 
    n14747 , 
    n14748 , 
    n14749 , 
    n14750 , 
    n14751 , 
    n14752 , 
    n14753 , 
    n14754 , 
    n14755 , 
    n14756 , 
    n14757 , 
    n14758 , 
    n14759 , 
    n14760 , 
    n14761 , 
    n14762 , 
    n14763 , 
    n14764 , 
    n14765 , 
    n14766 , 
    n14767 , 
    n14768 , 
    n14769 , 
    n14770 , 
    n14771 , 
    n14772 , 
    n14773 , 
    n14774 , 
    n14775 , 
    n14776 , 
    n14777 , 
    n14778 , 
    n14779 , 
    n14780 , 
    n14781 , 
    n14782 , 
    n14783 , 
    n14784 , 
    n14785 , 
    n14786 , 
    n14787 , 
    n14788 , 
    n14789 , 
    n14790 , 
    n14791 , 
    n14792 , 
    n14793 , 
    n14794 , 
    n14795 , 
    n14796 , 
    n14797 , 
    n14798 , 
    n14799 , 
    n14800 , 
    n14801 , 
    n14802 , 
    n14803 , 
    n14804 , 
    n14805 , 
    n14806 , 
    n14807 , 
    n14808 , 
    n14809 , 
    n14810 , 
    n14811 , 
    n14812 , 
    n14813 , 
    n14814 , 
    n14815 , 
    n14816 , 
    n14817 , 
    n14818 , 
    n14819 , 
    n14820 , 
    n14821 , 
    n14822 , 
    n14823 , 
    n14824 , 
    n14825 , 
    n14826 , 
    n14827 , 
    n14828 , 
    n14829 , 
    n14830 , 
    n14831 , 
    n14832 , 
    n14833 , 
    n14834 , 
    n14835 , 
    n14836 , 
    n14837 , 
    n14838 , 
    n14839 , 
    n14840 , 
    n14841 , 
    n14842 , 
    n14843 , 
    n14844 , 
    n14845 , 
    n14846 , 
    n14847 , 
    n14848 , 
    n14849 , 
    n14850 , 
    n14851 , 
    n14852 , 
    n14853 , 
    n14854 , 
    n14855 , 
    n14856 , 
    n14857 , 
    n14858 , 
    n14859 , 
    n14860 , 
    n14861 , 
    n14862 , 
    n14863 , 
    n14864 , 
    n14865 , 
    n14866 , 
    n14867 , 
    n14868 , 
    n14869 , 
    n14870 , 
    n14871 , 
    n14872 , 
    n14873 , 
    n14874 , 
    n14875 , 
    n14876 , 
    n14877 , 
    n14878 , 
    n14879 , 
    n14880 , 
    n14881 , 
    n14882 , 
    n14883 , 
    n14884 , 
    n14885 , 
    n14886 , 
    n14887 , 
    n14888 , 
    n14889 , 
    n14890 , 
    n14891 , 
    n14892 , 
    n14893 , 
    n14894 , 
    n14895 , 
    n14896 , 
    n14897 , 
    n14898 , 
    n14899 , 
    n14900 , 
    n14901 , 
    n14902 , 
    n14903 , 
    n14904 , 
    n14905 , 
    n14906 , 
    n14907 , 
    n14908 , 
    n14909 , 
    n14910 , 
    n14911 , 
    n14912 , 
    n14913 , 
    n14914 , 
    n14915 , 
    n14916 , 
    n14917 , 
    n14918 , 
    n14919 , 
    n14920 , 
    n14921 , 
    n14922 , 
    n14923 , 
    n14924 , 
    n14925 , 
    n14926 , 
    n14927 , 
    n14928 , 
    n14929 , 
    n14930 , 
    n14931 , 
    n14932 , 
    n14933 , 
    n14934 , 
    n14935 , 
    n14936 , 
    n14937 , 
    n14938 , 
    n14939 , 
    n14940 , 
    n14941 , 
    n14942 , 
    n14943 , 
    n14944 , 
    n14945 , 
    n14946 , 
    n14947 , 
    n14948 , 
    n14949 , 
    n14950 , 
    n14951 , 
    n14952 , 
    n14953 , 
    n14954 , 
    n14955 , 
    n14956 , 
    n14957 , 
    n14958 , 
    n14959 , 
    n14960 , 
    n14961 , 
    n14962 , 
    n14963 , 
    n14964 , 
    n14965 , 
    n14966 , 
    n14967 , 
    n14968 , 
    n14969 , 
    n14970 , 
    n14971 , 
    n14972 , 
    n14973 , 
    n14974 , 
    n14975 , 
    n14976 , 
    n14977 , 
    n14978 , 
    n14979 , 
    n14980 , 
    n14981 , 
    n14982 , 
    n14983 , 
    n14984 , 
    n14985 , 
    n14986 , 
    n14987 , 
    n14988 , 
    n14989 , 
    n14990 , 
    n14991 , 
    n14992 , 
    n14993 , 
    n14994 , 
    n14995 , 
    n14996 , 
    n14997 , 
    n14998 , 
    n14999 , 
    n15000 , 
    n15001 , 
    n15002 , 
    n15003 , 
    n15004 , 
    n15005 , 
    n15006 , 
    n15007 , 
    n15008 , 
    n15009 , 
    n15010 , 
    n15011 , 
    n15012 , 
    n15013 , 
    n15014 , 
    n15015 , 
    n15016 , 
    n15017 , 
    n15018 , 
    n15019 , 
    n15020 , 
    n15021 , 
    n15022 , 
    n15023 , 
    n15024 , 
    n15025 , 
    n15026 , 
    n15027 , 
    n15028 , 
    n15029 , 
    n15030 , 
    n15031 , 
    n15032 , 
    n15033 , 
    n15034 , 
    n15035 , 
    n15036 , 
    n15037 , 
    n15038 , 
    n15039 , 
    n15040 , 
    n15041 , 
    n15042 , 
    n15043 , 
    n15044 , 
    n15045 , 
    n15046 , 
    n15047 , 
    n15048 , 
    n15049 , 
    n15050 , 
    n15051 , 
    n15052 , 
    n15053 , 
    n15054 , 
    n15055 , 
    n15056 , 
    n15057 , 
    n15058 , 
    n15059 , 
    n15060 , 
    n15061 , 
    n15062 , 
    n15063 , 
    n15064 , 
    n15065 , 
    n15066 , 
    n15067 , 
    n15068 , 
    n15069 , 
    n15070 , 
    n15071 , 
    n15072 , 
    n15073 , 
    n15074 , 
    n15075 , 
    n15076 , 
    n15077 , 
    n15078 , 
    n15079 , 
    n15080 , 
    n15081 , 
    n15082 , 
    n15083 , 
    n15084 , 
    n15085 , 
    n15086 , 
    n15087 , 
    n15088 , 
    n15089 , 
    n15090 , 
    n15091 , 
    n15092 , 
    n15093 , 
    n15094 , 
    n15095 , 
    n15096 , 
    n15097 , 
    n15098 , 
    n15099 , 
    n15100 , 
    n15101 , 
    n15102 , 
    n15103 , 
    n15104 , 
    n15105 , 
    n15106 , 
    n15107 , 
    n15108 , 
    n15109 , 
    n15110 , 
    n15111 , 
    n15112 , 
    n15113 , 
    n15114 , 
    n15115 , 
    n15116 , 
    n15117 , 
    n15118 , 
    n15119 , 
    n15120 , 
    n15121 , 
    n15122 , 
    n15123 , 
    n15124 , 
    n15125 , 
    n15126 , 
    n15127 , 
    n15128 , 
    n15129 , 
    n15130 , 
    n15131 , 
    n15132 , 
    n15133 , 
    n15134 , 
    n15135 , 
    n15136 , 
    n15137 , 
    n15138 , 
    n15139 , 
    n15140 , 
    n15141 , 
    n15142 , 
    n15143 , 
    n15144 , 
    n15145 , 
    n15146 , 
    n15147 , 
    n15148 , 
    n15149 , 
    n15150 , 
    n15151 , 
    n15152 , 
    n15153 , 
    n15154 , 
    n15155 , 
    n15156 , 
    n15157 , 
    n15158 , 
    n15159 , 
    n15160 , 
    n15161 , 
    n15162 , 
    n15163 , 
    n15164 , 
    n15165 , 
    n15166 , 
    n15167 , 
    n15168 , 
    n15169 , 
    n15170 , 
    n15171 , 
    n15172 , 
    n15173 , 
    n15174 , 
    n15175 , 
    n15176 , 
    n15177 , 
    n15178 , 
    n15179 , 
    n15180 , 
    n15181 , 
    n15182 , 
    n15183 , 
    n15184 , 
    n15185 , 
    n15186 , 
    n15187 , 
    n15188 , 
    n15189 , 
    n15190 , 
    n15191 , 
    n15192 , 
    n15193 , 
    n15194 , 
    n15195 , 
    n15196 , 
    n15197 , 
    n15198 , 
    n15199 , 
    n15200 , 
    n15201 , 
    n15202 , 
    n15203 , 
    n15204 , 
    n15205 , 
    n15206 , 
    n15207 , 
    n15208 , 
    n15209 , 
    n15210 , 
    n15211 , 
    n15212 , 
    n15213 , 
    n15214 , 
    n15215 , 
    n15216 , 
    n15217 , 
    n15218 , 
    n15219 , 
    n15220 , 
    n15221 , 
    n15222 , 
    n15223 , 
    n15224 , 
    n15225 , 
    n15226 , 
    n15227 , 
    n15228 , 
    n15229 , 
    n15230 , 
    n15231 , 
    n15232 , 
    n15233 , 
    n15234 , 
    n15235 , 
    n15236 , 
    n15237 , 
    n15238 , 
    n15239 , 
    n15240 , 
    n15241 , 
    n15242 , 
    n15243 , 
    n15244 , 
    n15245 , 
    n15246 , 
    n15247 , 
    n15248 , 
    n15249 , 
    n15250 , 
    n15251 , 
    n15252 , 
    n15253 , 
    n15254 , 
    n15255 , 
    n15256 , 
    n15257 , 
    n15258 , 
    n15259 , 
    n15260 , 
    n15261 , 
    n15262 , 
    n15263 , 
    n15264 , 
    n15265 , 
    n15266 , 
    n15267 , 
    n15268 , 
    n15269 , 
    n15270 , 
    n15271 , 
    n15272 , 
    n15273 , 
    n15274 , 
    n15275 , 
    n15276 , 
    n15277 , 
    n15278 , 
    n15279 , 
    n15280 , 
    n15281 , 
    n15282 , 
    n15283 , 
    n15284 , 
    n15285 , 
    n15286 , 
    n15287 , 
    n15288 , 
    n15289 , 
    n15290 , 
    n15291 , 
    n15292 , 
    n15293 , 
    n15294 , 
    n15295 , 
    n15296 , 
    n15297 , 
    n15298 , 
    n15299 , 
    n15300 , 
    n15301 , 
    n15302 , 
    n15303 , 
    n15304 , 
    n15305 , 
    n15306 , 
    n15307 , 
    n15308 , 
    n15309 , 
    n15310 , 
    n15311 , 
    n15312 , 
    n15313 , 
    n15314 , 
    n15315 , 
    n15316 , 
    n15317 , 
    n15318 , 
    n15319 , 
    n15320 , 
    n15321 , 
    n15322 , 
    n15323 , 
    n15324 , 
    n15325 , 
    n15326 , 
    n15327 , 
    n15328 , 
    n15329 , 
    n15330 , 
    n15331 , 
    n15332 , 
    n15333 , 
    n15334 , 
    n15335 , 
    n15336 , 
    n15337 , 
    n15338 , 
    n15339 , 
    n15340 , 
    n15341 , 
    n15342 , 
    n15343 , 
    n15344 , 
    n15345 , 
    n15346 , 
    n15347 , 
    n15348 , 
    n15349 , 
    n15350 , 
    n15351 , 
    n15352 , 
    n15353 , 
    n15354 , 
    n15355 , 
    n15356 , 
    n15357 , 
    n15358 , 
    n15359 , 
    n15360 , 
    n15361 , 
    n15362 , 
    n15363 , 
    n15364 , 
    n15365 , 
    n15366 , 
    n15367 , 
    n15368 , 
    n15369 , 
    n15370 , 
    n15371 , 
    n15372 , 
    n15373 , 
    n15374 , 
    n15375 , 
    n15376 , 
    n15377 , 
    n15378 , 
    n15379 , 
    n15380 , 
    n15381 , 
    n15382 , 
    n15383 , 
    n15384 , 
    n15385 , 
    n15386 , 
    n15387 , 
    n15388 , 
    n15389 , 
    n15390 , 
    n15391 , 
    n15392 , 
    n15393 , 
    n15394 , 
    n15395 , 
    n15396 , 
    n15397 , 
    n15398 , 
    n15399 , 
    n15400 , 
    n15401 , 
    n15402 , 
    n15403 , 
    n15404 , 
    n15405 , 
    n15406 , 
    n15407 , 
    n15408 , 
    n15409 , 
    n15410 , 
    n15411 , 
    n15412 , 
    n15413 , 
    n15414 , 
    n15415 , 
    n15416 , 
    n15417 , 
    n15418 , 
    n15419 , 
    n15420 , 
    n15421 , 
    n15422 , 
    n15423 , 
    n15424 , 
    n15425 , 
    n15426 , 
    n15427 , 
    n15428 , 
    n15429 , 
    n15430 , 
    n15431 , 
    n15432 , 
    n15433 , 
    n15434 , 
    n15435 , 
    n15436 , 
    n15437 , 
    n15438 , 
    n15439 , 
    n15440 , 
    n15441 , 
    n15442 , 
    n15443 , 
    n15444 , 
    n15445 , 
    n15446 , 
    n15447 , 
    n15448 , 
    n15449 , 
    n15450 , 
    n15451 , 
    n15452 , 
    n15453 , 
    n15454 , 
    n15455 , 
    n15456 , 
    n15457 , 
    n15458 , 
    n15459 , 
    n15460 , 
    n15461 , 
    n15462 , 
    n15463 , 
    n15464 , 
    n15465 , 
    n15466 , 
    n15467 , 
    n15468 , 
    n15469 , 
    n15470 , 
    n15471 , 
    n15472 , 
    n15473 , 
    n15474 , 
    n15475 , 
    n15476 , 
    n15477 , 
    n15478 , 
    n15479 , 
    n15480 , 
    n15481 , 
    n15482 , 
    n15483 , 
    n15484 , 
    n15485 , 
    n15486 , 
    n15487 , 
    n15488 , 
    n15489 , 
    n15490 , 
    n15491 , 
    n15492 , 
    n15493 , 
    n15494 , 
    n15495 , 
    n15496 , 
    n15497 , 
    n15498 , 
    n15499 , 
    n15500 , 
    n15501 , 
    n15502 , 
    n15503 , 
    n15504 , 
    n15505 , 
    n15506 , 
    n15507 , 
    n15508 , 
    n15509 , 
    n15510 , 
    n15511 , 
    n15512 , 
    n15513 , 
    n15514 , 
    n15515 , 
    n15516 , 
    n15517 , 
    n15518 , 
    n15519 , 
    n15520 , 
    n15521 , 
    n15522 , 
    n15523 , 
    n15524 , 
    n15525 , 
    n15526 , 
    n15527 , 
    n15528 , 
    n15529 , 
    n15530 , 
    n15531 , 
    n15532 , 
    n15533 , 
    n15534 , 
    n15535 , 
    n15536 , 
    n15537 , 
    n15538 , 
    n15539 , 
    n15540 , 
    n15541 , 
    n15542 , 
    n15543 , 
    n15544 , 
    n15545 , 
    n15546 , 
    n15547 , 
    n15548 , 
    n15549 , 
    n15550 , 
    n15551 , 
    n15552 , 
    n15553 , 
    n15554 , 
    n15555 , 
    n15556 , 
    n15557 , 
    n15558 , 
    n15559 , 
    n15560 , 
    n15561 , 
    n15562 , 
    n15563 , 
    n15564 , 
    n15565 , 
    n15566 , 
    n15567 , 
    n15568 , 
    n15569 , 
    n15570 , 
    n15571 , 
    n15572 , 
    n15573 , 
    n15574 , 
    n15575 , 
    n15576 , 
    n15577 , 
    n15578 , 
    n15579 , 
    n15580 , 
    n15581 , 
    n15582 , 
    n15583 , 
    n15584 , 
    n15585 , 
    n15586 , 
    n15587 , 
    n15588 , 
    n15589 , 
    n15590 , 
    n15591 , 
    n15592 , 
    n15593 , 
    n15594 , 
    n15595 , 
    n15596 , 
    n15597 , 
    n15598 , 
    n15599 , 
    n15600 , 
    n15601 , 
    n15602 , 
    n15603 , 
    n15604 , 
    n15605 , 
    n15606 , 
    n15607 , 
    n15608 , 
    n15609 , 
    n15610 , 
    n15611 , 
    n15612 , 
    n15613 , 
    n15614 , 
    n15615 , 
    n15616 , 
    n15617 , 
    n15618 , 
    n15619 , 
    n15620 , 
    n15621 , 
    n15622 , 
    n15623 , 
    n15624 , 
    n15625 , 
    n15626 , 
    n15627 , 
    n15628 , 
    n15629 , 
    n15630 , 
    n15631 , 
    n15632 , 
    n15633 , 
    n15634 , 
    n15635 , 
    n15636 , 
    n15637 , 
    n15638 , 
    n15639 , 
    n15640 , 
    n15641 , 
    n15642 , 
    n15643 , 
    n15644 , 
    n15645 , 
    n15646 , 
    n15647 , 
    n15648 , 
    n15649 , 
    n15650 , 
    n15651 , 
    n15652 , 
    n15653 , 
    n15654 , 
    n15655 , 
    n15656 , 
    n15657 , 
    n15658 , 
    n15659 , 
    n15660 , 
    n15661 , 
    n15662 , 
    n15663 , 
    n15664 , 
    n15665 , 
    n15666 , 
    n15667 , 
    n15668 , 
    n15669 , 
    n15670 , 
    n15671 , 
    n15672 , 
    n15673 , 
    n15674 , 
    n15675 , 
    n15676 , 
    n15677 , 
    n15678 , 
    n15679 , 
    n15680 , 
    n15681 , 
    n15682 , 
    n15683 , 
    n15684 , 
    n15685 , 
    n15686 , 
    n15687 , 
    n15688 , 
    n15689 , 
    n15690 , 
    n15691 , 
    n15692 , 
    n15693 , 
    n15694 , 
    n15695 , 
    n15696 , 
    n15697 , 
    n15698 , 
    n15699 , 
    n15700 , 
    n15701 , 
    n15702 , 
    n15703 , 
    n15704 , 
    n15705 , 
    n15706 , 
    n15707 , 
    n15708 , 
    n15709 , 
    n15710 , 
    n15711 , 
    n15712 , 
    n15713 , 
    n15714 , 
    n15715 , 
    n15716 , 
    n15717 , 
    n15718 , 
    n15719 , 
    n15720 , 
    n15721 , 
    n15722 , 
    n15723 , 
    n15724 , 
    n15725 , 
    n15726 , 
    n15727 , 
    n15728 , 
    n15729 , 
    n15730 , 
    n15731 , 
    n15732 , 
    n15733 , 
    n15734 , 
    n15735 , 
    n15736 , 
    n15737 , 
    n15738 , 
    n15739 , 
    n15740 , 
    n15741 , 
    n15742 , 
    n15743 , 
    n15744 , 
    n15745 , 
    n15746 , 
    n15747 , 
    n15748 , 
    n15749 , 
    n15750 , 
    n15751 , 
    n15752 , 
    n15753 , 
    n15754 , 
    n15755 , 
    n15756 , 
    n15757 , 
    n15758 , 
    n15759 , 
    n15760 , 
    n15761 , 
    n15762 , 
    n15763 , 
    n15764 , 
    n15765 , 
    n15766 , 
    n15767 , 
    n15768 , 
    n15769 , 
    n15770 , 
    n15771 , 
    n15772 , 
    n15773 , 
    n15774 , 
    n15775 , 
    n15776 , 
    n15777 , 
    n15778 , 
    n15779 , 
    n15780 , 
    n15781 , 
    n15782 , 
    n15783 , 
    n15784 , 
    n15785 , 
    n15786 , 
    n15787 , 
    n15788 , 
    n15789 , 
    n15790 , 
    n15791 , 
    n15792 , 
    n15793 , 
    n15794 , 
    n15795 , 
    n15796 , 
    n15797 , 
    n15798 , 
    n15799 , 
    n15800 , 
    n15801 , 
    n15802 , 
    n15803 , 
    n15804 , 
    n15805 , 
    n15806 , 
    n15807 , 
    n15808 , 
    n15809 , 
    n15810 , 
    n15811 , 
    n15812 , 
    n15813 , 
    n15814 , 
    n15815 , 
    n15816 , 
    n15817 , 
    n15818 , 
    n15819 , 
    n15820 , 
    n15821 , 
    n15822 , 
    n15823 , 
    n15824 , 
    n15825 , 
    n15826 , 
    n15827 , 
    n15828 , 
    n15829 , 
    n15830 , 
    n15831 , 
    n15832 , 
    n15833 , 
    n15834 , 
    n15835 , 
    n15836 , 
    n15837 , 
    n15838 , 
    n15839 , 
    n15840 , 
    n15841 , 
    n15842 , 
    n15843 , 
    n15844 , 
    n15845 , 
    n15846 , 
    n15847 , 
    n15848 , 
    n15849 , 
    n15850 , 
    n15851 , 
    n15852 , 
    n15853 , 
    n15854 , 
    n15855 , 
    n15856 , 
    n15857 , 
    n15858 , 
    n15859 , 
    n15860 , 
    n15861 , 
    n15862 , 
    n15863 , 
    n15864 , 
    n15865 , 
    n15866 , 
    n15867 , 
    n15868 , 
    n15869 , 
    n15870 , 
    n15871 , 
    n15872 , 
    n15873 , 
    n15874 , 
    n15875 , 
    n15876 , 
    n15877 , 
    n15878 , 
    n15879 , 
    n15880 , 
    n15881 , 
    n15882 , 
    n15883 , 
    n15884 , 
    n15885 , 
    n15886 , 
    n15887 , 
    n15888 , 
    n15889 , 
    n15890 , 
    n15891 , 
    n15892 , 
    n15893 , 
    n15894 , 
    n15895 , 
    n15896 , 
    n15897 , 
    n15898 , 
    n15899 , 
    n15900 , 
    n15901 , 
    n15902 , 
    n15903 , 
    n15904 , 
    n15905 , 
    n15906 , 
    n15907 , 
    n15908 , 
    n15909 , 
    n15910 , 
    n15911 , 
    n15912 , 
    n15913 , 
    n15914 , 
    n15915 , 
    n15916 , 
    n15917 , 
    n15918 , 
    n15919 , 
    n15920 , 
    n15921 , 
    n15922 , 
    n15923 , 
    n15924 , 
    n15925 , 
    n15926 , 
    n15927 , 
    n15928 , 
    n15929 , 
    n15930 , 
    n15931 , 
    n15932 , 
    n15933 , 
    n15934 , 
    n15935 , 
    n15936 , 
    n15937 , 
    n15938 , 
    n15939 , 
    n15940 , 
    n15941 , 
    n15942 , 
    n15943 , 
    n15944 , 
    n15945 , 
    n15946 , 
    n15947 , 
    n15948 , 
    n15949 , 
    n15950 , 
    n15951 , 
    n15952 , 
    n15953 , 
    n15954 , 
    n15955 , 
    n15956 , 
    n15957 , 
    n15958 , 
    n15959 , 
    n15960 , 
    n15961 , 
    n15962 , 
    n15963 , 
    n15964 , 
    n15965 , 
    n15966 , 
    n15967 , 
    n15968 , 
    n15969 , 
    n15970 , 
    n15971 , 
    n15972 , 
    n15973 , 
    n15974 , 
    n15975 , 
    n15976 , 
    n15977 , 
    n15978 , 
    n15979 , 
    n15980 , 
    n15981 , 
    n15982 , 
    n15983 , 
    n15984 , 
    n15985 , 
    n15986 , 
    n15987 , 
    n15988 , 
    n15989 , 
    n15990 , 
    n15991 , 
    n15992 , 
    n15993 , 
    n15994 , 
    n15995 , 
    n15996 , 
    n15997 , 
    n15998 , 
    n15999 , 
    n16000 , 
    n16001 , 
    n16002 , 
    n16003 , 
    n16004 , 
    n16005 , 
    n16006 , 
    n16007 , 
    n16008 , 
    n16009 , 
    n16010 , 
    n16011 , 
    n16012 , 
    n16013 , 
    n16014 , 
    n16015 , 
    n16016 , 
    n16017 , 
    n16018 , 
    n16019 , 
    n16020 , 
    n16021 , 
    n16022 , 
    n16023 , 
    n16024 , 
    n16025 , 
    n16026 , 
    n16027 , 
    n16028 , 
    n16029 , 
    n16030 , 
    n16031 , 
    n16032 , 
    n16033 , 
    n16034 , 
    n16035 , 
    n16036 , 
    n16037 , 
    n16038 , 
    n16039 , 
    n16040 , 
    n16041 , 
    n16042 , 
    n16043 , 
    n16044 , 
    n16045 , 
    n16046 , 
    n16047 , 
    n16048 , 
    n16049 , 
    n16050 , 
    n16051 , 
    n16052 , 
    n16053 , 
    n16054 , 
    n16055 , 
    n16056 , 
    n16057 , 
    n16058 , 
    n16059 , 
    n16060 , 
    n16061 , 
    n16062 , 
    n16063 , 
    n16064 , 
    n16065 , 
    n16066 , 
    n16067 , 
    n16068 , 
    n16069 , 
    n16070 , 
    n16071 , 
    n16072 , 
    n16073 , 
    n16074 , 
    n16075 , 
    n16076 , 
    n16077 , 
    n16078 , 
    n16079 , 
    n16080 , 
    n16081 , 
    n16082 , 
    n16083 , 
    n16084 , 
    n16085 , 
    n16086 , 
    n16087 , 
    n16088 , 
    n16089 , 
    n16090 , 
    n16091 , 
    n16092 , 
    n16093 , 
    n16094 , 
    n16095 , 
    n16096 , 
    n16097 , 
    n16098 , 
    n16099 , 
    n16100 , 
    n16101 , 
    n16102 , 
    n16103 , 
    n16104 , 
    n16105 , 
    n16106 , 
    n16107 , 
    n16108 , 
    n16109 , 
    n16110 , 
    n16111 , 
    n16112 , 
    n16113 , 
    n16114 , 
    n16115 , 
    n16116 , 
    n16117 , 
    n16118 , 
    n16119 , 
    n16120 , 
    n16121 , 
    n16122 , 
    n16123 , 
    n16124 , 
    n16125 , 
    n16126 , 
    n16127 , 
    n16128 , 
    n16129 , 
    n16130 , 
    n16131 , 
    n16132 , 
    n16133 , 
    n16134 , 
    n16135 , 
    n16136 , 
    n16137 , 
    n16138 , 
    n16139 , 
    n16140 , 
    n16141 , 
    n16142 , 
    n16143 , 
    n16144 , 
    n16145 , 
    n16146 , 
    n16147 , 
    n16148 , 
    n16149 , 
    n16150 , 
    n16151 , 
    n16152 , 
    n16153 , 
    n16154 , 
    n16155 , 
    n16156 , 
    n16157 , 
    n16158 , 
    n16159 , 
    n16160 , 
    n16161 , 
    n16162 , 
    n16163 , 
    n16164 , 
    n16165 , 
    n16166 , 
    n16167 , 
    n16168 , 
    n16169 , 
    n16170 , 
    n16171 , 
    n16172 , 
    n16173 , 
    n16174 , 
    n16175 , 
    n16176 , 
    n16177 , 
    n16178 , 
    n16179 , 
    n16180 , 
    n16181 , 
    n16182 , 
    n16183 , 
    n16184 , 
    n16185 , 
    n16186 , 
    n16187 , 
    n16188 , 
    n16189 , 
    n16190 , 
    n16191 , 
    n16192 , 
    n16193 , 
    n16194 , 
    n16195 , 
    n16196 , 
    n16197 , 
    n16198 , 
    n16199 , 
    n16200 , 
    n16201 , 
    n16202 , 
    n16203 , 
    n16204 , 
    n16205 , 
    n16206 , 
    n16207 , 
    n16208 , 
    n16209 , 
    n16210 , 
    n16211 , 
    n16212 , 
    n16213 , 
    n16214 , 
    n16215 , 
    n16216 , 
    n16217 , 
    n16218 , 
    n16219 , 
    n16220 , 
    n16221 , 
    n16222 , 
    n16223 , 
    n16224 , 
    n16225 , 
    n16226 , 
    n16227 , 
    n16228 , 
    n16229 , 
    n16230 , 
    n16231 , 
    n16232 , 
    n16233 , 
    n16234 , 
    n16235 , 
    n16236 , 
    n16237 , 
    n16238 , 
    n16239 , 
    n16240 , 
    n16241 , 
    n16242 , 
    n16243 , 
    n16244 , 
    n16245 , 
    n16246 , 
    n16247 , 
    n16248 , 
    n16249 , 
    n16250 , 
    n16251 , 
    n16252 , 
    n16253 , 
    n16254 , 
    n16255 , 
    n16256 , 
    n16257 , 
    n16258 , 
    n16259 , 
    n16260 , 
    n16261 , 
    n16262 , 
    n16263 , 
    n16264 , 
    n16265 , 
    n16266 , 
    n16267 , 
    n16268 , 
    n16269 , 
    n16270 , 
    n16271 , 
    n16272 , 
    n16273 , 
    n16274 , 
    n16275 , 
    n16276 , 
    n16277 , 
    n16278 , 
    n16279 , 
    n16280 , 
    n16281 , 
    n16282 , 
    n16283 , 
    n16284 , 
    n16285 , 
    n16286 , 
    n16287 , 
    n16288 , 
    n16289 , 
    n16290 , 
    n16291 , 
    n16292 , 
    n16293 , 
    n16294 , 
    n16295 , 
    n16296 , 
    n16297 , 
    n16298 , 
    n16299 , 
    n16300 , 
    n16301 , 
    n16302 , 
    n16303 , 
    n16304 , 
    n16305 , 
    n16306 , 
    n16307 , 
    n16308 , 
    n16309 , 
    n16310 , 
    n16311 , 
    n16312 , 
    n16313 , 
    n16314 , 
    n16315 , 
    n16316 , 
    n16317 , 
    n16318 , 
    n16319 , 
    n16320 , 
    n16321 , 
    n16322 , 
    n16323 , 
    n16324 , 
    n16325 , 
    n16326 , 
    n16327 , 
    n16328 , 
    n16329 , 
    n16330 , 
    n16331 , 
    n16332 , 
    n16333 , 
    n16334 , 
    n16335 , 
    n16336 , 
    n16337 , 
    n16338 , 
    n16339 , 
    n16340 , 
    n16341 , 
    n16342 , 
    n16343 , 
    n16344 , 
    n16345 , 
    n16346 , 
    n16347 , 
    n16348 , 
    n16349 , 
    n16350 , 
    n16351 , 
    n16352 , 
    n16353 , 
    n16354 , 
    n16355 , 
    n16356 , 
    n16357 , 
    n16358 , 
    n16359 , 
    n16360 , 
    n16361 , 
    n16362 , 
    n16363 , 
    n16364 , 
    n16365 , 
    n16366 , 
    n16367 , 
    n16368 , 
    n16369 , 
    n16370 , 
    n16371 , 
    n16372 , 
    n16373 , 
    n16374 , 
    n16375 , 
    n16376 , 
    n16377 , 
    n16378 , 
    n16379 , 
    n16380 , 
    n16381 , 
    n16382 , 
    n16383 , 
    n16384 , 
    n16385 , 
    n16386 , 
    n16387 , 
    n16388 , 
    n16389 , 
    n16390 , 
    n16391 , 
    n16392 , 
    n16393 , 
    n16394 , 
    n16395 , 
    n16396 , 
    n16397 , 
    n16398 , 
    n16399 , 
    n16400 , 
    n16401 , 
    n16402 , 
    n16403 , 
    n16404 , 
    n16405 , 
    n16406 , 
    n16407 , 
    n16408 , 
    n16409 , 
    n16410 , 
    n16411 , 
    n16412 , 
    n16413 , 
    n16414 , 
    n16415 , 
    n16416 , 
    n16417 , 
    n16418 , 
    n16419 , 
    n16420 , 
    n16421 , 
    n16422 , 
    n16423 , 
    n16424 , 
    n16425 , 
    n16426 , 
    n16427 , 
    n16428 , 
    n16429 , 
    n16430 , 
    n16431 , 
    n16432 , 
    n16433 , 
    n16434 , 
    n16435 , 
    n16436 , 
    n16437 , 
    n16438 , 
    n16439 , 
    n16440 , 
    n16441 , 
    n16442 , 
    n16443 , 
    n16444 , 
    n16445 , 
    n16446 , 
    n16447 , 
    n16448 , 
    n16449 , 
    n16450 , 
    n16451 , 
    n16452 , 
    n16453 , 
    n16454 , 
    n16455 , 
    n16456 , 
    n16457 , 
    n16458 , 
    n16459 , 
    n16460 , 
    n16461 , 
    n16462 , 
    n16463 , 
    n16464 , 
    n16465 , 
    n16466 , 
    n16467 , 
    n16468 , 
    n16469 , 
    n16470 , 
    n16471 , 
    n16472 , 
    n16473 , 
    n16474 , 
    n16475 , 
    n16476 , 
    n16477 , 
    n16478 , 
    n16479 , 
    n16480 , 
    n16481 , 
    n16482 , 
    n16483 , 
    n16484 , 
    n16485 , 
    n16486 , 
    n16487 , 
    n16488 , 
    n16489 , 
    n16490 , 
    n16491 , 
    n16492 , 
    n16493 , 
    n16494 , 
    n16495 , 
    n16496 , 
    n16497 , 
    n16498 , 
    n16499 , 
    n16500 , 
    n16501 , 
    n16502 , 
    n16503 , 
    n16504 , 
    n16505 , 
    n16506 , 
    n16507 , 
    n16508 , 
    n16509 , 
    n16510 , 
    n16511 , 
    n16512 , 
    n16513 , 
    n16514 , 
    n16515 , 
    n16516 , 
    n16517 , 
    n16518 , 
    n16519 , 
    n16520 , 
    n16521 , 
    n16522 , 
    n16523 , 
    n16524 , 
    n16525 , 
    n16526 , 
    n16527 , 
    n16528 , 
    n16529 , 
    n16530 , 
    n16531 , 
    n16532 , 
    n16533 , 
    n16534 , 
    n16535 , 
    n16536 , 
    n16537 , 
    n16538 , 
    n16539 , 
    n16540 , 
    n16541 , 
    n16542 , 
    n16543 , 
    n16544 , 
    n16545 , 
    n16546 , 
    n16547 , 
    n16548 , 
    n16549 , 
    n16550 , 
    n16551 , 
    n16552 , 
    n16553 , 
    n16554 , 
    n16555 , 
    n16556 , 
    n16557 , 
    n16558 , 
    n16559 , 
    n16560 , 
    n16561 , 
    n16562 , 
    n16563 , 
    n16564 , 
    n16565 , 
    n16566 , 
    n16567 , 
    n16568 , 
    n16569 , 
    n16570 , 
    n16571 , 
    n16572 , 
    n16573 , 
    n16574 , 
    n16575 , 
    n16576 , 
    n16577 , 
    n16578 , 
    n16579 , 
    n16580 , 
    n16581 , 
    n16582 , 
    n16583 , 
    n16584 , 
    n16585 , 
    n16586 , 
    n16587 , 
    n16588 , 
    n16589 , 
    n16590 , 
    n16591 , 
    n16592 , 
    n16593 , 
    n16594 , 
    n16595 , 
    n16596 , 
    n16597 , 
    n16598 , 
    n16599 , 
    n16600 , 
    n16601 , 
    n16602 , 
    n16603 , 
    n16604 , 
    n16605 , 
    n16606 , 
    n16607 , 
    n16608 , 
    n16609 , 
    n16610 , 
    n16611 , 
    n16612 , 
    n16613 , 
    n16614 , 
    n16615 , 
    n16616 , 
    n16617 , 
    n16618 , 
    n16619 , 
    n16620 , 
    n16621 , 
    n16622 , 
    n16623 , 
    n16624 , 
    n16625 , 
    n16626 , 
    n16627 , 
    n16628 , 
    n16629 , 
    n16630 , 
    n16631 , 
    n16632 , 
    n16633 , 
    n16634 , 
    n16635 , 
    n16636 , 
    n16637 , 
    n16638 , 
    n16639 , 
    n16640 , 
    n16641 , 
    n16642 , 
    n16643 , 
    n16644 , 
    n16645 , 
    n16646 , 
    n16647 , 
    n16648 , 
    n16649 , 
    n16650 , 
    n16651 , 
    n16652 , 
    n16653 , 
    n16654 , 
    n16655 , 
    n16656 , 
    n16657 , 
    n16658 , 
    n16659 , 
    n16660 , 
    n16661 , 
    n16662 , 
    n16663 , 
    n16664 , 
    n16665 , 
    n16666 , 
    n16667 , 
    n16668 , 
    n16669 , 
    n16670 , 
    n16671 , 
    n16672 , 
    n16673 , 
    n16674 , 
    n16675 , 
    n16676 , 
    n16677 , 
    n16678 , 
    n16679 , 
    n16680 , 
    n16681 , 
    n16682 , 
    n16683 , 
    n16684 , 
    n16685 , 
    n16686 , 
    n16687 , 
    n16688 , 
    n16689 , 
    n16690 , 
    n16691 , 
    n16692 , 
    n16693 , 
    n16694 , 
    n16695 , 
    n16696 , 
    n16697 , 
    n16698 , 
    n16699 , 
    n16700 , 
    n16701 , 
    n16702 , 
    n16703 , 
    n16704 , 
    n16705 , 
    n16706 , 
    n16707 , 
    n16708 , 
    n16709 , 
    n16710 , 
    n16711 , 
    n16712 , 
    n16713 , 
    n16714 , 
    n16715 , 
    n16716 , 
    n16717 , 
    n16718 , 
    n16719 , 
    n16720 , 
    n16721 , 
    n16722 , 
    n16723 , 
    n16724 , 
    n16725 , 
    n16726 , 
    n16727 , 
    n16728 , 
    n16729 , 
    n16730 , 
    n16731 , 
    n16732 , 
    n16733 , 
    n16734 , 
    n16735 , 
    n16736 , 
    n16737 , 
    n16738 , 
    n16739 , 
    n16740 , 
    n16741 , 
    n16742 , 
    n16743 , 
    n16744 , 
    n16745 , 
    n16746 , 
    n16747 , 
    n16748 , 
    n16749 , 
    n16750 , 
    n16751 , 
    n16752 , 
    n16753 , 
    n16754 , 
    n16755 , 
    n16756 , 
    n16757 , 
    n16758 , 
    n16759 , 
    n16760 , 
    n16761 , 
    n16762 , 
    n16763 , 
    n16764 , 
    n16765 , 
    n16766 , 
    n16767 , 
    n16768 , 
    n16769 , 
    n16770 , 
    n16771 , 
    n16772 , 
    n16773 , 
    n16774 , 
    n16775 , 
    n16776 , 
    n16777 , 
    n16778 , 
    n16779 , 
    n16780 , 
    n16781 , 
    n16782 , 
    n16783 , 
    n16784 , 
    n16785 , 
    n16786 , 
    n16787 , 
    n16788 , 
    n16789 , 
    n16790 , 
    n16791 , 
    n16792 , 
    n16793 , 
    n16794 , 
    n16795 , 
    n16796 , 
    n16797 , 
    n16798 , 
    n16799 , 
    n16800 , 
    n16801 , 
    n16802 , 
    n16803 , 
    n16804 , 
    n16805 , 
    n16806 , 
    n16807 , 
    n16808 , 
    n16809 , 
    n16810 , 
    n16811 , 
    n16812 , 
    n16813 , 
    n16814 , 
    n16815 , 
    n16816 , 
    n16817 , 
    n16818 , 
    n16819 , 
    n16820 , 
    n16821 , 
    n16822 , 
    n16823 , 
    n16824 , 
    n16825 , 
    n16826 , 
    n16827 , 
    n16828 , 
    n16829 , 
    n16830 , 
    n16831 , 
    n16832 , 
    n16833 , 
    n16834 , 
    n16835 , 
    n16836 , 
    n16837 , 
    n16838 , 
    n16839 , 
    n16840 , 
    n16841 , 
    n16842 , 
    n16843 , 
    n16844 , 
    n16845 , 
    n16846 , 
    n16847 , 
    n16848 , 
    n16849 , 
    n16850 , 
    n16851 , 
    n16852 , 
    n16853 , 
    n16854 , 
    n16855 , 
    n16856 , 
    n16857 , 
    n16858 , 
    n16859 , 
    n16860 , 
    n16861 , 
    n16862 , 
    n16863 , 
    n16864 , 
    n16865 , 
    n16866 , 
    n16867 , 
    n16868 , 
    n16869 , 
    n16870 , 
    n16871 , 
    n16872 , 
    n16873 , 
    n16874 , 
    n16875 , 
    n16876 , 
    n16877 , 
    n16878 , 
    n16879 , 
    n16880 , 
    n16881 , 
    n16882 , 
    n16883 , 
    n16884 , 
    n16885 , 
    n16886 , 
    n16887 , 
    n16888 , 
    n16889 , 
    n16890 , 
    n16891 , 
    n16892 , 
    n16893 , 
    n16894 , 
    n16895 , 
    n16896 , 
    n16897 , 
    n16898 , 
    n16899 , 
    n16900 , 
    n16901 , 
    n16902 , 
    n16903 , 
    n16904 , 
    n16905 , 
    n16906 , 
    n16907 , 
    n16908 , 
    n16909 , 
    n16910 , 
    n16911 , 
    n16912 , 
    n16913 , 
    n16914 , 
    n16915 , 
    n16916 , 
    n16917 , 
    n16918 , 
    n16919 , 
    n16920 , 
    n16921 , 
    n16922 , 
    n16923 , 
    n16924 , 
    n16925 , 
    n16926 , 
    n16927 , 
    n16928 , 
    n16929 , 
    n16930 , 
    n16931 , 
    n16932 , 
    n16933 , 
    n16934 , 
    n16935 , 
    n16936 , 
    n16937 , 
    n16938 , 
    n16939 , 
    n16940 , 
    n16941 , 
    n16942 , 
    n16943 , 
    n16944 , 
    n16945 , 
    n16946 , 
    n16947 , 
    n16948 , 
    n16949 , 
    n16950 , 
    n16951 , 
    n16952 , 
    n16953 , 
    n16954 , 
    n16955 , 
    n16956 , 
    n16957 , 
    n16958 , 
    n16959 , 
    n16960 , 
    n16961 , 
    n16962 , 
    n16963 , 
    n16964 , 
    n16965 , 
    n16966 , 
    n16967 , 
    n16968 , 
    n16969 , 
    n16970 , 
    n16971 , 
    n16972 , 
    n16973 , 
    n16974 , 
    n16975 , 
    n16976 , 
    n16977 , 
    n16978 , 
    n16979 , 
    n16980 , 
    n16981 , 
    n16982 , 
    n16983 , 
    n16984 , 
    n16985 , 
    n16986 , 
    n16987 , 
    n16988 , 
    n16989 , 
    n16990 , 
    n16991 , 
    n16992 , 
    n16993 , 
    n16994 , 
    n16995 , 
    n16996 , 
    n16997 , 
    n16998 , 
    n16999 , 
    n17000 , 
    n17001 , 
    n17002 , 
    n17003 , 
    n17004 , 
    n17005 , 
    n17006 , 
    n17007 , 
    n17008 , 
    n17009 , 
    n17010 , 
    n17011 , 
    n17012 , 
    n17013 , 
    n17014 , 
    n17015 , 
    n17016 , 
    n17017 , 
    n17018 , 
    n17019 , 
    n17020 , 
    n17021 , 
    n17022 , 
    n17023 , 
    n17024 , 
    n17025 , 
    n17026 , 
    n17027 , 
    n17028 , 
    n17029 , 
    n17030 , 
    n17031 , 
    n17032 , 
    n17033 , 
    n17034 , 
    n17035 , 
    n17036 , 
    n17037 , 
    n17038 , 
    n17039 , 
    n17040 , 
    n17041 , 
    n17042 , 
    n17043 , 
    n17044 , 
    n17045 , 
    n17046 , 
    n17047 , 
    n17048 , 
    n17049 , 
    n17050 , 
    n17051 , 
    n17052 , 
    n17053 , 
    n17054 , 
    n17055 , 
    n17056 , 
    n17057 , 
    n17058 , 
    n17059 , 
    n17060 , 
    n17061 , 
    n17062 , 
    n17063 , 
    n17064 , 
    n17065 , 
    n17066 , 
    n17067 , 
    n17068 , 
    n17069 , 
    n17070 , 
    n17071 , 
    n17072 , 
    n17073 , 
    n17074 , 
    n17075 , 
    n17076 , 
    n17077 , 
    n17078 , 
    n17079 , 
    n17080 , 
    n17081 , 
    n17082 , 
    n17083 , 
    n17084 , 
    n17085 , 
    n17086 , 
    n17087 , 
    n17088 , 
    n17089 , 
    n17090 , 
    n17091 , 
    n17092 , 
    n17093 , 
    n17094 , 
    n17095 , 
    n17096 , 
    n17097 , 
    n17098 , 
    n17099 , 
    n17100 , 
    n17101 , 
    n17102 , 
    n17103 , 
    n17104 , 
    n17105 , 
    n17106 , 
    n17107 , 
    n17108 , 
    n17109 , 
    n17110 , 
    n17111 , 
    n17112 , 
    n17113 , 
    n17114 , 
    n17115 , 
    n17116 , 
    n17117 , 
    n17118 , 
    n17119 , 
    n17120 , 
    n17121 , 
    n17122 , 
    n17123 , 
    n17124 , 
    n17125 , 
    n17126 , 
    n17127 , 
    n17128 , 
    n17129 , 
    n17130 , 
    n17131 , 
    n17132 , 
    n17133 , 
    n17134 , 
    n17135 , 
    n17136 , 
    n17137 , 
    n17138 , 
    n17139 , 
    n17140 , 
    n17141 , 
    n17142 , 
    n17143 , 
    n17144 , 
    n17145 , 
    n17146 , 
    n17147 , 
    n17148 , 
    n17149 , 
    n17150 , 
    n17151 , 
    n17152 , 
    n17153 , 
    n17154 , 
    n17155 , 
    n17156 , 
    n17157 , 
    n17158 , 
    n17159 , 
    n17160 , 
    n17161 , 
    n17162 , 
    n17163 , 
    n17164 , 
    n17165 , 
    n17166 , 
    n17167 , 
    n17168 , 
    n17169 , 
    n17170 , 
    n17171 , 
    n17172 , 
    n17173 , 
    n17174 , 
    n17175 , 
    n17176 , 
    n17177 , 
    n17178 , 
    n17179 , 
    n17180 , 
    n17181 , 
    n17182 , 
    n17183 , 
    n17184 , 
    n17185 , 
    n17186 , 
    n17187 , 
    n17188 , 
    n17189 , 
    n17190 , 
    n17191 , 
    n17192 , 
    n17193 , 
    n17194 , 
    n17195 , 
    n17196 , 
    n17197 , 
    n17198 , 
    n17199 , 
    n17200 , 
    n17201 , 
    n17202 , 
    n17203 , 
    n17204 , 
    n17205 , 
    n17206 , 
    n17207 , 
    n17208 , 
    n17209 , 
    n17210 , 
    n17211 , 
    n17212 , 
    n17213 , 
    n17214 , 
    n17215 , 
    n17216 , 
    n17217 , 
    n17218 , 
    n17219 , 
    n17220 , 
    n17221 , 
    n17222 , 
    n17223 , 
    n17224 , 
    n17225 , 
    n17226 , 
    n17227 , 
    n17228 , 
    n17229 , 
    n17230 , 
    n17231 , 
    n17232 , 
    n17233 , 
    n17234 , 
    n17235 , 
    n17236 , 
    n17237 , 
    n17238 , 
    n17239 , 
    n17240 , 
    n17241 , 
    n17242 , 
    n17243 , 
    n17244 , 
    n17245 , 
    n17246 , 
    n17247 , 
    n17248 , 
    n17249 , 
    n17250 , 
    n17251 , 
    n17252 , 
    n17253 , 
    n17254 , 
    n17255 , 
    n17256 , 
    n17257 , 
    n17258 , 
    n17259 , 
    n17260 , 
    n17261 , 
    n17262 , 
    n17263 , 
    n17264 , 
    n17265 , 
    n17266 , 
    n17267 , 
    n17268 , 
    n17269 , 
    n17270 , 
    n17271 , 
    n17272 , 
    n17273 , 
    n17274 , 
    n17275 , 
    n17276 , 
    n17277 , 
    n17278 , 
    n17279 , 
    n17280 , 
    n17281 , 
    n17282 , 
    n17283 , 
    n17284 , 
    n17285 , 
    n17286 , 
    n17287 , 
    n17288 , 
    n17289 , 
    n17290 , 
    n17291 , 
    n17292 , 
    n17293 , 
    n17294 , 
    n17295 , 
    n17296 , 
    n17297 , 
    n17298 , 
    n17299 , 
    n17300 , 
    n17301 , 
    n17302 , 
    n17303 , 
    n17304 , 
    n17305 , 
    n17306 , 
    n17307 , 
    n17308 , 
    n17309 , 
    n17310 , 
    n17311 , 
    n17312 , 
    n17313 , 
    n17314 , 
    n17315 , 
    n17316 , 
    n17317 , 
    n17318 , 
    n17319 , 
    n17320 , 
    n17321 , 
    n17322 , 
    n17323 , 
    n17324 , 
    n17325 , 
    n17326 , 
    n17327 , 
    n17328 , 
    n17329 , 
    n17330 , 
    n17331 , 
    n17332 , 
    n17333 , 
    n17334 , 
    n17335 , 
    n17336 , 
    n17337 , 
    n17338 , 
    n17339 , 
    n17340 , 
    n17341 , 
    n17342 , 
    n17343 , 
    n17344 , 
    n17345 , 
    n17346 , 
    n17347 , 
    n17348 , 
    n17349 , 
    n17350 , 
    n17351 , 
    n17352 , 
    n17353 , 
    n17354 , 
    n17355 , 
    n17356 , 
    n17357 , 
    n17358 , 
    n17359 , 
    n17360 , 
    n17361 , 
    n17362 , 
    n17363 , 
    n17364 , 
    n17365 , 
    n17366 , 
    n17367 , 
    n17368 , 
    n17369 , 
    n17370 , 
    n17371 , 
    n17372 , 
    n17373 , 
    n17374 , 
    n17375 , 
    n17376 , 
    n17377 , 
    n17378 , 
    n17379 , 
    n17380 , 
    n17381 , 
    n17382 , 
    n17383 , 
    n17384 , 
    n17385 , 
    n17386 , 
    n17387 , 
    n17388 , 
    n17389 , 
    n17390 , 
    n17391 , 
    n17392 , 
    n17393 , 
    n17394 , 
    n17395 , 
    n17396 , 
    n17397 , 
    n17398 , 
    n17399 , 
    n17400 , 
    n17401 , 
    n17402 , 
    n17403 , 
    n17404 , 
    n17405 , 
    n17406 , 
    n17407 , 
    n17408 , 
    n17409 , 
    n17410 , 
    n17411 , 
    n17412 , 
    n17413 , 
    n17414 , 
    n17415 , 
    n17416 , 
    n17417 , 
    n17418 , 
    n17419 , 
    n17420 , 
    n17421 , 
    n17422 , 
    n17423 , 
    n17424 , 
    n17425 , 
    n17426 , 
    n17427 , 
    n17428 , 
    n17429 , 
    n17430 , 
    n17431 , 
    n17432 , 
    n17433 , 
    n17434 , 
    n17435 , 
    n17436 , 
    n17437 , 
    n17438 , 
    n17439 , 
    n17440 , 
    n17441 , 
    n17442 , 
    n17443 , 
    n17444 , 
    n17445 , 
    n17446 , 
    n17447 , 
    n17448 , 
    n17449 , 
    n17450 , 
    n17451 , 
    n17452 , 
    n17453 , 
    n17454 , 
    n17455 , 
    n17456 , 
    n17457 , 
    n17458 , 
    n17459 , 
    n17460 , 
    n17461 , 
    n17462 , 
    n17463 , 
    n17464 , 
    n17465 , 
    n17466 , 
    n17467 , 
    n17468 , 
    n17469 , 
    n17470 , 
    n17471 , 
    n17472 , 
    n17473 , 
    n17474 , 
    n17475 , 
    n17476 , 
    n17477 , 
    n17478 , 
    n17479 , 
    n17480 , 
    n17481 , 
    n17482 , 
    n17483 , 
    n17484 , 
    n17485 , 
    n17486 , 
    n17487 , 
    n17488 , 
    n17489 , 
    n17490 , 
    n17491 , 
    n17492 , 
    n17493 , 
    n17494 , 
    n17495 , 
    n17496 , 
    n17497 , 
    n17498 , 
    n17499 , 
    n17500 , 
    n17501 , 
    n17502 , 
    n17503 , 
    n17504 , 
    n17505 , 
    n17506 , 
    n17507 , 
    n17508 , 
    n17509 , 
    n17510 , 
    n17511 , 
    n17512 , 
    n17513 , 
    n17514 , 
    n17515 , 
    n17516 , 
    n17517 , 
    n17518 , 
    n17519 , 
    n17520 , 
    n17521 , 
    n17522 , 
    n17523 , 
    n17524 , 
    n17525 , 
    n17526 , 
    n17527 , 
    n17528 , 
    n17529 , 
    n17530 , 
    n17531 , 
    n17532 , 
    n17533 , 
    n17534 , 
    n17535 , 
    n17536 , 
    n17537 , 
    n17538 , 
    n17539 , 
    n17540 , 
    n17541 , 
    n17542 , 
    n17543 , 
    n17544 , 
    n17545 , 
    n17546 , 
    n17547 , 
    n17548 , 
    n17549 , 
    n17550 , 
    n17551 , 
    n17552 , 
    n17553 , 
    n17554 , 
    n17555 , 
    n17556 , 
    n17557 , 
    n17558 , 
    n17559 , 
    n17560 , 
    n17561 , 
    n17562 , 
    n17563 , 
    n17564 , 
    n17565 , 
    n17566 , 
    n17567 , 
    n17568 , 
    n17569 , 
    n17570 , 
    n17571 , 
    n17572 , 
    n17573 , 
    n17574 , 
    n17575 , 
    n17576 , 
    n17577 , 
    n17578 , 
    n17579 , 
    n17580 , 
    n17581 , 
    n17582 , 
    n17583 , 
    n17584 , 
    n17585 , 
    n17586 , 
    n17587 , 
    n17588 , 
    n17589 , 
    n17590 , 
    n17591 , 
    n17592 , 
    n17593 , 
    n17594 , 
    n17595 , 
    n17596 , 
    n17597 , 
    n17598 , 
    n17599 , 
    n17600 , 
    n17601 , 
    n17602 , 
    n17603 , 
    n17604 , 
    n17605 , 
    n17606 , 
    n17607 , 
    n17608 , 
    n17609 , 
    n17610 , 
    n17611 , 
    n17612 , 
    n17613 , 
    n17614 , 
    n17615 , 
    n17616 , 
    n17617 , 
    n17618 , 
    n17619 , 
    n17620 , 
    n17621 , 
    n17622 , 
    n17623 , 
    n17624 , 
    n17625 , 
    n17626 , 
    n17627 , 
    n17628 , 
    n17629 , 
    n17630 , 
    n17631 , 
    n17632 , 
    n17633 , 
    n17634 , 
    n17635 , 
    n17636 , 
    n17637 , 
    n17638 , 
    n17639 , 
    n17640 , 
    n17641 , 
    n17642 , 
    n17643 , 
    n17644 , 
    n17645 , 
    n17646 , 
    n17647 , 
    n17648 , 
    n17649 , 
    n17650 , 
    n17651 , 
    n17652 , 
    n17653 , 
    n17654 , 
    n17655 , 
    n17656 , 
    n17657 , 
    n17658 , 
    n17659 , 
    n17660 , 
    n17661 , 
    n17662 , 
    n17663 , 
    n17664 , 
    n17665 , 
    n17666 , 
    n17667 , 
    n17668 , 
    n17669 , 
    n17670 , 
    n17671 , 
    n17672 , 
    n17673 , 
    n17674 , 
    n17675 , 
    n17676 , 
    n17677 , 
    n17678 , 
    n17679 , 
    n17680 , 
    n17681 , 
    n17682 , 
    n17683 , 
    n17684 , 
    n17685 , 
    n17686 , 
    n17687 , 
    n17688 , 
    n17689 , 
    n17690 , 
    n17691 , 
    n17692 , 
    n17693 , 
    n17694 , 
    n17695 , 
    n17696 , 
    n17697 , 
    n17698 , 
    n17699 , 
    n17700 , 
    n17701 , 
    n17702 , 
    n17703 , 
    n17704 , 
    n17705 , 
    n17706 , 
    n17707 , 
    n17708 , 
    n17709 , 
    n17710 , 
    n17711 , 
    n17712 , 
    n17713 , 
    n17714 , 
    n17715 , 
    n17716 , 
    n17717 , 
    n17718 , 
    n17719 , 
    n17720 , 
    n17721 , 
    n17722 , 
    n17723 , 
    n17724 , 
    n17725 , 
    n17726 , 
    n17727 , 
    n17728 , 
    n17729 , 
    n17730 , 
    n17731 , 
    n17732 , 
    n17733 , 
    n17734 , 
    n17735 , 
    n17736 , 
    n17737 , 
    n17738 , 
    n17739 , 
    n17740 , 
    n17741 , 
    n17742 , 
    n17743 , 
    n17744 , 
    n17745 , 
    n17746 , 
    n17747 , 
    n17748 , 
    n17749 , 
    n17750 , 
    n17751 , 
    n17752 , 
    n17753 , 
    n17754 , 
    n17755 , 
    n17756 , 
    n17757 , 
    n17758 , 
    n17759 , 
    n17760 , 
    n17761 , 
    n17762 , 
    n17763 , 
    n17764 , 
    n17765 , 
    n17766 , 
    n17767 , 
    n17768 , 
    n17769 , 
    n17770 , 
    n17771 , 
    n17772 , 
    n17773 , 
    n17774 , 
    n17775 , 
    n17776 , 
    n17777 , 
    n17778 , 
    n17779 , 
    n17780 , 
    n17781 , 
    n17782 , 
    n17783 , 
    n17784 , 
    n17785 , 
    n17786 , 
    n17787 , 
    n17788 , 
    n17789 , 
    n17790 , 
    n17791 , 
    n17792 , 
    n17793 , 
    n17794 , 
    n17795 , 
    n17796 , 
    n17797 , 
    n17798 , 
    n17799 , 
    n17800 , 
    n17801 , 
    n17802 , 
    n17803 , 
    n17804 , 
    n17805 , 
    n17806 , 
    n17807 , 
    n17808 , 
    n17809 , 
    n17810 , 
    n17811 , 
    n17812 , 
    n17813 , 
    n17814 , 
    n17815 , 
    n17816 , 
    n17817 , 
    n17818 , 
    n17819 , 
    n17820 , 
    n17821 , 
    n17822 , 
    n17823 , 
    n17824 , 
    n17825 , 
    n17826 , 
    n17827 , 
    n17828 , 
    n17829 , 
    n17830 , 
    n17831 , 
    n17832 , 
    n17833 , 
    n17834 , 
    n17835 , 
    n17836 , 
    n17837 , 
    n17838 , 
    n17839 , 
    n17840 , 
    n17841 , 
    n17842 , 
    n17843 , 
    n17844 , 
    n17845 , 
    n17846 , 
    n17847 , 
    n17848 , 
    n17849 , 
    n17850 , 
    n17851 , 
    n17852 , 
    n17853 , 
    n17854 , 
    n17855 , 
    n17856 , 
    n17857 , 
    n17858 , 
    n17859 , 
    n17860 , 
    n17861 , 
    n17862 , 
    n17863 , 
    n17864 , 
    n17865 , 
    n17866 , 
    n17867 , 
    n17868 , 
    n17869 , 
    n17870 , 
    n17871 , 
    n17872 , 
    n17873 , 
    n17874 , 
    n17875 , 
    n17876 , 
    n17877 , 
    n17878 , 
    n17879 , 
    n17880 , 
    n17881 , 
    n17882 , 
    n17883 , 
    n17884 , 
    n17885 , 
    n17886 , 
    n17887 , 
    n17888 , 
    n17889 , 
    n17890 , 
    n17891 , 
    n17892 , 
    n17893 , 
    n17894 , 
    n17895 , 
    n17896 , 
    n17897 , 
    n17898 , 
    n17899 , 
    n17900 , 
    n17901 , 
    n17902 , 
    n17903 , 
    n17904 , 
    n17905 , 
    n17906 , 
    n17907 , 
    n17908 , 
    n17909 , 
    n17910 , 
    n17911 , 
    n17912 , 
    n17913 , 
    n17914 , 
    n17915 , 
    n17916 , 
    n17917 , 
    n17918 , 
    n17919 , 
    n17920 , 
    n17921 , 
    n17922 , 
    n17923 , 
    n17924 , 
    n17925 , 
    n17926 , 
    n17927 , 
    n17928 , 
    n17929 , 
    n17930 , 
    n17931 , 
    n17932 , 
    n17933 , 
    n17934 , 
    n17935 , 
    n17936 , 
    n17937 , 
    n17938 , 
    n17939 , 
    n17940 , 
    n17941 , 
    n17942 , 
    n17943 , 
    n17944 , 
    n17945 , 
    n17946 , 
    n17947 , 
    n17948 , 
    n17949 , 
    n17950 , 
    n17951 , 
    n17952 , 
    n17953 , 
    n17954 , 
    n17955 , 
    n17956 , 
    n17957 , 
    n17958 , 
    n17959 , 
    n17960 , 
    n17961 , 
    n17962 , 
    n17963 , 
    n17964 , 
    n17965 , 
    n17966 , 
    n17967 , 
    n17968 , 
    n17969 , 
    n17970 , 
    n17971 , 
    n17972 , 
    n17973 , 
    n17974 , 
    n17975 , 
    n17976 , 
    n17977 , 
    n17978 , 
    n17979 , 
    n17980 , 
    n17981 , 
    n17982 , 
    n17983 , 
    n17984 , 
    n17985 , 
    n17986 , 
    n17987 , 
    n17988 , 
    n17989 , 
    n17990 , 
    n17991 , 
    n17992 , 
    n17993 , 
    n17994 , 
    n17995 , 
    n17996 , 
    n17997 , 
    n17998 , 
    n17999 , 
    n18000 , 
    n18001 , 
    n18002 , 
    n18003 , 
    n18004 , 
    n18005 , 
    n18006 , 
    n18007 , 
    n18008 , 
    n18009 , 
    n18010 , 
    n18011 , 
    n18012 , 
    n18013 , 
    n18014 , 
    n18015 , 
    n18016 , 
    n18017 , 
    n18018 , 
    n18019 , 
    n18020 , 
    n18021 , 
    n18022 , 
    n18023 , 
    n18024 , 
    n18025 , 
    n18026 , 
    n18027 , 
    n18028 , 
    n18029 , 
    n18030 , 
    n18031 , 
    n18032 , 
    n18033 , 
    n18034 , 
    n18035 , 
    n18036 , 
    n18037 , 
    n18038 , 
    n18039 , 
    n18040 , 
    n18041 , 
    n18042 , 
    n18043 , 
    n18044 , 
    n18045 , 
    n18046 , 
    n18047 , 
    n18048 , 
    n18049 , 
    n18050 , 
    n18051 , 
    n18052 , 
    n18053 , 
    n18054 , 
    n18055 , 
    n18056 , 
    n18057 , 
    n18058 , 
    n18059 , 
    n18060 , 
    n18061 , 
    n18062 , 
    n18063 , 
    n18064 , 
    n18065 , 
    n18066 , 
    n18067 , 
    n18068 , 
    n18069 , 
    n18070 , 
    n18071 , 
    n18072 , 
    n18073 , 
    n18074 , 
    n18075 , 
    n18076 , 
    n18077 , 
    n18078 , 
    n18079 , 
    n18080 , 
    n18081 , 
    n18082 , 
    n18083 , 
    n18084 , 
    n18085 , 
    n18086 , 
    n18087 , 
    n18088 , 
    n18089 , 
    n18090 , 
    n18091 , 
    n18092 , 
    n18093 , 
    n18094 , 
    n18095 , 
    n18096 , 
    n18097 , 
    n18098 , 
    n18099 , 
    n18100 , 
    n18101 , 
    n18102 , 
    n18103 , 
    n18104 , 
    n18105 , 
    n18106 , 
    n18107 , 
    n18108 , 
    n18109 , 
    n18110 , 
    n18111 , 
    n18112 , 
    n18113 , 
    n18114 , 
    n18115 , 
    n18116 , 
    n18117 , 
    n18118 , 
    n18119 , 
    n18120 , 
    n18121 , 
    n18122 , 
    n18123 , 
    n18124 , 
    n18125 , 
    n18126 , 
    n18127 , 
    n18128 , 
    n18129 , 
    n18130 , 
    n18131 , 
    n18132 , 
    n18133 , 
    n18134 , 
    n18135 , 
    n18136 , 
    n18137 , 
    n18138 , 
    n18139 , 
    n18140 , 
    n18141 , 
    n18142 , 
    n18143 , 
    n18144 , 
    n18145 , 
    n18146 , 
    n18147 , 
    n18148 , 
    n18149 , 
    n18150 , 
    n18151 , 
    n18152 , 
    n18153 , 
    n18154 , 
    n18155 , 
    n18156 , 
    n18157 , 
    n18158 , 
    n18159 , 
    n18160 , 
    n18161 , 
    n18162 , 
    n18163 , 
    n18164 , 
    n18165 , 
    n18166 , 
    n18167 , 
    n18168 , 
    n18169 , 
    n18170 , 
    n18171 , 
    n18172 , 
    n18173 , 
    n18174 , 
    n18175 , 
    n18176 , 
    n18177 , 
    n18178 , 
    n18179 , 
    n18180 , 
    n18181 , 
    n18182 , 
    n18183 , 
    n18184 , 
    n18185 , 
    n18186 , 
    n18187 , 
    n18188 , 
    n18189 , 
    n18190 , 
    n18191 , 
    n18192 , 
    n18193 , 
    n18194 , 
    n18195 , 
    n18196 , 
    n18197 , 
    n18198 , 
    n18199 , 
    n18200 , 
    n18201 , 
    n18202 , 
    n18203 , 
    n18204 , 
    n18205 , 
    n18206 , 
    n18207 , 
    n18208 , 
    n18209 , 
    n18210 , 
    n18211 , 
    n18212 , 
    n18213 , 
    n18214 , 
    n18215 , 
    n18216 , 
    n18217 , 
    n18218 , 
    n18219 , 
    n18220 , 
    n18221 , 
    n18222 , 
    n18223 , 
    n18224 , 
    n18225 , 
    n18226 , 
    n18227 , 
    n18228 , 
    n18229 , 
    n18230 , 
    n18231 , 
    n18232 , 
    n18233 , 
    n18234 , 
    n18235 , 
    n18236 , 
    n18237 , 
    n18238 , 
    n18239 , 
    n18240 , 
    n18241 , 
    n18242 , 
    n18243 , 
    n18244 , 
    n18245 , 
    n18246 , 
    n18247 , 
    n18248 , 
    n18249 , 
    n18250 , 
    n18251 , 
    n18252 , 
    n18253 , 
    n18254 , 
    n18255 , 
    n18256 , 
    n18257 , 
    n18258 , 
    n18259 , 
    n18260 , 
    n18261 , 
    n18262 , 
    n18263 , 
    n18264 , 
    n18265 , 
    n18266 , 
    n18267 , 
    n18268 , 
    n18269 , 
    n18270 , 
    n18271 , 
    n18272 , 
    n18273 , 
    n18274 , 
    n18275 , 
    n18276 , 
    n18277 , 
    n18278 , 
    n18279 , 
    n18280 , 
    n18281 , 
    n18282 , 
    n18283 , 
    n18284 , 
    n18285 , 
    n18286 , 
    n18287 , 
    n18288 , 
    n18289 , 
    n18290 , 
    n18291 , 
    n18292 , 
    n18293 , 
    n18294 , 
    n18295 , 
    n18296 , 
    n18297 , 
    n18298 , 
    n18299 , 
    n18300 , 
    n18301 , 
    n18302 , 
    n18303 , 
    n18304 , 
    n18305 , 
    n18306 , 
    n18307 , 
    n18308 , 
    n18309 , 
    n18310 , 
    n18311 , 
    n18312 , 
    n18313 , 
    n18314 , 
    n18315 , 
    n18316 , 
    n18317 , 
    n18318 , 
    n18319 , 
    n18320 , 
    n18321 , 
    n18322 , 
    n18323 , 
    n18324 , 
    n18325 , 
    n18326 , 
    n18327 , 
    n18328 , 
    n18329 , 
    n18330 , 
    n18331 , 
    n18332 , 
    n18333 , 
    n18334 , 
    n18335 , 
    n18336 , 
    n18337 , 
    n18338 , 
    n18339 , 
    n18340 , 
    n18341 , 
    n18342 , 
    n18343 , 
    n18344 , 
    n18345 , 
    n18346 , 
    n18347 , 
    n18348 , 
    n18349 , 
    n18350 , 
    n18351 , 
    n18352 , 
    n18353 , 
    n18354 , 
    n18355 , 
    n18356 , 
    n18357 , 
    n18358 , 
    n18359 , 
    n18360 , 
    n18361 , 
    n18362 , 
    n18363 , 
    n18364 , 
    n18365 , 
    n18366 , 
    n18367 , 
    n18368 , 
    n18369 , 
    n18370 , 
    n18371 , 
    n18372 , 
    n18373 , 
    n18374 , 
    n18375 , 
    n18376 , 
    n18377 , 
    n18378 , 
    n18379 , 
    n18380 , 
    n18381 , 
    n18382 , 
    n18383 , 
    n18384 , 
    n18385 , 
    n18386 , 
    n18387 , 
    n18388 , 
    n18389 , 
    n18390 , 
    n18391 , 
    n18392 , 
    n18393 , 
    n18394 , 
    n18395 , 
    n18396 , 
    n18397 , 
    n18398 , 
    n18399 , 
    n18400 , 
    n18401 , 
    n18402 , 
    n18403 , 
    n18404 , 
    n18405 , 
    n18406 , 
    n18407 , 
    n18408 , 
    n18409 , 
    n18410 , 
    n18411 , 
    n18412 , 
    n18413 , 
    n18414 , 
    n18415 , 
    n18416 , 
    n18417 , 
    n18418 , 
    n18419 , 
    n18420 , 
    n18421 , 
    n18422 , 
    n18423 , 
    n18424 , 
    n18425 , 
    n18426 , 
    n18427 , 
    n18428 , 
    n18429 , 
    n18430 , 
    n18431 , 
    n18432 , 
    n18433 , 
    n18434 , 
    n18435 , 
    n18436 , 
    n18437 , 
    n18438 , 
    n18439 , 
    n18440 , 
    n18441 , 
    n18442 , 
    n18443 , 
    n18444 , 
    n18445 , 
    n18446 , 
    n18447 , 
    n18448 , 
    n18449 , 
    n18450 , 
    n18451 , 
    n18452 , 
    n18453 , 
    n18454 , 
    n18455 , 
    n18456 , 
    n18457 , 
    n18458 , 
    n18459 , 
    n18460 , 
    n18461 , 
    n18462 , 
    n18463 , 
    n18464 , 
    n18465 , 
    n18466 , 
    n18467 , 
    n18468 , 
    n18469 , 
    n18470 , 
    n18471 , 
    n18472 , 
    n18473 , 
    n18474 , 
    n18475 , 
    n18476 , 
    n18477 , 
    n18478 , 
    n18479 , 
    n18480 , 
    n18481 , 
    n18482 , 
    n18483 , 
    n18484 , 
    n18485 , 
    n18486 , 
    n18487 , 
    n18488 , 
    n18489 , 
    n18490 , 
    n18491 , 
    n18492 , 
    n18493 , 
    n18494 , 
    n18495 , 
    n18496 , 
    n18497 , 
    n18498 , 
    n18499 , 
    n18500 , 
    n18501 , 
    n18502 , 
    n18503 , 
    n18504 , 
    n18505 , 
    n18506 , 
    n18507 , 
    n18508 , 
    n18509 , 
    n18510 , 
    n18511 , 
    n18512 , 
    n18513 , 
    n18514 , 
    n18515 , 
    n18516 , 
    n18517 , 
    n18518 , 
    n18519 , 
    n18520 , 
    n18521 , 
    n18522 , 
    n18523 , 
    n18524 , 
    n18525 , 
    n18526 , 
    n18527 , 
    n18528 , 
    n18529 , 
    n18530 , 
    n18531 , 
    n18532 , 
    n18533 , 
    n18534 , 
    n18535 , 
    n18536 , 
    n18537 , 
    n18538 , 
    n18539 , 
    n18540 , 
    n18541 , 
    n18542 , 
    n18543 , 
    n18544 , 
    n18545 , 
    n18546 , 
    n18547 , 
    n18548 , 
    n18549 , 
    n18550 , 
    n18551 , 
    n18552 , 
    n18553 , 
    n18554 , 
    n18555 , 
    n18556 , 
    n18557 , 
    n18558 , 
    n18559 , 
    n18560 , 
    n18561 , 
    n18562 , 
    n18563 , 
    n18564 , 
    n18565 , 
    n18566 , 
    n18567 , 
    n18568 , 
    n18569 , 
    n18570 , 
    n18571 , 
    n18572 , 
    n18573 , 
    n18574 , 
    n18575 , 
    n18576 , 
    n18577 , 
    n18578 , 
    n18579 , 
    n18580 , 
    n18581 , 
    n18582 , 
    n18583 , 
    n18584 , 
    n18585 , 
    n18586 , 
    n18587 , 
    n18588 , 
    n18589 , 
    n18590 , 
    n18591 , 
    n18592 , 
    n18593 , 
    n18594 , 
    n18595 , 
    n18596 , 
    n18597 , 
    n18598 , 
    n18599 , 
    n18600 , 
    n18601 , 
    n18602 , 
    n18603 , 
    n18604 , 
    n18605 , 
    n18606 , 
    n18607 , 
    n18608 , 
    n18609 , 
    n18610 , 
    n18611 , 
    n18612 , 
    n18613 , 
    n18614 , 
    n18615 , 
    n18616 , 
    n18617 , 
    n18618 , 
    n18619 , 
    n18620 , 
    n18621 , 
    n18622 , 
    n18623 , 
    n18624 , 
    n18625 , 
    n18626 , 
    n18627 , 
    n18628 , 
    n18629 , 
    n18630 , 
    n18631 , 
    n18632 , 
    n18633 , 
    n18634 , 
    n18635 , 
    n18636 , 
    n18637 , 
    n18638 , 
    n18639 , 
    n18640 , 
    n18641 , 
    n18642 , 
    n18643 , 
    n18644 , 
    n18645 , 
    n18646 , 
    n18647 , 
    n18648 , 
    n18649 , 
    n18650 , 
    n18651 , 
    n18652 , 
    n18653 , 
    n18654 , 
    n18655 , 
    n18656 , 
    n18657 , 
    n18658 , 
    n18659 , 
    n18660 , 
    n18661 , 
    n18662 , 
    n18663 , 
    n18664 , 
    n18665 , 
    n18666 , 
    n18667 , 
    n18668 , 
    n18669 , 
    n18670 , 
    n18671 , 
    n18672 , 
    n18673 , 
    n18674 , 
    n18675 , 
    n18676 , 
    n18677 , 
    n18678 , 
    n18679 , 
    n18680 , 
    n18681 , 
    n18682 , 
    n18683 , 
    n18684 , 
    n18685 , 
    n18686 , 
    n18687 , 
    n18688 , 
    n18689 , 
    n18690 , 
    n18691 , 
    n18692 , 
    n18693 , 
    n18694 , 
    n18695 , 
    n18696 , 
    n18697 , 
    n18698 , 
    n18699 , 
    n18700 , 
    n18701 , 
    n18702 , 
    n18703 , 
    n18704 , 
    n18705 , 
    n18706 , 
    n18707 , 
    n18708 , 
    n18709 , 
    n18710 , 
    n18711 , 
    n18712 , 
    n18713 , 
    n18714 , 
    n18715 , 
    n18716 , 
    n18717 , 
    n18718 , 
    n18719 , 
    n18720 , 
    n18721 , 
    n18722 , 
    n18723 , 
    n18724 , 
    n18725 , 
    n18726 , 
    n18727 , 
    n18728 , 
    n18729 , 
    n18730 , 
    n18731 , 
    n18732 , 
    n18733 , 
    n18734 , 
    n18735 , 
    n18736 , 
    n18737 , 
    n18738 , 
    n18739 , 
    n18740 , 
    n18741 , 
    n18742 , 
    n18743 , 
    n18744 , 
    n18745 , 
    n18746 , 
    n18747 , 
    n18748 , 
    n18749 , 
    n18750 , 
    n18751 , 
    n18752 , 
    n18753 , 
    n18754 , 
    n18755 , 
    n18756 , 
    n18757 , 
    n18758 , 
    n18759 , 
    n18760 , 
    n18761 , 
    n18762 , 
    n18763 , 
    n18764 , 
    n18765 , 
    n18766 , 
    n18767 , 
    n18768 , 
    n18769 , 
    n18770 , 
    n18771 , 
    n18772 , 
    n18773 , 
    n18774 , 
    n18775 , 
    n18776 , 
    n18777 , 
    n18778 , 
    n18779 , 
    n18780 , 
    n18781 , 
    n18782 , 
    n18783 , 
    n18784 , 
    n18785 , 
    n18786 , 
    n18787 , 
    n18788 , 
    n18789 , 
    n18790 , 
    n18791 , 
    n18792 , 
    n18793 , 
    n18794 , 
    n18795 , 
    n18796 , 
    n18797 , 
    n18798 , 
    n18799 , 
    n18800 , 
    n18801 , 
    n18802 , 
    n18803 , 
    n18804 , 
    n18805 , 
    n18806 , 
    n18807 , 
    n18808 , 
    n18809 , 
    n18810 , 
    n18811 , 
    n18812 , 
    n18813 , 
    n18814 , 
    n18815 , 
    n18816 , 
    n18817 , 
    n18818 , 
    n18819 , 
    n18820 , 
    n18821 , 
    n18822 , 
    n18823 , 
    n18824 , 
    n18825 , 
    n18826 , 
    n18827 , 
    n18828 , 
    n18829 , 
    n18830 , 
    n18831 , 
    n18832 , 
    n18833 , 
    n18834 , 
    n18835 , 
    n18836 , 
    n18837 , 
    n18838 , 
    n18839 , 
    n18840 , 
    n18841 , 
    n18842 , 
    n18843 , 
    n18844 , 
    n18845 , 
    n18846 , 
    n18847 , 
    n18848 , 
    n18849 , 
    n18850 , 
    n18851 , 
    n18852 , 
    n18853 , 
    n18854 , 
    n18855 , 
    n18856 , 
    n18857 , 
    n18858 , 
    n18859 , 
    n18860 , 
    n18861 , 
    n18862 , 
    n18863 , 
    n18864 , 
    n18865 , 
    n18866 , 
    n18867 , 
    n18868 , 
    n18869 , 
    n18870 , 
    n18871 , 
    n18872 , 
    n18873 , 
    n18874 , 
    n18875 , 
    n18876 , 
    n18877 , 
    n18878 , 
    n18879 , 
    n18880 , 
    n18881 , 
    n18882 , 
    n18883 , 
    n18884 , 
    n18885 , 
    n18886 , 
    n18887 , 
    n18888 , 
    n18889 , 
    n18890 , 
    n18891 , 
    n18892 , 
    n18893 , 
    n18894 , 
    n18895 , 
    n18896 , 
    n18897 , 
    n18898 , 
    n18899 , 
    n18900 , 
    n18901 , 
    n18902 , 
    n18903 , 
    n18904 , 
    n18905 , 
    n18906 , 
    n18907 , 
    n18908 , 
    n18909 , 
    n18910 , 
    n18911 , 
    n18912 , 
    n18913 , 
    n18914 , 
    n18915 , 
    n18916 , 
    n18917 , 
    n18918 , 
    n18919 , 
    n18920 , 
    n18921 , 
    n18922 , 
    n18923 , 
    n18924 , 
    n18925 , 
    n18926 , 
    n18927 , 
    n18928 , 
    n18929 , 
    n18930 , 
    n18931 , 
    n18932 , 
    n18933 , 
    n18934 , 
    n18935 , 
    n18936 , 
    n18937 , 
    n18938 , 
    n18939 , 
    n18940 , 
    n18941 , 
    n18942 , 
    n18943 , 
    n18944 , 
    n18945 , 
    n18946 , 
    n18947 , 
    n18948 , 
    n18949 , 
    n18950 , 
    n18951 , 
    n18952 , 
    n18953 , 
    n18954 , 
    n18955 , 
    n18956 , 
    n18957 , 
    n18958 , 
    n18959 , 
    n18960 , 
    n18961 , 
    n18962 , 
    n18963 , 
    n18964 , 
    n18965 , 
    n18966 , 
    n18967 , 
    n18968 , 
    n18969 , 
    n18970 , 
    n18971 , 
    n18972 , 
    n18973 , 
    n18974 , 
    n18975 , 
    n18976 , 
    n18977 , 
    n18978 , 
    n18979 , 
    n18980 , 
    n18981 , 
    n18982 , 
    n18983 , 
    n18984 , 
    n18985 , 
    n18986 , 
    n18987 , 
    n18988 , 
    n18989 , 
    n18990 , 
    n18991 , 
    n18992 , 
    n18993 , 
    n18994 , 
    n18995 , 
    n18996 , 
    n18997 , 
    n18998 , 
    n18999 , 
    n19000 , 
    n19001 , 
    n19002 , 
    n19003 , 
    n19004 , 
    n19005 , 
    n19006 , 
    n19007 , 
    n19008 , 
    n19009 , 
    n19010 , 
    n19011 , 
    n19012 , 
    n19013 , 
    n19014 , 
    n19015 , 
    n19016 , 
    n19017 , 
    n19018 , 
    n19019 , 
    n19020 , 
    n19021 , 
    n19022 , 
    n19023 , 
    n19024 , 
    n19025 , 
    n19026 , 
    n19027 , 
    n19028 , 
    n19029 , 
    n19030 , 
    n19031 , 
    n19032 , 
    n19033 , 
    n19034 , 
    n19035 , 
    n19036 , 
    n19037 , 
    n19038 , 
    n19039 , 
    n19040 , 
    n19041 , 
    n19042 , 
    n19043 , 
    n19044 , 
    n19045 , 
    n19046 , 
    n19047 , 
    n19048 , 
    n19049 , 
    n19050 , 
    n19051 , 
    n19052 , 
    n19053 , 
    n19054 , 
    n19055 , 
    n19056 , 
    n19057 , 
    n19058 , 
    n19059 , 
    n19060 , 
    n19061 , 
    n19062 , 
    n19063 , 
    n19064 , 
    n19065 , 
    n19066 , 
    n19067 , 
    n19068 , 
    n19069 , 
    n19070 , 
    n19071 , 
    n19072 , 
    n19073 , 
    n19074 , 
    n19075 , 
    n19076 , 
    n19077 , 
    n19078 , 
    n19079 , 
    n19080 , 
    n19081 , 
    n19082 , 
    n19083 , 
    n19084 , 
    n19085 , 
    n19086 , 
    n19087 , 
    n19088 , 
    n19089 , 
    n19090 , 
    n19091 , 
    n19092 , 
    n19093 , 
    n19094 , 
    n19095 , 
    n19096 , 
    n19097 , 
    n19098 , 
    n19099 , 
    n19100 , 
    n19101 , 
    n19102 , 
    n19103 , 
    n19104 , 
    n19105 , 
    n19106 , 
    n19107 , 
    n19108 , 
    n19109 , 
    n19110 , 
    n19111 , 
    n19112 , 
    n19113 , 
    n19114 , 
    n19115 , 
    n19116 , 
    n19117 , 
    n19118 , 
    n19119 , 
    n19120 , 
    n19121 , 
    n19122 , 
    n19123 , 
    n19124 , 
    n19125 , 
    n19126 , 
    n19127 , 
    n19128 , 
    n19129 , 
    n19130 , 
    n19131 , 
    n19132 , 
    n19133 , 
    n19134 , 
    n19135 , 
    n19136 , 
    n19137 , 
    n19138 , 
    n19139 , 
    n19140 , 
    n19141 , 
    n19142 , 
    n19143 , 
    n19144 , 
    n19145 , 
    n19146 , 
    n19147 , 
    n19148 , 
    n19149 , 
    n19150 , 
    n19151 , 
    n19152 , 
    n19153 , 
    n19154 , 
    n19155 , 
    n19156 , 
    n19157 , 
    n19158 , 
    n19159 , 
    n19160 , 
    n19161 , 
    n19162 , 
    n19163 , 
    n19164 , 
    n19165 , 
    n19166 , 
    n19167 , 
    n19168 , 
    n19169 , 
    n19170 , 
    n19171 , 
    n19172 , 
    n19173 , 
    n19174 , 
    n19175 , 
    n19176 , 
    n19177 , 
    n19178 , 
    n19179 , 
    n19180 , 
    n19181 , 
    n19182 , 
    n19183 , 
    n19184 , 
    n19185 , 
    n19186 , 
    n19187 , 
    n19188 , 
    n19189 , 
    n19190 , 
    n19191 , 
    n19192 , 
    n19193 , 
    n19194 , 
    n19195 , 
    n19196 , 
    n19197 , 
    n19198 , 
    n19199 , 
    n19200 , 
    n19201 , 
    n19202 , 
    n19203 , 
    n19204 , 
    n19205 , 
    n19206 , 
    n19207 , 
    n19208 , 
    n19209 , 
    n19210 , 
    n19211 , 
    n19212 , 
    n19213 , 
    n19214 , 
    n19215 , 
    n19216 , 
    n19217 , 
    n19218 , 
    n19219 , 
    n19220 , 
    n19221 , 
    n19222 , 
    n19223 , 
    n19224 , 
    n19225 , 
    n19226 , 
    n19227 , 
    n19228 , 
    n19229 , 
    n19230 , 
    n19231 , 
    n19232 , 
    n19233 , 
    n19234 , 
    n19235 , 
    n19236 , 
    n19237 , 
    n19238 , 
    n19239 , 
    n19240 , 
    n19241 , 
    n19242 , 
    n19243 , 
    n19244 , 
    n19245 , 
    n19246 , 
    n19247 , 
    n19248 , 
    n19249 , 
    n19250 , 
    n19251 , 
    n19252 , 
    n19253 , 
    n19254 , 
    n19255 , 
    n19256 , 
    n19257 , 
    n19258 , 
    n19259 , 
    n19260 , 
    n19261 , 
    n19262 , 
    n19263 , 
    n19264 , 
    n19265 , 
    n19266 , 
    n19267 , 
    n19268 , 
    n19269 , 
    n19270 , 
    n19271 , 
    n19272 , 
    n19273 , 
    n19274 , 
    n19275 , 
    n19276 , 
    n19277 , 
    n19278 , 
    n19279 , 
    n19280 , 
    n19281 , 
    n19282 , 
    n19283 , 
    n19284 , 
    n19285 , 
    n19286 , 
    n19287 , 
    n19288 , 
    n19289 , 
    n19290 , 
    n19291 , 
    n19292 , 
    n19293 , 
    n19294 , 
    n19295 , 
    n19296 , 
    n19297 , 
    n19298 , 
    n19299 , 
    n19300 , 
    n19301 , 
    n19302 , 
    n19303 , 
    n19304 , 
    n19305 , 
    n19306 , 
    n19307 , 
    n19308 , 
    n19309 , 
    n19310 , 
    n19311 , 
    n19312 , 
    n19313 , 
    n19314 , 
    n19315 , 
    n19316 , 
    n19317 , 
    n19318 , 
    n19319 , 
    n19320 , 
    n19321 , 
    n19322 , 
    n19323 , 
    n19324 , 
    n19325 , 
    n19326 , 
    n19327 , 
    n19328 , 
    n19329 , 
    n19330 , 
    n19331 , 
    n19332 , 
    n19333 , 
    n19334 , 
    n19335 , 
    n19336 , 
    n19337 , 
    n19338 , 
    n19339 , 
    n19340 , 
    n19341 , 
    n19342 , 
    n19343 , 
    n19344 , 
    n19345 , 
    n19346 , 
    n19347 , 
    n19348 , 
    n19349 , 
    n19350 , 
    n19351 , 
    n19352 , 
    n19353 , 
    n19354 , 
    n19355 , 
    n19356 , 
    n19357 , 
    n19358 , 
    n19359 , 
    n19360 , 
    n19361 , 
    n19362 , 
    n19363 , 
    n19364 , 
    n19365 , 
    n19366 , 
    n19367 , 
    n19368 , 
    n19369 , 
    n19370 , 
    n19371 , 
    n19372 , 
    n19373 , 
    n19374 , 
    n19375 , 
    n19376 , 
    n19377 , 
    n19378 , 
    n19379 , 
    n19380 , 
    n19381 , 
    n19382 , 
    n19383 , 
    n19384 , 
    n19385 , 
    n19386 , 
    n19387 , 
    n19388 , 
    n19389 , 
    n19390 , 
    n19391 , 
    n19392 , 
    n19393 , 
    n19394 , 
    n19395 , 
    n19396 , 
    n19397 , 
    n19398 , 
    n19399 , 
    n19400 , 
    n19401 , 
    n19402 , 
    n19403 , 
    n19404 , 
    n19405 , 
    n19406 , 
    n19407 , 
    n19408 , 
    n19409 , 
    n19410 , 
    n19411 , 
    n19412 , 
    n19413 , 
    n19414 , 
    n19415 , 
    n19416 , 
    n19417 , 
    n19418 , 
    n19419 , 
    n19420 , 
    n19421 , 
    n19422 , 
    n19423 , 
    n19424 , 
    n19425 , 
    n19426 , 
    n19427 , 
    n19428 , 
    n19429 , 
    n19430 , 
    n19431 , 
    n19432 , 
    n19433 , 
    n19434 , 
    n19435 , 
    n19436 , 
    n19437 , 
    n19438 , 
    n19439 , 
    n19440 , 
    n19441 , 
    n19442 , 
    n19443 , 
    n19444 , 
    n19445 , 
    n19446 , 
    n19447 , 
    n19448 , 
    n19449 , 
    n19450 , 
    n19451 , 
    n19452 , 
    n19453 , 
    n19454 , 
    n19455 , 
    n19456 , 
    n19457 , 
    n19458 , 
    n19459 , 
    n19460 , 
    n19461 , 
    n19462 , 
    n19463 , 
    n19464 , 
    n19465 , 
    n19466 , 
    n19467 , 
    n19468 , 
    n19469 , 
    n19470 , 
    n19471 , 
    n19472 , 
    n19473 , 
    n19474 , 
    n19475 , 
    n19476 , 
    n19477 , 
    n19478 , 
    n19479 , 
    n19480 , 
    n19481 , 
    n19482 , 
    n19483 , 
    n19484 , 
    n19485 , 
    n19486 , 
    n19487 , 
    n19488 , 
    n19489 , 
    n19490 , 
    n19491 , 
    n19492 , 
    n19493 , 
    n19494 , 
    n19495 , 
    n19496 , 
    n19497 , 
    n19498 , 
    n19499 , 
    n19500 , 
    n19501 , 
    n19502 , 
    n19503 , 
    n19504 , 
    n19505 , 
    n19506 , 
    n19507 , 
    n19508 , 
    n19509 , 
    n19510 , 
    n19511 , 
    n19512 , 
    n19513 , 
    n19514 , 
    n19515 , 
    n19516 , 
    n19517 , 
    n19518 , 
    n19519 , 
    n19520 , 
    n19521 , 
    n19522 , 
    n19523 , 
    n19524 , 
    n19525 , 
    n19526 , 
    n19527 , 
    n19528 , 
    n19529 , 
    n19530 , 
    n19531 , 
    n19532 , 
    n19533 , 
    n19534 , 
    n19535 , 
    n19536 , 
    n19537 , 
    n19538 , 
    n19539 , 
    n19540 , 
    n19541 , 
    n19542 , 
    n19543 , 
    n19544 , 
    n19545 , 
    n19546 , 
    n19547 , 
    n19548 , 
    n19549 , 
    n19550 , 
    n19551 , 
    n19552 , 
    n19553 , 
    n19554 , 
    n19555 , 
    n19556 , 
    n19557 , 
    n19558 , 
    n19559 , 
    n19560 , 
    n19561 , 
    n19562 , 
    n19563 , 
    n19564 , 
    n19565 , 
    n19566 , 
    n19567 , 
    n19568 , 
    n19569 , 
    n19570 , 
    n19571 , 
    n19572 , 
    n19573 , 
    n19574 , 
    n19575 , 
    n19576 , 
    n19577 , 
    n19578 , 
    n19579 , 
    n19580 , 
    n19581 , 
    n19582 , 
    n19583 , 
    n19584 , 
    n19585 , 
    n19586 , 
    n19587 , 
    n19588 , 
    n19589 , 
    n19590 , 
    n19591 , 
    n19592 , 
    n19593 , 
    n19594 , 
    n19595 , 
    n19596 , 
    n19597 , 
    n19598 , 
    n19599 , 
    n19600 , 
    n19601 , 
    n19602 , 
    n19603 , 
    n19604 , 
    n19605 , 
    n19606 , 
    n19607 , 
    n19608 , 
    n19609 , 
    n19610 , 
    n19611 , 
    n19612 , 
    n19613 , 
    n19614 , 
    n19615 , 
    n19616 , 
    n19617 , 
    n19618 , 
    n19619 , 
    n19620 , 
    n19621 , 
    n19622 , 
    n19623 , 
    n19624 , 
    n19625 , 
    n19626 , 
    n19627 , 
    n19628 , 
    n19629 , 
    n19630 , 
    n19631 , 
    n19632 , 
    n19633 , 
    n19634 , 
    n19635 , 
    n19636 , 
    n19637 , 
    n19638 , 
    n19639 , 
    n19640 , 
    n19641 , 
    n19642 , 
    n19643 , 
    n19644 , 
    n19645 , 
    n19646 , 
    n19647 , 
    n19648 , 
    n19649 , 
    n19650 , 
    n19651 , 
    n19652 , 
    n19653 , 
    n19654 , 
    n19655 , 
    n19656 , 
    n19657 , 
    n19658 , 
    n19659 , 
    n19660 , 
    n19661 , 
    n19662 , 
    n19663 , 
    n19664 , 
    n19665 , 
    n19666 , 
    n19667 , 
    n19668 , 
    n19669 , 
    n19670 , 
    n19671 , 
    n19672 , 
    n19673 , 
    n19674 , 
    n19675 , 
    n19676 , 
    n19677 , 
    n19678 , 
    n19679 , 
    n19680 , 
    n19681 , 
    n19682 , 
    n19683 , 
    n19684 , 
    n19685 , 
    n19686 , 
    n19687 , 
    n19688 , 
    n19689 , 
    n19690 , 
    n19691 , 
    n19692 , 
    n19693 , 
    n19694 , 
    n19695 , 
    n19696 , 
    n19697 , 
    n19698 , 
    n19699 , 
    n19700 , 
    n19701 , 
    n19702 , 
    n19703 , 
    n19704 , 
    n19705 , 
    n19706 , 
    n19707 , 
    n19708 , 
    n19709 , 
    n19710 , 
    n19711 , 
    n19712 , 
    n19713 , 
    n19714 , 
    n19715 , 
    n19716 , 
    n19717 , 
    n19718 , 
    n19719 , 
    n19720 , 
    n19721 , 
    n19722 , 
    n19723 , 
    n19724 , 
    n19725 , 
    n19726 , 
    n19727 , 
    n19728 , 
    n19729 , 
    n19730 , 
    n19731 , 
    n19732 , 
    n19733 , 
    n19734 , 
    n19735 , 
    n19736 , 
    n19737 , 
    n19738 , 
    n19739 , 
    n19740 , 
    n19741 , 
    n19742 , 
    n19743 , 
    n19744 , 
    n19745 , 
    n19746 , 
    n19747 , 
    n19748 , 
    n19749 , 
    n19750 , 
    n19751 , 
    n19752 , 
    n19753 , 
    n19754 , 
    n19755 , 
    n19756 , 
    n19757 , 
    n19758 , 
    n19759 , 
    n19760 , 
    n19761 , 
    n19762 , 
    n19763 , 
    n19764 , 
    n19765 , 
    n19766 , 
    n19767 , 
    n19768 , 
    n19769 , 
    n19770 , 
    n19771 , 
    n19772 , 
    n19773 , 
    n19774 , 
    n19775 , 
    n19776 , 
    n19777 , 
    n19778 , 
    n19779 , 
    n19780 , 
    n19781 , 
    n19782 , 
    n19783 , 
    n19784 , 
    n19785 , 
    n19786 , 
    n19787 , 
    n19788 , 
    n19789 , 
    n19790 , 
    n19791 , 
    n19792 , 
    n19793 , 
    n19794 , 
    n19795 , 
    n19796 , 
    n19797 , 
    n19798 , 
    n19799 , 
    n19800 , 
    n19801 , 
    n19802 , 
    n19803 , 
    n19804 , 
    n19805 , 
    n19806 , 
    n19807 , 
    n19808 , 
    n19809 , 
    n19810 , 
    n19811 , 
    n19812 , 
    n19813 , 
    n19814 , 
    n19815 , 
    n19816 , 
    n19817 , 
    n19818 , 
    n19819 , 
    n19820 , 
    n19821 , 
    n19822 , 
    n19823 , 
    n19824 , 
    n19825 , 
    n19826 , 
    n19827 , 
    n19828 , 
    n19829 , 
    n19830 , 
    n19831 , 
    n19832 , 
    n19833 , 
    n19834 , 
    n19835 , 
    n19836 , 
    n19837 , 
    n19838 , 
    n19839 , 
    n19840 , 
    n19841 , 
    n19842 , 
    n19843 , 
    n19844 , 
    n19845 , 
    n19846 , 
    n19847 , 
    n19848 , 
    n19849 , 
    n19850 , 
    n19851 , 
    n19852 , 
    n19853 , 
    n19854 , 
    n19855 , 
    n19856 , 
    n19857 , 
    n19858 , 
    n19859 , 
    n19860 , 
    n19861 , 
    n19862 , 
    n19863 , 
    n19864 , 
    n19865 , 
    n19866 , 
    n19867 , 
    n19868 , 
    n19869 , 
    n19870 , 
    n19871 , 
    n19872 , 
    n19873 , 
    n19874 , 
    n19875 , 
    n19876 , 
    n19877 , 
    n19878 , 
    n19879 , 
    n19880 , 
    n19881 , 
    n19882 , 
    n19883 , 
    n19884 , 
    n19885 , 
    n19886 , 
    n19887 , 
    n19888 , 
    n19889 , 
    n19890 , 
    n19891 , 
    n19892 , 
    n19893 , 
    n19894 , 
    n19895 , 
    n19896 , 
    n19897 , 
    n19898 , 
    n19899 , 
    n19900 , 
    n19901 , 
    n19902 , 
    n19903 , 
    n19904 , 
    n19905 , 
    n19906 , 
    n19907 , 
    n19908 , 
    n19909 , 
    n19910 , 
    n19911 , 
    n19912 , 
    n19913 , 
    n19914 , 
    n19915 , 
    n19916 , 
    n19917 , 
    n19918 , 
    n19919 , 
    n19920 , 
    n19921 , 
    n19922 , 
    n19923 , 
    n19924 , 
    n19925 , 
    n19926 , 
    n19927 , 
    n19928 , 
    n19929 , 
    n19930 , 
    n19931 , 
    n19932 , 
    n19933 , 
    n19934 , 
    n19935 , 
    n19936 , 
    n19937 , 
    n19938 , 
    n19939 , 
    n19940 , 
    n19941 , 
    n19942 , 
    n19943 , 
    n19944 , 
    n19945 , 
    n19946 , 
    n19947 , 
    n19948 , 
    n19949 , 
    n19950 , 
    n19951 , 
    n19952 , 
    n19953 , 
    n19954 , 
    n19955 , 
    n19956 , 
    n19957 , 
    n19958 , 
    n19959 , 
    n19960 , 
    n19961 , 
    n19962 , 
    n19963 , 
    n19964 , 
    n19965 , 
    n19966 , 
    n19967 , 
    n19968 , 
    n19969 , 
    n19970 , 
    n19971 , 
    n19972 , 
    n19973 , 
    n19974 , 
    n19975 , 
    n19976 , 
    n19977 , 
    n19978 , 
    n19979 , 
    n19980 , 
    n19981 , 
    n19982 , 
    n19983 , 
    n19984 , 
    n19985 , 
    n19986 , 
    n19987 , 
    n19988 , 
    n19989 , 
    n19990 , 
    n19991 , 
    n19992 , 
    n19993 , 
    n19994 , 
    n19995 , 
    n19996 , 
    n19997 , 
    n19998 , 
    n19999 , 
    n20000 , 
    n20001 , 
    n20002 , 
    n20003 , 
    n20004 , 
    n20005 , 
    n20006 , 
    n20007 , 
    n20008 , 
    n20009 , 
    n20010 , 
    n20011 , 
    n20012 , 
    n20013 , 
    n20014 , 
    n20015 , 
    n20016 , 
    n20017 , 
    n20018 , 
    n20019 , 
    n20020 , 
    n20021 , 
    n20022 , 
    n20023 , 
    n20024 , 
    n20025 , 
    n20026 , 
    n20027 , 
    n20028 , 
    n20029 , 
    n20030 , 
    n20031 , 
    n20032 , 
    n20033 , 
    n20034 , 
    n20035 , 
    n20036 , 
    n20037 , 
    n20038 , 
    n20039 , 
    n20040 , 
    n20041 , 
    n20042 , 
    n20043 , 
    n20044 , 
    n20045 , 
    n20046 , 
    n20047 , 
    n20048 , 
    n20049 , 
    n20050 , 
    n20051 , 
    n20052 , 
    n20053 , 
    n20054 , 
    n20055 , 
    n20056 , 
    n20057 , 
    n20058 , 
    n20059 , 
    n20060 , 
    n20061 , 
    n20062 , 
    n20063 , 
    n20064 , 
    n20065 , 
    n20066 , 
    n20067 , 
    n20068 , 
    n20069 , 
    n20070 , 
    n20071 , 
    n20072 , 
    n20073 , 
    n20074 , 
    n20075 , 
    n20076 , 
    n20077 , 
    n20078 , 
    n20079 , 
    n20080 , 
    n20081 , 
    n20082 , 
    n20083 , 
    n20084 , 
    n20085 , 
    n20086 , 
    n20087 , 
    n20088 , 
    n20089 , 
    n20090 , 
    n20091 , 
    n20092 , 
    n20093 , 
    n20094 , 
    n20095 , 
    n20096 , 
    n20097 , 
    n20098 , 
    n20099 , 
    n20100 , 
    n20101 , 
    n20102 , 
    n20103 , 
    n20104 , 
    n20105 , 
    n20106 , 
    n20107 , 
    n20108 , 
    n20109 , 
    n20110 , 
    n20111 , 
    n20112 , 
    n20113 , 
    n20114 , 
    n20115 , 
    n20116 , 
    n20117 , 
    n20118 , 
    n20119 , 
    n20120 , 
    n20121 , 
    n20122 , 
    n20123 , 
    n20124 , 
    n20125 , 
    n20126 , 
    n20127 , 
    n20128 , 
    n20129 , 
    n20130 , 
    n20131 , 
    n20132 , 
    n20133 , 
    n20134 , 
    n20135 , 
    n20136 , 
    n20137 , 
    n20138 , 
    n20139 , 
    n20140 , 
    n20141 , 
    n20142 , 
    n20143 , 
    n20144 , 
    n20145 , 
    n20146 , 
    n20147 , 
    n20148 , 
    n20149 , 
    n20150 , 
    n20151 , 
    n20152 , 
    n20153 , 
    n20154 , 
    n20155 , 
    n20156 , 
    n20157 , 
    n20158 , 
    n20159 , 
    n20160 , 
    n20161 , 
    n20162 , 
    n20163 , 
    n20164 , 
    n20165 , 
    n20166 , 
    n20167 , 
    n20168 , 
    n20169 , 
    n20170 , 
    n20171 , 
    n20172 , 
    n20173 , 
    n20174 , 
    n20175 , 
    n20176 , 
    n20177 , 
    n20178 , 
    n20179 , 
    n20180 , 
    n20181 , 
    n20182 , 
    n20183 , 
    n20184 , 
    n20185 , 
    n20186 , 
    n20187 , 
    n20188 , 
    n20189 , 
    n20190 , 
    n20191 , 
    n20192 , 
    n20193 , 
    n20194 , 
    n20195 , 
    n20196 , 
    n20197 , 
    n20198 , 
    n20199 , 
    n20200 , 
    n20201 , 
    n20202 , 
    n20203 , 
    n20204 , 
    n20205 , 
    n20206 , 
    n20207 , 
    n20208 , 
    n20209 , 
    n20210 , 
    n20211 , 
    n20212 , 
    n20213 , 
    n20214 , 
    n20215 , 
    n20216 , 
    n20217 , 
    n20218 , 
    n20219 , 
    n20220 , 
    n20221 , 
    n20222 , 
    n20223 , 
    n20224 , 
    n20225 , 
    n20226 , 
    n20227 , 
    n20228 , 
    n20229 , 
    n20230 , 
    n20231 , 
    n20232 , 
    n20233 , 
    n20234 , 
    n20235 , 
    n20236 , 
    n20237 , 
    n20238 , 
    n20239 , 
    n20240 , 
    n20241 , 
    n20242 , 
    n20243 , 
    n20244 , 
    n20245 , 
    n20246 , 
    n20247 , 
    n20248 , 
    n20249 , 
    n20250 , 
    n20251 , 
    n20252 , 
    n20253 , 
    n20254 , 
    n20255 , 
    n20256 , 
    n20257 , 
    n20258 , 
    n20259 , 
    n20260 , 
    n20261 , 
    n20262 , 
    n20263 , 
    n20264 , 
    n20265 , 
    n20266 , 
    n20267 , 
    n20268 , 
    n20269 , 
    n20270 , 
    n20271 , 
    n20272 , 
    n20273 , 
    n20274 , 
    n20275 , 
    n20276 , 
    n20277 , 
    n20278 , 
    n20279 , 
    n20280 , 
    n20281 , 
    n20282 , 
    n20283 , 
    n20284 , 
    n20285 , 
    n20286 , 
    n20287 , 
    n20288 , 
    n20289 , 
    n20290 , 
    n20291 , 
    n20292 , 
    n20293 , 
    n20294 , 
    n20295 , 
    n20296 , 
    n20297 , 
    n20298 , 
    n20299 , 
    n20300 , 
    n20301 , 
    n20302 , 
    n20303 , 
    n20304 , 
    n20305 , 
    n20306 , 
    n20307 , 
    n20308 , 
    n20309 , 
    n20310 , 
    n20311 , 
    n20312 , 
    n20313 , 
    n20314 , 
    n20315 , 
    n20316 , 
    n20317 , 
    n20318 , 
    n20319 , 
    n20320 , 
    n20321 , 
    n20322 , 
    n20323 , 
    n20324 , 
    n20325 , 
    n20326 , 
    n20327 , 
    n20328 , 
    n20329 , 
    n20330 , 
    n20331 , 
    n20332 , 
    n20333 , 
    n20334 , 
    n20335 , 
    n20336 , 
    n20337 , 
    n20338 , 
    n20339 , 
    n20340 , 
    n20341 , 
    n20342 , 
    n20343 , 
    n20344 , 
    n20345 , 
    n20346 , 
    n20347 , 
    n20348 , 
    n20349 , 
    n20350 , 
    n20351 , 
    n20352 , 
    n20353 , 
    n20354 , 
    n20355 , 
    n20356 , 
    n20357 , 
    n20358 , 
    n20359 , 
    n20360 , 
    n20361 , 
    n20362 , 
    n20363 , 
    n20364 , 
    n20365 , 
    n20366 , 
    n20367 , 
    n20368 , 
    n20369 , 
    n20370 , 
    n20371 , 
    n20372 , 
    n20373 , 
    n20374 , 
    n20375 , 
    n20376 , 
    n20377 , 
    n20378 , 
    n20379 , 
    n20380 , 
    n20381 , 
    n20382 , 
    n20383 , 
    n20384 , 
    n20385 , 
    n20386 , 
    n20387 , 
    n20388 , 
    n20389 , 
    n20390 , 
    n20391 , 
    n20392 , 
    n20393 , 
    n20394 , 
    n20395 , 
    n20396 , 
    n20397 , 
    n20398 , 
    n20399 , 
    n20400 , 
    n20401 , 
    n20402 , 
    n20403 , 
    n20404 , 
    n20405 , 
    n20406 , 
    n20407 , 
    n20408 , 
    n20409 , 
    n20410 , 
    n20411 , 
    n20412 , 
    n20413 , 
    n20414 , 
    n20415 , 
    n20416 , 
    n20417 , 
    n20418 , 
    n20419 , 
    n20420 , 
    n20421 , 
    n20422 , 
    n20423 , 
    n20424 , 
    n20425 , 
    n20426 , 
    n20427 , 
    n20428 , 
    n20429 , 
    n20430 , 
    n20431 , 
    n20432 , 
    n20433 , 
    n20434 , 
    n20435 , 
    n20436 , 
    n20437 , 
    n20438 , 
    n20439 , 
    n20440 , 
    n20441 , 
    n20442 , 
    n20443 , 
    n20444 , 
    n20445 , 
    n20446 , 
    n20447 , 
    n20448 , 
    n20449 , 
    n20450 , 
    n20451 , 
    n20452 , 
    n20453 , 
    n20454 , 
    n20455 , 
    n20456 , 
    n20457 , 
    n20458 , 
    n20459 , 
    n20460 , 
    n20461 , 
    n20462 , 
    n20463 , 
    n20464 , 
    n20465 , 
    n20466 , 
    n20467 , 
    n20468 , 
    n20469 , 
    n20470 , 
    n20471 , 
    n20472 , 
    n20473 , 
    n20474 , 
    n20475 , 
    n20476 , 
    n20477 , 
    n20478 , 
    n20479 , 
    n20480 , 
    n20481 , 
    n20482 , 
    n20483 , 
    n20484 , 
    n20485 , 
    n20486 , 
    n20487 , 
    n20488 , 
    n20489 , 
    n20490 , 
    n20491 , 
    n20492 , 
    n20493 , 
    n20494 , 
    n20495 , 
    n20496 , 
    n20497 , 
    n20498 , 
    n20499 , 
    n20500 , 
    n20501 , 
    n20502 , 
    n20503 , 
    n20504 , 
    n20505 , 
    n20506 , 
    n20507 , 
    n20508 , 
    n20509 , 
    n20510 , 
    n20511 , 
    n20512 , 
    n20513 , 
    n20514 , 
    n20515 , 
    n20516 , 
    n20517 , 
    n20518 , 
    n20519 , 
    n20520 , 
    n20521 , 
    n20522 , 
    n20523 , 
    n20524 , 
    n20525 , 
    n20526 , 
    n20527 , 
    n20528 , 
    n20529 , 
    n20530 , 
    n20531 , 
    n20532 , 
    n20533 , 
    n20534 , 
    n20535 , 
    n20536 , 
    n20537 , 
    n20538 , 
    n20539 , 
    n20540 , 
    n20541 , 
    n20542 , 
    n20543 , 
    n20544 , 
    n20545 , 
    n20546 , 
    n20547 , 
    n20548 , 
    n20549 , 
    n20550 , 
    n20551 , 
    n20552 , 
    n20553 , 
    n20554 , 
    n20555 , 
    n20556 , 
    n20557 , 
    n20558 , 
    n20559 , 
    n20560 , 
    n20561 , 
    n20562 , 
    n20563 , 
    n20564 , 
    n20565 , 
    n20566 , 
    n20567 , 
    n20568 , 
    n20569 , 
    n20570 , 
    n20571 , 
    n20572 , 
    n20573 , 
    n20574 , 
    n20575 , 
    n20576 , 
    n20577 , 
    n20578 , 
    n20579 , 
    n20580 , 
    n20581 , 
    n20582 , 
    n20583 , 
    n20584 , 
    n20585 , 
    n20586 , 
    n20587 , 
    n20588 , 
    n20589 , 
    n20590 , 
    n20591 , 
    n20592 , 
    n20593 , 
    n20594 , 
    n20595 , 
    n20596 , 
    n20597 , 
    n20598 , 
    n20599 , 
    n20600 , 
    n20601 , 
    n20602 , 
    n20603 , 
    n20604 , 
    n20605 , 
    n20606 , 
    n20607 , 
    n20608 , 
    n20609 , 
    n20610 , 
    n20611 , 
    n20612 , 
    n20613 , 
    n20614 , 
    n20615 , 
    n20616 , 
    n20617 , 
    n20618 , 
    n20619 , 
    n20620 , 
    n20621 , 
    n20622 , 
    n20623 , 
    n20624 , 
    n20625 , 
    n20626 , 
    n20627 , 
    n20628 , 
    n20629 , 
    n20630 , 
    n20631 , 
    n20632 , 
    n20633 , 
    n20634 , 
    n20635 , 
    n20636 , 
    n20637 , 
    n20638 , 
    n20639 , 
    n20640 , 
    n20641 , 
    n20642 , 
    n20643 , 
    n20644 , 
    n20645 , 
    n20646 , 
    n20647 , 
    n20648 , 
    n20649 , 
    n20650 , 
    n20651 , 
    n20652 , 
    n20653 , 
    n20654 , 
    n20655 , 
    n20656 , 
    n20657 , 
    n20658 , 
    n20659 , 
    n20660 , 
    n20661 , 
    n20662 , 
    n20663 , 
    n20664 , 
    n20665 , 
    n20666 , 
    n20667 , 
    n20668 , 
    n20669 , 
    n20670 , 
    n20671 , 
    n20672 , 
    n20673 , 
    n20674 , 
    n20675 , 
    n20676 , 
    n20677 , 
    n20678 , 
    n20679 , 
    n20680 , 
    n20681 , 
    n20682 , 
    n20683 , 
    n20684 , 
    n20685 , 
    n20686 , 
    n20687 , 
    n20688 , 
    n20689 , 
    n20690 , 
    n20691 , 
    n20692 , 
    n20693 , 
    n20694 , 
    n20695 , 
    n20696 , 
    n20697 , 
    n20698 , 
    n20699 , 
    n20700 , 
    n20701 , 
    n20702 , 
    n20703 , 
    n20704 , 
    n20705 , 
    n20706 , 
    n20707 , 
    n20708 , 
    n20709 , 
    n20710 , 
    n20711 , 
    n20712 , 
    n20713 , 
    n20714 , 
    n20715 , 
    n20716 , 
    n20717 , 
    n20718 , 
    n20719 , 
    n20720 , 
    n20721 , 
    n20722 , 
    n20723 , 
    n20724 , 
    n20725 , 
    n20726 , 
    n20727 , 
    n20728 , 
    n20729 , 
    n20730 , 
    n20731 , 
    n20732 , 
    n20733 , 
    n20734 , 
    n20735 , 
    n20736 , 
    n20737 , 
    n20738 , 
    n20739 , 
    n20740 , 
    n20741 , 
    n20742 , 
    n20743 , 
    n20744 , 
    n20745 , 
    n20746 , 
    n20747 , 
    n20748 , 
    n20749 , 
    n20750 , 
    n20751 , 
    n20752 , 
    n20753 , 
    n20754 , 
    n20755 , 
    n20756 , 
    n20757 , 
    n20758 , 
    n20759 , 
    n20760 , 
    n20761 , 
    n20762 , 
    n20763 , 
    n20764 , 
    n20765 , 
    n20766 , 
    n20767 , 
    n20768 , 
    n20769 , 
    n20770 , 
    n20771 , 
    n20772 , 
    n20773 , 
    n20774 , 
    n20775 , 
    n20776 , 
    n20777 , 
    n20778 , 
    n20779 , 
    n20780 , 
    n20781 , 
    n20782 , 
    n20783 , 
    n20784 , 
    n20785 , 
    n20786 , 
    n20787 , 
    n20788 , 
    n20789 , 
    n20790 , 
    n20791 , 
    n20792 , 
    n20793 , 
    n20794 , 
    n20795 , 
    n20796 , 
    n20797 , 
    n20798 , 
    n20799 , 
    n20800 , 
    n20801 , 
    n20802 , 
    n20803 , 
    n20804 , 
    n20805 , 
    n20806 , 
    n20807 , 
    n20808 , 
    n20809 , 
    n20810 , 
    n20811 , 
    n20812 , 
    n20813 , 
    n20814 , 
    n20815 , 
    n20816 , 
    n20817 , 
    n20818 , 
    n20819 , 
    n20820 , 
    n20821 , 
    n20822 , 
    n20823 , 
    n20824 , 
    n20825 , 
    n20826 , 
    n20827 , 
    n20828 , 
    n20829 , 
    n20830 , 
    n20831 , 
    n20832 , 
    n20833 , 
    n20834 , 
    n20835 , 
    n20836 , 
    n20837 , 
    n20838 , 
    n20839 , 
    n20840 , 
    n20841 , 
    n20842 , 
    n20843 , 
    n20844 , 
    n20845 , 
    n20846 , 
    n20847 , 
    n20848 , 
    n20849 , 
    n20850 , 
    n20851 , 
    n20852 , 
    n20853 , 
    n20854 , 
    n20855 , 
    n20856 , 
    n20857 , 
    n20858 , 
    n20859 , 
    n20860 , 
    n20861 , 
    n20862 , 
    n20863 , 
    n20864 , 
    n20865 , 
    n20866 , 
    n20867 , 
    n20868 , 
    n20869 , 
    n20870 , 
    n20871 , 
    n20872 , 
    n20873 , 
    n20874 , 
    n20875 , 
    n20876 , 
    n20877 , 
    n20878 , 
    n20879 , 
    n20880 , 
    n20881 , 
    n20882 , 
    n20883 , 
    n20884 , 
    n20885 , 
    n20886 , 
    n20887 , 
    n20888 , 
    n20889 , 
    n20890 , 
    n20891 , 
    n20892 , 
    n20893 , 
    n20894 , 
    n20895 , 
    n20896 , 
    n20897 , 
    n20898 , 
    n20899 , 
    n20900 , 
    n20901 , 
    n20902 , 
    n20903 , 
    n20904 , 
    n20905 , 
    n20906 , 
    n20907 , 
    n20908 , 
    n20909 , 
    n20910 , 
    n20911 , 
    n20912 , 
    n20913 , 
    n20914 , 
    n20915 , 
    n20916 , 
    n20917 , 
    n20918 , 
    n20919 , 
    n20920 , 
    n20921 , 
    n20922 , 
    n20923 , 
    n20924 , 
    n20925 , 
    n20926 , 
    n20927 , 
    n20928 , 
    n20929 , 
    n20930 , 
    n20931 , 
    n20932 , 
    n20933 , 
    n20934 , 
    n20935 , 
    n20936 , 
    n20937 , 
    n20938 , 
    n20939 , 
    n20940 , 
    n20941 , 
    n20942 , 
    n20943 , 
    n20944 , 
    n20945 , 
    n20946 , 
    n20947 , 
    n20948 , 
    n20949 , 
    n20950 , 
    n20951 , 
    n20952 , 
    n20953 , 
    n20954 , 
    n20955 , 
    n20956 , 
    n20957 , 
    n20958 , 
    n20959 , 
    n20960 , 
    n20961 , 
    n20962 , 
    n20963 , 
    n20964 , 
    n20965 , 
    n20966 , 
    n20967 , 
    n20968 , 
    n20969 , 
    n20970 , 
    n20971 , 
    n20972 , 
    n20973 , 
    n20974 , 
    n20975 , 
    n20976 , 
    n20977 , 
    n20978 , 
    n20979 , 
    n20980 , 
    n20981 , 
    n20982 , 
    n20983 , 
    n20984 , 
    n20985 , 
    n20986 , 
    n20987 , 
    n20988 , 
    n20989 , 
    n20990 , 
    n20991 , 
    n20992 , 
    n20993 , 
    n20994 , 
    n20995 , 
    n20996 , 
    n20997 , 
    n20998 , 
    n20999 , 
    n21000 , 
    n21001 , 
    n21002 , 
    n21003 , 
    n21004 , 
    n21005 , 
    n21006 , 
    n21007 , 
    n21008 , 
    n21009 , 
    n21010 , 
    n21011 , 
    n21012 , 
    n21013 , 
    n21014 , 
    n21015 , 
    n21016 , 
    n21017 , 
    n21018 , 
    n21019 , 
    n21020 , 
    n21021 , 
    n21022 , 
    n21023 , 
    n21024 , 
    n21025 , 
    n21026 , 
    n21027 , 
    n21028 , 
    n21029 , 
    n21030 , 
    n21031 , 
    n21032 , 
    n21033 , 
    n21034 , 
    n21035 , 
    n21036 , 
    n21037 , 
    n21038 , 
    n21039 , 
    n21040 , 
    n21041 , 
    n21042 , 
    n21043 , 
    n21044 , 
    n21045 , 
    n21046 , 
    n21047 , 
    n21048 , 
    n21049 , 
    n21050 , 
    n21051 , 
    n21052 , 
    n21053 , 
    n21054 , 
    n21055 , 
    n21056 , 
    n21057 , 
    n21058 , 
    n21059 , 
    n21060 , 
    n21061 , 
    n21062 , 
    n21063 , 
    n21064 , 
    n21065 , 
    n21066 , 
    n21067 , 
    n21068 , 
    n21069 , 
    n21070 , 
    n21071 , 
    n21072 , 
    n21073 , 
    n21074 , 
    n21075 , 
    n21076 , 
    n21077 , 
    n21078 , 
    n21079 , 
    n21080 , 
    n21081 , 
    n21082 , 
    n21083 , 
    n21084 , 
    n21085 , 
    n21086 , 
    n21087 , 
    n21088 , 
    n21089 , 
    n21090 , 
    n21091 , 
    n21092 , 
    n21093 , 
    n21094 , 
    n21095 , 
    n21096 , 
    n21097 , 
    n21098 , 
    n21099 , 
    n21100 , 
    n21101 , 
    n21102 , 
    n21103 , 
    n21104 , 
    n21105 , 
    n21106 , 
    n21107 , 
    n21108 , 
    n21109 , 
    n21110 , 
    n21111 , 
    n21112 , 
    n21113 , 
    n21114 , 
    n21115 , 
    n21116 , 
    n21117 , 
    n21118 , 
    n21119 , 
    n21120 , 
    n21121 , 
    n21122 , 
    n21123 , 
    n21124 , 
    n21125 , 
    n21126 , 
    n21127 , 
    n21128 , 
    n21129 , 
    n21130 , 
    n21131 , 
    n21132 , 
    n21133 , 
    n21134 , 
    n21135 , 
    n21136 , 
    n21137 , 
    n21138 , 
    n21139 , 
    n21140 , 
    n21141 , 
    n21142 , 
    n21143 , 
    n21144 , 
    n21145 , 
    n21146 , 
    n21147 , 
    n21148 , 
    n21149 , 
    n21150 , 
    n21151 , 
    n21152 , 
    n21153 , 
    n21154 , 
    n21155 , 
    n21156 , 
    n21157 , 
    n21158 , 
    n21159 , 
    n21160 , 
    n21161 , 
    n21162 , 
    n21163 , 
    n21164 , 
    n21165 , 
    n21166 , 
    n21167 , 
    n21168 , 
    n21169 , 
    n21170 , 
    n21171 , 
    n21172 , 
    n21173 , 
    n21174 , 
    n21175 , 
    n21176 , 
    n21177 , 
    n21178 , 
    n21179 , 
    n21180 , 
    n21181 , 
    n21182 , 
    n21183 , 
    n21184 , 
    n21185 , 
    n21186 , 
    n21187 , 
    n21188 , 
    n21189 , 
    n21190 , 
    n21191 , 
    n21192 , 
    n21193 , 
    n21194 , 
    n21195 , 
    n21196 , 
    n21197 , 
    n21198 , 
    n21199 , 
    n21200 , 
    n21201 , 
    n21202 , 
    n21203 , 
    n21204 , 
    n21205 , 
    n21206 , 
    n21207 , 
    n21208 , 
    n21209 , 
    n21210 , 
    n21211 , 
    n21212 , 
    n21213 , 
    n21214 , 
    n21215 , 
    n21216 , 
    n21217 , 
    n21218 , 
    n21219 , 
    n21220 , 
    n21221 , 
    n21222 , 
    n21223 , 
    n21224 , 
    n21225 , 
    n21226 , 
    n21227 , 
    n21228 , 
    n21229 , 
    n21230 , 
    n21231 , 
    n21232 , 
    n21233 , 
    n21234 , 
    n21235 , 
    n21236 , 
    n21237 , 
    n21238 , 
    n21239 , 
    n21240 , 
    n21241 , 
    n21242 , 
    n21243 , 
    n21244 , 
    n21245 , 
    n21246 , 
    n21247 , 
    n21248 , 
    n21249 , 
    n21250 , 
    n21251 , 
    n21252 , 
    n21253 , 
    n21254 , 
    n21255 , 
    n21256 , 
    n21257 , 
    n21258 , 
    n21259 , 
    n21260 , 
    n21261 , 
    n21262 , 
    n21263 , 
    n21264 , 
    n21265 , 
    n21266 , 
    n21267 , 
    n21268 , 
    n21269 , 
    n21270 , 
    n21271 , 
    n21272 , 
    n21273 , 
    n21274 , 
    n21275 , 
    n21276 , 
    n21277 , 
    n21278 , 
    n21279 , 
    n21280 , 
    n21281 , 
    n21282 , 
    n21283 , 
    n21284 , 
    n21285 , 
    n21286 , 
    n21287 , 
    n21288 , 
    n21289 , 
    n21290 , 
    n21291 , 
    n21292 , 
    n21293 , 
    n21294 , 
    n21295 , 
    n21296 , 
    n21297 , 
    n21298 , 
    n21299 , 
    n21300 , 
    n21301 , 
    n21302 , 
    n21303 , 
    n21304 , 
    n21305 , 
    n21306 , 
    n21307 , 
    n21308 , 
    n21309 , 
    n21310 , 
    n21311 , 
    n21312 , 
    n21313 , 
    n21314 , 
    n21315 , 
    n21316 , 
    n21317 , 
    n21318 , 
    n21319 , 
    n21320 , 
    n21321 , 
    n21322 , 
    n21323 , 
    n21324 , 
    n21325 , 
    n21326 , 
    n21327 , 
    n21328 , 
    n21329 , 
    n21330 , 
    n21331 , 
    n21332 , 
    n21333 , 
    n21334 , 
    n21335 , 
    n21336 , 
    n21337 , 
    n21338 , 
    n21339 , 
    n21340 , 
    n21341 , 
    n21342 , 
    n21343 , 
    n21344 , 
    n21345 , 
    n21346 , 
    n21347 , 
    n21348 , 
    n21349 , 
    n21350 , 
    n21351 , 
    n21352 , 
    n21353 , 
    n21354 , 
    n21355 , 
    n21356 , 
    n21357 , 
    n21358 , 
    n21359 , 
    n21360 , 
    n21361 , 
    n21362 , 
    n21363 , 
    n21364 , 
    n21365 , 
    n21366 , 
    n21367 , 
    n21368 , 
    n21369 , 
    n21370 , 
    n21371 , 
    n21372 , 
    n21373 , 
    n21374 , 
    n21375 , 
    n21376 , 
    n21377 , 
    n21378 , 
    n21379 , 
    n21380 , 
    n21381 , 
    n21382 , 
    n21383 , 
    n21384 , 
    n21385 , 
    n21386 , 
    n21387 , 
    n21388 , 
    n21389 , 
    n21390 , 
    n21391 , 
    n21392 , 
    n21393 , 
    n21394 , 
    n21395 , 
    n21396 , 
    n21397 , 
    n21398 , 
    n21399 , 
    n21400 , 
    n21401 , 
    n21402 , 
    n21403 , 
    n21404 , 
    n21405 , 
    n21406 , 
    n21407 , 
    n21408 , 
    n21409 , 
    n21410 , 
    n21411 , 
    n21412 , 
    n21413 , 
    n21414 , 
    n21415 , 
    n21416 , 
    n21417 , 
    n21418 , 
    n21419 , 
    n21420 , 
    n21421 , 
    n21422 , 
    n21423 , 
    n21424 , 
    n21425 , 
    n21426 , 
    n21427 , 
    n21428 , 
    n21429 , 
    n21430 , 
    n21431 , 
    n21432 , 
    n21433 , 
    n21434 , 
    n21435 , 
    n21436 , 
    n21437 , 
    n21438 , 
    n21439 , 
    n21440 , 
    n21441 , 
    n21442 , 
    n21443 , 
    n21444 , 
    n21445 , 
    n21446 , 
    n21447 , 
    n21448 , 
    n21449 , 
    n21450 , 
    n21451 , 
    n21452 , 
    n21453 , 
    n21454 , 
    n21455 , 
    n21456 , 
    n21457 , 
    n21458 , 
    n21459 , 
    n21460 , 
    n21461 , 
    n21462 , 
    n21463 , 
    n21464 , 
    n21465 , 
    n21466 , 
    n21467 , 
    n21468 , 
    n21469 , 
    n21470 , 
    n21471 , 
    n21472 , 
    n21473 , 
    n21474 , 
    n21475 , 
    n21476 , 
    n21477 , 
    n21478 , 
    n21479 , 
    n21480 , 
    n21481 , 
    n21482 , 
    n21483 , 
    n21484 , 
    n21485 , 
    n21486 , 
    n21487 , 
    n21488 , 
    n21489 , 
    n21490 , 
    n21491 , 
    n21492 , 
    n21493 , 
    n21494 , 
    n21495 , 
    n21496 , 
    n21497 , 
    n21498 , 
    n21499 , 
    n21500 , 
    n21501 , 
    n21502 , 
    n21503 , 
    n21504 , 
    n21505 , 
    n21506 , 
    n21507 , 
    n21508 , 
    n21509 , 
    n21510 , 
    n21511 , 
    n21512 , 
    n21513 , 
    n21514 , 
    n21515 , 
    n21516 , 
    n21517 , 
    n21518 , 
    n21519 , 
    n21520 , 
    n21521 , 
    n21522 , 
    n21523 , 
    n21524 , 
    n21525 , 
    n21526 , 
    n21527 , 
    n21528 , 
    n21529 , 
    n21530 , 
    n21531 , 
    n21532 , 
    n21533 , 
    n21534 , 
    n21535 , 
    n21536 , 
    n21537 , 
    n21538 , 
    n21539 , 
    n21540 , 
    n21541 , 
    n21542 , 
    n21543 , 
    n21544 , 
    n21545 , 
    n21546 , 
    n21547 , 
    n21548 , 
    n21549 , 
    n21550 , 
    n21551 , 
    n21552 , 
    n21553 , 
    n21554 , 
    n21555 , 
    n21556 , 
    n21557 , 
    n21558 , 
    n21559 , 
    n21560 , 
    n21561 , 
    n21562 , 
    n21563 , 
    n21564 , 
    n21565 , 
    n21566 , 
    n21567 , 
    n21568 , 
    n21569 , 
    n21570 , 
    n21571 , 
    n21572 , 
    n21573 , 
    n21574 , 
    n21575 , 
    n21576 , 
    n21577 , 
    n21578 , 
    n21579 , 
    n21580 , 
    n21581 , 
    n21582 , 
    n21583 , 
    n21584 , 
    n21585 , 
    n21586 , 
    n21587 , 
    n21588 , 
    n21589 , 
    n21590 , 
    n21591 , 
    n21592 , 
    n21593 , 
    n21594 , 
    n21595 , 
    n21596 , 
    n21597 , 
    n21598 , 
    n21599 , 
    n21600 , 
    n21601 , 
    n21602 , 
    n21603 , 
    n21604 , 
    n21605 , 
    n21606 , 
    n21607 , 
    n21608 , 
    n21609 , 
    n21610 , 
    n21611 , 
    n21612 , 
    n21613 , 
    n21614 , 
    n21615 , 
    n21616 , 
    n21617 , 
    n21618 , 
    n21619 , 
    n21620 , 
    n21621 , 
    n21622 , 
    n21623 , 
    n21624 , 
    n21625 , 
    n21626 , 
    n21627 , 
    n21628 , 
    n21629 , 
    n21630 , 
    n21631 , 
    n21632 , 
    n21633 , 
    n21634 , 
    n21635 , 
    n21636 , 
    n21637 , 
    n21638 , 
    n21639 , 
    n21640 , 
    n21641 , 
    n21642 , 
    n21643 , 
    n21644 , 
    n21645 , 
    n21646 , 
    n21647 , 
    n21648 , 
    n21649 , 
    n21650 , 
    n21651 , 
    n21652 , 
    n21653 , 
    n21654 , 
    n21655 , 
    n21656 , 
    n21657 , 
    n21658 , 
    n21659 , 
    n21660 , 
    n21661 , 
    n21662 , 
    n21663 , 
    n21664 , 
    n21665 , 
    n21666 , 
    n21667 , 
    n21668 , 
    n21669 , 
    n21670 , 
    n21671 , 
    n21672 , 
    n21673 , 
    n21674 , 
    n21675 , 
    n21676 , 
    n21677 , 
    n21678 , 
    n21679 , 
    n21680 , 
    n21681 , 
    n21682 , 
    n21683 , 
    n21684 , 
    n21685 , 
    n21686 , 
    n21687 , 
    n21688 , 
    n21689 , 
    n21690 , 
    n21691 , 
    n21692 , 
    n21693 , 
    n21694 , 
    n21695 , 
    n21696 , 
    n21697 , 
    n21698 , 
    n21699 , 
    n21700 , 
    n21701 , 
    n21702 , 
    n21703 , 
    n21704 , 
    n21705 , 
    n21706 , 
    n21707 , 
    n21708 , 
    n21709 , 
    n21710 , 
    n21711 , 
    n21712 , 
    n21713 , 
    n21714 , 
    n21715 , 
    n21716 , 
    n21717 , 
    n21718 , 
    n21719 , 
    n21720 , 
    n21721 , 
    n21722 , 
    n21723 , 
    n21724 , 
    n21725 , 
    n21726 , 
    n21727 , 
    n21728 , 
    n21729 , 
    n21730 , 
    n21731 , 
    n21732 , 
    n21733 , 
    n21734 , 
    n21735 , 
    n21736 , 
    n21737 , 
    n21738 , 
    n21739 , 
    n21740 , 
    n21741 , 
    n21742 , 
    n21743 , 
    n21744 , 
    n21745 , 
    n21746 , 
    n21747 , 
    n21748 , 
    n21749 , 
    n21750 , 
    n21751 , 
    n21752 , 
    n21753 , 
    n21754 , 
    n21755 , 
    n21756 , 
    n21757 , 
    n21758 , 
    n21759 , 
    n21760 , 
    n21761 , 
    n21762 , 
    n21763 , 
    n21764 , 
    n21765 , 
    n21766 , 
    n21767 , 
    n21768 , 
    n21769 , 
    n21770 , 
    n21771 , 
    n21772 , 
    n21773 , 
    n21774 , 
    n21775 , 
    n21776 , 
    n21777 , 
    n21778 , 
    n21779 , 
    n21780 , 
    n21781 , 
    n21782 , 
    n21783 , 
    n21784 , 
    n21785 , 
    n21786 , 
    n21787 , 
    n21788 , 
    n21789 , 
    n21790 , 
    n21791 , 
    n21792 , 
    n21793 , 
    n21794 , 
    n21795 , 
    n21796 , 
    n21797 , 
    n21798 , 
    n21799 , 
    n21800 , 
    n21801 , 
    n21802 , 
    n21803 , 
    n21804 , 
    n21805 , 
    n21806 , 
    n21807 , 
    n21808 , 
    n21809 , 
    n21810 , 
    n21811 , 
    n21812 , 
    n21813 , 
    n21814 , 
    n21815 , 
    n21816 , 
    n21817 , 
    n21818 , 
    n21819 , 
    n21820 , 
    n21821 , 
    n21822 , 
    n21823 , 
    n21824 , 
    n21825 , 
    n21826 , 
    n21827 , 
    n21828 , 
    n21829 , 
    n21830 , 
    n21831 , 
    n21832 , 
    n21833 , 
    n21834 , 
    n21835 , 
    n21836 , 
    n21837 , 
    n21838 , 
    n21839 , 
    n21840 , 
    n21841 , 
    n21842 , 
    n21843 , 
    n21844 , 
    n21845 , 
    n21846 , 
    n21847 , 
    n21848 , 
    n21849 , 
    n21850 , 
    n21851 , 
    n21852 , 
    n21853 , 
    n21854 , 
    n21855 , 
    n21856 , 
    n21857 , 
    n21858 , 
    n21859 , 
    n21860 , 
    n21861 , 
    n21862 , 
    n21863 , 
    n21864 , 
    n21865 , 
    n21866 , 
    n21867 , 
    n21868 , 
    n21869 , 
    n21870 , 
    n21871 , 
    n21872 , 
    n21873 , 
    n21874 , 
    n21875 , 
    n21876 , 
    n21877 , 
    n21878 , 
    n21879 , 
    n21880 , 
    n21881 , 
    n21882 , 
    n21883 , 
    n21884 , 
    n21885 , 
    n21886 , 
    n21887 , 
    n21888 , 
    n21889 , 
    n21890 , 
    n21891 , 
    n21892 , 
    n21893 , 
    n21894 , 
    n21895 , 
    n21896 , 
    n21897 , 
    n21898 , 
    n21899 , 
    n21900 , 
    n21901 , 
    n21902 , 
    n21903 , 
    n21904 , 
    n21905 , 
    n21906 , 
    n21907 , 
    n21908 , 
    n21909 , 
    n21910 , 
    n21911 , 
    n21912 , 
    n21913 , 
    n21914 , 
    n21915 , 
    n21916 , 
    n21917 , 
    n21918 , 
    n21919 , 
    n21920 , 
    n21921 , 
    n21922 , 
    n21923 , 
    n21924 , 
    n21925 , 
    n21926 , 
    n21927 , 
    n21928 , 
    n21929 , 
    n21930 , 
    n21931 , 
    n21932 , 
    n21933 , 
    n21934 , 
    n21935 , 
    n21936 , 
    n21937 , 
    n21938 , 
    n21939 , 
    n21940 , 
    n21941 , 
    n21942 , 
    n21943 , 
    n21944 , 
    n21945 , 
    n21946 , 
    n21947 , 
    n21948 , 
    n21949 , 
    n21950 , 
    n21951 , 
    n21952 , 
    n21953 , 
    n21954 , 
    n21955 , 
    n21956 , 
    n21957 , 
    n21958 , 
    n21959 , 
    n21960 , 
    n21961 , 
    n21962 , 
    n21963 , 
    n21964 , 
    n21965 , 
    n21966 , 
    n21967 , 
    n21968 , 
    n21969 , 
    n21970 , 
    n21971 , 
    n21972 , 
    n21973 , 
    n21974 , 
    n21975 , 
    n21976 , 
    n21977 , 
    n21978 , 
    n21979 , 
    n21980 , 
    n21981 , 
    n21982 , 
    n21983 , 
    n21984 , 
    n21985 , 
    n21986 , 
    n21987 , 
    n21988 , 
    n21989 , 
    n21990 , 
    n21991 , 
    n21992 , 
    n21993 , 
    n21994 , 
    n21995 , 
    n21996 , 
    n21997 , 
    n21998 , 
    n21999 , 
    n22000 , 
    n22001 , 
    n22002 , 
    n22003 , 
    n22004 , 
    n22005 , 
    n22006 , 
    n22007 , 
    n22008 , 
    n22009 , 
    n22010 , 
    n22011 , 
    n22012 , 
    n22013 , 
    n22014 , 
    n22015 , 
    n22016 , 
    n22017 , 
    n22018 , 
    n22019 , 
    n22020 , 
    n22021 , 
    n22022 , 
    n22023 , 
    n22024 , 
    n22025 , 
    n22026 , 
    n22027 , 
    n22028 , 
    n22029 , 
    n22030 , 
    n22031 , 
    n22032 , 
    n22033 , 
    n22034 , 
    n22035 , 
    n22036 , 
    n22037 , 
    n22038 , 
    n22039 , 
    n22040 , 
    n22041 , 
    n22042 , 
    n22043 , 
    n22044 , 
    n22045 , 
    n22046 , 
    n22047 , 
    n22048 , 
    n22049 , 
    n22050 , 
    n22051 , 
    n22052 , 
    n22053 , 
    n22054 , 
    n22055 , 
    n22056 , 
    n22057 , 
    n22058 , 
    n22059 , 
    n22060 , 
    n22061 , 
    n22062 , 
    n22063 , 
    n22064 , 
    n22065 , 
    n22066 , 
    n22067 , 
    n22068 , 
    n22069 , 
    n22070 , 
    n22071 , 
    n22072 , 
    n22073 , 
    n22074 , 
    n22075 , 
    n22076 , 
    n22077 , 
    n22078 , 
    n22079 , 
    n22080 , 
    n22081 , 
    n22082 , 
    n22083 , 
    n22084 , 
    n22085 , 
    n22086 , 
    n22087 , 
    n22088 , 
    n22089 , 
    n22090 , 
    n22091 , 
    n22092 , 
    n22093 , 
    n22094 , 
    n22095 , 
    n22096 , 
    n22097 , 
    n22098 , 
    n22099 , 
    n22100 , 
    n22101 , 
    n22102 , 
    n22103 , 
    n22104 , 
    n22105 , 
    n22106 , 
    n22107 , 
    n22108 , 
    n22109 , 
    n22110 , 
    n22111 , 
    n22112 , 
    n22113 , 
    n22114 , 
    n22115 , 
    n22116 , 
    n22117 , 
    n22118 , 
    n22119 , 
    n22120 , 
    n22121 , 
    n22122 , 
    n22123 , 
    n22124 , 
    n22125 , 
    n22126 , 
    n22127 , 
    n22128 , 
    n22129 , 
    n22130 , 
    n22131 , 
    n22132 , 
    n22133 , 
    n22134 , 
    n22135 , 
    n22136 , 
    n22137 , 
    n22138 , 
    n22139 , 
    n22140 , 
    n22141 , 
    n22142 , 
    n22143 , 
    n22144 , 
    n22145 , 
    n22146 , 
    n22147 , 
    n22148 , 
    n22149 , 
    n22150 , 
    n22151 , 
    n22152 , 
    n22153 , 
    n22154 , 
    n22155 , 
    n22156 , 
    n22157 , 
    n22158 , 
    n22159 , 
    n22160 , 
    n22161 , 
    n22162 , 
    n22163 , 
    n22164 , 
    n22165 , 
    n22166 , 
    n22167 , 
    n22168 , 
    n22169 , 
    n22170 , 
    n22171 , 
    n22172 , 
    n22173 , 
    n22174 , 
    n22175 , 
    n22176 , 
    n22177 , 
    n22178 , 
    n22179 , 
    n22180 , 
    n22181 , 
    n22182 , 
    n22183 , 
    n22184 , 
    n22185 , 
    n22186 , 
    n22187 , 
    n22188 , 
    n22189 , 
    n22190 , 
    n22191 , 
    n22192 , 
    n22193 , 
    n22194 , 
    n22195 , 
    n22196 , 
    n22197 , 
    n22198 , 
    n22199 , 
    n22200 , 
    n22201 , 
    n22202 , 
    n22203 , 
    n22204 , 
    n22205 , 
    n22206 , 
    n22207 , 
    n22208 , 
    n22209 , 
    n22210 , 
    n22211 , 
    n22212 , 
    n22213 , 
    n22214 , 
    n22215 , 
    n22216 , 
    n22217 , 
    n22218 , 
    n22219 , 
    n22220 , 
    n22221 , 
    n22222 , 
    n22223 , 
    n22224 , 
    n22225 , 
    n22226 , 
    n22227 , 
    n22228 , 
    n22229 , 
    n22230 , 
    n22231 , 
    n22232 , 
    n22233 , 
    n22234 , 
    n22235 , 
    n22236 , 
    n22237 , 
    n22238 , 
    n22239 , 
    n22240 , 
    n22241 , 
    n22242 , 
    n22243 , 
    n22244 , 
    n22245 , 
    n22246 , 
    n22247 , 
    n22248 , 
    n22249 , 
    n22250 , 
    n22251 , 
    n22252 , 
    n22253 , 
    n22254 , 
    n22255 , 
    n22256 , 
    n22257 , 
    n22258 , 
    n22259 , 
    n22260 , 
    n22261 , 
    n22262 , 
    n22263 , 
    n22264 , 
    n22265 , 
    n22266 , 
    n22267 , 
    n22268 , 
    n22269 , 
    n22270 , 
    n22271 , 
    n22272 , 
    n22273 , 
    n22274 , 
    n22275 , 
    n22276 , 
    n22277 , 
    n22278 , 
    n22279 , 
    n22280 , 
    n22281 , 
    n22282 , 
    n22283 , 
    n22284 , 
    n22285 , 
    n22286 , 
    n22287 , 
    n22288 , 
    n22289 , 
    n22290 , 
    n22291 , 
    n22292 , 
    n22293 , 
    n22294 , 
    n22295 , 
    n22296 , 
    n22297 , 
    n22298 , 
    n22299 , 
    n22300 , 
    n22301 , 
    n22302 , 
    n22303 , 
    n22304 , 
    n22305 , 
    n22306 , 
    n22307 , 
    n22308 , 
    n22309 , 
    n22310 , 
    n22311 , 
    n22312 , 
    n22313 , 
    n22314 , 
    n22315 , 
    n22316 , 
    n22317 , 
    n22318 , 
    n22319 , 
    n22320 , 
    n22321 , 
    n22322 , 
    n22323 , 
    n22324 , 
    n22325 , 
    n22326 , 
    n22327 , 
    n22328 , 
    n22329 , 
    n22330 , 
    n22331 , 
    n22332 , 
    n22333 , 
    n22334 , 
    n22335 , 
    n22336 , 
    n22337 , 
    n22338 , 
    n22339 , 
    n22340 , 
    n22341 , 
    n22342 , 
    n22343 , 
    n22344 , 
    n22345 , 
    n22346 , 
    n22347 , 
    n22348 , 
    n22349 , 
    n22350 , 
    n22351 , 
    n22352 , 
    n22353 , 
    n22354 , 
    n22355 , 
    n22356 , 
    n22357 , 
    n22358 , 
    n22359 , 
    n22360 , 
    n22361 , 
    n22362 , 
    n22363 , 
    n22364 , 
    n22365 , 
    n22366 , 
    n22367 , 
    n22368 , 
    n22369 , 
    n22370 , 
    n22371 , 
    n22372 , 
    n22373 , 
    n22374 , 
    n22375 , 
    n22376 , 
    n22377 , 
    n22378 , 
    n22379 , 
    n22380 , 
    n22381 , 
    n22382 , 
    n22383 , 
    n22384 , 
    n22385 , 
    n22386 , 
    n22387 , 
    n22388 , 
    n22389 , 
    n22390 , 
    n22391 , 
    n22392 , 
    n22393 , 
    n22394 , 
    n22395 , 
    n22396 , 
    n22397 , 
    n22398 , 
    n22399 , 
    n22400 , 
    n22401 , 
    n22402 , 
    n22403 , 
    n22404 , 
    n22405 , 
    n22406 , 
    n22407 , 
    n22408 , 
    n22409 , 
    n22410 , 
    n22411 , 
    n22412 , 
    n22413 , 
    n22414 , 
    n22415 , 
    n22416 , 
    n22417 , 
    n22418 , 
    n22419 , 
    n22420 , 
    n22421 , 
    n22422 , 
    n22423 , 
    n22424 , 
    n22425 , 
    n22426 , 
    n22427 , 
    n22428 , 
    n22429 , 
    n22430 , 
    n22431 , 
    n22432 , 
    n22433 , 
    n22434 , 
    n22435 , 
    n22436 , 
    n22437 , 
    n22438 , 
    n22439 , 
    n22440 , 
    n22441 , 
    n22442 , 
    n22443 , 
    n22444 , 
    n22445 , 
    n22446 , 
    n22447 , 
    n22448 , 
    n22449 , 
    n22450 , 
    n22451 , 
    n22452 , 
    n22453 , 
    n22454 , 
    n22455 , 
    n22456 , 
    n22457 , 
    n22458 , 
    n22459 , 
    n22460 , 
    n22461 , 
    n22462 , 
    n22463 , 
    n22464 , 
    n22465 , 
    n22466 , 
    n22467 , 
    n22468 , 
    n22469 , 
    n22470 , 
    n22471 , 
    n22472 , 
    n22473 , 
    n22474 , 
    n22475 , 
    n22476 , 
    n22477 , 
    n22478 , 
    n22479 , 
    n22480 , 
    n22481 , 
    n22482 , 
    n22483 , 
    n22484 , 
    n22485 , 
    n22486 , 
    n22487 , 
    n22488 , 
    n22489 , 
    n22490 , 
    n22491 , 
    n22492 , 
    n22493 , 
    n22494 , 
    n22495 , 
    n22496 , 
    n22497 , 
    n22498 , 
    n22499 , 
    n22500 , 
    n22501 , 
    n22502 , 
    n22503 , 
    n22504 , 
    n22505 , 
    n22506 , 
    n22507 , 
    n22508 , 
    n22509 , 
    n22510 , 
    n22511 , 
    n22512 , 
    n22513 , 
    n22514 , 
    n22515 , 
    n22516 , 
    n22517 , 
    n22518 , 
    n22519 , 
    n22520 , 
    n22521 , 
    n22522 , 
    n22523 , 
    n22524 , 
    n22525 , 
    n22526 , 
    n22527 , 
    n22528 , 
    n22529 , 
    n22530 , 
    n22531 , 
    n22532 , 
    n22533 , 
    n22534 , 
    n22535 , 
    n22536 , 
    n22537 , 
    n22538 , 
    n22539 , 
    n22540 , 
    n22541 , 
    n22542 , 
    n22543 , 
    n22544 , 
    n22545 , 
    n22546 , 
    n22547 , 
    n22548 , 
    n22549 , 
    n22550 , 
    n22551 , 
    n22552 , 
    n22553 , 
    n22554 , 
    n22555 , 
    n22556 , 
    n22557 , 
    n22558 , 
    n22559 , 
    n22560 , 
    n22561 , 
    n22562 , 
    n22563 , 
    n22564 , 
    n22565 , 
    n22566 , 
    n22567 , 
    n22568 , 
    n22569 , 
    n22570 , 
    n22571 , 
    n22572 , 
    n22573 , 
    n22574 , 
    n22575 , 
    n22576 , 
    n22577 , 
    n22578 , 
    n22579 , 
    n22580 , 
    n22581 , 
    n22582 , 
    n22583 , 
    n22584 , 
    n22585 , 
    n22586 , 
    n22587 , 
    n22588 , 
    n22589 , 
    n22590 , 
    n22591 , 
    n22592 , 
    n22593 , 
    n22594 , 
    n22595 , 
    n22596 , 
    n22597 , 
    n22598 , 
    n22599 , 
    n22600 , 
    n22601 , 
    n22602 , 
    n22603 , 
    n22604 , 
    n22605 , 
    n22606 , 
    n22607 , 
    n22608 , 
    n22609 , 
    n22610 , 
    n22611 , 
    n22612 , 
    n22613 , 
    n22614 , 
    n22615 , 
    n22616 , 
    n22617 , 
    n22618 , 
    n22619 , 
    n22620 , 
    n22621 , 
    n22622 , 
    n22623 , 
    n22624 , 
    n22625 , 
    n22626 , 
    n22627 , 
    n22628 , 
    n22629 , 
    n22630 , 
    n22631 , 
    n22632 , 
    n22633 , 
    n22634 , 
    n22635 , 
    n22636 , 
    n22637 , 
    n22638 , 
    n22639 , 
    n22640 , 
    n22641 , 
    n22642 , 
    n22643 , 
    n22644 , 
    n22645 , 
    n22646 , 
    n22647 , 
    n22648 , 
    n22649 , 
    n22650 , 
    n22651 , 
    n22652 , 
    n22653 , 
    n22654 , 
    n22655 , 
    n22656 , 
    n22657 , 
    n22658 , 
    n22659 , 
    n22660 , 
    n22661 , 
    n22662 , 
    n22663 , 
    n22664 , 
    n22665 , 
    n22666 , 
    n22667 , 
    n22668 , 
    n22669 , 
    n22670 , 
    n22671 , 
    n22672 , 
    n22673 , 
    n22674 , 
    n22675 , 
    n22676 , 
    n22677 , 
    n22678 , 
    n22679 , 
    n22680 , 
    n22681 , 
    n22682 , 
    n22683 , 
    n22684 , 
    n22685 , 
    n22686 , 
    n22687 , 
    n22688 , 
    n22689 , 
    n22690 , 
    n22691 , 
    n22692 , 
    n22693 , 
    n22694 , 
    n22695 , 
    n22696 , 
    n22697 , 
    n22698 , 
    n22699 , 
    n22700 , 
    n22701 , 
    n22702 , 
    n22703 , 
    n22704 , 
    n22705 , 
    n22706 , 
    n22707 , 
    n22708 , 
    n22709 , 
    n22710 , 
    n22711 , 
    n22712 , 
    n22713 , 
    n22714 , 
    n22715 , 
    n22716 , 
    n22717 , 
    n22718 , 
    n22719 , 
    n22720 , 
    n22721 , 
    n22722 , 
    n22723 , 
    n22724 , 
    n22725 , 
    n22726 , 
    n22727 , 
    n22728 , 
    n22729 , 
    n22730 , 
    n22731 , 
    n22732 , 
    n22733 , 
    n22734 , 
    n22735 , 
    n22736 , 
    n22737 , 
    n22738 , 
    n22739 , 
    n22740 , 
    n22741 , 
    n22742 , 
    n22743 , 
    n22744 , 
    n22745 , 
    n22746 , 
    n22747 , 
    n22748 , 
    n22749 , 
    n22750 , 
    n22751 , 
    n22752 , 
    n22753 , 
    n22754 , 
    n22755 , 
    n22756 , 
    n22757 , 
    n22758 , 
    n22759 , 
    n22760 , 
    n22761 , 
    n22762 , 
    n22763 , 
    n22764 , 
    n22765 , 
    n22766 , 
    n22767 , 
    n22768 , 
    n22769 , 
    n22770 , 
    n22771 , 
    n22772 , 
    n22773 , 
    n22774 , 
    n22775 , 
    n22776 , 
    n22777 , 
    n22778 , 
    n22779 , 
    n22780 , 
    n22781 , 
    n22782 , 
    n22783 , 
    n22784 , 
    n22785 , 
    n22786 , 
    n22787 , 
    n22788 , 
    n22789 , 
    n22790 , 
    n22791 , 
    n22792 , 
    n22793 , 
    n22794 , 
    n22795 , 
    n22796 , 
    n22797 , 
    n22798 , 
    n22799 , 
    n22800 , 
    n22801 , 
    n22802 , 
    n22803 , 
    n22804 , 
    n22805 , 
    n22806 , 
    n22807 , 
    n22808 , 
    n22809 , 
    n22810 , 
    n22811 , 
    n22812 , 
    n22813 , 
    n22814 , 
    n22815 , 
    n22816 , 
    n22817 , 
    n22818 , 
    n22819 , 
    n22820 , 
    n22821 , 
    n22822 , 
    n22823 , 
    n22824 , 
    n22825 , 
    n22826 , 
    n22827 , 
    n22828 , 
    n22829 , 
    n22830 , 
    n22831 , 
    n22832 , 
    n22833 , 
    n22834 , 
    n22835 , 
    n22836 , 
    n22837 , 
    n22838 , 
    n22839 , 
    n22840 , 
    n22841 , 
    n22842 , 
    n22843 , 
    n22844 , 
    n22845 , 
    n22846 , 
    n22847 , 
    n22848 , 
    n22849 , 
    n22850 , 
    n22851 , 
    n22852 , 
    n22853 , 
    n22854 , 
    n22855 , 
    n22856 , 
    n22857 , 
    n22858 , 
    n22859 , 
    n22860 , 
    n22861 , 
    n22862 , 
    n22863 , 
    n22864 , 
    n22865 , 
    n22866 , 
    n22867 , 
    n22868 , 
    n22869 , 
    n22870 , 
    n22871 , 
    n22872 , 
    n22873 , 
    n22874 , 
    n22875 , 
    n22876 , 
    n22877 , 
    n22878 , 
    n22879 , 
    n22880 , 
    n22881 , 
    n22882 , 
    n22883 , 
    n22884 , 
    n22885 , 
    n22886 , 
    n22887 , 
    n22888 , 
    n22889 , 
    n22890 , 
    n22891 , 
    n22892 , 
    n22893 , 
    n22894 , 
    n22895 , 
    n22896 , 
    n22897 , 
    n22898 , 
    n22899 , 
    n22900 , 
    n22901 , 
    n22902 , 
    n22903 , 
    n22904 , 
    n22905 , 
    n22906 , 
    n22907 , 
    n22908 , 
    n22909 , 
    n22910 , 
    n22911 , 
    n22912 , 
    n22913 , 
    n22914 , 
    n22915 , 
    n22916 , 
    n22917 , 
    n22918 , 
    n22919 , 
    n22920 , 
    n22921 , 
    n22922 , 
    n22923 , 
    n22924 , 
    n22925 , 
    n22926 , 
    n22927 , 
    n22928 , 
    n22929 , 
    n22930 , 
    n22931 , 
    n22932 , 
    n22933 , 
    n22934 , 
    n22935 , 
    n22936 , 
    n22937 , 
    n22938 , 
    n22939 , 
    n22940 , 
    n22941 , 
    n22942 , 
    n22943 , 
    n22944 , 
    n22945 , 
    n22946 , 
    n22947 , 
    n22948 , 
    n22949 , 
    n22950 , 
    n22951 , 
    n22952 , 
    n22953 , 
    n22954 , 
    n22955 , 
    n22956 , 
    n22957 , 
    n22958 , 
    n22959 , 
    n22960 , 
    n22961 , 
    n22962 , 
    n22963 , 
    n22964 , 
    n22965 , 
    n22966 , 
    n22967 , 
    n22968 , 
    n22969 , 
    n22970 , 
    n22971 , 
    n22972 , 
    n22973 , 
    n22974 , 
    n22975 , 
    n22976 , 
    n22977 , 
    n22978 , 
    n22979 , 
    n22980 , 
    n22981 , 
    n22982 , 
    n22983 , 
    n22984 , 
    n22985 , 
    n22986 , 
    n22987 , 
    n22988 , 
    n22989 , 
    n22990 , 
    n22991 , 
    n22992 , 
    n22993 , 
    n22994 , 
    n22995 , 
    n22996 , 
    n22997 , 
    n22998 , 
    n22999 , 
    n23000 , 
    n23001 , 
    n23002 , 
    n23003 , 
    n23004 , 
    n23005 , 
    n23006 , 
    n23007 , 
    n23008 , 
    n23009 , 
    n23010 , 
    n23011 , 
    n23012 , 
    n23013 , 
    n23014 , 
    n23015 , 
    n23016 , 
    n23017 , 
    n23018 , 
    n23019 , 
    n23020 , 
    n23021 , 
    n23022 , 
    n23023 , 
    n23024 , 
    n23025 , 
    n23026 , 
    n23027 , 
    n23028 , 
    n23029 , 
    n23030 , 
    n23031 , 
    n23032 , 
    n23033 , 
    n23034 , 
    n23035 , 
    n23036 , 
    n23037 , 
    n23038 , 
    n23039 , 
    n23040 , 
    n23041 , 
    n23042 , 
    n23043 , 
    n23044 , 
    n23045 , 
    n23046 , 
    n23047 , 
    n23048 , 
    n23049 , 
    n23050 , 
    n23051 , 
    n23052 , 
    n23053 , 
    n23054 , 
    n23055 , 
    n23056 , 
    n23057 , 
    n23058 , 
    n23059 , 
    n23060 , 
    n23061 , 
    n23062 , 
    n23063 , 
    n23064 , 
    n23065 , 
    n23066 , 
    n23067 , 
    n23068 , 
    n23069 , 
    n23070 , 
    n23071 , 
    n23072 , 
    n23073 , 
    n23074 , 
    n23075 , 
    n23076 , 
    n23077 , 
    n23078 , 
    n23079 , 
    n23080 , 
    n23081 , 
    n23082 , 
    n23083 , 
    n23084 , 
    n23085 , 
    n23086 , 
    n23087 , 
    n23088 , 
    n23089 , 
    n23090 , 
    n23091 , 
    n23092 , 
    n23093 , 
    n23094 , 
    n23095 , 
    n23096 , 
    n23097 , 
    n23098 , 
    n23099 , 
    n23100 , 
    n23101 , 
    n23102 , 
    n23103 , 
    n23104 , 
    n23105 , 
    n23106 , 
    n23107 , 
    n23108 , 
    n23109 , 
    n23110 , 
    n23111 , 
    n23112 , 
    n23113 , 
    n23114 , 
    n23115 , 
    n23116 , 
    n23117 , 
    n23118 , 
    n23119 , 
    n23120 , 
    n23121 , 
    n23122 , 
    n23123 , 
    n23124 , 
    n23125 , 
    n23126 , 
    n23127 , 
    n23128 , 
    n23129 , 
    n23130 , 
    n23131 , 
    n23132 , 
    n23133 , 
    n23134 , 
    n23135 , 
    n23136 , 
    n23137 , 
    n23138 , 
    n23139 , 
    n23140 , 
    n23141 , 
    n23142 , 
    n23143 , 
    n23144 , 
    n23145 , 
    n23146 , 
    n23147 , 
    n23148 , 
    n23149 , 
    n23150 , 
    n23151 , 
    n23152 , 
    n23153 , 
    n23154 , 
    n23155 , 
    n23156 , 
    n23157 , 
    n23158 , 
    n23159 , 
    n23160 , 
    n23161 , 
    n23162 , 
    n23163 , 
    n23164 , 
    n23165 , 
    n23166 , 
    n23167 , 
    n23168 , 
    n23169 , 
    n23170 , 
    n23171 , 
    n23172 , 
    n23173 , 
    n23174 , 
    n23175 , 
    n23176 , 
    n23177 , 
    n23178 , 
    n23179 , 
    n23180 , 
    n23181 , 
    n23182 , 
    n23183 , 
    n23184 , 
    n23185 , 
    n23186 , 
    n23187 , 
    n23188 , 
    n23189 , 
    n23190 , 
    n23191 , 
    n23192 , 
    n23193 , 
    n23194 , 
    n23195 , 
    n23196 , 
    n23197 , 
    n23198 , 
    n23199 , 
    n23200 , 
    n23201 , 
    n23202 , 
    n23203 , 
    n23204 , 
    n23205 , 
    n23206 , 
    n23207 , 
    n23208 , 
    n23209 , 
    n23210 , 
    n23211 , 
    n23212 , 
    n23213 , 
    n23214 , 
    n23215 , 
    n23216 , 
    n23217 , 
    n23218 , 
    n23219 , 
    n23220 , 
    n23221 , 
    n23222 , 
    n23223 , 
    n23224 , 
    n23225 , 
    n23226 , 
    n23227 , 
    n23228 , 
    n23229 , 
    n23230 , 
    n23231 , 
    n23232 , 
    n23233 , 
    n23234 , 
    n23235 , 
    n23236 , 
    n23237 , 
    n23238 , 
    n23239 , 
    n23240 , 
    n23241 , 
    n23242 , 
    n23243 , 
    n23244 , 
    n23245 , 
    n23246 , 
    n23247 , 
    n23248 , 
    n23249 , 
    n23250 , 
    n23251 , 
    n23252 , 
    n23253 , 
    n23254 , 
    n23255 , 
    n23256 , 
    n23257 , 
    n23258 , 
    n23259 , 
    n23260 , 
    n23261 , 
    n23262 , 
    n23263 , 
    n23264 , 
    n23265 , 
    n23266 , 
    n23267 , 
    n23268 , 
    n23269 , 
    n23270 , 
    n23271 , 
    n23272 , 
    n23273 , 
    n23274 , 
    n23275 , 
    n23276 , 
    n23277 , 
    n23278 , 
    n23279 , 
    n23280 , 
    n23281 , 
    n23282 , 
    n23283 , 
    n23284 , 
    n23285 , 
    n23286 , 
    n23287 , 
    n23288 , 
    n23289 , 
    n23290 , 
    n23291 , 
    n23292 , 
    n23293 , 
    n23294 , 
    n23295 , 
    n23296 , 
    n23297 , 
    n23298 , 
    n23299 , 
    n23300 , 
    n23301 , 
    n23302 , 
    n23303 , 
    n23304 , 
    n23305 , 
    n23306 , 
    n23307 , 
    n23308 , 
    n23309 , 
    n23310 , 
    n23311 , 
    n23312 , 
    n23313 , 
    n23314 , 
    n23315 , 
    n23316 , 
    n23317 , 
    n23318 , 
    n23319 , 
    n23320 , 
    n23321 , 
    n23322 , 
    n23323 , 
    n23324 , 
    n23325 , 
    n23326 , 
    n23327 , 
    n23328 , 
    n23329 , 
    n23330 , 
    n23331 , 
    n23332 , 
    n23333 , 
    n23334 , 
    n23335 , 
    n23336 , 
    n23337 , 
    n23338 , 
    n23339 , 
    n23340 , 
    n23341 , 
    n23342 , 
    n23343 , 
    n23344 , 
    n23345 , 
    n23346 , 
    n23347 , 
    n23348 , 
    n23349 , 
    n23350 , 
    n23351 , 
    n23352 , 
    n23353 , 
    n23354 , 
    n23355 , 
    n23356 , 
    n23357 , 
    n23358 , 
    n23359 , 
    n23360 , 
    n23361 , 
    n23362 , 
    n23363 , 
    n23364 , 
    n23365 , 
    n23366 , 
    n23367 , 
    n23368 , 
    n23369 , 
    n23370 , 
    n23371 , 
    n23372 , 
    n23373 , 
    n23374 , 
    n23375 , 
    n23376 , 
    n23377 , 
    n23378 , 
    n23379 , 
    n23380 , 
    n23381 , 
    n23382 , 
    n23383 , 
    n23384 , 
    n23385 , 
    n23386 , 
    n23387 , 
    n23388 , 
    n23389 , 
    n23390 , 
    n23391 , 
    n23392 , 
    n23393 , 
    n23394 , 
    n23395 , 
    n23396 , 
    n23397 , 
    n23398 , 
    n23399 , 
    n23400 , 
    n23401 , 
    n23402 , 
    n23403 , 
    n23404 , 
    n23405 , 
    n23406 , 
    n23407 , 
    n23408 , 
    n23409 , 
    n23410 , 
    n23411 , 
    n23412 , 
    n23413 , 
    n23414 , 
    n23415 , 
    n23416 , 
    n23417 , 
    n23418 , 
    n23419 , 
    n23420 , 
    n23421 , 
    n23422 , 
    n23423 , 
    n23424 , 
    n23425 , 
    n23426 , 
    n23427 , 
    n23428 , 
    n23429 , 
    n23430 , 
    n23431 , 
    n23432 , 
    n23433 , 
    n23434 , 
    n23435 , 
    n23436 , 
    n23437 , 
    n23438 , 
    n23439 , 
    n23440 , 
    n23441 , 
    n23442 , 
    n23443 , 
    n23444 , 
    n23445 , 
    n23446 , 
    n23447 , 
    n23448 , 
    n23449 , 
    n23450 , 
    n23451 , 
    n23452 , 
    n23453 , 
    n23454 , 
    n23455 , 
    n23456 , 
    n23457 , 
    n23458 , 
    n23459 , 
    n23460 , 
    n23461 , 
    n23462 , 
    n23463 , 
    n23464 , 
    n23465 , 
    n23466 , 
    n23467 , 
    n23468 , 
    n23469 , 
    n23470 , 
    n23471 , 
    n23472 , 
    n23473 , 
    n23474 , 
    n23475 , 
    n23476 , 
    n23477 , 
    n23478 , 
    n23479 , 
    n23480 , 
    n23481 , 
    n23482 , 
    n23483 , 
    n23484 , 
    n23485 , 
    n23486 , 
    n23487 , 
    n23488 , 
    n23489 , 
    n23490 , 
    n23491 , 
    n23492 , 
    n23493 , 
    n23494 , 
    n23495 , 
    n23496 , 
    n23497 , 
    n23498 , 
    n23499 , 
    n23500 , 
    n23501 , 
    n23502 , 
    n23503 , 
    n23504 , 
    n23505 , 
    n23506 , 
    n23507 , 
    n23508 , 
    n23509 , 
    n23510 , 
    n23511 , 
    n23512 , 
    n23513 , 
    n23514 , 
    n23515 , 
    n23516 , 
    n23517 , 
    n23518 , 
    n23519 , 
    n23520 , 
    n23521 , 
    n23522 , 
    n23523 , 
    n23524 , 
    n23525 , 
    n23526 , 
    n23527 , 
    n23528 , 
    n23529 , 
    n23530 , 
    n23531 , 
    n23532 , 
    n23533 , 
    n23534 , 
    n23535 , 
    n23536 , 
    n23537 , 
    n23538 , 
    n23539 , 
    n23540 , 
    n23541 , 
    n23542 , 
    n23543 , 
    n23544 , 
    n23545 , 
    n23546 , 
    n23547 , 
    n23548 , 
    n23549 , 
    n23550 , 
    n23551 , 
    n23552 , 
    n23553 , 
    n23554 , 
    n23555 , 
    n23556 , 
    n23557 , 
    n23558 , 
    n23559 , 
    n23560 , 
    n23561 , 
    n23562 , 
    n23563 , 
    n23564 , 
    n23565 , 
    n23566 , 
    n23567 , 
    n23568 , 
    n23569 , 
    n23570 , 
    n23571 , 
    n23572 , 
    n23573 , 
    n23574 , 
    n23575 , 
    n23576 , 
    n23577 , 
    n23578 , 
    n23579 , 
    n23580 , 
    n23581 , 
    n23582 , 
    n23583 , 
    n23584 , 
    n23585 , 
    n23586 , 
    n23587 , 
    n23588 , 
    n23589 , 
    n23590 , 
    n23591 , 
    n23592 , 
    n23593 , 
    n23594 , 
    n23595 , 
    n23596 , 
    n23597 , 
    n23598 , 
    n23599 , 
    n23600 , 
    n23601 , 
    n23602 , 
    n23603 , 
    n23604 , 
    n23605 , 
    n23606 , 
    n23607 , 
    n23608 , 
    n23609 , 
    n23610 , 
    n23611 , 
    n23612 , 
    n23613 , 
    n23614 , 
    n23615 , 
    n23616 , 
    n23617 , 
    n23618 , 
    n23619 , 
    n23620 , 
    n23621 , 
    n23622 , 
    n23623 , 
    n23624 , 
    n23625 , 
    n23626 , 
    n23627 , 
    n23628 , 
    n23629 , 
    n23630 , 
    n23631 , 
    n23632 , 
    n23633 , 
    n23634 , 
    n23635 , 
    n23636 , 
    n23637 , 
    n23638 , 
    n23639 , 
    n23640 , 
    n23641 , 
    n23642 , 
    n23643 , 
    n23644 , 
    n23645 , 
    n23646 , 
    n23647 , 
    n23648 , 
    n23649 , 
    n23650 , 
    n23651 , 
    n23652 , 
    n23653 , 
    n23654 , 
    n23655 , 
    n23656 , 
    n23657 , 
    n23658 , 
    n23659 , 
    n23660 , 
    n23661 , 
    n23662 , 
    n23663 , 
    n23664 , 
    n23665 , 
    n23666 , 
    n23667 , 
    n23668 , 
    n23669 , 
    n23670 , 
    n23671 , 
    n23672 , 
    n23673 , 
    n23674 , 
    n23675 , 
    n23676 , 
    n23677 , 
    n23678 , 
    n23679 , 
    n23680 , 
    n23681 , 
    n23682 , 
    n23683 , 
    n23684 , 
    n23685 , 
    n23686 , 
    n23687 , 
    n23688 , 
    n23689 , 
    n23690 , 
    n23691 , 
    n23692 , 
    n23693 , 
    n23694 , 
    n23695 , 
    n23696 , 
    n23697 , 
    n23698 , 
    n23699 , 
    n23700 , 
    n23701 , 
    n23702 , 
    n23703 , 
    n23704 , 
    n23705 , 
    n23706 , 
    n23707 , 
    n23708 , 
    n23709 , 
    n23710 , 
    n23711 , 
    n23712 , 
    n23713 , 
    n23714 , 
    n23715 , 
    n23716 , 
    n23717 , 
    n23718 , 
    n23719 , 
    n23720 , 
    n23721 , 
    n23722 , 
    n23723 , 
    n23724 , 
    n23725 , 
    n23726 , 
    n23727 , 
    n23728 , 
    n23729 , 
    n23730 , 
    n23731 , 
    n23732 , 
    n23733 , 
    n23734 , 
    n23735 , 
    n23736 , 
    n23737 , 
    n23738 , 
    n23739 , 
    n23740 , 
    n23741 , 
    n23742 , 
    n23743 , 
    n23744 , 
    n23745 , 
    n23746 , 
    n23747 , 
    n23748 , 
    n23749 , 
    n23750 , 
    n23751 , 
    n23752 , 
    n23753 , 
    n23754 , 
    n23755 , 
    n23756 , 
    n23757 , 
    n23758 , 
    n23759 , 
    n23760 , 
    n23761 , 
    n23762 , 
    n23763 , 
    n23764 , 
    n23765 , 
    n23766 , 
    n23767 , 
    n23768 , 
    n23769 , 
    n23770 , 
    n23771 , 
    n23772 , 
    n23773 , 
    n23774 , 
    n23775 , 
    n23776 , 
    n23777 , 
    n23778 , 
    n23779 , 
    n23780 , 
    n23781 , 
    n23782 , 
    n23783 , 
    n23784 , 
    n23785 , 
    n23786 , 
    n23787 , 
    n23788 , 
    n23789 , 
    n23790 , 
    n23791 , 
    n23792 , 
    n23793 , 
    n23794 , 
    n23795 , 
    n23796 , 
    n23797 , 
    n23798 , 
    n23799 , 
    n23800 , 
    n23801 , 
    n23802 , 
    n23803 , 
    n23804 , 
    n23805 , 
    n23806 , 
    n23807 , 
    n23808 , 
    n23809 , 
    n23810 , 
    n23811 , 
    n23812 , 
    n23813 , 
    n23814 , 
    n23815 , 
    n23816 , 
    n23817 , 
    n23818 , 
    n23819 , 
    n23820 , 
    n23821 , 
    n23822 , 
    n23823 , 
    n23824 , 
    n23825 , 
    n23826 , 
    n23827 , 
    n23828 , 
    n23829 , 
    n23830 , 
    n23831 , 
    n23832 , 
    n23833 , 
    n23834 , 
    n23835 , 
    n23836 , 
    n23837 , 
    n23838 , 
    n23839 , 
    n23840 , 
    n23841 , 
    n23842 , 
    n23843 , 
    n23844 , 
    n23845 , 
    n23846 , 
    n23847 , 
    n23848 , 
    n23849 , 
    n23850 , 
    n23851 , 
    n23852 , 
    n23853 , 
    n23854 , 
    n23855 , 
    n23856 , 
    n23857 , 
    n23858 , 
    n23859 , 
    n23860 , 
    n23861 , 
    n23862 , 
    n23863 , 
    n23864 , 
    n23865 , 
    n23866 , 
    n23867 , 
    n23868 , 
    n23869 , 
    n23870 , 
    n23871 , 
    n23872 , 
    n23873 , 
    n23874 , 
    n23875 , 
    n23876 , 
    n23877 , 
    n23878 , 
    n23879 , 
    n23880 , 
    n23881 , 
    n23882 , 
    n23883 , 
    n23884 , 
    n23885 , 
    n23886 , 
    n23887 , 
    n23888 , 
    n23889 , 
    n23890 , 
    n23891 , 
    n23892 , 
    n23893 , 
    n23894 , 
    n23895 , 
    n23896 , 
    n23897 , 
    n23898 , 
    n23899 , 
    n23900 , 
    n23901 , 
    n23902 , 
    n23903 , 
    n23904 , 
    n23905 , 
    n23906 , 
    n23907 , 
    n23908 , 
    n23909 , 
    n23910 , 
    n23911 , 
    n23912 , 
    n23913 , 
    n23914 , 
    n23915 , 
    n23916 , 
    n23917 , 
    n23918 , 
    n23919 , 
    n23920 , 
    n23921 , 
    n23922 , 
    n23923 , 
    n23924 , 
    n23925 , 
    n23926 , 
    n23927 , 
    n23928 , 
    n23929 , 
    n23930 , 
    n23931 , 
    n23932 , 
    n23933 , 
    n23934 , 
    n23935 , 
    n23936 , 
    n23937 , 
    n23938 , 
    n23939 , 
    n23940 , 
    n23941 , 
    n23942 , 
    n23943 , 
    n23944 , 
    n23945 , 
    n23946 , 
    n23947 , 
    n23948 , 
    n23949 , 
    n23950 , 
    n23951 , 
    n23952 , 
    n23953 , 
    n23954 , 
    n23955 , 
    n23956 , 
    n23957 , 
    n23958 , 
    n23959 , 
    n23960 , 
    n23961 , 
    n23962 , 
    n23963 , 
    n23964 , 
    n23965 , 
    n23966 , 
    n23967 , 
    n23968 , 
    n23969 , 
    n23970 , 
    n23971 , 
    n23972 , 
    n23973 , 
    n23974 , 
    n23975 , 
    n23976 , 
    n23977 , 
    n23978 , 
    n23979 , 
    n23980 , 
    n23981 , 
    n23982 , 
    n23983 , 
    n23984 , 
    n23985 , 
    n23986 , 
    n23987 , 
    n23988 , 
    n23989 , 
    n23990 , 
    n23991 , 
    n23992 , 
    n23993 , 
    n23994 , 
    n23995 , 
    n23996 , 
    n23997 , 
    n23998 , 
    n23999 , 
    n24000 , 
    n24001 , 
    n24002 , 
    n24003 , 
    n24004 , 
    n24005 , 
    n24006 , 
    n24007 , 
    n24008 , 
    n24009 , 
    n24010 , 
    n24011 , 
    n24012 , 
    n24013 , 
    n24014 , 
    n24015 , 
    n24016 , 
    n24017 , 
    n24018 , 
    n24019 , 
    n24020 , 
    n24021 , 
    n24022 , 
    n24023 , 
    n24024 , 
    n24025 , 
    n24026 , 
    n24027 , 
    n24028 , 
    n24029 , 
    n24030 , 
    n24031 , 
    n24032 , 
    n24033 , 
    n24034 , 
    n24035 , 
    n24036 , 
    n24037 , 
    n24038 , 
    n24039 , 
    n24040 , 
    n24041 , 
    n24042 , 
    n24043 , 
    n24044 , 
    n24045 , 
    n24046 , 
    n24047 , 
    n24048 , 
    n24049 , 
    n24050 , 
    n24051 , 
    n24052 , 
    n24053 , 
    n24054 , 
    n24055 , 
    n24056 , 
    n24057 , 
    n24058 , 
    n24059 , 
    n24060 , 
    n24061 , 
    n24062 , 
    n24063 , 
    n24064 , 
    n24065 , 
    n24066 , 
    n24067 , 
    n24068 , 
    n24069 , 
    n24070 , 
    n24071 , 
    n24072 , 
    n24073 , 
    n24074 , 
    n24075 , 
    n24076 , 
    n24077 , 
    n24078 , 
    n24079 , 
    n24080 , 
    n24081 , 
    n24082 , 
    n24083 , 
    n24084 , 
    n24085 , 
    n24086 , 
    n24087 , 
    n24088 , 
    n24089 , 
    n24090 , 
    n24091 , 
    n24092 , 
    n24093 , 
    n24094 , 
    n24095 , 
    n24096 , 
    n24097 , 
    n24098 , 
    n24099 , 
    n24100 , 
    n24101 , 
    n24102 , 
    n24103 , 
    n24104 , 
    n24105 , 
    n24106 , 
    n24107 , 
    n24108 , 
    n24109 , 
    n24110 , 
    n24111 , 
    n24112 , 
    n24113 , 
    n24114 , 
    n24115 , 
    n24116 , 
    n24117 , 
    n24118 , 
    n24119 , 
    n24120 , 
    n24121 , 
    n24122 , 
    n24123 , 
    n24124 , 
    n24125 , 
    n24126 , 
    n24127 , 
    n24128 , 
    n24129 , 
    n24130 , 
    n24131 , 
    n24132 , 
    n24133 , 
    n24134 , 
    n24135 , 
    n24136 , 
    n24137 , 
    n24138 , 
    n24139 , 
    n24140 , 
    n24141 , 
    n24142 , 
    n24143 , 
    n24144 , 
    n24145 , 
    n24146 , 
    n24147 , 
    n24148 , 
    n24149 , 
    n24150 , 
    n24151 , 
    n24152 , 
    n24153 , 
    n24154 , 
    n24155 , 
    n24156 , 
    n24157 , 
    n24158 , 
    n24159 , 
    n24160 , 
    n24161 , 
    n24162 , 
    n24163 , 
    n24164 , 
    n24165 , 
    n24166 , 
    n24167 , 
    n24168 , 
    n24169 , 
    n24170 , 
    n24171 , 
    n24172 , 
    n24173 , 
    n24174 , 
    n24175 , 
    n24176 , 
    n24177 , 
    n24178 , 
    n24179 , 
    n24180 , 
    n24181 , 
    n24182 , 
    n24183 , 
    n24184 , 
    n24185 , 
    n24186 , 
    n24187 , 
    n24188 , 
    n24189 , 
    n24190 , 
    n24191 , 
    n24192 , 
    n24193 , 
    n24194 , 
    n24195 , 
    n24196 , 
    n24197 , 
    n24198 , 
    n24199 , 
    n24200 , 
    n24201 , 
    n24202 , 
    n24203 , 
    n24204 , 
    n24205 , 
    n24206 , 
    n24207 , 
    n24208 , 
    n24209 , 
    n24210 , 
    n24211 , 
    n24212 , 
    n24213 , 
    n24214 , 
    n24215 , 
    n24216 , 
    n24217 , 
    n24218 , 
    n24219 , 
    n24220 , 
    n24221 , 
    n24222 , 
    n24223 , 
    n24224 , 
    n24225 , 
    n24226 , 
    n24227 , 
    n24228 , 
    n24229 , 
    n24230 , 
    n24231 , 
    n24232 , 
    n24233 , 
    n24234 , 
    n24235 , 
    n24236 , 
    n24237 , 
    n24238 , 
    n24239 , 
    n24240 , 
    n24241 , 
    n24242 , 
    n24243 , 
    n24244 , 
    n24245 , 
    n24246 , 
    n24247 , 
    n24248 , 
    n24249 , 
    n24250 , 
    n24251 , 
    n24252 , 
    n24253 , 
    n24254 , 
    n24255 , 
    n24256 , 
    n24257 , 
    n24258 , 
    n24259 , 
    n24260 , 
    n24261 , 
    n24262 , 
    n24263 , 
    n24264 , 
    n24265 , 
    n24266 , 
    n24267 , 
    n24268 , 
    n24269 , 
    n24270 , 
    n24271 , 
    n24272 , 
    n24273 , 
    n24274 , 
    n24275 , 
    n24276 , 
    n24277 , 
    n24278 , 
    n24279 , 
    n24280 , 
    n24281 , 
    n24282 , 
    n24283 , 
    n24284 , 
    n24285 , 
    n24286 , 
    n24287 , 
    n24288 , 
    n24289 , 
    n24290 , 
    n24291 , 
    n24292 , 
    n24293 , 
    n24294 , 
    n24295 , 
    n24296 , 
    n24297 , 
    n24298 , 
    n24299 , 
    n24300 , 
    n24301 , 
    n24302 , 
    n24303 , 
    n24304 , 
    n24305 , 
    n24306 , 
    n24307 , 
    n24308 , 
    n24309 , 
    n24310 , 
    n24311 , 
    n24312 , 
    n24313 , 
    n24314 , 
    n24315 , 
    n24316 , 
    n24317 , 
    n24318 , 
    n24319 , 
    n24320 , 
    n24321 , 
    n24322 , 
    n24323 , 
    n24324 , 
    n24325 , 
    n24326 , 
    n24327 , 
    n24328 , 
    n24329 , 
    n24330 , 
    n24331 , 
    n24332 , 
    n24333 , 
    n24334 , 
    n24335 , 
    n24336 , 
    n24337 , 
    n24338 , 
    n24339 , 
    n24340 , 
    n24341 , 
    n24342 , 
    n24343 , 
    n24344 , 
    n24345 , 
    n24346 , 
    n24347 , 
    n24348 , 
    n24349 , 
    n24350 , 
    n24351 , 
    n24352 , 
    n24353 , 
    n24354 , 
    n24355 , 
    n24356 , 
    n24357 , 
    n24358 , 
    n24359 , 
    n24360 , 
    n24361 , 
    n24362 , 
    n24363 , 
    n24364 , 
    n24365 , 
    n24366 , 
    n24367 , 
    n24368 , 
    n24369 , 
    n24370 , 
    n24371 , 
    n24372 , 
    n24373 , 
    n24374 , 
    n24375 , 
    n24376 , 
    n24377 , 
    n24378 , 
    n24379 , 
    n24380 , 
    n24381 , 
    n24382 , 
    n24383 , 
    n24384 , 
    n24385 , 
    n24386 , 
    n24387 , 
    n24388 , 
    n24389 , 
    n24390 , 
    n24391 , 
    n24392 , 
    n24393 , 
    n24394 , 
    n24395 , 
    n24396 , 
    n24397 , 
    n24398 , 
    n24399 , 
    n24400 , 
    n24401 , 
    n24402 , 
    n24403 , 
    n24404 , 
    n24405 , 
    n24406 , 
    n24407 , 
    n24408 , 
    n24409 , 
    n24410 , 
    n24411 , 
    n24412 , 
    n24413 , 
    n24414 , 
    n24415 , 
    n24416 , 
    n24417 , 
    n24418 , 
    n24419 , 
    n24420 , 
    n24421 , 
    n24422 , 
    n24423 , 
    n24424 , 
    n24425 , 
    n24426 , 
    n24427 , 
    n24428 , 
    n24429 , 
    n24430 , 
    n24431 , 
    n24432 , 
    n24433 , 
    n24434 , 
    n24435 , 
    n24436 , 
    n24437 , 
    n24438 , 
    n24439 , 
    n24440 , 
    n24441 , 
    n24442 , 
    n24443 , 
    n24444 , 
    n24445 , 
    n24446 , 
    n24447 , 
    n24448 , 
    n24449 , 
    n24450 , 
    n24451 , 
    n24452 , 
    n24453 , 
    n24454 , 
    n24455 , 
    n24456 , 
    n24457 , 
    n24458 , 
    n24459 , 
    n24460 , 
    n24461 , 
    n24462 , 
    n24463 , 
    n24464 , 
    n24465 , 
    n24466 , 
    n24467 , 
    n24468 , 
    n24469 , 
    n24470 , 
    n24471 , 
    n24472 , 
    n24473 , 
    n24474 , 
    n24475 , 
    n24476 , 
    n24477 , 
    n24478 , 
    n24479 , 
    n24480 , 
    n24481 , 
    n24482 , 
    n24483 , 
    n24484 , 
    n24485 , 
    n24486 , 
    n24487 , 
    n24488 , 
    n24489 , 
    n24490 , 
    n24491 , 
    n24492 , 
    n24493 , 
    n24494 , 
    n24495 , 
    n24496 , 
    n24497 , 
    n24498 , 
    n24499 , 
    n24500 , 
    n24501 , 
    n24502 , 
    n24503 , 
    n24504 , 
    n24505 , 
    n24506 , 
    n24507 , 
    n24508 , 
    n24509 , 
    n24510 , 
    n24511 , 
    n24512 , 
    n24513 , 
    n24514 , 
    n24515 , 
    n24516 , 
    n24517 , 
    n24518 , 
    n24519 , 
    n24520 , 
    n24521 , 
    n24522 , 
    n24523 , 
    n24524 , 
    n24525 , 
    n24526 , 
    n24527 , 
    n24528 , 
    n24529 , 
    n24530 , 
    n24531 , 
    n24532 , 
    n24533 , 
    n24534 , 
    n24535 , 
    n24536 , 
    n24537 , 
    n24538 , 
    n24539 , 
    n24540 , 
    n24541 , 
    n24542 , 
    n24543 , 
    n24544 , 
    n24545 , 
    n24546 , 
    n24547 , 
    n24548 , 
    n24549 , 
    n24550 , 
    n24551 , 
    n24552 , 
    n24553 , 
    n24554 , 
    n24555 , 
    n24556 , 
    n24557 , 
    n24558 , 
    n24559 , 
    n24560 , 
    n24561 , 
    n24562 , 
    n24563 , 
    n24564 , 
    n24565 , 
    n24566 , 
    n24567 , 
    n24568 , 
    n24569 , 
    n24570 , 
    n24571 , 
    n24572 , 
    n24573 , 
    n24574 , 
    n24575 , 
    n24576 , 
    n24577 , 
    n24578 , 
    n24579 , 
    n24580 , 
    n24581 , 
    n24582 , 
    n24583 , 
    n24584 , 
    n24585 , 
    n24586 , 
    n24587 , 
    n24588 , 
    n24589 , 
    n24590 , 
    n24591 , 
    n24592 , 
    n24593 , 
    n24594 , 
    n24595 , 
    n24596 , 
    n24597 , 
    n24598 , 
    n24599 , 
    n24600 , 
    n24601 , 
    n24602 , 
    n24603 , 
    n24604 , 
    n24605 , 
    n24606 , 
    n24607 , 
    n24608 , 
    n24609 , 
    n24610 , 
    n24611 , 
    n24612 , 
    n24613 , 
    n24614 , 
    n24615 , 
    n24616 , 
    n24617 , 
    n24618 , 
    n24619 , 
    n24620 , 
    n24621 , 
    n24622 , 
    n24623 , 
    n24624 , 
    n24625 , 
    n24626 , 
    n24627 , 
    n24628 , 
    n24629 , 
    n24630 , 
    n24631 , 
    n24632 , 
    n24633 , 
    n24634 , 
    n24635 , 
    n24636 , 
    n24637 , 
    n24638 , 
    n24639 , 
    n24640 , 
    n24641 , 
    n24642 , 
    n24643 , 
    n24644 , 
    n24645 , 
    n24646 , 
    n24647 , 
    n24648 , 
    n24649 , 
    n24650 , 
    n24651 , 
    n24652 , 
    n24653 , 
    n24654 , 
    n24655 , 
    n24656 , 
    n24657 , 
    n24658 , 
    n24659 , 
    n24660 , 
    n24661 , 
    n24662 , 
    n24663 , 
    n24664 , 
    n24665 , 
    n24666 , 
    n24667 , 
    n24668 , 
    n24669 , 
    n24670 , 
    n24671 , 
    n24672 , 
    n24673 , 
    n24674 , 
    n24675 , 
    n24676 , 
    n24677 , 
    n24678 , 
    n24679 , 
    n24680 , 
    n24681 , 
    n24682 , 
    n24683 , 
    n24684 , 
    n24685 , 
    n24686 , 
    n24687 , 
    n24688 , 
    n24689 , 
    n24690 , 
    n24691 , 
    n24692 , 
    n24693 , 
    n24694 , 
    n24695 , 
    n24696 , 
    n24697 , 
    n24698 , 
    n24699 , 
    n24700 , 
    n24701 , 
    n24702 , 
    n24703 , 
    n24704 , 
    n24705 , 
    n24706 , 
    n24707 , 
    n24708 , 
    n24709 , 
    n24710 , 
    n24711 , 
    n24712 , 
    n24713 , 
    n24714 , 
    n24715 , 
    n24716 , 
    n24717 , 
    n24718 , 
    n24719 , 
    n24720 , 
    n24721 , 
    n24722 , 
    n24723 , 
    n24724 , 
    n24725 , 
    n24726 , 
    n24727 , 
    n24728 , 
    n24729 , 
    n24730 , 
    n24731 , 
    n24732 , 
    n24733 , 
    n24734 , 
    n24735 , 
    n24736 , 
    n24737 , 
    n24738 , 
    n24739 , 
    n24740 , 
    n24741 , 
    n24742 , 
    n24743 , 
    n24744 , 
    n24745 , 
    n24746 , 
    n24747 , 
    n24748 , 
    n24749 , 
    n24750 , 
    n24751 , 
    n24752 , 
    n24753 , 
    n24754 , 
    n24755 , 
    n24756 , 
    n24757 , 
    n24758 , 
    n24759 , 
    n24760 , 
    n24761 , 
    n24762 , 
    n24763 , 
    n24764 , 
    n24765 , 
    n24766 , 
    n24767 , 
    n24768 , 
    n24769 , 
    n24770 , 
    n24771 , 
    n24772 , 
    n24773 , 
    n24774 , 
    n24775 , 
    n24776 , 
    n24777 , 
    n24778 , 
    n24779 , 
    n24780 , 
    n24781 , 
    n24782 , 
    n24783 , 
    n24784 , 
    n24785 , 
    n24786 , 
    n24787 , 
    n24788 , 
    n24789 , 
    n24790 , 
    n24791 , 
    n24792 , 
    n24793 , 
    n24794 , 
    n24795 , 
    n24796 , 
    n24797 , 
    n24798 , 
    n24799 , 
    n24800 , 
    n24801 , 
    n24802 , 
    n24803 , 
    n24804 , 
    n24805 , 
    n24806 , 
    n24807 , 
    n24808 , 
    n24809 , 
    n24810 , 
    n24811 , 
    n24812 , 
    n24813 , 
    n24814 , 
    n24815 , 
    n24816 , 
    n24817 , 
    n24818 , 
    n24819 , 
    n24820 , 
    n24821 , 
    n24822 , 
    n24823 , 
    n24824 , 
    n24825 , 
    n24826 , 
    n24827 , 
    n24828 , 
    n24829 , 
    n24830 , 
    n24831 , 
    n24832 , 
    n24833 , 
    n24834 , 
    n24835 , 
    n24836 , 
    n24837 , 
    n24838 , 
    n24839 , 
    n24840 , 
    n24841 , 
    n24842 , 
    n24843 , 
    n24844 , 
    n24845 , 
    n24846 , 
    n24847 , 
    n24848 , 
    n24849 , 
    n24850 , 
    n24851 , 
    n24852 , 
    n24853 , 
    n24854 , 
    n24855 , 
    n24856 , 
    n24857 , 
    n24858 , 
    n24859 , 
    n24860 , 
    n24861 , 
    n24862 , 
    n24863 , 
    n24864 , 
    n24865 , 
    n24866 , 
    n24867 , 
    n24868 , 
    n24869 , 
    n24870 , 
    n24871 , 
    n24872 , 
    n24873 , 
    n24874 , 
    n24875 , 
    n24876 , 
    n24877 , 
    n24878 , 
    n24879 , 
    n24880 , 
    n24881 , 
    n24882 , 
    n24883 , 
    n24884 , 
    n24885 , 
    n24886 , 
    n24887 , 
    n24888 , 
    n24889 , 
    n24890 , 
    n24891 , 
    n24892 , 
    n24893 , 
    n24894 , 
    n24895 , 
    n24896 , 
    n24897 , 
    n24898 , 
    n24899 , 
    n24900 , 
    n24901 , 
    n24902 , 
    n24903 , 
    n24904 , 
    n24905 , 
    n24906 , 
    n24907 , 
    n24908 , 
    n24909 , 
    n24910 , 
    n24911 , 
    n24912 , 
    n24913 , 
    n24914 , 
    n24915 , 
    n24916 , 
    n24917 , 
    n24918 , 
    n24919 , 
    n24920 , 
    n24921 , 
    n24922 , 
    n24923 , 
    n24924 , 
    n24925 , 
    n24926 , 
    n24927 , 
    n24928 , 
    n24929 , 
    n24930 , 
    n24931 , 
    n24932 , 
    n24933 , 
    n24934 , 
    n24935 , 
    n24936 , 
    n24937 , 
    n24938 , 
    n24939 , 
    n24940 , 
    n24941 , 
    n24942 , 
    n24943 , 
    n24944 , 
    n24945 , 
    n24946 , 
    n24947 , 
    n24948 , 
    n24949 , 
    n24950 , 
    n24951 , 
    n24952 , 
    n24953 , 
    n24954 , 
    n24955 , 
    n24956 , 
    n24957 , 
    n24958 , 
    n24959 , 
    n24960 , 
    n24961 , 
    n24962 , 
    n24963 , 
    n24964 , 
    n24965 , 
    n24966 , 
    n24967 , 
    n24968 , 
    n24969 , 
    n24970 , 
    n24971 , 
    n24972 , 
    n24973 , 
    n24974 , 
    n24975 , 
    n24976 , 
    n24977 , 
    n24978 , 
    n24979 , 
    n24980 , 
    n24981 , 
    n24982 , 
    n24983 , 
    n24984 , 
    n24985 , 
    n24986 , 
    n24987 , 
    n24988 , 
    n24989 , 
    n24990 , 
    n24991 , 
    n24992 , 
    n24993 , 
    n24994 , 
    n24995 , 
    n24996 , 
    n24997 , 
    n24998 , 
    n24999 , 
    n25000 , 
    n25001 , 
    n25002 , 
    n25003 , 
    n25004 , 
    n25005 , 
    n25006 , 
    n25007 , 
    n25008 , 
    n25009 , 
    n25010 , 
    n25011 , 
    n25012 , 
    n25013 , 
    n25014 , 
    n25015 , 
    n25016 , 
    n25017 , 
    n25018 , 
    n25019 , 
    n25020 , 
    n25021 , 
    n25022 , 
    n25023 , 
    n25024 , 
    n25025 , 
    n25026 , 
    n25027 , 
    n25028 , 
    n25029 , 
    n25030 , 
    n25031 , 
    n25032 , 
    n25033 , 
    n25034 , 
    n25035 , 
    n25036 , 
    n25037 , 
    n25038 , 
    n25039 , 
    n25040 , 
    n25041 , 
    n25042 , 
    n25043 , 
    n25044 , 
    n25045 , 
    n25046 , 
    n25047 , 
    n25048 , 
    n25049 , 
    n25050 , 
    n25051 , 
    n25052 , 
    n25053 , 
    n25054 , 
    n25055 , 
    n25056 , 
    n25057 , 
    n25058 , 
    n25059 , 
    n25060 , 
    n25061 , 
    n25062 , 
    n25063 , 
    n25064 , 
    n25065 , 
    n25066 , 
    n25067 , 
    n25068 , 
    n25069 , 
    n25070 , 
    n25071 , 
    n25072 , 
    n25073 , 
    n25074 , 
    n25075 , 
    n25076 , 
    n25077 , 
    n25078 , 
    n25079 , 
    n25080 , 
    n25081 , 
    n25082 , 
    n25083 , 
    n25084 , 
    n25085 , 
    n25086 , 
    n25087 , 
    n25088 , 
    n25089 , 
    n25090 , 
    n25091 , 
    n25092 , 
    n25093 , 
    n25094 , 
    n25095 , 
    n25096 , 
    n25097 , 
    n25098 , 
    n25099 , 
    n25100 , 
    n25101 , 
    n25102 , 
    n25103 , 
    n25104 , 
    n25105 , 
    n25106 , 
    n25107 , 
    n25108 , 
    n25109 , 
    n25110 , 
    n25111 , 
    n25112 , 
    n25113 , 
    n25114 , 
    n25115 , 
    n25116 , 
    n25117 , 
    n25118 , 
    n25119 , 
    n25120 , 
    n25121 , 
    n25122 , 
    n25123 , 
    n25124 , 
    n25125 , 
    n25126 , 
    n25127 , 
    n25128 , 
    n25129 , 
    n25130 , 
    n25131 , 
    n25132 , 
    n25133 , 
    n25134 , 
    n25135 , 
    n25136 , 
    n25137 , 
    n25138 , 
    n25139 , 
    n25140 , 
    n25141 , 
    n25142 , 
    n25143 , 
    n25144 , 
    n25145 , 
    n25146 , 
    n25147 , 
    n25148 , 
    n25149 , 
    n25150 , 
    n25151 , 
    n25152 , 
    n25153 , 
    n25154 , 
    n25155 , 
    n25156 , 
    n25157 , 
    n25158 , 
    n25159 , 
    n25160 , 
    n25161 , 
    n25162 , 
    n25163 , 
    n25164 , 
    n25165 , 
    n25166 , 
    n25167 , 
    n25168 , 
    n25169 , 
    n25170 , 
    n25171 , 
    n25172 , 
    n25173 , 
    n25174 , 
    n25175 , 
    n25176 , 
    n25177 , 
    n25178 , 
    n25179 , 
    n25180 , 
    n25181 , 
    n25182 , 
    n25183 , 
    n25184 , 
    n25185 , 
    n25186 , 
    n25187 , 
    n25188 , 
    n25189 , 
    n25190 , 
    n25191 , 
    n25192 , 
    n25193 , 
    n25194 , 
    n25195 , 
    n25196 , 
    n25197 , 
    n25198 , 
    n25199 , 
    n25200 , 
    n25201 , 
    n25202 , 
    n25203 , 
    n25204 , 
    n25205 , 
    n25206 , 
    n25207 , 
    n25208 , 
    n25209 , 
    n25210 , 
    n25211 , 
    n25212 , 
    n25213 , 
    n25214 , 
    n25215 , 
    n25216 , 
    n25217 , 
    n25218 , 
    n25219 , 
    n25220 , 
    n25221 , 
    n25222 , 
    n25223 , 
    n25224 , 
    n25225 , 
    n25226 , 
    n25227 , 
    n25228 , 
    n25229 , 
    n25230 , 
    n25231 , 
    n25232 , 
    n25233 , 
    n25234 , 
    n25235 , 
    n25236 , 
    n25237 , 
    n25238 , 
    n25239 , 
    n25240 , 
    n25241 , 
    n25242 , 
    n25243 , 
    n25244 , 
    n25245 , 
    n25246 , 
    n25247 , 
    n25248 , 
    n25249 , 
    n25250 , 
    n25251 , 
    n25252 , 
    n25253 , 
    n25254 , 
    n25255 , 
    n25256 , 
    n25257 , 
    n25258 , 
    n25259 , 
    n25260 , 
    n25261 , 
    n25262 , 
    n25263 , 
    n25264 , 
    n25265 , 
    n25266 , 
    n25267 , 
    n25268 , 
    n25269 , 
    n25270 , 
    n25271 , 
    n25272 , 
    n25273 , 
    n25274 , 
    n25275 , 
    n25276 , 
    n25277 , 
    n25278 , 
    n25279 , 
    n25280 , 
    n25281 , 
    n25282 , 
    n25283 , 
    n25284 , 
    n25285 , 
    n25286 , 
    n25287 , 
    n25288 , 
    n25289 , 
    n25290 , 
    n25291 , 
    n25292 , 
    n25293 , 
    n25294 , 
    n25295 , 
    n25296 , 
    n25297 , 
    n25298 , 
    n25299 , 
    n25300 , 
    n25301 , 
    n25302 , 
    n25303 , 
    n25304 , 
    n25305 , 
    n25306 , 
    n25307 , 
    n25308 , 
    n25309 , 
    n25310 , 
    n25311 , 
    n25312 , 
    n25313 , 
    n25314 , 
    n25315 ;
wire n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , 
     n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , 
     n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , 
     n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , 
     n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , 
     n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , 
     n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , 
     n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , 
     n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , 
     n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , 
     n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , 
     n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , 
     n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , 
     n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , 
     n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , 
     n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , 
     n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , 
     n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , 
     n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , 
     n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , 
     n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , 
     n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , 
     n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , 
     n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , 
     n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , 
     n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , 
     n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , 
     n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , 
     n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , 
     n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , 
     n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , 
     n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , 
     n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , 
     n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , 
     n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , 
     n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , 
     n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , 
     n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
     n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
     n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
     n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
     n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
     n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
     n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
     n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
     n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , 
     n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , 
     n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , 
     n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , 
     n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , 
     n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , 
     n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , 
     n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , 
     n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , 
     n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , 
     n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , 
     n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
     n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , 
     n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , 
     n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , 
     n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , 
     n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , 
     n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , 
     n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , 
     n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , 
     n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , 
     n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , 
     n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , 
     n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , 
     n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , 
     n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , 
     n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , 
     n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , 
     n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , 
     n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , 
     n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , 
     n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , 
     n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , 
     n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , 
     n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , 
     n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , 
     n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , 
     n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , 
     n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , 
     n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , 
     n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , 
     n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , 
     n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , 
     n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , 
     n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , 
     n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , 
     n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , 
     n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , 
     n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , 
     n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , 
     n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , 
     n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , 
     n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , 
     n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , 
     n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , 
     n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , 
     n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , 
     n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , 
     n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , 
     n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , 
     n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , 
     n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , 
     n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , 
     n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , 
     n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , 
     n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , 
     n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , 
     n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , 
     n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , 
     n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , 
     n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , 
     n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , 
     n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , 
     n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , 
     n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , 
     n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , 
     n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , 
     n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , 
     n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , 
     n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , 
     n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , 
     n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , 
     n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , 
     n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , 
     n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , 
     n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , 
     n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , 
     n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , 
     n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , 
     n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , 
     n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , 
     n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , 
     n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , 
     n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , 
     n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , 
     n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , 
     n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , 
     n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , 
     n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , 
     n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , 
     n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , 
     n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , 
     n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , 
     n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , 
     n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , 
     n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , 
     n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , 
     n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , 
     n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , 
     n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , 
     n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , 
     n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , 
     n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , 
     n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , 
     n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , 
     n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , 
     n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , 
     n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , 
     n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , 
     n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , 
     n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , 
     n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , 
     n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , 
     n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , 
     n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , 
     n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , 
     n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , 
     n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , 
     n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , 
     n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , 
     n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , 
     n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , 
     n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , 
     n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , 
     n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , 
     n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , 
     n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , 
     n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , 
     n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , 
     n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , 
     n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , 
     n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , 
     n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , 
     n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , 
     n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , 
     n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , 
     n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , 
     n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , 
     n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , 
     n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , 
     n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , 
     n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , 
     n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , 
     n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , 
     n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , 
     n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , 
     n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , 
     n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , 
     n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , 
     n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , 
     n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , 
     n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , 
     n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , 
     n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , 
     n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , 
     n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , 
     n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , 
     n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , 
     n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , 
     n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , 
     n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , 
     n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , 
     n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , 
     n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , 
     n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , 
     n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , 
     n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , 
     n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , 
     n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , 
     n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , 
     n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , 
     n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , 
     n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , 
     n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , 
     n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , 
     n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , 
     n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , 
     n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , 
     n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , 
     n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , 
     n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , 
     n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , 
     n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , 
     n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , 
     n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , 
     n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , 
     n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , 
     n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , 
     n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , 
     n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , 
     n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , 
     n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , 
     n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , 
     n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , 
     n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , 
     n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , 
     n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , 
     n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , 
     n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , 
     n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , 
     n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , 
     n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , 
     n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , 
     n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , 
     n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , 
     n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , 
     n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , 
     n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , 
     n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , 
     n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , 
     n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , 
     n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , 
     n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , 
     n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , 
     n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , 
     n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , 
     n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , 
     n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , 
     n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , 
     n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , 
     n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , 
     n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , 
     n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , 
     n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , 
     n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , 
     n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , 
     n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , 
     n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , 
     n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , 
     n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , 
     n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , 
     n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , 
     n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , 
     n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , 
     n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , 
     n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , 
     n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , 
     n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , 
     n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , 
     n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , 
     n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , 
     n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , 
     n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , 
     n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , 
     n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , 
     n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , 
     n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , 
     n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , 
     n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , 
     n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , 
     n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , 
     n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , 
     n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , 
     n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , 
     n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , 
     n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , 
     n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , 
     n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , 
     n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , 
     n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , 
     n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , 
     n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , 
     n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , 
     n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , 
     n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , 
     n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , 
     n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , 
     n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , 
     n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , 
     n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , 
     n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , 
     n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , 
     n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , 
     n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , 
     n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , 
     n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , 
     n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , 
     n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , 
     n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , 
     n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , 
     n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , 
     n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , 
     n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , 
     n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , 
     n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , 
     n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , 
     n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , 
     n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , 
     n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , 
     n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , 
     n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , 
     n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , 
     n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , 
     n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , 
     n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , 
     n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , 
     n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , 
     n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , 
     n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , 
     n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , 
     n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , 
     n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , 
     n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , 
     n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
     n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , 
     n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , 
     n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , 
     n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , 
     n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , 
     n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , 
     n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , 
     n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , 
     n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , 
     n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , 
     n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , 
     n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , 
     n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , 
     n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , 
     n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , 
     n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , 
     n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , 
     n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , 
     n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , 
     n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , 
     n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , 
     n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , 
     n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , 
     n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , 
     n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , 
     n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , 
     n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , 
     n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , 
     n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , 
     n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , 
     n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , 
     n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , 
     n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , 
     n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , 
     n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , 
     n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , 
     n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , 
     n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , 
     n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , 
     n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , 
     n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , 
     n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , 
     n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , 
     n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , 
     n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , 
     n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , 
     n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , 
     n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , 
     n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , 
     n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , 
     n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , 
     n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , 
     n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , 
     n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , 
     n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , 
     n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , 
     n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , 
     n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , 
     n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , 
     n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , 
     n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , 
     n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , 
     n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , 
     n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , 
     n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , 
     n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , 
     n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , 
     n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , 
     n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , 
     n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , 
     n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , 
     n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , 
     n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , 
     n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , 
     n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , 
     n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , 
     n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , 
     n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , 
     n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , 
     n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , 
     n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , 
     n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , 
     n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , 
     n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , 
     n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , 
     n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , 
     n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , 
     n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , 
     n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , 
     n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , 
     n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , 
     n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , 
     n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , 
     n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , 
     n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , 
     n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , 
     n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , 
     n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , 
     n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , 
     n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , 
     n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , 
     n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , 
     n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , 
     n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , 
     n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , 
     n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , 
     n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , 
     n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , 
     n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , 
     n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , 
     n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , 
     n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , 
     n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , 
     n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , 
     n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , 
     n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , 
     n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , 
     n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , 
     n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , 
     n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , 
     n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , 
     n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , 
     n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , 
     n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , 
     n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , 
     n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , 
     n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , 
     n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , 
     n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , 
     n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , 
     n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , 
     n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , 
     n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , 
     n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , 
     n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , 
     n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , 
     n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , 
     n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , 
     n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , 
     n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , 
     n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , 
     n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , 
     n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , 
     n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , 
     n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , 
     n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , 
     n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , 
     n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , 
     n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , 
     n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , 
     n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , 
     n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , 
     n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , 
     n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , 
     n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , 
     n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , 
     n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , 
     n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , 
     n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , 
     n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , 
     n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , 
     n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , 
     n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , 
     n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , 
     n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , 
     n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , 
     n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , 
     n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , 
     n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , 
     n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , 
     n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , 
     n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , 
     n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , 
     n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , 
     n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , 
     n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , 
     n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , 
     n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , 
     n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , 
     n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , 
     n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , 
     n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , 
     n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , 
     n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , 
     n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , 
     n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , 
     n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , 
     n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , 
     n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , 
     n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , 
     n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , 
     n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , 
     n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , 
     n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , 
     n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , 
     n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , 
     n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , 
     n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , 
     n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , 
     n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , 
     n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , 
     n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , 
     n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , 
     n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , 
     n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , 
     n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , 
     n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , 
     n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , 
     n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , 
     n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , 
     n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , 
     n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , 
     n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , 
     n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , 
     n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , 
     n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , 
     n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , 
     n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , 
     n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , 
     n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , 
     n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , 
     n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , 
     n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , 
     n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , 
     n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , 
     n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , 
     n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , 
     n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , 
     n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , 
     n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , 
     n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , 
     n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , 
     n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , 
     n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , 
     n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , 
     n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , 
     n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , 
     n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , 
     n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , 
     n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , 
     n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , 
     n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , 
     n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , 
     n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , 
     n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , 
     n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , 
     n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , 
     n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , 
     n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , 
     n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , 
     n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , 
     n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , 
     n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , 
     n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , 
     n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , 
     n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , 
     n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , 
     n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , 
     n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , 
     n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , 
     n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , 
     n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , 
     n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , 
     n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , 
     n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , 
     n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , 
     n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , 
     n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , 
     n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , 
     n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , 
     n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , 
     n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , 
     n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , 
     n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , 
     n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , 
     n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , 
     n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , 
     n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , 
     n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , 
     n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , 
     n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , 
     n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , 
     n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , 
     n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , 
     n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , 
     n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , 
     n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , 
     n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , 
     n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , 
     n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , 
     n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , 
     n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , 
     n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , 
     n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , 
     n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , 
     n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , 
     n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , 
     n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , 
     n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , 
     n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , 
     n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , 
     n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , 
     n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , 
     n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , 
     n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , 
     n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , 
     n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , 
     n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , 
     n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , 
     n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , 
     n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , 
     n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , 
     n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , 
     n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , 
     n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , 
     n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , 
     n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , 
     n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , 
     n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , 
     n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , 
     n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , 
     n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , 
     n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , 
     n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , 
     n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , 
     n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , 
     n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , 
     n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , 
     n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , 
     n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , 
     n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , 
     n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , 
     n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , 
     n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , 
     n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , 
     n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , 
     n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , 
     n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , 
     n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , 
     n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , 
     n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , 
     n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , 
     n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , 
     n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , 
     n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , 
     n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , 
     n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , 
     n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , 
     n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , 
     n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , 
     n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , 
     n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , 
     n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , 
     n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , 
     n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , 
     n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , 
     n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , 
     n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , 
     n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , 
     n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , 
     n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , 
     n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , 
     n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , 
     n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , 
     n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , 
     n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , 
     n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , 
     n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , 
     n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , 
     n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , 
     n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , 
     n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , 
     n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , 
     n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , 
     n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , 
     n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , 
     n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , 
     n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , 
     n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , 
     n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , 
     n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , 
     n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , 
     n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , 
     n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , 
     n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , 
     n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , 
     n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , 
     n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , 
     n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , 
     n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , 
     n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , 
     n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , 
     n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , 
     n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , 
     n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , 
     n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , 
     n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , 
     n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , 
     n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , 
     n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , 
     n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , 
     n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , 
     n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , 
     n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , 
     n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , 
     n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , 
     n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , 
     n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , 
     n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , 
     n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , 
     n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , 
     n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , 
     n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , 
     n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , 
     n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , 
     n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , 
     n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , 
     n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , 
     n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , 
     n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , 
     n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , 
     n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , 
     n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , 
     n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , 
     n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , 
     n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , 
     n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , 
     n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , 
     n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , 
     n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , 
     n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , 
     n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , 
     n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , 
     n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , 
     n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , 
     n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , 
     n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , 
     n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , 
     n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , 
     n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , 
     n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , 
     n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , 
     n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , 
     n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , 
     n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , 
     n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , 
     n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , 
     n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , 
     n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , 
     n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , 
     n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , 
     n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , 
     n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , 
     n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , 
     n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , 
     n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , 
     n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , 
     n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , 
     n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , 
     n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , 
     n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , 
     n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , 
     n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , 
     n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , 
     n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , 
     n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , 
     n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , 
     n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , 
     n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , 
     n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , 
     n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , 
     n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , 
     n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , 
     n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , 
     n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , 
     n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , 
     n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , 
     n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , 
     n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , 
     n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , 
     n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , 
     n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , 
     n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , 
     n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , 
     n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , 
     n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , 
     n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , 
     n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , 
     n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , 
     n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , 
     n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , 
     n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , 
     n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , 
     n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , 
     n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , 
     n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , 
     n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , 
     n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , 
     n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , 
     n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , 
     n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , 
     n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , 
     n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , 
     n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , 
     n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , 
     n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , 
     n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , 
     n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , 
     n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , 
     n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , 
     n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , 
     n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , 
     n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , 
     n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , 
     n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , 
     n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , 
     n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , 
     n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , 
     n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , 
     n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , 
     n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , 
     n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , 
     n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , 
     n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , 
     n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , 
     n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , 
     n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , 
     n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , 
     n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , 
     n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , 
     n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , 
     n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , 
     n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , 
     n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , 
     n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , 
     n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , 
     n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , 
     n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , 
     n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , 
     n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , 
     n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , 
     n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , 
     n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , 
     n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , 
     n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , 
     n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , 
     n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , 
     n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , 
     n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , 
     n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , 
     n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , 
     n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , 
     n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , 
     n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , 
     n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , 
     n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , 
     n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , 
     n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , 
     n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , 
     n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , 
     n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , 
     n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , 
     n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , 
     n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , 
     n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , 
     n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , 
     n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , 
     n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , 
     n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , 
     n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , 
     n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , 
     n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , 
     n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , 
     n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , 
     n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , 
     n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , 
     n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , 
     n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , 
     n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , 
     n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , 
     n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , 
     n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , 
     n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , 
     n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , 
     n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , 
     n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , 
     n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , 
     n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , 
     n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , 
     n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , 
     n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , 
     n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , 
     n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , 
     n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , 
     n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , 
     n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , 
     n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , 
     n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , 
     n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , 
     n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , 
     n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , 
     n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , 
     n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , 
     n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , 
     n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , 
     n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , 
     n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , 
     n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , 
     n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , 
     n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , 
     n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , 
     n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , 
     n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , 
     n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , 
     n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , 
     n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , 
     n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , 
     n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , 
     n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , 
     n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , 
     n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , 
     n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , 
     n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , 
     n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , 
     n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , 
     n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , 
     n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , 
     n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , 
     n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , 
     n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , 
     n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , 
     n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , 
     n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , 
     n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , 
     n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , 
     n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , 
     n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , 
     n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , 
     n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , 
     n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , 
     n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , 
     n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , 
     n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , 
     n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , 
     n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , 
     n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , 
     n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , 
     n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , 
     n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , 
     n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , 
     n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , 
     n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , 
     n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , 
     n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , 
     n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , 
     n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , 
     n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , 
     n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , 
     n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , 
     n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , 
     n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , 
     n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , 
     n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , 
     n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , 
     n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , 
     n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , 
     n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , 
     n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , 
     n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , 
     n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , 
     n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , 
     n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , 
     n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , 
     n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , 
     n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , 
     n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , 
     n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , 
     n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , 
     n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , 
     n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , 
     n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , 
     n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , 
     n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , 
     n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , 
     n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , 
     n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , 
     n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , 
     n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , 
     n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , 
     n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , 
     n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , 
     n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , 
     n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , 
     n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , 
     n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , 
     n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , 
     n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , 
     n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , 
     n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , 
     n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , 
     n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , 
     n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , 
     n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , 
     n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , 
     n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , 
     n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , 
     n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , 
     n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , 
     n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , 
     n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , 
     n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , 
     n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , 
     n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , 
     n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , 
     n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , 
     n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , 
     n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , 
     n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , 
     n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , 
     n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , 
     n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , 
     n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , 
     n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , 
     n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , 
     n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , 
     n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , 
     n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , 
     n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , 
     n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , 
     n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , 
     n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , 
     n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , 
     n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , 
     n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , 
     n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , 
     n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , 
     n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , 
     n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , 
     n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , 
     n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , 
     n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , 
     n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , 
     n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , 
     n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , 
     n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , 
     n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , 
     n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , 
     n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , 
     n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , 
     n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , 
     n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , 
     n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , 
     n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , 
     n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , 
     n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , 
     n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , 
     n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , 
     n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , 
     n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , 
     n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , 
     n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , 
     n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , 
     n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , 
     n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , 
     n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , 
     n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , 
     n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , 
     n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , 
     n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , 
     n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , 
     n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , 
     n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , 
     n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , 
     n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , 
     n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , 
     n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , 
     n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , 
     n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , 
     n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , 
     n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , 
     n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , 
     n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , 
     n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , 
     n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , 
     n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , 
     n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , 
     n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , 
     n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , 
     n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , 
     n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , 
     n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , 
     n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , 
     n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , 
     n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , 
     n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , 
     n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , 
     n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , 
     n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , 
     n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , 
     n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , 
     n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , 
     n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , 
     n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , 
     n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , 
     n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , 
     n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , 
     n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , 
     n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , 
     n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , 
     n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , 
     n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , 
     n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , 
     n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , 
     n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , 
     n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , 
     n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , 
     n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , 
     n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , 
     n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , 
     n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , 
     n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , 
     n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , 
     n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , 
     n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , 
     n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , 
     n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , 
     n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , 
     n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , 
     n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , 
     n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , 
     n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , 
     n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , 
     n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , 
     n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , 
     n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , 
     n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , 
     n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , 
     n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , 
     n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , 
     n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , 
     n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , 
     n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , 
     n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , 
     n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , 
     n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , 
     n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , 
     n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , 
     n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , 
     n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , 
     n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , 
     n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , 
     n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , 
     n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , 
     n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , 
     n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , 
     n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , 
     n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , 
     n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , 
     n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , 
     n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , 
     n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , 
     n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , 
     n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , 
     n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , 
     n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , 
     n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , 
     n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , 
     n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , 
     n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , 
     n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , 
     n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , 
     n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , 
     n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , 
     n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , 
     n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , 
     n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , 
     n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , 
     n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , 
     n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , 
     n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , 
     n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , 
     n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , 
     n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , 
     n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , 
     n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , 
     n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , 
     n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , 
     n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , 
     n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , 
     n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , 
     n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , 
     n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , 
     n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , 
     n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , 
     n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , 
     n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , 
     n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , 
     n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , 
     n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , 
     n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , 
     n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , 
     n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , 
     n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , 
     n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , 
     n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , 
     n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , 
     n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , 
     n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , 
     n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , 
     n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , 
     n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , 
     n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , 
     n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , 
     n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , 
     n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , 
     n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , 
     n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , 
     n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , 
     n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , 
     n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , 
     n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , 
     n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , 
     n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , 
     n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , 
     n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , 
     n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , 
     n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , 
     n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , 
     n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , 
     n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , 
     n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , 
     n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , 
     n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , 
     n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , 
     n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , 
     n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , 
     n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , 
     n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , 
     n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , 
     n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , 
     n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , 
     n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , 
     n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , 
     n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , 
     n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , 
     n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , 
     n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , 
     n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , 
     n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , 
     n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , 
     n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , 
     n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , 
     n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , 
     n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , 
     n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , 
     n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , 
     n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , 
     n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , 
     n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , 
     n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , 
     n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , 
     n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , 
     n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , 
     n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , 
     n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , 
     n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , 
     n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , 
     n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , 
     n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , 
     n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , 
     n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , 
     n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , 
     n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , 
     n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , 
     n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , 
     n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , 
     n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , 
     n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , 
     n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , 
     n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , 
     n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , 
     n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , 
     n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , 
     n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , 
     n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , 
     n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , 
     n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , 
     n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , 
     n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , 
     n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , 
     n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , 
     n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , 
     n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , 
     n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , 
     n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , 
     n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , 
     n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , 
     n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , 
     n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , 
     n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , 
     n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , 
     n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , 
     n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , 
     n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , 
     n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , 
     n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , 
     n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , 
     n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , 
     n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , 
     n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , 
     n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , 
     n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , 
     n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , 
     n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , 
     n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , 
     n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , 
     n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , 
     n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , 
     n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , 
     n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , 
     n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , 
     n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , 
     n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , 
     n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , 
     n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , 
     n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , 
     n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , 
     n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , 
     n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , 
     n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , 
     n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , 
     n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , 
     n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , 
     n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , 
     n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , 
     n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , 
     n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , 
     n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , 
     n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , 
     n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , 
     n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , 
     n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , 
     n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , 
     n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , 
     n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , 
     n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , 
     n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , 
     n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , 
     n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , 
     n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , 
     n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , 
     n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , 
     n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , 
     n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , 
     n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , 
     n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , 
     n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , 
     n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , 
     n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , 
     n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , 
     n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , 
     n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , 
     n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , 
     n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , 
     n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , 
     n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , 
     n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , 
     n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , 
     n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , 
     n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , 
     n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , 
     n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , 
     n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , 
     n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , 
     n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , 
     n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , 
     n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , 
     n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , 
     n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , 
     n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , 
     n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , 
     n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , 
     n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , 
     n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , 
     n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , 
     n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , 
     n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , 
     n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , 
     n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , 
     n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , 
     n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , 
     n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , 
     n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , 
     n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , 
     n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , 
     n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , 
     n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , 
     n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , 
     n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , 
     n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , 
     n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , 
     n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , 
     n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , 
     n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , 
     n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , 
     n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , 
     n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , 
     n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , 
     n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , 
     n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , 
     n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , 
     n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , 
     n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , 
     n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , 
     n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , 
     n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , 
     n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , 
     n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , 
     n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , 
     n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , 
     n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , 
     n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , 
     n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , 
     n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , 
     n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , 
     n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , 
     n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , 
     n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , 
     n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , 
     n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , 
     n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , 
     n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , 
     n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , 
     n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , 
     n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , 
     n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , 
     n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , 
     n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , 
     n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , 
     n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , 
     n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , 
     n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , 
     n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , 
     n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , 
     n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , 
     n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , 
     n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , 
     n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , 
     n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , 
     n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , 
     n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , 
     n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , 
     n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , 
     n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , 
     n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , 
     n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , 
     n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , 
     n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , 
     n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , 
     n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , 
     n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , 
     n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , 
     n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , 
     n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , 
     n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , 
     n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , 
     n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , 
     n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , 
     n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , 
     n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , 
     n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , 
     n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , 
     n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , 
     n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , 
     n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , 
     n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , 
     n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , 
     n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , 
     n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , 
     n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , 
     n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , 
     n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , 
     n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , 
     n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , 
     n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , 
     n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , 
     n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , 
     n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , 
     n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , 
     n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , 
     n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , 
     n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , 
     n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , 
     n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , 
     n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , 
     n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , 
     n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , 
     n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , 
     n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , 
     n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , 
     n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , 
     n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , 
     n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , 
     n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , 
     n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , 
     n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , 
     n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , 
     n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , 
     n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , 
     n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , 
     n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , 
     n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , 
     n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , 
     n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , 
     n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , 
     n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , 
     n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , 
     n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , 
     n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , 
     n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , 
     n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , 
     n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , 
     n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , 
     n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , 
     n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , 
     n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , 
     n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , 
     n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , 
     n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , 
     n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , 
     n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , 
     n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , 
     n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , 
     n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , 
     n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , 
     n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , 
     n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , 
     n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , 
     n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , 
     n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , 
     n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , 
     n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , 
     n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , 
     n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , 
     n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , 
     n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , 
     n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , 
     n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , 
     n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , 
     n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , 
     n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , 
     n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , 
     n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , 
     n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , 
     n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , 
     n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , 
     n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , 
     n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , 
     n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , 
     n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , 
     n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , 
     n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , 
     n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , 
     n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , 
     n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , 
     n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , 
     n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , 
     n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , 
     n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , 
     n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , 
     n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , 
     n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , 
     n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , 
     n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , 
     n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , 
     n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , 
     n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , 
     n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , 
     n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , 
     n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , 
     n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , 
     n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , 
     n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , 
     n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , 
     n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , 
     n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , 
     n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , 
     n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , 
     n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , 
     n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , 
     n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , 
     n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , 
     n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , 
     n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , 
     n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , 
     n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , 
     n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , 
     n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , 
     n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , 
     n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , 
     n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , 
     n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , 
     n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , 
     n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , 
     n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , 
     n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , 
     n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , 
     n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , 
     n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , 
     n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , 
     n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , 
     n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , 
     n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , 
     n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , 
     n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , 
     n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , 
     n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , 
     n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , 
     n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , 
     n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , 
     n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , 
     n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , 
     n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , 
     n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , 
     n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , 
     n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , 
     n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , 
     n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , 
     n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , 
     n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , 
     n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , 
     n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , 
     n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , 
     n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , 
     n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , 
     n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , 
     n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , 
     n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , 
     n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , 
     n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , 
     n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , 
     n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , 
     n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , 
     n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , 
     n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , 
     n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , 
     n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , 
     n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , 
     n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , 
     n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , 
     n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , 
     n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , 
     n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , 
     n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , 
     n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , 
     n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , 
     n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , 
     n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , 
     n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , 
     n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , 
     n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , 
     n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , 
     n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , 
     n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , 
     n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , 
     n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , 
     n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , 
     n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , 
     n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , 
     n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , 
     n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , 
     n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , 
     n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , 
     n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , 
     n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , 
     n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , 
     n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , 
     n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , 
     n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , 
     n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , 
     n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , 
     n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , 
     n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , 
     n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , 
     n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , 
     n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , 
     n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , 
     n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , 
     n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , 
     n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , 
     n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , 
     n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , 
     n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , 
     n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , 
     n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , 
     n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , 
     n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , 
     n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , 
     n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , 
     n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , 
     n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , 
     n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , 
     n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , 
     n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , 
     n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , 
     n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , 
     n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , 
     n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , 
     n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , 
     n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , 
     n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , 
     n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , 
     n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , 
     n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , 
     n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , 
     n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , 
     n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , 
     n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , 
     n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , 
     n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , 
     n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , 
     n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , 
     n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , 
     n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , 
     n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , 
     n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , 
     n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , 
     n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , 
     n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , 
     n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , 
     n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , 
     n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , 
     n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , 
     n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , 
     n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , 
     n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , 
     n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , 
     n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , 
     n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , 
     n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , 
     n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , 
     n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , 
     n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , 
     n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , 
     n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , 
     n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , 
     n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , 
     n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , 
     n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , 
     n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , 
     n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , 
     n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , 
     n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , 
     n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , 
     n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , 
     n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , 
     n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , 
     n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , 
     n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , 
     n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , 
     n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , 
     n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , 
     n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , 
     n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , 
     n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , 
     n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , 
     n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , 
     n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , 
     n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , 
     n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , 
     n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , 
     n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , 
     n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , 
     n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , 
     n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , 
     n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , 
     n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , 
     n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , 
     n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , 
     n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , 
     n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , 
     n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , 
     n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , 
     n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , 
     n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , 
     n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , 
     n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , 
     n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , 
     n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , 
     n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , 
     n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , 
     n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , 
     n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , 
     n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , 
     n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , 
     n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , 
     n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , 
     n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , 
     n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , 
     n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , 
     n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , 
     n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , 
     n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , 
     n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , 
     n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , 
     n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , 
     n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , 
     n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , 
     n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , 
     n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , 
     n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , 
     n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , 
     n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , 
     n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , 
     n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , 
     n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , 
     n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , 
     n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , 
     n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , 
     n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , 
     n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , 
     n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , 
     n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , 
     n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , 
     n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , 
     n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , 
     n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , 
     n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , 
     n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , 
     n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , 
     n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , 
     n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , 
     n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , 
     n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , 
     n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , 
     n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , 
     n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , 
     n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , 
     n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , 
     n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , 
     n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , 
     n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , 
     n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , 
     n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , 
     n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , 
     n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , 
     n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , 
     n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , 
     n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , 
     n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , 
     n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , 
     n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , 
     n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , 
     n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , 
     n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , 
     n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , 
     n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , 
     n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , 
     n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , 
     n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , 
     n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , 
     n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , 
     n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , 
     n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , 
     n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , 
     n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , 
     n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , 
     n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , 
     n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , 
     n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , 
     n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , 
     n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , 
     n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , 
     n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , 
     n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , 
     n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , 
     n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , 
     n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , 
     n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , 
     n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , 
     n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , 
     n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , 
     n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , 
     n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , 
     n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , 
     n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , 
     n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , 
     n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , 
     n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , 
     n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , 
     n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , 
     n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , 
     n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , 
     n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , 
     n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , 
     n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , 
     n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , 
     n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , 
     n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , 
     n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , 
     n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , 
     n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , 
     n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , 
     n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , 
     n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , 
     n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , 
     n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , 
     n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , 
     n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , 
     n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , 
     n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , 
     n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , 
     n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , 
     n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , 
     n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , 
     n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , 
     n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , 
     n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , 
     n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , 
     n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , 
     n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , 
     n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , 
     n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , 
     n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , 
     n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , 
     n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , 
     n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , 
     n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , 
     n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , 
     n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , 
     n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , 
     n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , 
     n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , 
     n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , 
     n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , 
     n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , 
     n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , 
     n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , 
     n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , 
     n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , 
     n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , 
     n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , 
     n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , 
     n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , 
     n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , 
     n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , 
     n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , 
     n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , 
     n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , 
     n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , 
     n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , 
     n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , 
     n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , 
     n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , 
     n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , 
     n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , 
     n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , 
     n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , 
     n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , 
     n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , 
     n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , 
     n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , 
     n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , 
     n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , 
     n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , 
     n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , 
     n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , 
     n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , 
     n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , 
     n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , 
     n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , 
     n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , 
     n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , 
     n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , 
     n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , 
     n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , 
     n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , 
     n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , 
     n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , 
     n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , 
     n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , 
     n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , 
     n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , 
     n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , 
     n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , 
     n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , 
     n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , 
     n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , 
     n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , 
     n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , 
     n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , 
     n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , 
     n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , 
     n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , 
     n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , 
     n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , 
     n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , 
     n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , 
     n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , 
     n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , 
     n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , 
     n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , 
     n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , 
     n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , 
     n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , 
     n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , 
     n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , 
     n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , 
     n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , 
     n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , 
     n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , 
     n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , 
     n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , 
     n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , 
     n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , 
     n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , 
     n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , 
     n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , 
     n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , 
     n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , 
     n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , 
     n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , 
     n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , 
     n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , 
     n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , 
     n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , 
     n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , 
     n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , 
     n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , 
     n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , 
     n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , 
     n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , 
     n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , 
     n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , 
     n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , 
     n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , 
     n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , 
     n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , 
     n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , 
     n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , 
     n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , 
     n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , 
     n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , 
     n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , 
     n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , 
     n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , 
     n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , 
     n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , 
     n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , 
     n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , 
     n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , 
     n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , 
     n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , 
     n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , 
     n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , 
     n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , 
     n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , 
     n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , 
     n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , 
     n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , 
     n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , 
     n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , 
     n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , 
     n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , 
     n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , 
     n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , 
     n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , 
     n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , 
     n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , 
     n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , 
     n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , 
     n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , 
     n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , 
     n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , 
     n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , 
     n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , 
     n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , 
     n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , 
     n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , 
     n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , 
     n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , 
     n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , 
     n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , 
     n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , 
     n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , 
     n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , 
     n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , 
     n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , 
     n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , 
     n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , 
     n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , 
     n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , 
     n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , 
     n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , 
     n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , 
     n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , 
     n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , 
     n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , 
     n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , 
     n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , 
     n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , 
     n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , 
     n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , 
     n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , 
     n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , 
     n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , 
     n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , 
     n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , 
     n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , 
     n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , 
     n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , 
     n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , 
     n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , 
     n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , 
     n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , 
     n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , 
     n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , 
     n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , 
     n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , 
     n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , 
     n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , 
     n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , 
     n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , 
     n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , 
     n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , 
     n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , 
     n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , 
     n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , 
     n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , 
     n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , 
     n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , 
     n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , 
     n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , 
     n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , 
     n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , 
     n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , 
     n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , 
     n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , 
     n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , 
     n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , 
     n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , 
     n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , 
     n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , 
     n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , 
     n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , 
     n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , 
     n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , 
     n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , 
     n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , 
     n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , 
     n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , 
     n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , 
     n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , 
     n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , 
     n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , 
     n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , 
     n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , 
     n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , 
     n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , 
     n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , 
     n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , 
     n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , 
     n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , 
     n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , 
     n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , 
     n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , 
     n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , 
     n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , 
     n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , 
     n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , 
     n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , 
     n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , 
     n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , 
     n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , 
     n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , 
     n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , 
     n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , 
     n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , 
     n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , 
     n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , 
     n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , 
     n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , 
     n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , 
     n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , 
     n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , 
     n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , 
     n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , 
     n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , 
     n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , 
     n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , 
     n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , 
     n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , 
     n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , 
     n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , 
     n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , 
     n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , 
     n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , 
     n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , 
     n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , 
     n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , 
     n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , 
     n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , 
     n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , 
     n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , 
     n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , 
     n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , 
     n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , 
     n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , 
     n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , 
     n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , 
     n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , 
     n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , 
     n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , 
     n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , 
     n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , 
     n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , 
     n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , 
     n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , 
     n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , 
     n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , 
     n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , 
     n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , 
     n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , 
     n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , 
     n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , 
     n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , 
     n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , 
     n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , 
     n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , 
     n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , 
     n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , 
     n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , 
     n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , 
     n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , 
     n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , 
     n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , 
     n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , 
     n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , 
     n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , 
     n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , 
     n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , 
     n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , 
     n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , 
     n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , 
     n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , 
     n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , 
     n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , 
     n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , 
     n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , 
     n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , 
     n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , 
     n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , 
     n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , 
     n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , 
     n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , 
     n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , 
     n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , 
     n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , 
     n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , 
     n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , 
     n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , 
     n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , 
     n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , 
     n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , 
     n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , 
     n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , 
     n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , 
     n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , 
     n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , 
     n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , 
     n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , 
     n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , 
     n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , 
     n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , 
     n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , 
     n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , 
     n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , 
     n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , 
     n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , 
     n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , 
     n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , 
     n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , 
     n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , 
     n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , 
     n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , 
     n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , 
     n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , 
     n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , 
     n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , 
     n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , 
     n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , 
     n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , 
     n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , 
     n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , 
     n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , 
     n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , 
     n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , 
     n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , 
     n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , 
     n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , 
     n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , 
     n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , 
     n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , 
     n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , 
     n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , 
     n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , 
     n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , 
     n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , 
     n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , 
     n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , 
     n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , 
     n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , 
     n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , 
     n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , 
     n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , 
     n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , 
     n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , 
     n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , 
     n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , 
     n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , 
     n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , 
     n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , 
     n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , 
     n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , 
     n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , 
     n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , 
     n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , 
     n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , 
     n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , 
     n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , 
     n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , 
     n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , 
     n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , 
     n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , 
     n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , 
     n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , 
     n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , 
     n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , 
     n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , 
     n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , 
     n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , 
     n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , 
     n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , 
     n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , 
     n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , 
     n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , 
     n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , 
     n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , 
     n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , 
     n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , 
     n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , 
     n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , 
     n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , 
     n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , 
     n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , 
     n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , 
     n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , 
     n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , 
     n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , 
     n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , 
     n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , 
     n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , 
     n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , 
     n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , 
     n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , 
     n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , 
     n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , 
     n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , 
     n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , 
     n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , 
     n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , 
     n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , 
     n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , 
     n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , 
     n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , 
     n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , 
     n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , 
     n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , 
     n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , 
     n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , 
     n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , 
     n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , 
     n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , 
     n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , 
     n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , 
     n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , 
     n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , 
     n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , 
     n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , 
     n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , 
     n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , 
     n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , 
     n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , 
     n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , 
     n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , 
     n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , 
     n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , 
     n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , 
     n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , 
     n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , 
     n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , 
     n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , 
     n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , 
     n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , 
     n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , 
     n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , 
     n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , 
     n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , 
     n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , 
     n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , 
     n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , 
     n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , 
     n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , 
     n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , 
     n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , 
     n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , 
     n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , 
     n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , 
     n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , 
     n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , 
     n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , 
     n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , 
     n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , 
     n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , 
     n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , 
     n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , 
     n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , 
     n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , 
     n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , 
     n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , 
     n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , 
     n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , 
     n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , 
     n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , 
     n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , 
     n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , 
     n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , 
     n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , 
     n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , 
     n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , 
     n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , 
     n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , 
     n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , 
     n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , 
     n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , 
     n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , 
     n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , 
     n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , 
     n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , 
     n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , 
     n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , 
     n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , 
     n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , 
     n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , 
     n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , 
     n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , 
     n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , 
     n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , 
     n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , 
     n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , 
     n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , 
     n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , 
     n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , 
     n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , 
     n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , 
     n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , 
     n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , 
     n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , 
     n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , 
     n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , 
     n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , 
     n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , 
     n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , 
     n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , 
     n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , 
     n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , 
     n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , 
     n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , 
     n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , 
     n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , 
     n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , 
     n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , 
     n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , 
     n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , 
     n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , 
     n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , 
     n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , 
     n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , 
     n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , 
     n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , 
     n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , 
     n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , 
     n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , 
     n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , 
     n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , 
     n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , 
     n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , 
     n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , 
     n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , 
     n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , 
     n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , 
     n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , 
     n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , 
     n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , 
     n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , 
     n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , 
     n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , 
     n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , 
     n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , 
     n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , 
     n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , 
     n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , 
     n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , 
     n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , 
     n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , 
     n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , 
     n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , 
     n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , 
     n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , 
     n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , 
     n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , 
     n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , 
     n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , 
     n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , 
     n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , 
     n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , 
     n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , 
     n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , 
     n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , 
     n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , 
     n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , 
     n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , 
     n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , 
     n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , 
     n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , 
     n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , 
     n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , 
     n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , 
     n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , 
     n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , 
     n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , 
     n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , 
     n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , 
     n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , 
     n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , 
     n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , 
     n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , 
     n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , 
     n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , 
     n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , 
     n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , 
     n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , 
     n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , 
     n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , 
     n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , 
     n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , 
     n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , 
     n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , 
     n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , 
     n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , 
     n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , 
     n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , 
     n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , 
     n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , 
     n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , 
     n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , 
     n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , 
     n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , 
     n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , 
     n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , 
     n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , 
     n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , 
     n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , 
     n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , 
     n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , 
     n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , 
     n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , 
     n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , 
     n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , 
     n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , 
     n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , 
     n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , 
     n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , 
     n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , 
     n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , 
     n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , 
     n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , 
     n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , 
     n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , 
     n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , 
     n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , 
     n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , 
     n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , 
     n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , 
     n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , 
     n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , 
     n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , 
     n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , 
     n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , 
     n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , 
     n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , 
     n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , 
     n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , 
     n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , 
     n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , 
     n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , 
     n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , 
     n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , 
     n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , 
     n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , 
     n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , 
     n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , 
     n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , 
     n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , 
     n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , 
     n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , 
     n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , 
     n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , 
     n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , 
     n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , 
     n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , 
     n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , 
     n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , 
     n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , 
     n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , 
     n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , 
     n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , 
     n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , 
     n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , 
     n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , 
     n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , 
     n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , 
     n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , 
     n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , 
     n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , 
     n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , 
     n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , 
     n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , 
     n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , 
     n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , 
     n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , 
     n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , 
     n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , 
     n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , 
     n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , 
     n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , 
     n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , 
     n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , 
     n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , 
     n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , 
     n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , 
     n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , 
     n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , 
     n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , 
     n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , 
     n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , 
     n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , 
     n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , 
     n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , 
     n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , 
     n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , 
     n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , 
     n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , 
     n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , 
     n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , 
     n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , 
     n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , 
     n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , 
     n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , 
     n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , 
     n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , 
     n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , 
     n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , 
     n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , 
     n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , 
     n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , 
     n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , 
     n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , 
     n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , 
     n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , 
     n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , 
     n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , 
     n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , 
     n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , 
     n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , 
     n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , 
     n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , 
     n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , 
     n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , 
     n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , 
     n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , 
     n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , 
     n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , 
     n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , 
     n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , 
     n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , 
     n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , 
     n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , 
     n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , 
     n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , 
     n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , 
     n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , 
     n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , 
     n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , 
     n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , 
     n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , 
     n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , 
     n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , 
     n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , 
     n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , 
     n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , 
     n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , 
     n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , 
     n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , 
     n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , 
     n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , 
     n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , 
     n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , 
     n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , 
     n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , 
     n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , 
     n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , 
     n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , 
     n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , 
     n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , 
     n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , 
     n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , 
     n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , 
     n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , 
     n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , 
     n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , 
     n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , 
     n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , 
     n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , 
     n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , 
     n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , 
     n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , 
     n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , 
     n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , 
     n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , 
     n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , 
     n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , 
     n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , 
     n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , 
     n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , 
     n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , 
     n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , 
     n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , 
     n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , 
     n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , 
     n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , 
     n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , 
     n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , 
     n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , 
     n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , 
     n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , 
     n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , 
     n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , 
     n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , 
     n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , 
     n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , 
     n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , 
     n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , 
     n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , 
     n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , 
     n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , 
     n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , 
     n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , 
     n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , 
     n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , 
     n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , 
     n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , 
     n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , 
     n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , 
     n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , 
     n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , 
     n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , 
     n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , 
     n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , 
     n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , 
     n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , 
     n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , 
     n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , 
     n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , 
     n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , 
     n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , 
     n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , 
     n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , 
     n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , 
     n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , 
     n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , 
     n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , 
     n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , 
     n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , 
     n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , 
     n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , 
     n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , 
     n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , 
     n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , 
     n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , 
     n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , 
     n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , 
     n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , 
     n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , 
     n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , 
     n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , 
     n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , 
     n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , 
     n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , 
     n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , 
     n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , 
     n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , 
     n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , 
     n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , 
     n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , 
     n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , 
     n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , 
     n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , 
     n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , 
     n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , 
     n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , 
     n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , 
     n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , 
     n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , 
     n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , 
     n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , 
     n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , 
     n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , 
     n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , 
     n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , 
     n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , 
     n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , 
     n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , 
     n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , 
     n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , 
     n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , 
     n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , 
     n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , 
     n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , 
     n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , 
     n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , 
     n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , 
     n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , 
     n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , 
     n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , 
     n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , 
     n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , 
     n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , 
     n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , 
     n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , 
     n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , 
     n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , 
     n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , 
     n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , 
     n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , 
     n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , 
     n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , 
     n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , 
     n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , 
     n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , 
     n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , 
     n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , 
     n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , 
     n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , 
     n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , 
     n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , 
     n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , 
     n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , 
     n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , 
     n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , 
     n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , 
     n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , 
     n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , 
     n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , 
     n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , 
     n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , 
     n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , 
     n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , 
     n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , 
     n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , 
     n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , 
     n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , 
     n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , 
     n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , 
     n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , 
     n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , 
     n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , 
     n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , 
     n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , 
     n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , 
     n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , 
     n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , 
     n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , 
     n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , 
     n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , 
     n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , 
     n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , 
     n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , 
     n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , 
     n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , 
     n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , 
     n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , 
     n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , 
     n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , 
     n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , 
     n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , 
     n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , 
     n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , 
     n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , 
     n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , 
     n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , 
     n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , 
     n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , 
     n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , 
     n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , 
     n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , 
     n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , 
     n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , 
     n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , 
     n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , 
     n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , 
     n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , 
     n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , 
     n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , 
     n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , 
     n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , 
     n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , 
     n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , 
     n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , 
     n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , 
     n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , 
     n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , 
     n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , 
     n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , 
     n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , 
     n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , 
     n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , 
     n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , 
     n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , 
     n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , 
     n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , 
     n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , 
     n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , 
     n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , 
     n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , 
     n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , 
     n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , 
     n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , 
     n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , 
     n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , 
     n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , 
     n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , 
     n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , 
     n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , 
     n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , 
     n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , 
     n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , 
     n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , 
     n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , 
     n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , 
     n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , 
     n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , 
     n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , 
     n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , 
     n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , 
     n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , 
     n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , 
     n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , 
     n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , 
     n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , 
     n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , 
     n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , 
     n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , 
     n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , 
     n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , 
     n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , 
     n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , 
     n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , 
     n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , 
     n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , 
     n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , 
     n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , 
     n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , 
     n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , 
     n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , 
     n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , 
     n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , 
     n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , 
     n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , 
     n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , 
     n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , 
     n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , 
     n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , 
     n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , 
     n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , 
     n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , 
     n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , 
     n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , 
     n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , 
     n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , 
     n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , 
     n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , 
     n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , 
     n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , 
     n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , 
     n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , 
     n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , 
     n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , 
     n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , 
     n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , 
     n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , 
     n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , 
     n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , 
     n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , 
     n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , 
     n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , 
     n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , 
     n56075 , n56076 , n56077 , n56078 ;
buf ( RI19a859b8_2755 , n0 );
buf ( RI19a23510_2794 , n1 );
buf ( RI19a22f70_2797 , n2 );
buf ( RI1754a798_67 , n3 );
buf ( RI19a23e70_2789 , n4 );
buf ( RI19ad04a8_2209 , n5 );
buf ( RI1754c610_2 , n6 );
buf ( RI17465568_1242 , n7 );
buf ( RI19a8fd50_2684 , n8 );
buf ( RI1753aa78_586 , n9 );
buf ( RI1749f948_958 , n10 );
buf ( RI19ab7530_2399 , n11 );
buf ( RI17534808_603 , n12 );
buf ( RI173ba970_1846 , n13 );
buf ( RI17403660_1491 , n14 );
buf ( RI173efea8_1586 , n15 );
buf ( RI174741a8_1170 , n16 );
buf ( RI19a9a160_2611 , n17 );
buf ( RI174bfb80_814 , n18 );
buf ( RI19ac9938_2258 , n19 );
buf ( RI1738f1d0_2058 , n20 );
buf ( RI173d7ec0_1703 , n21 );
buf ( RI1744f998_1348 , n22 );
buf ( RI174cedd8_767 , n23 );
buf ( RI19ac4460_2297 , n24 );
buf ( RI1746f630_1193 , n25 );
buf ( RI19a8a2d8_2723 , n26 );
buf ( RI174b8308_838 , n27 );
buf ( RI19abbe50_2368 , n28 );
buf ( RI1738a658_2081 , n29 );
buf ( RI173d3348_1726 , n30 );
buf ( RI1744ae20_1371 , n31 );
buf ( RI1747e270_1121 , n32 );
buf ( RI19aa5560_2527 , n33 );
buf ( RI174cf300_766 , n34 );
buf ( RI19a869a8_2748 , n35 );
buf ( RI17398f50_2010 , n36 );
buf ( RI173e1c40_1655 , n37 );
buf ( RI17459a60_1299 , n38 );
buf ( RI173a7500_1940 , n39 );
buf ( RI1747dbe0_1123 , n40 );
buf ( RI19a93fe0_2654 , n41 );
buf ( RI174ce8b0_768 , n42 );
buf ( RI19ac4280_2298 , n43 );
buf ( RI173988c0_2012 , n44 );
buf ( RI173e15b0_1657 , n45 );
buf ( RI174593d0_1301 , n46 );
buf ( RI1749b118_980 , n47 );
buf ( RI19aa7e28_2510 , n48 );
buf ( RI1752d698_625 , n49 );
buf ( RI19a89e28_2725 , n50 );
buf ( RI173b5df8_1869 , n51 );
buf ( RI173fee30_1513 , n52 );
buf ( RI173c2620_1808 , n53 );
buf ( RI1740fb40_1431 , n54 );
buf ( RI174944d0_1013 , n55 );
buf ( RI19aaac18_2490 , n56 );
buf ( RI17522c70_658 , n57 );
buf ( RI19aa5a88_2525 , n58 );
buf ( RI173af1b0_1902 , n59 );
buf ( RI173f7ea0_1547 , n60 );
buf ( RI1733d8d0_2141 , n61 );
buf ( RI17468d30_1225 , n62 );
buf ( RI19a8d410_2702 , n63 );
buf ( RI174b1a08_870 , n64 );
buf ( RI19abe4c0_2347 , n65 );
buf ( RI17343168_2114 , n66 );
buf ( RI173cc6e8_1759 , n67 );
buf ( RI17415720_1403 , n68 );
buf ( RI1745d570_1281 , n69 );
buf ( RI17473488_1174 , n70 );
buf ( RI19a99698_2616 , n71 );
buf ( RI174be6e0_818 , n72 );
buf ( RI19ac90c8_2262 , n73 );
buf ( RI1738e4b0_2062 , n74 );
buf ( RI173d71a0_1707 , n75 );
buf ( RI1744ec78_1352 , n76 );
buf ( RI174909c0_1031 , n77 );
buf ( RI19aad468_2473 , n78 );
buf ( RI1751cfa0_676 , n79 );
buf ( RI19abe2e0_2348 , n80 );
buf ( RI173ab6a0_1920 , n81 );
buf ( RI173f4390_1565 , n82 );
buf ( RI1750ecc0_720 , n83 );
buf ( RI17497608_998 , n84 );
buf ( RI19aaa510_2493 , n85 );
buf ( RI17488d10_1069 , n86 );
buf ( RI19aa0970_2564 , n87 );
buf ( RI17510bb0_714 , n88 );
buf ( RI19acf680_2215 , n89 );
buf ( RI173a3d38_1957 , n90 );
buf ( RI173eca28_1602 , n91 );
buf ( RI17483130_1097 , n92 );
buf ( RI174a6590_925 , n93 );
buf ( RI19ab2148_2439 , n94 );
buf ( RI17337cf0_2169 , n95 );
buf ( RI173c1270_1814 , n96 );
buf ( RI17409f60_1459 , n97 );
buf ( RI17460d38_1264 , n98 );
buf ( RI17335c20_2179 , n99 );
buf ( RI17495bc8_1006 , n100 );
buf ( RI19aabb90_2484 , n101 );
buf ( RI17525088_651 , n102 );
buf ( RI19aaf448_2459 , n103 );
buf ( RI173b08a8_1895 , n104 );
buf ( RI173f9598_1540 , n105 );
buf ( RI1738bd50_2074 , n106 );
buf ( RI1746a428_1218 , n107 );
buf ( RI19a8bbb0_2713 , n108 );
buf ( RI174b3100_863 , n109 );
buf ( RI19abd188_2358 , n110 );
buf ( RI17344860_2107 , n111 );
buf ( RI173ce128_1751 , n112 );
buf ( RI17445c18_1396 , n113 );
buf ( RI17444ef8_1400 , n114 );
buf ( RI174a3ae8_938 , n115 );
buf ( RI19ab52f8_2415 , n116 );
buf ( RI17335590_2181 , n117 );
buf ( RI173beb10_1826 , n118 );
buf ( RI17407800_1471 , n119 );
buf ( RI17447ce8_1386 , n120 );
buf ( RI17478690_1149 , n121 );
buf ( RI19a97dc0_2627 , n122 );
buf ( RI174c62a0_794 , n123 );
buf ( RI19ac7b38_2272 , n124 );
buf ( RI17393370_2038 , n125 );
buf ( RI173dc060_1683 , n126 );
buf ( RI17453b38_1328 , n127 );
buf ( RI17465bf8_1240 , n128 );
buf ( RI19a8ffa8_2683 , n129 );
buf ( RI174ae8d0_885 , n130 );
buf ( RI19ac0680_2328 , n131 );
buf ( RI17340030_2129 , n132 );
buf ( RI173c95b0_1774 , n133 );
buf ( RI174125e8_1418 , n134 );
buf ( RI17482de8_1098 , n135 );
buf ( RI19aa3aa8_2540 , n136 );
buf ( RI17507628_743 , n137 );
buf ( RI19a84e00_2760 , n138 );
buf ( RI1739dac8_1987 , n139 );
buf ( RI173e6b00_1631 , n140 );
buf ( RI1745e5d8_1276 , n141 );
buf ( RI17508ff0_738 , n142 );
buf ( RI19a82f88_2773 , n143 );
buf ( RI17475210_1165 , n144 );
buf ( RI19a98630_2623 , n145 );
buf ( RI174c1548_809 , n146 );
buf ( RI19ac81c8_2269 , n147 );
buf ( RI17390238_2053 , n148 );
buf ( RI173d8f28_1698 , n149 );
buf ( RI17450a00_1343 , n150 );
buf ( RI17492a90_1021 , n151 );
buf ( RI19aac6d0_2480 , n152 );
buf ( RI17520330_666 , n153 );
buf ( RI19ab3c00_2425 , n154 );
buf ( RI173ad770_1910 , n155 );
buf ( RI173f6460_1555 , n156 );
buf ( RI1752f060_620 , n157 );
buf ( RI174c8be0_786 , n158 );
buf ( RI174809d0_1109 , n159 );
buf ( RI19aa4a98_2532 , n160 );
buf ( RI17501ef8_754 , n161 );
buf ( RI19a85e68_2753 , n162 );
buf ( RI1739b6b0_1998 , n163 );
buf ( RI173e43a0_1643 , n164 );
buf ( RI1745c1c0_1287 , n165 );
buf ( RI1749df08_966 , n166 );
buf ( RI19ab8d90_2389 , n167 );
buf ( RI17531ec8_611 , n168 );
buf ( RI173b8f30_1854 , n169 );
buf ( RI17401c20_1499 , n170 );
buf ( RI173dfeb8_1664 , n171 );
buf ( RI174a5f00_927 , n172 );
buf ( RI19ab4380_2422 , n173 );
buf ( RI174972c0_999 , n174 );
buf ( RI19aaa330_2494 , n175 );
buf ( RI175274a0_644 , n176 );
buf ( RI19aa12d0_2559 , n177 );
buf ( RI173b1fa0_1888 , n178 );
buf ( RI173fac90_1533 , n179 );
buf ( RI1739b9f8_1997 , n180 );
buf ( RI1746bb20_1211 , n181 );
buf ( RI19a8cb28_2706 , n182 );
buf ( RI174b47f8_856 , n183 );
buf ( RI19abddb8_2351 , n184 );
buf ( RI17345f58_2100 , n185 );
buf ( RI173cf820_1744 , n186 );
buf ( RI17447310_1389 , n187 );
buf ( RI174b6580_847 , n188 );
buf ( RI19abcdc8_2360 , n189 );
buf ( RI174a7fd0_917 , n190 );
buf ( RI19ab3138_2431 , n191 );
buf ( RI17339730_2161 , n192 );
buf ( RI173c2cb0_1806 , n193 );
buf ( RI1740b9a0_1451 , n194 );
buf ( RI173895f0_2086 , n195 );
buf ( RI1747c830_1129 , n196 );
buf ( RI19a93068_2661 , n197 );
buf ( RI174cc9c0_774 , n198 );
buf ( RI19ac3290_2305 , n199 );
buf ( RI17397510_2018 , n200 );
buf ( RI173e0200_1663 , n201 );
buf ( RI17458020_1307 , n202 );
buf ( RI1744fce0_1347 , n203 );
buf ( RI17465f40_1239 , n204 );
buf ( RI19a90188_2682 , n205 );
buf ( RI174aec18_884 , n206 );
buf ( RI19ac0860_2327 , n207 );
buf ( RI17340378_2128 , n208 );
buf ( RI173c98f8_1773 , n209 );
buf ( RI17412930_1417 , n210 );
buf ( RI17483478_1096 , n211 );
buf ( RI19aa3c88_2539 , n212 );
buf ( RI17508078_741 , n213 );
buf ( RI19a85058_2759 , n214 );
buf ( RI1739e158_1985 , n215 );
buf ( RI173e7190_1629 , n216 );
buf ( RI1745ec68_1274 , n217 );
buf ( RI174820c8_1102 , n218 );
buf ( RI19aa3238_2544 , n219 );
buf ( RI174737d0_1173 , n220 );
buf ( RI19a998f0_2615 , n221 );
buf ( RI174bec08_817 , n222 );
buf ( RI19ac92a8_2261 , n223 );
buf ( RI1738e7f8_2061 , n224 );
buf ( RI173d74e8_1706 , n225 );
buf ( RI1744efc0_1351 , n226 );
buf ( RI17491050_1029 , n227 );
buf ( RI19aad648_2472 , n228 );
buf ( RI1751d9f0_674 , n229 );
buf ( RI19abf690_2337 , n230 );
buf ( RI173abd30_1918 , n231 );
buf ( RI173f4a20_1563 , n232 );
buf ( RI17512aa0_708 , n233 );
buf ( RI1751ab88_683 , n234 );
buf ( RI19a23678_2793 , n235 );
buf ( RI17480688_1110 , n236 );
buf ( RI19aa48b8_2533 , n237 );
buf ( RI175019d0_755 , n238 );
buf ( RI19a85c10_2754 , n239 );
buf ( RI1739b368_1999 , n240 );
buf ( RI173e4058_1644 , n241 );
buf ( RI1745be78_1288 , n242 );
buf ( RI1749dbc0_967 , n243 );
buf ( RI19ab8b38_2390 , n244 );
buf ( RI175319a0_612 , n245 );
buf ( RI173b8be8_1855 , n246 );
buf ( RI174018d8_1500 , n247 );
buf ( RI173ddaa0_1675 , n248 );
buf ( RI174b8650_837 , n249 );
buf ( RI19acb300_2246 , n250 );
buf ( RI174613c8_1262 , n251 );
buf ( RI19a91e98_2669 , n252 );
buf ( RI174aa0a0_907 , n253 );
buf ( RI19ac21b0_2313 , n254 );
buf ( RI1733b800_2151 , n255 );
buf ( RI173c4d80_1796 , n256 );
buf ( RI1740da70_1441 , n257 );
buf ( RI1747e5b8_1120 , n258 );
buf ( RI19aa5740_2526 , n259 );
buf ( RI174cf828_765 , n260 );
buf ( RI19a86c00_2747 , n261 );
buf ( RI17399298_2009 , n262 );
buf ( RI173e1f88_1654 , n263 );
buf ( RI17459da8_1298 , n264 );
buf ( RI173a7848_1939 , n265 );
buf ( RI1747df28_1122 , n266 );
buf ( RI19a94238_2653 , n267 );
buf ( RI17398c08_2011 , n268 );
buf ( RI173e18f8_1656 , n269 );
buf ( RI17459718_1300 , n270 );
buf ( RI1748cb68_1050 , n271 );
buf ( RI19aafad8_2456 , n272 );
buf ( RI175172d0_694 , n273 );
buf ( RI19a85508_2757 , n274 );
buf ( RI173a7b90_1938 , n275 );
buf ( RI173f0880_1583 , n276 );
buf ( RI174a9d58_908 , n277 );
buf ( RI173f9c28_1538 , n278 );
buf ( RI17487618_1076 , n279 );
buf ( RI19a9fae8_2571 , n280 );
buf ( RI1750e798_721 , n281 );
buf ( RI19ace870_2221 , n282 );
buf ( RI173a2640_1964 , n283 );
buf ( RI173eb330_1609 , n284 );
buf ( RI17475558_1164 , n285 );
buf ( RI174a4b50_933 , n286 );
buf ( RI19ab36d8_2428 , n287 );
buf ( RI173365f8_2176 , n288 );
buf ( RI173bfb78_1821 , n289 );
buf ( RI17408868_1466 , n290 );
buf ( RI17453160_1331 , n291 );
buf ( RI17335f68_2178 , n292 );
buf ( RI17495f10_1005 , n293 );
buf ( RI19aa9688_2500 , n294 );
buf ( RI175255b0_650 , n295 );
buf ( RI19a981f8_2625 , n296 );
buf ( RI173b0bf0_1894 , n297 );
buf ( RI173f98e0_1539 , n298 );
buf ( RI1738e168_2063 , n299 );
buf ( RI1746a770_1217 , n300 );
buf ( RI19a8be08_2712 , n301 );
buf ( RI174b3448_862 , n302 );
buf ( RI19abd2f0_2357 , n303 );
buf ( RI17344ba8_2106 , n304 );
buf ( RI173ce470_1750 , n305 );
buf ( RI17445f60_1395 , n306 );
buf ( RI17340a08_2126 , n307 );
buf ( RI174a0668_954 , n308 );
buf ( RI19ab7f80_2395 , n309 );
buf ( RI17535ca8_599 , n310 );
buf ( RI173bb690_1842 , n311 );
buf ( RI17404380_1487 , n312 );
buf ( RI173f8f08_1542 , n313 );
buf ( RI17474ec8_1166 , n314 );
buf ( RI19a983d8_2624 , n315 );
buf ( RI174c1020_810 , n316 );
buf ( RI19ac7f70_2270 , n317 );
buf ( RI1738fef0_2054 , n318 );
buf ( RI173d8be0_1699 , n319 );
buf ( RI174506b8_1344 , n320 );
buf ( RI173d39d8_1724 , n321 );
buf ( RI17461710_1261 , n322 );
buf ( RI19a920f0_2668 , n323 );
buf ( RI174aa3e8_906 , n324 );
buf ( RI19ac2390_2312 , n325 );
buf ( RI1733bb48_2150 , n326 );
buf ( RI173c50c8_1795 , n327 );
buf ( RI1740ddb8_1440 , n328 );
buf ( RI1747ec48_1118 , n329 );
buf ( RI19aa5dd0_2524 , n330 );
buf ( RI174d0278_763 , n331 );
buf ( RI19a86fc0_2745 , n332 );
buf ( RI17399928_2007 , n333 );
buf ( RI173e2618_1652 , n334 );
buf ( RI1745a438_1296 , n335 );
buf ( RI17509518_737 , n336 );
buf ( RI19a831e0_2772 , n337 );
buf ( RI174758a0_1163 , n338 );
buf ( RI19a98888_2622 , n339 );
buf ( RI174c1f98_807 , n340 );
buf ( RI19ac8330_2268 , n341 );
buf ( RI173908c8_2051 , n342 );
buf ( RI173d95b8_1696 , n343 );
buf ( RI17451090_1341 , n344 );
buf ( RI17492dd8_1020 , n345 );
buf ( RI19aac838_2479 , n346 );
buf ( RI17520858_665 , n347 );
buf ( RI19ab54d8_2414 , n348 );
buf ( RI173adab8_1909 , n349 );
buf ( RI173f67a8_1554 , n350 );
buf ( RI17532918_609 , n351 );
buf ( RI173b1c58_1889 , n352 );
buf ( RI17488680_1071 , n353 );
buf ( RI19aa05b0_2566 , n354 );
buf ( RI17510160_716 , n355 );
buf ( RI19acf1d0_2217 , n356 );
buf ( RI173a36a8_1959 , n357 );
buf ( RI173ec398_1604 , n358 );
buf ( RI1747e900_1119 , n359 );
buf ( RI17337660_2171 , n360 );
buf ( RI173c0be0_1816 , n361 );
buf ( RI174098d0_1461 , n362 );
buf ( RI1745c508_1286 , n363 );
buf ( RI17405730_1481 , n364 );
buf ( RI17493468_1018 , n365 );
buf ( RI19aaca18_2478 , n366 );
buf ( RI175212a8_663 , n367 );
buf ( RI19ab6cc0_2403 , n368 );
buf ( RI173ae148_1907 , n369 );
buf ( RI173f6e38_1552 , n370 );
buf ( RI17332458_2196 , n371 );
buf ( RI17467980_1231 , n372 );
buf ( RI19a8efb8_2690 , n373 );
buf ( RI174b0658_876 , n374 );
buf ( RI19abfa50_2335 , n375 );
buf ( RI17341db8_2120 , n376 );
buf ( RI173cb338_1765 , n377 );
buf ( RI17414370_1409 , n378 );
buf ( RI174b68c8_846 , n379 );
buf ( RI19abaa28_2376 , n380 );
buf ( RI174a8318_916 , n381 );
buf ( RI19ab0e10_2447 , n382 );
buf ( RI17339a78_2160 , n383 );
buf ( RI173c2ff8_1805 , n384 );
buf ( RI1740bce8_1450 , n385 );
buf ( RI173a0228_1975 , n386 );
buf ( RI1747cb78_1128 , n387 );
buf ( RI19a932c0_2660 , n388 );
buf ( RI174ccee8_773 , n389 );
buf ( RI19ac34e8_2304 , n390 );
buf ( RI17397858_2017 , n391 );
buf ( RI173e0548_1662 , n392 );
buf ( RI17458368_1306 , n393 );
buf ( RI173915e8_2047 , n394 );
buf ( RI17468010_1229 , n395 );
buf ( RI19a8f210_2689 , n396 );
buf ( RI174b0ce8_874 , n397 );
buf ( RI19abfc30_2334 , n398 );
buf ( RI17342448_2118 , n399 );
buf ( RI173cb9c8_1763 , n400 );
buf ( RI17414a00_1407 , n401 );
buf ( RI17485200_1087 , n402 );
buf ( RI19aa2e78_2546 , n403 );
buf ( RI1750aee0_732 , n404 );
buf ( RI19a83f78_2766 , n405 );
buf ( RI1739fee0_1976 , n406 );
buf ( RI173e8f18_1620 , n407 );
buf ( RI174609f0_1265 , n408 );
buf ( RI173e9f80_1615 , n409 );
buf ( RI17477628_1154 , n410 );
buf ( RI19a976b8_2630 , n411 );
buf ( RI174c4e00_798 , n412 );
buf ( RI19ac74a8_2275 , n413 );
buf ( RI17392650_2042 , n414 );
buf ( RI173db340_1687 , n415 );
buf ( RI17452e18_1332 , n416 );
buf ( RI17494ea8_1010 , n417 );
buf ( RI19aab410_2487 , n418 );
buf ( RI17523be8_655 , n419 );
buf ( RI19aaa858_2492 , n420 );
buf ( RI173afb88_1899 , n421 );
buf ( RI173f8878_1544 , n422 );
buf ( RI17344518_2108 , n423 );
buf ( RI1751b0b0_682 , n424 );
buf ( RI19a23858_2792 , n425 );
buf ( RI173c39d0_1802 , n426 );
buf ( RI1749a3f8_984 , n427 );
buf ( RI19aa71f8_2515 , n428 );
buf ( RI1752c1f8_629 , n429 );
buf ( RI19a88460_2736 , n430 );
buf ( RI173b50d8_1873 , n431 );
buf ( RI173fe110_1517 , n432 );
buf ( RI173b95c0_1852 , n433 );
buf ( RI1746ec58_1196 , n434 );
buf ( RI19a89888_2727 , n435 );
buf ( RI174b7930_841 , n436 );
buf ( RI19abb5e0_2372 , n437 );
buf ( RI17389c80_2084 , n438 );
buf ( RI173d2970_1729 , n439 );
buf ( RI1744a448_1374 , n440 );
buf ( RI173d2cb8_1728 , n441 );
buf ( RI174a9380_911 , n442 );
buf ( RI19ab1860_2442 , n443 );
buf ( RI1733aae0_2155 , n444 );
buf ( RI173c4060_1800 , n445 );
buf ( RI1740cd50_1445 , n446 );
buf ( RI17411f58_1420 , n447 );
buf ( RI17491398_1028 , n448 );
buf ( RI19aad828_2471 , n449 );
buf ( RI1751df18_673 , n450 );
buf ( RI19ac0a40_2326 , n451 );
buf ( RI173ac078_1917 , n452 );
buf ( RI173f4d68_1562 , n453 );
buf ( RI17516358_697 , n454 );
buf ( RI1733be90_2149 , n455 );
buf ( RI1749baf0_977 , n456 );
buf ( RI19ab9a38_2383 , n457 );
buf ( RI1752e610_622 , n458 );
buf ( RI173b67d0_1866 , n459 );
buf ( RI173ff808_1510 , n460 );
buf ( RI173c9268_1775 , n461 );
buf ( RI17470350_1189 , n462 );
buf ( RI19a9c5f0_2595 , n463 );
buf ( RI174b9460_834 , n464 );
buf ( RI19acb828_2243 , n465 );
buf ( RI1738b378_2077 , n466 );
buf ( RI173d4068_1722 , n467 );
buf ( RI1744bb40_1367 , n468 );
buf ( RI173dd410_1677 , n469 );
buf ( RI1746b148_1214 , n470 );
buf ( RI19a8c498_2709 , n471 );
buf ( RI174b3e20_859 , n472 );
buf ( RI19abd890_2354 , n473 );
buf ( RI17345580_2103 , n474 );
buf ( RI173cee48_1747 , n475 );
buf ( RI17446938_1392 , n476 );
buf ( RI174a9a10_909 , n477 );
buf ( RI19ab1ef0_2440 , n478 );
buf ( RI1733b170_2153 , n479 );
buf ( RI173c46f0_1798 , n480 );
buf ( RI1740d3e0_1443 , n481 );
buf ( RI175361d0_598 , n482 );
buf ( RI1746f978_1192 , n483 );
buf ( RI19a9bfd8_2598 , n484 );
buf ( RI1738a9a0_2080 , n485 );
buf ( RI173d3690_1725 , n486 );
buf ( RI1744b168_1370 , n487 );
buf ( RI174c7c68_789 , n488 );
buf ( RI19ac6080_2284 , n489 );
buf ( RI1746ae00_1215 , n490 );
buf ( RI19a8c240_2710 , n491 );
buf ( RI174b3ad8_860 , n492 );
buf ( RI19abd6b0_2355 , n493 );
buf ( RI17345238_2104 , n494 );
buf ( RI173ceb00_1748 , n495 );
buf ( RI174465f0_1393 , n496 );
buf ( RI17488338_1072 , n497 );
buf ( RI19aa0358_2567 , n498 );
buf ( RI1750fc38_717 , n499 );
buf ( RI19acef78_2218 , n500 );
buf ( RI173a3360_1960 , n501 );
buf ( RI173ec050_1605 , n502 );
buf ( RI1747c4e8_1130 , n503 );
buf ( RI173a2cd0_1962 , n504 );
buf ( RI174793b0_1145 , n505 );
buf ( RI19a96038_2640 , n506 );
buf ( RI174c7740_790 , n507 );
buf ( RI19ac5e28_2285 , n508 );
buf ( RI17394090_2034 , n509 );
buf ( RI173dcd80_1679 , n510 );
buf ( RI17454858_1324 , n511 );
buf ( RI174968e8_1002 , n512 );
buf ( RI19aa9d90_2497 , n513 );
buf ( RI17526528_647 , n514 );
buf ( RI19a9cc08_2592 , n515 );
buf ( RI173b15c8_1891 , n516 );
buf ( RI173fa2b8_1536 , n517 );
buf ( RI17394db0_2030 , n518 );
buf ( RI17539830_589 , n519 );
buf ( RI17539218_590 , n520 );
buf ( RI175385e8_592 , n521 );
buf ( RI17537fd0_593 , n522 );
buf ( RI175379b8_594 , n523 );
buf ( RI17536770_597 , n524 );
buf ( RI17539e48_588 , n525 );
buf ( RI174844e0_1091 , n526 );
buf ( RI19aa2248_2551 , n527 );
buf ( RI17509a40_736 , n528 );
buf ( RI19a83438_2771 , n529 );
buf ( RI1739f1c0_1980 , n530 );
buf ( RI173e81f8_1624 , n531 );
buf ( RI1745fcd0_1269 , n532 );
buf ( RI174a1a18_948 , n533 );
buf ( RI19ab63d8_2407 , n534 );
buf ( RI173334c0_2191 , n535 );
buf ( RI173bca40_1836 , n536 );
buf ( RI174046c8_1486 , n537 );
buf ( RI174d1208_760 , n538 );
buf ( RI19a876c8_2742 , n539 );
buf ( RI174709e0_1187 , n540 );
buf ( RI19a9ca28_2593 , n541 );
buf ( RI174b9eb0_832 , n542 );
buf ( RI19acbc60_2241 , n543 );
buf ( RI1738ba08_2075 , n544 );
buf ( RI173d46f8_1720 , n545 );
buf ( RI1744c1d0_1365 , n546 );
buf ( RI1748df18_1044 , n547 );
buf ( RI19ab0870_2450 , n548 );
buf ( RI175191c0_688 , n549 );
buf ( RI19ac1d78_2315 , n550 );
buf ( RI173a8f40_1932 , n551 );
buf ( RI173f1c30_1577 , n552 );
buf ( RI174b75e8_842 , n553 );
buf ( RI173ad0e0_1912 , n554 );
buf ( RI17483b08_1094 , n555 );
buf ( RI19aa1d20_2554 , n556 );
buf ( RI17508ac8_739 , n557 );
buf ( RI19a82d30_2774 , n558 );
buf ( RI1739e7e8_1983 , n559 );
buf ( RI173e7820_1627 , n560 );
buf ( RI1745f2f8_1272 , n561 );
buf ( RI174a1040_951 , n562 );
buf ( RI19ab5d48_2410 , n563 );
buf ( RI17332ae8_2194 , n564 );
buf ( RI173bc068_1839 , n565 );
buf ( RI17404d58_1484 , n566 );
buf ( RI173fda80_1519 , n567 );
buf ( RI174a1388_950 , n568 );
buf ( RI19ab5f28_2409 , n569 );
buf ( RI174672f0_1233 , n570 );
buf ( RI19a8e8b0_2693 , n571 );
buf ( RI174affc8_878 , n572 );
buf ( RI19abf4b0_2338 , n573 );
buf ( RI17341728_2122 , n574 );
buf ( RI173caca8_1767 , n575 );
buf ( RI17413ce0_1411 , n576 );
buf ( RI174b1d50_869 , n577 );
buf ( RI19abe6a0_2346 , n578 );
buf ( RI174a3458_940 , n579 );
buf ( RI19ab4dd0_2417 , n580 );
buf ( RI17334f00_2183 , n581 );
buf ( RI173be480_1828 , n582 );
buf ( RI17407170_1473 , n583 );
buf ( RI174146b8_1408 , n584 );
buf ( RI17478000_1151 , n585 );
buf ( RI19a97820_2629 , n586 );
buf ( RI174c5850_796 , n587 );
buf ( RI19ac7700_2274 , n588 );
buf ( RI17392ce0_2040 , n589 );
buf ( RI173db9d0_1685 , n590 );
buf ( RI174534a8_1330 , n591 );
buf ( RI1738ca70_2070 , n592 );
buf ( RI17463150_1253 , n593 );
buf ( RI19a90cc8_2677 , n594 );
buf ( RI174abe28_898 , n595 );
buf ( RI19ac1148_2322 , n596 );
buf ( RI1733d588_2142 , n597 );
buf ( RI173c6b08_1787 , n598 );
buf ( RI1740f7f8_1432 , n599 );
buf ( RI1748be48_1054 , n600 );
buf ( RI19a9e030_2584 , n601 );
buf ( RI1747d898_1124 , n602 );
buf ( RI19a93d88_2655 , n603 );
buf ( RI174ce388_769 , n604 );
buf ( RI19ac40a0_2299 , n605 );
buf ( RI17398578_2013 , n606 );
buf ( RI173e1268_1658 , n607 );
buf ( RI17459088_1302 , n608 );
buf ( RI1749add0_981 , n609 );
buf ( RI19aa7c48_2511 , n610 );
buf ( RI1752d170_626 , n611 );
buf ( RI19a88e38_2732 , n612 );
buf ( RI173b5ab0_1870 , n613 );
buf ( RI173feae8_1514 , n614 );
buf ( RI173c0208_1819 , n615 );
buf ( RI1752a308_635 , n616 );
buf ( RI19a95048_2647 , n617 );
buf ( RI1748a750_1061 , n618 );
buf ( RI19a9f548_2574 , n619 );
buf ( RI17513a18_705 , n620 );
buf ( RI19ace168_2224 , n621 );
buf ( RI173a5778_1949 , n622 );
buf ( RI173ee468_1594 , n623 );
buf ( RI17493120_1019 , n624 );
buf ( RI173bee58_1825 , n625 );
buf ( RI17495880_1007 , n626 );
buf ( RI19aab938_2485 , n627 );
buf ( RI17524b60_652 , n628 );
buf ( RI19aadb70_2470 , n629 );
buf ( RI173b0560_1896 , n630 );
buf ( RI173f9250_1541 , n631 );
buf ( RI17389938_2085 , n632 );
buf ( RI17469d98_1220 , n633 );
buf ( RI19a8dfc8_2697 , n634 );
buf ( RI174b2a70_865 , n635 );
buf ( RI19abeda8_2342 , n636 );
buf ( RI173441d0_2109 , n637 );
buf ( RI173cd750_1754 , n638 );
buf ( RI17445588_1398 , n639 );
buf ( RI173a3018_1961 , n640 );
buf ( RI174796f8_1144 , n641 );
buf ( RI19a96290_2639 , n642 );
buf ( RI173943d8_2033 , n643 );
buf ( RI173dd0c8_1678 , n644 );
buf ( RI17454ba0_1323 , n645 );
buf ( RI17496c30_1001 , n646 );
buf ( RI19aa9f70_2496 , n647 );
buf ( RI17526a50_646 , n648 );
buf ( RI19a9e6c0_2581 , n649 );
buf ( RI173b1910_1890 , n650 );
buf ( RI173fa600_1535 , n651 );
buf ( RI173971c8_2019 , n652 );
buf ( RI173f53f8_1560 , n653 );
buf ( RI174a0320_955 , n654 );
buf ( RI19ab7da0_2396 , n655 );
buf ( RI17535780_600 , n656 );
buf ( RI173bb348_1843 , n657 );
buf ( RI17404038_1488 , n658 );
buf ( RI173f6af0_1553 , n659 );
buf ( RI173e4a30_1641 , n660 );
buf ( RI1748ffe8_1034 , n661 );
buf ( RI19aaf628_2458 , n662 );
buf ( RI1751c028_679 , n663 );
buf ( RI19a23150_2796 , n664 );
buf ( RI173aacc8_1923 , n665 );
buf ( RI173f39b8_1568 , n666 );
buf ( RI17502420_753 , n667 );
buf ( RI17464848_1246 , n668 );
buf ( RI19a919e8_2671 , n669 );
buf ( RI174ad520_891 , n670 );
buf ( RI19ac1b98_2316 , n671 );
buf ( RI1733ec80_2135 , n672 );
buf ( RI173c8200_1780 , n673 );
buf ( RI17410ef0_1425 , n674 );
buf ( RI1733c1d8_2148 , n675 );
buf ( RI1749be38_976 , n676 );
buf ( RI19ab9c18_2382 , n677 );
buf ( RI1752eb38_621 , n678 );
buf ( RI173b6b18_1865 , n679 );
buf ( RI173ffb50_1509 , n680 );
buf ( RI173cb680_1764 , n681 );
buf ( RI17470698_1188 , n682 );
buf ( RI19a9c848_2594 , n683 );
buf ( RI174b9988_833 , n684 );
buf ( RI19acba08_2242 , n685 );
buf ( RI1738b6c0_2076 , n686 );
buf ( RI173d43b0_1721 , n687 );
buf ( RI1744be88_1366 , n688 );
buf ( RI173dd758_1676 , n689 );
buf ( RI1746b490_1213 , n690 );
buf ( RI19a8c6f0_2708 , n691 );
buf ( RI174b4168_858 , n692 );
buf ( RI19abd9f8_2353 , n693 );
buf ( RI173458c8_2102 , n694 );
buf ( RI173cf190_1746 , n695 );
buf ( RI17446c80_1391 , n696 );
buf ( RI174889c8_1070 , n697 );
buf ( RI19aa0790_2565 , n698 );
buf ( RI17510688_715 , n699 );
buf ( RI19acf428_2216 , n700 );
buf ( RI173a39f0_1958 , n701 );
buf ( RI173ec6e0_1603 , n702 );
buf ( RI17480d18_1108 , n703 );
buf ( RI174a2dc8_942 , n704 );
buf ( RI173ad428_1911 , n705 );
buf ( RI17483e50_1093 , n706 );
buf ( RI19aa1f00_2553 , n707 );
buf ( RI1739eb30_1982 , n708 );
buf ( RI173e7b68_1626 , n709 );
buf ( RI1745f640_1271 , n710 );
buf ( RI17332e30_2193 , n711 );
buf ( RI173bc3b0_1838 , n712 );
buf ( RI174050a0_1483 , n713 );
buf ( RI173ffe98_1508 , n714 );
buf ( RI17400f00_1503 , n715 );
buf ( RI1748ec38_1040 , n716 );
buf ( RI19aae7a0_2465 , n717 );
buf ( RI1751a138_685 , n718 );
buf ( RI19a23330_2795 , n719 );
buf ( RI173a9918_1929 , n720 );
buf ( RI173f2608_1574 , n721 );
buf ( RI174be1b8_819 , n722 );
buf ( RI174118c8_1422 , n723 );
buf ( RI1749f600_959 , n724 );
buf ( RI19ab73c8_2400 , n725 );
buf ( RI175342e0_604 , n726 );
buf ( RI173ba628_1847 , n727 );
buf ( RI17403318_1492 , n728 );
buf ( RI173eda90_1597 , n729 );
buf ( RI17473e60_1171 , n730 );
buf ( RI19a99f80_2612 , n731 );
buf ( RI174bf658_815 , n732 );
buf ( RI19ac96e0_2259 , n733 );
buf ( RI1738ee88_2059 , n734 );
buf ( RI173d7b78_1704 , n735 );
buf ( RI1744f650_1349 , n736 );
buf ( RI1738cdb8_2069 , n737 );
buf ( RI174637e0_1251 , n738 );
buf ( RI19a90f20_2676 , n739 );
buf ( RI174ac4b8_896 , n740 );
buf ( RI19ac12b0_2321 , n741 );
buf ( RI1733dc18_2140 , n742 );
buf ( RI173c7198_1785 , n743 );
buf ( RI1740fe88_1430 , n744 );
buf ( RI173e5750_1637 , n745 );
buf ( RI17472df8_1176 , n746 );
buf ( RI19a9bd80_2599 , n747 );
buf ( RI174bd768_821 , n748 );
buf ( RI19acb120_2247 , n749 );
buf ( RI1738de20_2064 , n750 );
buf ( RI173d6b10_1709 , n751 );
buf ( RI1744e5e8_1354 , n752 );
buf ( RI17490678_1032 , n753 );
buf ( RI19aad300_2474 , n754 );
buf ( RI1751ca78_677 , n755 );
buf ( RI19abcfa8_2359 , n756 );
buf ( RI173ab358_1921 , n757 );
buf ( RI173f4048_1566 , n758 );
buf ( RI1750b408_731 , n759 );
buf ( RI173b2630_1886 , n760 );
buf ( RI1748ade0_1059 , n761 );
buf ( RI19a9d400_2589 , n762 );
buf ( RI17514468_703 , n763 );
buf ( RI19acc200_2238 , n764 );
buf ( RI173a5e08_1947 , n765 );
buf ( RI173eeaf8_1592 , n766 );
buf ( RI17497950_997 , n767 );
buf ( RI174a8660_915 , n768 );
buf ( RI19ab0ff0_2446 , n769 );
buf ( RI17339dc0_2159 , n770 );
buf ( RI173c3340_1804 , n771 );
buf ( RI1740c030_1449 , n772 );
buf ( RI173b6e60_1864 , n773 );
buf ( RI173bf1a0_1824 , n774 );
buf ( RI174a4808_934 , n775 );
buf ( RI19ab34f8_2429 , n776 );
buf ( RI173362b0_2177 , n777 );
buf ( RI173bf830_1822 , n778 );
buf ( RI17408520_1467 , n779 );
buf ( RI17450d48_1342 , n780 );
buf ( RI1744b7f8_1368 , n781 );
buf ( RI17461a58_1260 , n782 );
buf ( RI19a922d0_2667 , n783 );
buf ( RI174aa730_905 , n784 );
buf ( RI19ac25e8_2311 , n785 );
buf ( RI173c5410_1794 , n786 );
buf ( RI1740e100_1439 , n787 );
buf ( RI1747ef90_1117 , n788 );
buf ( RI19aa5fb0_2523 , n789 );
buf ( RI174d07a0_762 , n790 );
buf ( RI19a87218_2744 , n791 );
buf ( RI17399c70_2006 , n792 );
buf ( RI173e2960_1651 , n793 );
buf ( RI1745a780_1295 , n794 );
buf ( RI173acd98_1913 , n795 );
buf ( RI174837c0_1095 , n796 );
buf ( RI19aa3ee0_2538 , n797 );
buf ( RI175085a0_740 , n798 );
buf ( RI19a852b0_2758 , n799 );
buf ( RI1739e4a0_1984 , n800 );
buf ( RI173e74d8_1628 , n801 );
buf ( RI1745efb0_1273 , n802 );
buf ( RI174a0cf8_952 , n803 );
buf ( RI19ab5a00_2411 , n804 );
buf ( RI173327a0_2195 , n805 );
buf ( RI173bbd20_1840 , n806 );
buf ( RI17404a10_1485 , n807 );
buf ( RI173fb668_1530 , n808 );
buf ( RI17400870_1505 , n809 );
buf ( RI17462ac0_1255 , n810 );
buf ( RI19a92e10_2662 , n811 );
buf ( RI174ab798_900 , n812 );
buf ( RI19ac30b0_2306 , n813 );
buf ( RI1733cef8_2144 , n814 );
buf ( RI173c6478_1789 , n815 );
buf ( RI1740f168_1434 , n816 );
buf ( RI17411238_1424 , n817 );
buf ( RI1749ef70_961 , n818 );
buf ( RI19ab7008_2402 , n819 );
buf ( RI17533890_606 , n820 );
buf ( RI173b9f98_1849 , n821 );
buf ( RI17402c88_1494 , n822 );
buf ( RI173e9260_1619 , n823 );
buf ( RI1746aab8_1216 , n824 );
buf ( RI19a8bfe8_2711 , n825 );
buf ( RI174b3790_861 , n826 );
buf ( RI19abd4d0_2356 , n827 );
buf ( RI17344ef0_2105 , n828 );
buf ( RI173ce7b8_1749 , n829 );
buf ( RI174462a8_1394 , n830 );
buf ( RI17487ff0_1073 , n831 );
buf ( RI19aa0100_2568 , n832 );
buf ( RI1750f710_718 , n833 );
buf ( RI19aced20_2219 , n834 );
buf ( RI173ebd08_1606 , n835 );
buf ( RI1747a0d0_1141 , n836 );
buf ( RI17479068_1146 , n837 );
buf ( RI19a95de0_2641 , n838 );
buf ( RI174c7218_791 , n839 );
buf ( RI19ac5bd0_2286 , n840 );
buf ( RI17393d48_2035 , n841 );
buf ( RI173dca38_1680 , n842 );
buf ( RI17454510_1325 , n843 );
buf ( RI174965a0_1003 , n844 );
buf ( RI19aa9bb0_2498 , n845 );
buf ( RI17526000_648 , n846 );
buf ( RI19a9b420_2603 , n847 );
buf ( RI173b1280_1892 , n848 );
buf ( RI173f9f70_1537 , n849 );
buf ( RI17392998_2041 , n850 );
buf ( RI17482758_1100 , n851 );
buf ( RI19aa3580_2542 , n852 );
buf ( RI17506bd8_745 , n853 );
buf ( RI19a84950_2762 , n854 );
buf ( RI1739d438_1989 , n855 );
buf ( RI173e6470_1633 , n856 );
buf ( RI1745df48_1278 , n857 );
buf ( RI1749fc90_957 , n858 );
buf ( RI19ab7878_2398 , n859 );
buf ( RI17534d30_602 , n860 );
buf ( RI173bacb8_1845 , n861 );
buf ( RI174039a8_1490 , n862 );
buf ( RI173f22c0_1575 , n863 );
buf ( RI174ae240_887 , n864 );
buf ( RI19ac04a0_2329 , n865 );
buf ( RI1733f9a0_2131 , n866 );
buf ( RI173c8f20_1776 , n867 );
buf ( RI17411c10_1421 , n868 );
buf ( RI1749b7a8_978 , n869 );
buf ( RI19ab98d0_2384 , n870 );
buf ( RI1752e0e8_623 , n871 );
buf ( RI173b6488_1867 , n872 );
buf ( RI173ff4c0_1511 , n873 );
buf ( RI173c6e50_1786 , n874 );
buf ( RI17470008_1190 , n875 );
buf ( RI19a9c398_2596 , n876 );
buf ( RI174b8f38_835 , n877 );
buf ( RI19acb648_2244 , n878 );
buf ( RI1738b030_2078 , n879 );
buf ( RI173d3d20_1723 , n880 );
buf ( RI174d0cc8_761 , n881 );
buf ( RI19a87470_2743 , n882 );
buf ( RI1748dbd0_1045 , n883 );
buf ( RI19ab0528_2451 , n884 );
buf ( RI17518c98_689 , n885 );
buf ( RI19ab3a20_2426 , n886 );
buf ( RI173a8bf8_1933 , n887 );
buf ( RI173f18e8_1578 , n888 );
buf ( RI174b51d0_853 , n889 );
buf ( RI174a3110_941 , n890 );
buf ( RI19ab4bf0_2418 , n891 );
buf ( RI17334bb8_2184 , n892 );
buf ( RI173be138_1829 , n893 );
buf ( RI17406e28_1474 , n894 );
buf ( RI174122a0_1419 , n895 );
buf ( RI1738c728_2071 , n896 );
buf ( RI17462e08_1254 , n897 );
buf ( RI19a90a70_2678 , n898 );
buf ( RI174abae0_899 , n899 );
buf ( RI19ac0f68_2323 , n900 );
buf ( RI1733d240_2143 , n901 );
buf ( RI173c67c0_1788 , n902 );
buf ( RI1740f4b0_1433 , n903 );
buf ( RI17480340_1111 , n904 );
buf ( RI19aa46d8_2534 , n905 );
buf ( RI175014a8_756 , n906 );
buf ( RI1739b020_2000 , n907 );
buf ( RI173e3d10_1645 , n908 );
buf ( RI1745bb30_1289 , n909 );
buf ( RI173e50c0_1639 , n910 );
buf ( RI17472768_1178 , n911 );
buf ( RI19a9b8d0_2601 , n912 );
buf ( RI174bcd18_823 , n913 );
buf ( RI19acadd8_2249 , n914 );
buf ( RI1738d790_2066 , n915 );
buf ( RI173d6480_1711 , n916 );
buf ( RI1744df58_1356 , n917 );
buf ( RI17529de0_636 , n918 );
buf ( RI19a93518_2659 , n919 );
buf ( RI1748a408_1062 , n920 );
buf ( RI19a9f368_2575 , n921 );
buf ( RI175134f0_706 , n922 );
buf ( RI19acdf10_2225 , n923 );
buf ( RI173a5430_1950 , n924 );
buf ( RI173ee120_1595 , n925 );
buf ( RI17490d08_1030 , n926 );
buf ( RI174a7c88_918 , n927 );
buf ( RI19ab2f58_2432 , n928 );
buf ( RI173393e8_2162 , n929 );
buf ( RI173c2968_1807 , n930 );
buf ( RI1740b658_1452 , n931 );
buf ( RI17332110_2197 , n932 );
buf ( RI174951f0_1009 , n933 );
buf ( RI19aab5f0_2486 , n934 );
buf ( RI17524110_654 , n935 );
buf ( RI19aac388_2481 , n936 );
buf ( RI173afed0_1898 , n937 );
buf ( RI173f8bc0_1543 , n938 );
buf ( RI17346930_2097 , n939 );
buf ( RI17469a50_1221 , n940 );
buf ( RI19a8dd70_2698 , n941 );
buf ( RI174b2728_866 , n942 );
buf ( RI19abebc8_2343 , n943 );
buf ( RI17343e88_2110 , n944 );
buf ( RI173cd408_1755 , n945 );
buf ( RI17445240_1399 , n946 );
buf ( RI174a4178_936 , n947 );
buf ( RI19ab5820_2412 , n948 );
buf ( RI17407e90_1469 , n949 );
buf ( RI1744c518_1364 , n950 );
buf ( RI17478d20_1147 , n951 );
buf ( RI19a95b88_2642 , n952 );
buf ( RI174c6cf0_792 , n953 );
buf ( RI19ac5978_2287 , n954 );
buf ( RI17393a00_2036 , n955 );
buf ( RI173dc6f0_1681 , n956 );
buf ( RI174541c8_1326 , n957 );
buf ( RI173f50b0_1561 , n958 );
buf ( RI17482aa0_1099 , n959 );
buf ( RI19aa38c8_2541 , n960 );
buf ( RI17507100_744 , n961 );
buf ( RI19a84ba8_2761 , n962 );
buf ( RI1739d780_1988 , n963 );
buf ( RI173e67b8_1632 , n964 );
buf ( RI1745e290_1277 , n965 );
buf ( RI1749ffd8_956 , n966 );
buf ( RI19ab7a58_2397 , n967 );
buf ( RI17535258_601 , n968 );
buf ( RI173bb000_1844 , n969 );
buf ( RI17403cf0_1489 , n970 );
buf ( RI173f46d8_1564 , n971 );
buf ( RI173e22d0_1653 , n972 );
buf ( RI1748fca0_1035 , n973 );
buf ( RI19aaf268_2460 , n974 );
buf ( RI1751bb00_680 , n975 );
buf ( RI19a23c18_2790 , n976 );
buf ( RI173aa980_1924 , n977 );
buf ( RI173f3670_1569 , n978 );
buf ( RI174cfd50_764 , n979 );
buf ( RI17464500_1247 , n980 );
buf ( RI19a91808_2672 , n981 );
buf ( RI174ad1d8_892 , n982 );
buf ( RI19ac1a30_2317 , n983 );
buf ( RI1733e938_2136 , n984 );
buf ( RI173c7eb8_1781 , n985 );
buf ( RI17410ba8_1426 , n986 );
buf ( RI174a09b0_953 , n987 );
buf ( RI1747d550_1125 , n988 );
buf ( RI19a93ba8_2656 , n989 );
buf ( RI174cde60_770 , n990 );
buf ( RI19ac3d58_2300 , n991 );
buf ( RI17398230_2014 , n992 );
buf ( RI173e0f20_1659 , n993 );
buf ( RI17458d40_1303 , n994 );
buf ( RI1749aa88_982 , n995 );
buf ( RI19aa7a68_2512 , n996 );
buf ( RI1752cc48_627 , n997 );
buf ( RI19a88be0_2733 , n998 );
buf ( RI173b5768_1871 , n999 );
buf ( RI173fe7a0_1515 , n1000 );
buf ( RI173bddf0_1830 , n1001 );
buf ( RI17400bb8_1504 , n1002 );
buf ( RI1748e260_1043 , n1003 );
buf ( RI19ab0a50_2449 , n1004 );
buf ( RI175196e8_687 , n1005 );
buf ( RI19ad0238_2210 , n1006 );
buf ( RI173a9288_1931 , n1007 );
buf ( RI173f1f78_1576 , n1008 );
buf ( RI174ba3d8_831 , n1009 );
buf ( RI17411580_1423 , n1010 );
buf ( RI1749f2b8_960 , n1011 );
buf ( RI19ab71e8_2401 , n1012 );
buf ( RI17533db8_605 , n1013 );
buf ( RI173ba2e0_1848 , n1014 );
buf ( RI17402fd0_1493 , n1015 );
buf ( RI173eb678_1608 , n1016 );
buf ( RI17473b18_1172 , n1017 );
buf ( RI19a99d28_2613 , n1018 );
buf ( RI174bf130_816 , n1019 );
buf ( RI19ac9500_2260 , n1020 );
buf ( RI1738eb40_2060 , n1021 );
buf ( RI173d7830_1705 , n1022 );
buf ( RI1744f308_1350 , n1023 );
buf ( RI173e5408_1638 , n1024 );
buf ( RI17472ab0_1177 , n1025 );
buf ( RI19a9bb28_2600 , n1026 );
buf ( RI174bd240_822 , n1027 );
buf ( RI19acaf40_2248 , n1028 );
buf ( RI1738dad8_2065 , n1029 );
buf ( RI173d67c8_1710 , n1030 );
buf ( RI1744e2a0_1355 , n1031 );
buf ( RI17490330_1033 , n1032 );
buf ( RI19aaf790_2457 , n1033 );
buf ( RI1751c550_678 , n1034 );
buf ( RI19a83b40_2768 , n1035 );
buf ( RI173ab010_1922 , n1036 );
buf ( RI173f3d00_1567 , n1037 );
buf ( RI17507b50_742 , n1038 );
buf ( RI173b0218_1897 , n1039 );
buf ( RI1748aa98_1060 , n1040 );
buf ( RI19a9f728_2573 , n1041 );
buf ( RI17513f40_704 , n1042 );
buf ( RI19ace3c0_2223 , n1043 );
buf ( RI173a5ac0_1948 , n1044 );
buf ( RI173ee7b0_1593 , n1045 );
buf ( RI17495538_1008 , n1046 );
buf ( RI174a44c0_935 , n1047 );
buf ( RI19ab3318_2430 , n1048 );
buf ( RI173bf4e8_1823 , n1049 );
buf ( RI174081d8_1468 , n1050 );
buf ( RI1744e930_1353 , n1051 );
buf ( RI1744b4b0_1369 , n1052 );
buf ( RI1733f310_2133 , n1053 );
buf ( RI1746f2e8_1194 , n1054 );
buf ( RI19a8a080_2724 , n1055 );
buf ( RI174b7fc0_839 , n1056 );
buf ( RI19abbc70_2369 , n1057 );
buf ( RI1738a310_2082 , n1058 );
buf ( RI173d3000_1727 , n1059 );
buf ( RI1744aad8_1372 , n1060 );
buf ( RI1748c820_1051 , n1061 );
buf ( RI19a9e468_2582 , n1062 );
buf ( RI17516da8_695 , n1063 );
buf ( RI19acd100_2231 , n1064 );
buf ( RI173f0538_1584 , n1065 );
buf ( RI174a7940_919 , n1066 );
buf ( RI173a6e70_1942 , n1067 );
buf ( RI17486f88_1078 , n1068 );
buf ( RI19aa19d8_2555 , n1069 );
buf ( RI1750dd48_723 , n1070 );
buf ( RI19a82b50_2775 , n1071 );
buf ( RI173a1fb0_1966 , n1072 );
buf ( RI173eaca0_1611 , n1073 );
buf ( RI17470d28_1186 , n1074 );
buf ( RI17465220_1243 , n1075 );
buf ( RI19a8faf8_2685 , n1076 );
buf ( RI174a6248_926 , n1077 );
buf ( RI19ab4560_2421 , n1078 );
buf ( RI173379a8_2170 , n1079 );
buf ( RI173c0f28_1815 , n1080 );
buf ( RI17409c18_1460 , n1081 );
buf ( RI1745e920_1275 , n1082 );
buf ( RI173358d8_2180 , n1083 );
buf ( RI17474838_1168 , n1084 );
buf ( RI19a9a610_2609 , n1085 );
buf ( RI174c05d0_812 , n1086 );
buf ( RI19ac9de8_2256 , n1087 );
buf ( RI1738f860_2056 , n1088 );
buf ( RI173d8550_1701 , n1089 );
buf ( RI17450028_1346 , n1090 );
buf ( RI17492748_1022 , n1091 );
buf ( RI19aac040_2482 , n1092 );
buf ( RI1751fe08_667 , n1093 );
buf ( RI19ab2508_2437 , n1094 );
buf ( RI173f6118_1556 , n1095 );
buf ( RI1752b7a8_631 , n1096 );
buf ( RI174a5870_929 , n1097 );
buf ( RI19ab3de0_2424 , n1098 );
buf ( RI17336fd0_2173 , n1099 );
buf ( RI173c0550_1818 , n1100 );
buf ( RI17409240_1463 , n1101 );
buf ( RI17457cd8_1308 , n1102 );
buf ( RI174a5bb8_928 , n1103 );
buf ( RI19ab4038_2423 , n1104 );
buf ( RI17496f78_1000 , n1105 );
buf ( RI19aaa150_2495 , n1106 );
buf ( RI17526f78_645 , n1107 );
buf ( RI19a9fcc8_2570 , n1108 );
buf ( RI173fa948_1534 , n1109 );
buf ( RI173995e0_2008 , n1110 );
buf ( RI1746b7d8_1212 , n1111 );
buf ( RI19a8c948_2707 , n1112 );
buf ( RI174b44b0_857 , n1113 );
buf ( RI19abdbd8_2352 , n1114 );
buf ( RI17345c10_2101 , n1115 );
buf ( RI173cf4d8_1745 , n1116 );
buf ( RI17446fc8_1390 , n1117 );
buf ( RI174b6238_848 , n1118 );
buf ( RI19abcbe8_2361 , n1119 );
buf ( RI1747c1a0_1131 , n1120 );
buf ( RI19a95930_2643 , n1121 );
buf ( RI174cbf70_776 , n1122 );
buf ( RI19ac5720_2288 , n1123 );
buf ( RI17396e80_2020 , n1124 );
buf ( RI173dfb70_1665 , n1125 );
buf ( RI17457648_1310 , n1126 );
buf ( RI17390f58_2049 , n1127 );
buf ( RI17467638_1232 , n1128 );
buf ( RI19a8ed60_2691 , n1129 );
buf ( RI174b0310_877 , n1130 );
buf ( RI19abf870_2336 , n1131 );
buf ( RI17341a70_2121 , n1132 );
buf ( RI173caff0_1766 , n1133 );
buf ( RI17414028_1410 , n1134 );
buf ( RI17484b70_1089 , n1135 );
buf ( RI19aa27e8_2549 , n1136 );
buf ( RI1750a490_734 , n1137 );
buf ( RI19a838e8_2769 , n1138 );
buf ( RI1739f850_1978 , n1139 );
buf ( RI173e8888_1622 , n1140 );
buf ( RI17460360_1267 , n1141 );
buf ( RI17481d80_1103 , n1142 );
buf ( RI19aa3058_2545 , n1143 );
buf ( RI1751a660_684 , n1144 );
buf ( RI1749d878_968 , n1145 );
buf ( RI19ab8958_2391 , n1146 );
buf ( RI17531478_613 , n1147 );
buf ( RI173b88a0_1856 , n1148 );
buf ( RI17401590_1501 , n1149 );
buf ( RI173db688_1686 , n1150 );
buf ( RI17499a20_987 , n1151 );
buf ( RI19aa6d48_2517 , n1152 );
buf ( RI1752b280_632 , n1153 );
buf ( RI19a88028_2738 , n1154 );
buf ( RI173b4700_1876 , n1155 );
buf ( RI173fd738_1520 , n1156 );
buf ( RI173b4a48_1875 , n1157 );
buf ( RI1746e280_1199 , n1158 );
buf ( RI19a894c8_2729 , n1159 );
buf ( RI174b6f58_844 , n1160 );
buf ( RI19abaf50_2374 , n1161 );
buf ( RI173599e0_2088 , n1162 );
buf ( RI173d1f98_1732 , n1163 );
buf ( RI17449a70_1377 , n1164 );
buf ( RI174872d0_1077 , n1165 );
buf ( RI19a9f908_2572 , n1166 );
buf ( RI1750e270_722 , n1167 );
buf ( RI19ace618_2222 , n1168 );
buf ( RI173a22f8_1965 , n1169 );
buf ( RI173eafe8_1610 , n1170 );
buf ( RI17473140_1175 , n1171 );
buf ( RI173406c0_2127 , n1172 );
buf ( RI17474b80_1167 , n1173 );
buf ( RI19a9a868_2608 , n1174 );
buf ( RI174c0af8_811 , n1175 );
buf ( RI19aca040_2255 , n1176 );
buf ( RI1738fba8_2055 , n1177 );
buf ( RI173d8898_1700 , n1178 );
buf ( RI17450370_1345 , n1179 );
buf ( RI17337318_2172 , n1180 );
buf ( RI173c0898_1817 , n1181 );
buf ( RI17409588_1462 , n1182 );
buf ( RI1745a0f0_1297 , n1183 );
buf ( RI174053e8_1482 , n1184 );
buf ( RI173912a0_2048 , n1185 );
buf ( RI17484eb8_1088 , n1186 );
buf ( RI19aa2c20_2547 , n1187 );
buf ( RI1750a9b8_733 , n1188 );
buf ( RI19a83d20_2767 , n1189 );
buf ( RI1739fb98_1977 , n1190 );
buf ( RI173e8bd0_1621 , n1191 );
buf ( RI174606a8_1266 , n1192 );
buf ( RI173e9c38_1616 , n1193 );
buf ( RI174772e0_1155 , n1194 );
buf ( RI19a97460_2631 , n1195 );
buf ( RI174c48d8_799 , n1196 );
buf ( RI19ac7250_2276 , n1197 );
buf ( RI17392308_2043 , n1198 );
buf ( RI173daff8_1688 , n1199 );
buf ( RI17452ad0_1333 , n1200 );
buf ( RI17494b60_1011 , n1201 );
buf ( RI19aab0c8_2488 , n1202 );
buf ( RI175236c0_656 , n1203 );
buf ( RI19aa8f80_2503 , n1204 );
buf ( RI173af840_1900 , n1205 );
buf ( RI173f8530_1545 , n1206 );
buf ( RI17342100_2119 , n1207 );
buf ( RI173c3688_1803 , n1208 );
buf ( RI1749a0b0_985 , n1209 );
buf ( RI19aa7090_2516 , n1210 );
buf ( RI1752bcd0_630 , n1211 );
buf ( RI19a88208_2737 , n1212 );
buf ( RI173b4d90_1874 , n1213 );
buf ( RI173fddc8_1518 , n1214 );
buf ( RI173b71a8_1863 , n1215 );
buf ( RI1746e5c8_1198 , n1216 );
buf ( RI19a89720_2728 , n1217 );
buf ( RI174b72a0_843 , n1218 );
buf ( RI19abb298_2373 , n1219 );
buf ( RI173892a8_2087 , n1220 );
buf ( RI173d22e0_1731 , n1221 );
buf ( RI17449db8_1376 , n1222 );
buf ( RI174a9038_912 , n1223 );
buf ( RI19ab16f8_2443 , n1224 );
buf ( RI1733a798_2156 , n1225 );
buf ( RI173c3d18_1801 , n1226 );
buf ( RI1740ca08_1446 , n1227 );
buf ( RI173fb320_1531 , n1228 );
buf ( RI173413e0_2123 , n1229 );
buf ( RI17475be8_1162 , n1230 );
buf ( RI19a98ae0_2621 , n1231 );
buf ( RI174c24c0_806 , n1232 );
buf ( RI19ac8510_2267 , n1233 );
buf ( RI17390c10_2050 , n1234 );
buf ( RI173d9900_1695 , n1235 );
buf ( RI174513d8_1340 , n1236 );
buf ( RI174620e8_1258 , n1237 );
buf ( RI19a92708_2665 , n1238 );
buf ( RI174aadc0_903 , n1239 );
buf ( RI19ac2a98_2309 , n1240 );
buf ( RI1733c520_2147 , n1241 );
buf ( RI173c5aa0_1792 , n1242 );
buf ( RI1740e790_1437 , n1243 );
buf ( RI1747f620_1115 , n1244 );
buf ( RI19aa62f8_2521 , n1245 );
buf ( RI1739a300_2004 , n1246 );
buf ( RI173e2ff0_1649 , n1247 );
buf ( RI1745ae10_1293 , n1248 );
buf ( RI17491a28_1026 , n1249 );
buf ( RI19aadfa8_2468 , n1250 );
buf ( RI1751e968_671 , n1251 );
buf ( RI19ac36c8_2303 , n1252 );
buf ( RI173ac708_1915 , n1253 );
buf ( RI1751d4c8_675 , n1254 );
buf ( RI17461da0_1259 , n1255 );
buf ( RI19a92528_2666 , n1256 );
buf ( RI174aaa78_904 , n1257 );
buf ( RI19ac2840_2310 , n1258 );
buf ( RI173c5758_1793 , n1259 );
buf ( RI1740e448_1438 , n1260 );
buf ( RI1747f2d8_1116 , n1261 );
buf ( RI19aa6190_2522 , n1262 );
buf ( RI17399fb8_2005 , n1263 );
buf ( RI173e2ca8_1650 , n1264 );
buf ( RI1745aac8_1294 , n1265 );
buf ( RI1748d540_1047 , n1266 );
buf ( RI19ab01e0_2453 , n1267 );
buf ( RI17518248_691 , n1268 );
buf ( RI19a94df0_2648 , n1269 );
buf ( RI173a8568_1935 , n1270 );
buf ( RI173f1258_1580 , n1271 );
buf ( RI174b09a0_875 , n1272 );
buf ( RI17336940_2175 , n1273 );
buf ( RI17476278_1160 , n1274 );
buf ( RI19a98f90_2619 , n1275 );
buf ( RI174c2f10_804 , n1276 );
buf ( RI19ac89c0_2265 , n1277 );
buf ( RI173d9f90_1693 , n1278 );
buf ( RI17451a68_1338 , n1279 );
buf ( RI17493af8_1016 , n1280 );
buf ( RI19aacdd8_2476 , n1281 );
buf ( RI17521cf8_661 , n1282 );
buf ( RI19ab9df8_2381 , n1283 );
buf ( RI173ae7d8_1905 , n1284 );
buf ( RI173f74c8_1550 , n1285 );
buf ( RI17336c88_2174 , n1286 );
buf ( RI173b2978_1885 , n1287 );
buf ( RI17489058_1068 , n1288 );
buf ( RI19a9e8a0_2580 , n1289 );
buf ( RI175110d8_713 , n1290 );
buf ( RI19acd358_2230 , n1291 );
buf ( RI173a4080_1956 , n1292 );
buf ( RI173ecd70_1601 , n1293 );
buf ( RI17485548_1086 , n1294 );
buf ( RI174a68d8_924 , n1295 );
buf ( RI19ab2328_2438 , n1296 );
buf ( RI17338038_2168 , n1297 );
buf ( RI173c15b8_1813 , n1298 );
buf ( RI1740a2a8_1458 , n1299 );
buf ( RI17477970_1153 , n1300 );
buf ( RI17406108_1478 , n1301 );
buf ( RI17493e40_1015 , n1302 );
buf ( RI19aad120_2475 , n1303 );
buf ( RI17522220_660 , n1304 );
buf ( RI19abba90_2370 , n1305 );
buf ( RI173aeb20_1904 , n1306 );
buf ( RI173f7810_1549 , n1307 );
buf ( RI173390a0_2163 , n1308 );
buf ( RI174686a0_1227 , n1309 );
buf ( RI19a8cd80_2705 , n1310 );
buf ( RI174b1378_872 , n1311 );
buf ( RI19abdf98_2350 , n1312 );
buf ( RI17342ad8_2116 , n1313 );
buf ( RI173cc058_1761 , n1314 );
buf ( RI17415090_1405 , n1315 );
buf ( RI174a8cf0_913 , n1316 );
buf ( RI19ab1518_2444 , n1317 );
buf ( RI1733a450_2157 , n1318 );
buf ( RI1740c6c0_1447 , n1319 );
buf ( RI173e46e8_1642 , n1320 );
buf ( RI17391fc0_2044 , n1321 );
buf ( RI174689e8_1226 , n1322 );
buf ( RI19a8cfd8_2704 , n1323 );
buf ( RI174b16c0_871 , n1324 );
buf ( RI19abe100_2349 , n1325 );
buf ( RI17342e20_2115 , n1326 );
buf ( RI173cc3a0_1760 , n1327 );
buf ( RI174153d8_1404 , n1328 );
buf ( RI17485f20_1083 , n1329 );
buf ( RI19aa0f10_2561 , n1330 );
buf ( RI1750c380_728 , n1331 );
buf ( RI19acfd88_2212 , n1332 );
buf ( RI173a0f48_1971 , n1333 );
buf ( RI174658b0_1241 , n1334 );
buf ( RI173ea958_1612 , n1335 );
buf ( RI174816f0_1105 , n1336 );
buf ( RI19aa5218_2529 , n1337 );
buf ( RI17503398_750 , n1338 );
buf ( RI19a864f8_2750 , n1339 );
buf ( RI1739c3d0_1994 , n1340 );
buf ( RI1745cee0_1283 , n1341 );
buf ( RI1749ec28_962 , n1342 );
buf ( RI19ab9498_2386 , n1343 );
buf ( RI17533368_607 , n1344 );
buf ( RI173b9c50_1850 , n1345 );
buf ( RI17402940_1495 , n1346 );
buf ( RI173e6e48_1630 , n1347 );
buf ( RI173c43a8_1799 , n1348 );
buf ( RI1749b460_979 , n1349 );
buf ( RI19ab96f0_2385 , n1350 );
buf ( RI1752dbc0_624 , n1351 );
buf ( RI173b6140_1868 , n1352 );
buf ( RI173ff178_1512 , n1353 );
buf ( RI173c4a38_1797 , n1354 );
buf ( RI1746fcc0_1191 , n1355 );
buf ( RI19a9c1b8_2597 , n1356 );
buf ( RI174b8a10_836 , n1357 );
buf ( RI19acb4e0_2245 , n1358 );
buf ( RI1738ace8_2079 , n1359 );
buf ( RI1744a100_1375 , n1360 );
buf ( RI17466918_1236 , n1361 );
buf ( RI19a8e220_2696 , n1362 );
buf ( RI17462430_1257 , n1363 );
buf ( RI19a92960_2664 , n1364 );
buf ( RI174ab108_902 , n1365 );
buf ( RI19ac2cf0_2308 , n1366 );
buf ( RI1733c868_2146 , n1367 );
buf ( RI173c5de8_1791 , n1368 );
buf ( RI1740ead8_1436 , n1369 );
buf ( RI1747f968_1114 , n1370 );
buf ( RI19aa6640_2520 , n1371 );
buf ( RI17500530_759 , n1372 );
buf ( RI19a87920_2741 , n1373 );
buf ( RI1739a648_2003 , n1374 );
buf ( RI173e3338_1648 , n1375 );
buf ( RI1745b158_1292 , n1376 );
buf ( RI174744f0_1169 , n1377 );
buf ( RI19a9a3b8_2610 , n1378 );
buf ( RI174c00a8_813 , n1379 );
buf ( RI19ac9b90_2257 , n1380 );
buf ( RI1738f518_2057 , n1381 );
buf ( RI173d8208_1702 , n1382 );
buf ( RI17491d70_1025 , n1383 );
buf ( RI19aae110_2467 , n1384 );
buf ( RI1751ee90_670 , n1385 );
buf ( RI19ac4f28_2292 , n1386 );
buf ( RI173aca50_1914 , n1387 );
buf ( RI173f5740_1559 , n1388 );
buf ( RI17520d80_664 , n1389 );
buf ( RI174989b8_992 , n1390 );
buf ( RI19aa8bc0_2505 , n1391 );
buf ( RI1748a0c0_1063 , n1392 );
buf ( RI19a9f188_2576 , n1393 );
buf ( RI17512fc8_707 , n1394 );
buf ( RI19acdcb8_2226 , n1395 );
buf ( RI173a50e8_1951 , n1396 );
buf ( RI173eddd8_1596 , n1397 );
buf ( RI1748e8f0_1041 , n1398 );
buf ( RI174a75f8_920 , n1399 );
buf ( RI19ab2d78_2433 , n1400 );
buf ( RI17338d58_2164 , n1401 );
buf ( RI173c22d8_1809 , n1402 );
buf ( RI1740afc8_1454 , n1403 );
buf ( RI17512578_709 , n1404 );
buf ( RI17406450_1477 , n1405 );
buf ( RI17494188_1014 , n1406 );
buf ( RI19aaaa38_2491 , n1407 );
buf ( RI17522748_659 , n1408 );
buf ( RI19aa4318_2536 , n1409 );
buf ( RI173aee68_1903 , n1410 );
buf ( RI173f7b58_1548 , n1411 );
buf ( RI1733b4b8_2152 , n1412 );
buf ( RI17466c60_1235 , n1413 );
buf ( RI19a8e478_2695 , n1414 );
buf ( RI174af938_880 , n1415 );
buf ( RI19abf0f0_2340 , n1416 );
buf ( RI17341098_2124 , n1417 );
buf ( RI173ca618_1769 , n1418 );
buf ( RI17413650_1413 , n1419 );
buf ( RI17484198_1092 , n1420 );
buf ( RI19aa2068_2552 , n1421 );
buf ( RI1739ee78_1981 , n1422 );
buf ( RI173e7eb0_1625 , n1423 );
buf ( RI1745f988_1270 , n1424 );
buf ( RI174789d8_1148 , n1425 );
buf ( RI19a98018_2626 , n1426 );
buf ( RI174c67c8_793 , n1427 );
buf ( RI19ac7d90_2271 , n1428 );
buf ( RI173936b8_2037 , n1429 );
buf ( RI173dc3a8_1682 , n1430 );
buf ( RI17453e80_1327 , n1431 );
buf ( RI17503de8_748 , n1432 );
buf ( RI19a841d0_2765 , n1433 );
buf ( RI1739ca60_1992 , n1434 );
buf ( RI173e5a98_1636 , n1435 );
buf ( RI174a6f68_922 , n1436 );
buf ( RI19ab29b8_2435 , n1437 );
buf ( RI17498670_993 , n1438 );
buf ( RI19aa8878_2506 , n1439 );
buf ( RI17529390_638 , n1440 );
buf ( RI19a90368_2681 , n1441 );
buf ( RI173b3350_1882 , n1442 );
buf ( RI173fc388_1526 , n1443 );
buf ( RI173a71b8_1941 , n1444 );
buf ( RI1746ced0_1205 , n1445 );
buf ( RI19a8af08_2718 , n1446 );
buf ( RI174b5ba8_850 , n1447 );
buf ( RI19abc8a0_2363 , n1448 );
buf ( RI17347308_2094 , n1449 );
buf ( RI173d0bd0_1738 , n1450 );
buf ( RI174486c0_1383 , n1451 );
buf ( RI17466fa8_1234 , n1452 );
buf ( RI19a8e6d0_2694 , n1453 );
buf ( RI174afc80_879 , n1454 );
buf ( RI19abf2d0_2339 , n1455 );
buf ( RI173ca960_1768 , n1456 );
buf ( RI17413998_1412 , n1457 );
buf ( RI174920b8_1024 , n1458 );
buf ( RI19aae458_2466 , n1459 );
buf ( RI1751f3b8_669 , n1460 );
buf ( RI19ac6878_2281 , n1461 );
buf ( RI173f5a88_1558 , n1462 );
buf ( RI17524638_653 , n1463 );
buf ( RI1740a5f0_1457 , n1464 );
buf ( RI17498328_994 , n1465 );
buf ( RI19aa8530_2507 , n1466 );
buf ( RI17528e68_639 , n1467 );
buf ( RI19a8eb08_2692 , n1468 );
buf ( RI173b3008_1883 , n1469 );
buf ( RI173fc040_1527 , n1470 );
buf ( RI173a4da0_1952 , n1471 );
buf ( RI1746cb88_1206 , n1472 );
buf ( RI19a8acb0_2719 , n1473 );
buf ( RI174b5860_851 , n1474 );
buf ( RI19abc6c0_2364 , n1475 );
buf ( RI17346fc0_2095 , n1476 );
buf ( RI173d0888_1739 , n1477 );
buf ( RI17448378_1384 , n1478 );
buf ( RI174996d8_988 , n1479 );
buf ( RI19aa6b68_2518 , n1480 );
buf ( RI1752ad58_633 , n1481 );
buf ( RI19a87dd0_2739 , n1482 );
buf ( RI173b43b8_1877 , n1483 );
buf ( RI173fd3f0_1521 , n1484 );
buf ( RI1746df38_1200 , n1485 );
buf ( RI19a89270_2730 , n1486 );
buf ( RI174b6c10_845 , n1487 );
buf ( RI19abad70_2375 , n1488 );
buf ( RI17359698_2089 , n1489 );
buf ( RI173d1c50_1733 , n1490 );
buf ( RI17449728_1378 , n1491 );
buf ( RI1747a418_1140 , n1492 );
buf ( RI19a96bf0_2635 , n1493 );
buf ( RI174c9108_785 , n1494 );
buf ( RI19ac69e0_2280 , n1495 );
buf ( RI173950f8_2029 , n1496 );
buf ( RI173ddde8_1674 , n1497 );
buf ( RI174558c0_1319 , n1498 );
buf ( RI174665d0_1237 , n1499 );
buf ( RI19a90818_2679 , n1500 );
buf ( RI174af2a8_882 , n1501 );
buf ( RI19ac0d88_2324 , n1502 );
buf ( RI173c9f88_1771 , n1503 );
buf ( RI17412fc0_1415 , n1504 );
buf ( RI1749c4c8_974 , n1505 );
buf ( RI19aba050_2380 , n1506 );
buf ( RI1752f588_619 , n1507 );
buf ( RI173b74f0_1862 , n1508 );
buf ( RI174001e0_1507 , n1509 );
buf ( RI173cdde0_1752 , n1510 );
buf ( RI173964a8_2023 , n1511 );
buf ( RI173eee40_1591 , n1512 );
buf ( RI1733fce8_2130 , n1513 );
buf ( RI174adef8_888 , n1514 );
buf ( RI19ac0338_2330 , n1515 );
buf ( RI1733f658_2132 , n1516 );
buf ( RI173c8bd8_1777 , n1517 );
buf ( RI17454ee8_1322 , n1518 );
buf ( RI174a4e98_932 , n1519 );
buf ( RI19ab3840_2427 , n1520 );
buf ( RI173bfec0_1820 , n1521 );
buf ( RI17408bb0_1465 , n1522 );
buf ( RI17455578_1320 , n1523 );
buf ( RI17479a40_1143 , n1524 );
buf ( RI19a964e8_2638 , n1525 );
buf ( RI174c8190_788 , n1526 );
buf ( RI19ac63c8_2283 , n1527 );
buf ( RI17394720_2032 , n1528 );
buf ( RI17496258_1004 , n1529 );
buf ( RI19aa9868_2499 , n1530 );
buf ( RI17525ad8_649 , n1531 );
buf ( RI19a99ad0_2614 , n1532 );
buf ( RI173b0f38_1893 , n1533 );
buf ( RI17390580_2052 , n1534 );
buf ( RI1747fcb0_1113 , n1535 );
buf ( RI19aa6988_2519 , n1536 );
buf ( RI17500a58_758 , n1537 );
buf ( RI19a87b78_2740 , n1538 );
buf ( RI1739a990_2002 , n1539 );
buf ( RI173e3680_1647 , n1540 );
buf ( RI1745b4a0_1291 , n1541 );
buf ( RI1749d1e8_970 , n1542 );
buf ( RI19ab82c8_2394 , n1543 );
buf ( RI17530a28_615 , n1544 );
buf ( RI173b8210_1858 , n1545 );
buf ( RI173d6e58_1708 , n1546 );
buf ( RI1744a790_1373 , n1547 );
buf ( RI17511600_712 , n1548 );
buf ( RI19acd5b0_2229 , n1549 );
buf ( RI1747adf0_1137 , n1550 );
buf ( RI19a946e8_2651 , n1551 );
buf ( RI174ca080_782 , n1552 );
buf ( RI19ac4910_2295 , n1553 );
buf ( RI17395ad0_2026 , n1554 );
buf ( RI173de7c0_1671 , n1555 );
buf ( RI17456298_1316 , n1556 );
buf ( RI17486268_1082 , n1557 );
buf ( RI19aa10f0_2560 , n1558 );
buf ( RI1750c8a8_727 , n1559 );
buf ( RI19acffe0_2211 , n1560 );
buf ( RI173a1290_1970 , n1561 );
buf ( RI17467cc8_1230 , n1562 );
buf ( RI174a37a0_939 , n1563 );
buf ( RI19ab5118_2416 , n1564 );
buf ( RI17335248_2182 , n1565 );
buf ( RI173be7c8_1827 , n1566 );
buf ( RI174074b8_1472 , n1567 );
buf ( RI174458d0_1397 , n1568 );
buf ( RI1749cb58_972 , n1569 );
buf ( RI19aba578_2378 , n1570 );
buf ( RI17455230_1321 , n1571 );
buf ( RI17523198_657 , n1572 );
buf ( RI19aa7540_2514 , n1573 );
buf ( RI17464b90_1245 , n1574 );
buf ( RI19a8f648_2687 , n1575 );
buf ( RI174ad868_890 , n1576 );
buf ( RI19abff78_2332 , n1577 );
buf ( RI1733efc8_2134 , n1578 );
buf ( RI173c8548_1779 , n1579 );
buf ( RI173c8890_1778 , n1580 );
buf ( RI174916e0_1027 , n1581 );
buf ( RI19aadd50_2469 , n1582 );
buf ( RI1751e440_672 , n1583 );
buf ( RI19ac1f58_2314 , n1584 );
buf ( RI173ac3c0_1916 , n1585 );
buf ( RI17519c10_686 , n1586 );
buf ( RI17515e30_698 , n1587 );
buf ( RI19accc50_2233 , n1588 );
buf ( RI173efb60_1587 , n1589 );
buf ( RI174a96c8_910 , n1590 );
buf ( RI19ab1ba8_2441 , n1591 );
buf ( RI1733ae28_2154 , n1592 );
buf ( RI1740d098_1444 , n1593 );
buf ( RI17457990_1309 , n1594 );
buf ( RI1749a740_983 , n1595 );
buf ( RI19aa7888_2513 , n1596 );
buf ( RI1752c720_628 , n1597 );
buf ( RI19a88a00_2734 , n1598 );
buf ( RI173b5420_1872 , n1599 );
buf ( RI173fe458_1516 , n1600 );
buf ( RI173bb9d8_1841 , n1601 );
buf ( RI1746efa0_1195 , n1602 );
buf ( RI19a89bd0_2726 , n1603 );
buf ( RI174b7c78_840 , n1604 );
buf ( RI19abb748_2371 , n1605 );
buf ( RI17389fc8_2083 , n1606 );
buf ( RI175279c8_643 , n1607 );
buf ( RI19aa29c8_2548 , n1608 );
buf ( RI173b22e8_1887 , n1609 );
buf ( RI173fafd8_1532 , n1610 );
buf ( RI1739de10_1986 , n1611 );
buf ( RI173a7ed8_1937 , n1612 );
buf ( RI17497c98_996 , n1613 );
buf ( RI19aa8080_2509 , n1614 );
buf ( RI17528418_641 , n1615 );
buf ( RI19a8b958_2714 , n1616 );
buf ( RI173fb9b0_1529 , n1617 );
buf ( RI173a0570_1974 , n1618 );
buf ( RI1746c1b0_1209 , n1619 );
buf ( RI19a8a878_2721 , n1620 );
buf ( RI174b4e88_854 , n1621 );
buf ( RI19abc378_2366 , n1622 );
buf ( RI173465e8_2098 , n1623 );
buf ( RI173cfeb0_1742 , n1624 );
buf ( RI174479a0_1387 , n1625 );
buf ( RI174acb48_894 , n1626 );
buf ( RI19ac1670_2319 , n1627 );
buf ( RI17395e18_2025 , n1628 );
buf ( RI1746c840_1207 , n1629 );
buf ( RI19a8aad0_2720 , n1630 );
buf ( RI174b5518_852 , n1631 );
buf ( RI19abc4e0_2365 , n1632 );
buf ( RI17346c78_2096 , n1633 );
buf ( RI173d0540_1740 , n1634 );
buf ( RI17448030_1385 , n1635 );
buf ( RI17489a30_1065 , n1636 );
buf ( RI19a9efa8_2577 , n1637 );
buf ( RI17512050_710 , n1638 );
buf ( RI19acda60_2227 , n1639 );
buf ( RI173a4a58_1953 , n1640 );
buf ( RI173ed748_1598 , n1641 );
buf ( RI1748c190_1053 , n1642 );
buf ( RI174a2738_944 , n1643 );
buf ( RI19ab4740_2420 , n1644 );
buf ( RI173341e0_2187 , n1645 );
buf ( RI173bd760_1832 , n1646 );
buf ( RI1740d728_1442 , n1647 );
buf ( RI1748c4d8_1052 , n1648 );
buf ( RI19a9e288_2583 , n1649 );
buf ( RI17516880_696 , n1650 );
buf ( RI19accea8_2232 , n1651 );
buf ( RI173f01f0_1585 , n1652 );
buf ( RI174a5528_930 , n1653 );
buf ( RI17499390_989 , n1654 );
buf ( RI19aa9430_2501 , n1655 );
buf ( RI1752a830_634 , n1656 );
buf ( RI19a96998_2636 , n1657 );
buf ( RI173b4070_1878 , n1658 );
buf ( RI173fd0a8_1522 , n1659 );
buf ( RI1746dbf0_1201 , n1660 );
buf ( RI19a89018_2731 , n1661 );
buf ( RI17359350_2090 , n1662 );
buf ( RI173d1908_1734 , n1663 );
buf ( RI174493e0_1379 , n1664 );
buf ( RI17466288_1238 , n1665 );
buf ( RI19a905c0_2680 , n1666 );
buf ( RI174aef60_883 , n1667 );
buf ( RI19ac0ba8_2325 , n1668 );
buf ( RI173c9c40_1772 , n1669 );
buf ( RI17412c78_1416 , n1670 );
buf ( RI1746e910_1197 , n1671 );
buf ( RI1752ffd8_617 , n1672 );
buf ( RI173b7b80_1860 , n1673 );
buf ( RI173d2628_1730 , n1674 );
buf ( RI17497fe0_995 , n1675 );
buf ( RI19aa81e8_2508 , n1676 );
buf ( RI17528940_640 , n1677 );
buf ( RI19a8d230_2703 , n1678 );
buf ( RI173b2cc0_1884 , n1679 );
buf ( RI173fbcf8_1528 , n1680 );
buf ( RI173a2988_1963 , n1681 );
buf ( RI17485bd8_1084 , n1682 );
buf ( RI19aa0d30_2562 , n1683 );
buf ( RI1750be58_729 , n1684 );
buf ( RI19acfb30_2213 , n1685 );
buf ( RI173a0c00_1972 , n1686 );
buf ( RI173e98f0_1617 , n1687 );
buf ( RI17463498_1252 , n1688 );
buf ( RI1748d888_1046 , n1689 );
buf ( RI19ab03c0_2452 , n1690 );
buf ( RI17518770_690 , n1691 );
buf ( RI19aa40c0_2537 , n1692 );
buf ( RI173a88b0_1934 , n1693 );
buf ( RI173f15a0_1579 , n1694 );
buf ( RI174b2db8_864 , n1695 );
buf ( RI17484828_1090 , n1696 );
buf ( RI19aa24a0_2550 , n1697 );
buf ( RI17509f68_735 , n1698 );
buf ( RI19a83690_2770 , n1699 );
buf ( RI1739f508_1979 , n1700 );
buf ( RI173e8540_1623 , n1701 );
buf ( RI17460018_1268 , n1702 );
buf ( RI174a1d60_947 , n1703 );
buf ( RI19ab65b8_2406 , n1704 );
buf ( RI17333808_2190 , n1705 );
buf ( RI173bcd88_1835 , n1706 );
buf ( RI17405a78_1480 , n1707 );
buf ( RI17406ae0_1475 , n1708 );
buf ( RI1749cea0_971 , n1709 );
buf ( RI19aba8c0_2377 , n1710 );
buf ( RI17530500_616 , n1711 );
buf ( RI173b7ec8_1859 , n1712 );
buf ( RI173d4a40_1719 , n1713 );
buf ( RI17471700_1183 , n1714 );
buf ( RI19a9aac0_2607 , n1715 );
buf ( RI174bb350_828 , n1716 );
buf ( RI19aca298_2254 , n1717 );
buf ( RI173d5418_1716 , n1718 );
buf ( RI1744cef0_1361 , n1719 );
buf ( RI173a4710_1954 , n1720 );
buf ( RI1747b138_1136 , n1721 );
buf ( RI19a94940_2650 , n1722 );
buf ( RI174ca5a8_781 , n1723 );
buf ( RI19ac4b68_2294 , n1724 );
buf ( RI173deb08_1670 , n1725 );
buf ( RI174565e0_1315 , n1726 );
buf ( RI174720d8_1180 , n1727 );
buf ( RI19a9b1c8_2604 , n1728 );
buf ( RI174bc2c8_825 , n1729 );
buf ( RI19aca9a0_2251 , n1730 );
buf ( RI1738d100_2068 , n1731 );
buf ( RI173d5df0_1713 , n1732 );
buf ( RI1744d8c8_1358 , n1733 );
buf ( RI173df198_1668 , n1734 );
buf ( RI17485890_1085 , n1735 );
buf ( RI19aa0b50_2563 , n1736 );
buf ( RI1750b930_730 , n1737 );
buf ( RI19acf8d8_2214 , n1738 );
buf ( RI173a08b8_1973 , n1739 );
buf ( RI173e95a8_1618 , n1740 );
buf ( RI17461080_1263 , n1741 );
buf ( RI174a2a80_943 , n1742 );
buf ( RI19ab48a8_2419 , n1743 );
buf ( RI17334528_2186 , n1744 );
buf ( RI173bdaa8_1831 , n1745 );
buf ( RI17406798_1476 , n1746 );
buf ( RI17464ed8_1244 , n1747 );
buf ( RI19a8f8a0_2686 , n1748 );
buf ( RI174adbb0_889 , n1749 );
buf ( RI19ac0158_2331 , n1750 );
buf ( RI17482410_1101 , n1751 );
buf ( RI19aa3418_2543 , n1752 );
buf ( RI175066b0_746 , n1753 );
buf ( RI19a846f8_2763 , n1754 );
buf ( RI1739d0f0_1990 , n1755 );
buf ( RI173e6128_1634 , n1756 );
buf ( RI1745dc00_1279 , n1757 );
buf ( RI173cfb68_1743 , n1758 );
buf ( RI1744d238_1360 , n1759 );
buf ( RI17471a48_1182 , n1760 );
buf ( RI19a9ad18_2606 , n1761 );
buf ( RI174bb878_827 , n1762 );
buf ( RI19aca4f0_2253 , n1763 );
buf ( RI173d5760_1715 , n1764 );
buf ( RI174caff8_779 , n1765 );
buf ( RI19ac5108_2291 , n1766 );
buf ( RI174865b0_1081 , n1767 );
buf ( RI19aa1438_2558 , n1768 );
buf ( RI1750cdd0_726 , n1769 );
buf ( RI19a82538_2778 , n1770 );
buf ( RI173a15d8_1969 , n1771 );
buf ( RI173ea2c8_1614 , n1772 );
buf ( RI1746a0e0_1219 , n1773 );
buf ( RI174693c0_1223 , n1774 );
buf ( RI19a8d8c0_2700 , n1775 );
buf ( RI174b2098_868 , n1776 );
buf ( RI19abe808_2345 , n1777 );
buf ( RI173437f8_2112 , n1778 );
buf ( RI173ccd78_1757 , n1779 );
buf ( RI17444bb0_1401 , n1780 );
buf ( RI17479d88_1142 , n1781 );
buf ( RI19a96740_2637 , n1782 );
buf ( RI174c86b8_787 , n1783 );
buf ( RI19ac6620_2282 , n1784 );
buf ( RI17394a68_2031 , n1785 );
buf ( RI1744d580_1359 , n1786 );
buf ( RI17471070_1185 , n1787 );
buf ( RI19a9ce60_2591 , n1788 );
buf ( RI174ba900_830 , n1789 );
buf ( RI19acbe40_2240 , n1790 );
buf ( RI1738c098_2073 , n1791 );
buf ( RI173d4d88_1718 , n1792 );
buf ( RI1744c860_1363 , n1793 );
buf ( RI1753a460_587 , n1794 );
buf ( RI175373a0_595 , n1795 );
buf ( RI174a16d0_949 , n1796 );
buf ( RI19ab6090_2408 , n1797 );
buf ( RI17478348_1150 , n1798 );
buf ( RI19a97b68_2628 , n1799 );
buf ( RI174c5d78_795 , n1800 );
buf ( RI19ac7958_2273 , n1801 );
buf ( RI17393028_2039 , n1802 );
buf ( RI173dbd18_1684 , n1803 );
buf ( RI174537f0_1329 , n1804 );
buf ( RI17514990_702 , n1805 );
buf ( RI17410860_1427 , n1806 );
buf ( RI1749e250_965 , n1807 );
buf ( RI19ab8f70_2388 , n1808 );
buf ( RI175323f0_610 , n1809 );
buf ( RI173b9278_1853 , n1810 );
buf ( RI17401f68_1498 , n1811 );
buf ( RI173a1c68_1967 , n1812 );
buf ( RI173d9270_1697 , n1813 );
buf ( RI1748ef80_1039 , n1814 );
buf ( RI19aae980_2464 , n1815 );
buf ( RI173a9c60_1928 , n1816 );
buf ( RI173f2950_1573 , n1817 );
buf ( RI174c1a70_808 , n1818 );
buf ( RI17471d90_1181 , n1819 );
buf ( RI19a9af70_2605 , n1820 );
buf ( RI174bbda0_826 , n1821 );
buf ( RI19aca748_2252 , n1822 );
buf ( RI173d5aa8_1714 , n1823 );
buf ( RI1748f610_1037 , n1824 );
buf ( RI19aaeea8_2462 , n1825 );
buf ( RI173aa2f0_1926 , n1826 );
buf ( RI173f2fe0_1571 , n1827 );
buf ( RI174a72b0_921 , n1828 );
buf ( RI19ab2b98_2434 , n1829 );
buf ( RI17338a10_2165 , n1830 );
buf ( RI173c1f90_1810 , n1831 );
buf ( RI1740ac80_1455 , n1832 );
buf ( RI174bdc90_820 , n1833 );
buf ( RI17494818_1012 , n1834 );
buf ( RI19aaad80_2489 , n1835 );
buf ( RI173af4f8_1901 , n1836 );
buf ( RI173f81e8_1546 , n1837 );
buf ( RI17469078_1224 , n1838 );
buf ( RI19a8d668_2701 , n1839 );
buf ( RI173434b0_2113 , n1840 );
buf ( RI173cca30_1758 , n1841 );
buf ( RI17415a68_1402 , n1842 );
buf ( RI1748f2c8_1038 , n1843 );
buf ( RI19aaeb60_2463 , n1844 );
buf ( RI173a9fa8_1927 , n1845 );
buf ( RI173f2c98_1572 , n1846 );
buf ( RI174c5328_797 , n1847 );
buf ( RI17463b28_1250 , n1848 );
buf ( RI19a91100_2675 , n1849 );
buf ( RI174ac800_895 , n1850 );
buf ( RI19ac1490_2320 , n1851 );
buf ( RI1733df60_2139 , n1852 );
buf ( RI173c74e0_1784 , n1853 );
buf ( RI174101d0_1429 , n1854 );
buf ( RI17499d68_986 , n1855 );
buf ( RI17492400_1023 , n1856 );
buf ( RI19aabcf8_2483 , n1857 );
buf ( RI1749e8e0_963 , n1858 );
buf ( RI19ab92b8_2387 , n1859 );
buf ( RI17532e40_608 , n1860 );
buf ( RI173b9908_1851 , n1861 );
buf ( RI174025f8_1496 , n1862 );
buf ( RI173a95d0_1930 , n1863 );
buf ( RI174af5f0_881 , n1864 );
buf ( RI19abef88_2341 , n1865 );
buf ( RI17340d50_2125 , n1866 );
buf ( RI173ca2d0_1770 , n1867 );
buf ( RI17413308_1414 , n1868 );
buf ( RI17476f98_1156 , n1869 );
buf ( RI19a97208_2632 , n1870 );
buf ( RI174c43b0_800 , n1871 );
buf ( RI19ac6ff8_2277 , n1872 );
buf ( RI173dacb0_1689 , n1873 );
buf ( RI17452788_1334 , n1874 );
buf ( RI1748b470_1057 , n1875 );
buf ( RI19a9d9a0_2587 , n1876 );
buf ( RI1747cec0_1127 , n1877 );
buf ( RI19a936f8_2658 , n1878 );
buf ( RI174cd410_772 , n1879 );
buf ( RI19ac3920_2302 , n1880 );
buf ( RI17397ba0_2016 , n1881 );
buf ( RI173e0890_1661 , n1882 );
buf ( RI174586b0_1305 , n1883 );
buf ( RI1749c810_973 , n1884 );
buf ( RI19aba398_2379 , n1885 );
buf ( RI17462778_1256 , n1886 );
buf ( RI19a92bb8_2663 , n1887 );
buf ( RI174ab450_901 , n1888 );
buf ( RI19ac2f48_2307 , n1889 );
buf ( RI1733cbb0_2145 , n1890 );
buf ( RI173c6130_1790 , n1891 );
buf ( RI1740ee20_1435 , n1892 );
buf ( RI1747a760_1139 , n1893 );
buf ( RI19a96e48_2634 , n1894 );
buf ( RI174c9630_784 , n1895 );
buf ( RI19ac6bc0_2279 , n1896 );
buf ( RI17395440_2028 , n1897 );
buf ( RI173de130_1673 , n1898 );
buf ( RI17455c08_1318 , n1899 );
buf ( RI1752fab0_618 , n1900 );
buf ( RI173b7838_1861 , n1901 );
buf ( RI17400528_1506 , n1902 );
buf ( RI173d01f8_1741 , n1903 );
buf ( RI173967f0_2022 , n1904 );
buf ( RI1746d218_1204 , n1905 );
buf ( RI19a8b250_2717 , n1906 );
buf ( RI174b5ef0_849 , n1907 );
buf ( RI19abca80_2362 , n1908 );
buf ( RI17347650_2093 , n1909 );
buf ( RI173d0f18_1737 , n1910 );
buf ( RI17448a08_1382 , n1911 );
buf ( RI174896e8_1066 , n1912 );
buf ( RI19a9ed50_2578 , n1913 );
buf ( RI173bc6f8_1837 , n1914 );
buf ( RI1748d1f8_1048 , n1915 );
buf ( RI19ab0000_2454 , n1916 );
buf ( RI17517d20_692 , n1917 );
buf ( RI19a887a8_2735 , n1918 );
buf ( RI173a8220_1936 , n1919 );
buf ( RI173f0f10_1581 , n1920 );
buf ( RI174ae588_886 , n1921 );
buf ( RI1747bb10_1133 , n1922 );
buf ( RI19a954f8_2645 , n1923 );
buf ( RI174cb520_778 , n1924 );
buf ( RI19ac52e8_2290 , n1925 );
buf ( RI173df4e0_1667 , n1926 );
buf ( RI17456fb8_1312 , n1927 );
buf ( RI174c3e88_801 , n1928 );
buf ( RI19ac6e18_2278 , n1929 );
buf ( RI17487960_1075 , n1930 );
buf ( RI174713b8_1184 , n1931 );
buf ( RI19a9d1a8_2590 , n1932 );
buf ( RI174bae28_829 , n1933 );
buf ( RI19acc020_2239 , n1934 );
buf ( RI1738c3e0_2072 , n1935 );
buf ( RI173d50d0_1717 , n1936 );
buf ( RI1744cba8_1362 , n1937 );
buf ( RI17514eb8_701 , n1938 );
buf ( RI19acc5c0_2236 , n1939 );
buf ( RI17457300_1311 , n1940 );
buf ( RI1746d560_1203 , n1941 );
buf ( RI19a8b4a8_2716 , n1942 );
buf ( RI17358cc0_2092 , n1943 );
buf ( RI173d1278_1736 , n1944 );
buf ( RI17448d50_1381 , n1945 );
buf ( RI17476c50_1157 , n1946 );
buf ( RI19a97028_2633 , n1947 );
buf ( RI17391c78_2045 , n1948 );
buf ( RI173da968_1690 , n1949 );
buf ( RI17452440_1335 , n1950 );
buf ( RI17530f50_614 , n1951 );
buf ( RI175153e0_700 , n1952 );
buf ( RI19acc818_2235 , n1953 );
buf ( RI1747d208_1126 , n1954 );
buf ( RI19a93950_2657 , n1955 );
buf ( RI174cd938_771 , n1956 );
buf ( RI19ac3b00_2301 , n1957 );
buf ( RI17397ee8_2015 , n1958 );
buf ( RI173e0bd8_1660 , n1959 );
buf ( RI174589f8_1304 , n1960 );
buf ( RI174a20a8_946 , n1961 );
buf ( RI19ab6900_2405 , n1962 );
buf ( RI17333b50_2189 , n1963 );
buf ( RI173bd0d0_1834 , n1964 );
buf ( RI17405dc0_1479 , n1965 );
buf ( RI17408ef8_1464 , n1966 );
buf ( RI17476908_1158 , n1967 );
buf ( RI19a99440_2617 , n1968 );
buf ( RI174c3960_802 , n1969 );
buf ( RI19ac8e70_2263 , n1970 );
buf ( RI17391930_2046 , n1971 );
buf ( RI173da620_1691 , n1972 );
buf ( RI174520f8_1336 , n1973 );
buf ( RI174813a8_1106 , n1974 );
buf ( RI19aa4ed0_2530 , n1975 );
buf ( RI17502e70_751 , n1976 );
buf ( RI19a86318_2751 , n1977 );
buf ( RI1739c088_1995 , n1978 );
buf ( RI1745cb98_1284 , n1979 );
buf ( RI17469708_1222 , n1980 );
buf ( RI19a8db18_2699 , n1981 );
buf ( RI174b23e0_867 , n1982 );
buf ( RI19abe9e8_2344 , n1983 );
buf ( RI17343b40_2111 , n1984 );
buf ( RI173cd0c0_1756 , n1985 );
buf ( RI17486c40_1079 , n1986 );
buf ( RI19aa17f8_2556 , n1987 );
buf ( RI1750d820_724 , n1988 );
buf ( RI19a82970_2776 , n1989 );
buf ( RI17499048_990 , n1990 );
buf ( RI19aa90e8_2502 , n1991 );
buf ( RI173b3d28_1879 , n1992 );
buf ( RI173fcd60_1523 , n1993 );
buf ( RI173ade00_1908 , n1994 );
buf ( RI173a6498_1945 , n1995 );
buf ( RI173ef188_1590 , n1996 );
buf ( RI1749c180_975 , n1997 );
buf ( RI1748b7b8_1056 , n1998 );
buf ( RI19a9dbf8_2586 , n1999 );
buf ( RI173a67e0_1944 , n2000 );
buf ( RI173ef4d0_1589 , n2001 );
buf ( RI1749e598_964 , n2002 );
buf ( RI1747be58_1132 , n2003 );
buf ( RI19a95750_2644 , n2004 );
buf ( RI174cba48_777 , n2005 );
buf ( RI19ac5540_2289 , n2006 );
buf ( RI17396b38_2021 , n2007 );
buf ( RI173df828_1666 , n2008 );
buf ( RI174765c0_1159 , n2009 );
buf ( RI19a991e8_2618 , n2010 );
buf ( RI174c3438_803 , n2011 );
buf ( RI19ac8c18_2264 , n2012 );
buf ( RI173da2d8_1692 , n2013 );
buf ( RI17451db0_1337 , n2014 );
buf ( RI1748ceb0_1049 , n2015 );
buf ( RI19aafcb8_2455 , n2016 );
buf ( RI175177f8_693 , n2017 );
buf ( RI19a86de0_2746 , n2018 );
buf ( RI173f0bc8_1582 , n2019 );
buf ( RI174ac170_897 , n2020 );
buf ( RI1748b128_1058 , n2021 );
buf ( RI19a9d658_2588 , n2022 );
buf ( RI19acc3e0_2237 , n2023 );
buf ( RI173a6150_1946 , n2024 );
buf ( RI174a89a8_914 , n2025 );
buf ( RI19ab11d0_2445 , n2026 );
buf ( RI1733a108_2158 , n2027 );
buf ( RI1740c378_1448 , n2028 );
buf ( RI173cda98_1753 , n2029 );
buf ( RI174a23f0_945 , n2030 );
buf ( RI19ab6ae0_2404 , n2031 );
buf ( RI17333e98_2188 , n2032 );
buf ( RI173bd418_1833 , n2033 );
buf ( RI1740b310_1453 , n2034 );
buf ( RI17500f80_757 , n2035 );
buf ( RI19a85760_2756 , n2036 );
buf ( RI174937b0_1017 , n2037 );
buf ( RI19aacbf8_2477 , n2038 );
buf ( RI175217d0_662 , n2039 );
buf ( RI19ab8778_2392 , n2040 );
buf ( RI173ae490_1906 , n2041 );
buf ( RI173f7180_1551 , n2042 );
buf ( RI17334870_2185 , n2043 );
buf ( RI174a3e30_937 , n2044 );
buf ( RI19ab5640_2413 , n2045 );
buf ( RI17407b48_1470 , n2046 );
buf ( RI173f5dd0_1557 , n2047 );
buf ( RI173de478_1672 , n2048 );
buf ( RI1746be68_1210 , n2049 );
buf ( RI19a8a530_2722 , n2050 );
buf ( RI174b4b40_855 , n2051 );
buf ( RI19abc198_2367 , n2052 );
buf ( RI173462a0_2099 , n2053 );
buf ( RI17447658_1388 , n2054 );
buf ( RI174893a0_1067 , n2055 );
buf ( RI19a9eaf8_2579 , n2056 );
buf ( RI173a43c8_1955 , n2057 );
buf ( RI173ed0b8_1600 , n2058 );
buf ( RI17463e70_1249 , n2059 );
buf ( RI19a91358_2674 , n2060 );
buf ( RI1733e2a8_2138 , n2061 );
buf ( RI173c7828_1783 , n2062 );
buf ( RI17410518_1428 , n2063 );
buf ( RI174641b8_1248 , n2064 );
buf ( RI19a915b0_2673 , n2065 );
buf ( RI174ace90_893 , n2066 );
buf ( RI19ac1850_2318 , n2067 );
buf ( RI1733e5f0_2137 , n2068 );
buf ( RI173c7b70_1782 , n2069 );
buf ( RI17475f30_1161 , n2070 );
buf ( RI19a98d38_2620 , n2071 );
buf ( RI174c29e8_805 , n2072 );
buf ( RI19ac8768_2266 , n2073 );
buf ( RI173d9c48_1694 , n2074 );
buf ( RI17451720_1339 , n2075 );
buf ( RI1748f958_1036 , n2076 );
buf ( RI19aaf088_2461 , n2077 );
buf ( RI1751b5d8_681 , n2078 );
buf ( RI19a23a38_2791 , n2079 );
buf ( RI173aa638_1925 , n2080 );
buf ( RI173f3328_1570 , n2081 );
buf ( RI174cc498_775 , n2082 );
buf ( RI1748bb00_1055 , n2083 );
buf ( RI19a9de50_2585 , n2084 );
buf ( RI17515908_699 , n2085 );
buf ( RI19acc9f8_2234 , n2086 );
buf ( RI173a6b28_1943 , n2087 );
buf ( RI173ef818_1588 , n2088 );
buf ( RI1751f8e0_668 , n2089 );
buf ( RI19ab0c30_2448 , n2090 );
buf ( RI17527ef0_642 , n2091 );
buf ( RI17468358_1228 , n2092 );
buf ( RI19a8f3f0_2688 , n2093 );
buf ( RI174b1030_873 , n2094 );
buf ( RI19abfd98_2333 , n2095 );
buf ( RI17342790_2117 , n2096 );
buf ( RI173cbd10_1762 , n2097 );
buf ( RI17414d48_1406 , n2098 );
buf ( RI17487ca8_1074 , n2099 );
buf ( RI19a9ff20_2569 , n2100 );
buf ( RI1750f1e8_719 , n2101 );
buf ( RI19aceac8_2220 , n2102 );
buf ( RI173eb9c0_1607 , n2103 );
buf ( RI17477cb8_1152 , n2104 );
buf ( RI17333178_2192 , n2105 );
buf ( RI174022b0_1497 , n2106 );
buf ( RI17456c70_1313 , n2107 );
buf ( RI17472420_1179 , n2108 );
buf ( RI19a9b678_2602 , n2109 );
buf ( RI174bc7f0_824 , n2110 );
buf ( RI19acabf8_2250 , n2111 );
buf ( RI1738d448_2067 , n2112 );
buf ( RI173d6138_1712 , n2113 );
buf ( RI1744dc10_1357 , n2114 );
buf ( RI1745b7e8_1290 , n2115 );
buf ( RI173c1900_1812 , n2116 );
buf ( RI17481a38_1104 , n2117 );
buf ( RI19aa53f8_2528 , n2118 );
buf ( RI175038c0_749 , n2119 );
buf ( RI19a86750_2749 , n2120 );
buf ( RI1739c718_1993 , n2121 );
buf ( RI1745d228_1282 , n2122 );
buf ( RI174c9b58_783 , n2123 );
buf ( RI19ac46b8_2296 , n2124 );
buf ( RI1747b480_1135 , n2125 );
buf ( RI19a94b98_2649 , n2126 );
buf ( RI174a6c20_923 , n2127 );
buf ( RI19ab2670_2436 , n2128 );
buf ( RI17338380_2167 , n2129 );
buf ( RI1748e5a8_1042 , n2130 );
buf ( RI174caad0_780 , n2131 );
buf ( RI19ac4dc0_2293 , n2132 );
buf ( RI17396160_2024 , n2133 );
buf ( RI173dee50_1669 , n2134 );
buf ( RI17456928_1314 , n2135 );
buf ( RI1747aaa8_1138 , n2136 );
buf ( RI19a94490_2652 , n2137 );
buf ( RI17395788_2027 , n2138 );
buf ( RI17455f50_1317 , n2139 );
buf ( RI1747fff8_1112 , n2140 );
buf ( RI19aa44f8_2535 , n2141 );
buf ( RI1739acd8_2001 , n2142 );
buf ( RI173e39c8_1646 , n2143 );
buf ( RI1749d530_969 , n2144 );
buf ( RI19ab8430_2393 , n2145 );
buf ( RI173b8558_1857 , n2146 );
buf ( RI17401248_1502 , n2147 );
buf ( RI17481060_1107 , n2148 );
buf ( RI19aa4cf0_2531 , n2149 );
buf ( RI17502948_752 , n2150 );
buf ( RI19a860c0_2752 , n2151 );
buf ( RI1739bd40_1996 , n2152 );
buf ( RI173e4d78_1640 , n2153 );
buf ( RI1745c850_1285 , n2154 );
buf ( RI17511b28_711 , n2155 );
buf ( RI19acd808_2228 , n2156 );
buf ( RI173ed400_1599 , n2157 );
buf ( RI17489d78_1064 , n2158 );
buf ( RI1747b7c8_1134 , n2159 );
buf ( RI19a952a0_2646 , n2160 );
buf ( RI173386c8_2166 , n2161 );
buf ( RI173c1c48_1811 , n2162 );
buf ( RI1740a938_1456 , n2163 );
buf ( RI174a51e0_931 , n2164 );
buf ( RI17359008_2091 , n2165 );
buf ( RI175298b8_637 , n2166 );
buf ( RI19a91c40_2670 , n2167 );
buf ( RI173b3698_1881 , n2168 );
buf ( RI173fc6d0_1525 , n2169 );
buf ( RI17498d00_991 , n2170 );
buf ( RI19aa8da0_2504 , n2171 );
buf ( RI173b39e0_1880 , n2172 );
buf ( RI173fca18_1524 , n2173 );
buf ( RI173ab9e8_1919 , n2174 );
buf ( RI173d15c0_1735 , n2175 );
buf ( RI17506188_747 , n2176 );
buf ( RI19a843b0_2764 , n2177 );
buf ( RI1739cda8_1991 , n2178 );
buf ( RI173e5de0_1635 , n2179 );
buf ( RI1745d8b8_1280 , n2180 );
buf ( RI1746d8a8_1202 , n2181 );
buf ( RI19a8b700_2715 , n2182 );
buf ( RI1750d2f8_725 , n2183 );
buf ( RI19a82790_2777 , n2184 );
buf ( RI174868f8_1080 , n2185 );
buf ( RI19aa1618_2557 , n2186 );
buf ( RI173a1920_1968 , n2187 );
buf ( RI173ea610_1613 , n2188 );
buf ( RI1746c4f8_1208 , n2189 );
buf ( RI17449098_1380 , n2190 );
buf ( RI1754bad0_26 , n2191 );
buf ( RI1754a5b8_71 , n2192 );
buf ( RI1754a630_70 , n2193 );
buf ( RI1754a6a8_69 , n2194 );
buf ( RI1754a720_68 , n2195 );
buf ( RI17538c00_591 , n2196 );
buf ( RI19a25298_2780 , n2197 );
buf ( RI1754b788_33 , n2198 );
buf ( RI1754b878_31 , n2199 );
buf ( RI1754c430_6 , n2200 );
buf ( RI17536d88_596 , n2201 );
buf ( RI1754b800_32 , n2202 );
buf ( RI1754b530_38 , n2203 );
buf ( RI19a822e0_2779 , n2204 );
buf ( RI19ad0700_2208 , n2205 );
buf ( RI1754bcb0_22 , n2206 );
buf ( RI19a24ed8_2782 , n2207 );
buf ( RI19a250b8_2781 , n2208 );
buf ( RI1754be18_19 , n2209 );
buf ( RI1754b350_42 , n2210 );
buf ( RI1754c250_10 , n2211 );
buf ( RI1754b1e8_45 , n2212 );
buf ( RI19a24320_2787 , n2213 );
buf ( RI19a24578_2786 , n2214 );
buf ( RI1754b5a8_37 , n2215 );
buf ( RI19ad21b8_2198 , n2216 );
buf ( RI1754c160_12 , n2217 );
buf ( RI1754a900_64 , n2218 );
buf ( RI19a24c80_2783 , n2219 );
buf ( RI1754bf08_17 , n2220 );
buf ( RI1754ac48_57 , n2221 );
buf ( RI1754bf80_16 , n2222 );
buf ( RI1754bc38_23 , n2223 );
buf ( RI19a240c8_2788 , n2224 );
buf ( RI1754c070_14 , n2225 );
buf ( RI1754b3c8_41 , n2226 );
buf ( RI1754af18_51 , n2227 );
buf ( RI1754b080_48 , n2228 );
buf ( RI1754af90_50 , n2229 );
buf ( RI1754bda0_20 , n2230 );
buf ( RI1754aea0_52 , n2231 );
buf ( RI1754b260_44 , n2232 );
buf ( RI19ad0bb0_2206 , n2233 );
buf ( RI19a24a28_2784 , n2234 );
buf ( RI1754ae28_53 , n2235 );
buf ( RI1754a888_65 , n2236 );
buf ( RI1754bbc0_24 , n2237 );
buf ( RI19ad0e08_2205 , n2238 );
buf ( RI1754a810_66 , n2239 );
buf ( RI1754b440_40 , n2240 );
buf ( RI1754adb0_54 , n2241 );
buf ( RI1754c3b8_7 , n2242 );
buf ( RI19ad1060_2204 , n2243 );
buf ( RI1754ba58_27 , n2244 );
buf ( RI1754c340_8 , n2245 );
buf ( RI1754aa68_61 , n2246 );
buf ( RI1754ad38_55 , n2247 );
buf ( RI19ad12b8_2203 , n2248 );
buf ( RI1754be90_18 , n2249 );
buf ( RI1754c2c8_9 , n2250 );
buf ( RI1754c1d8_11 , n2251 );
buf ( RI19a247d0_2785 , n2252 );
buf ( RI1754b170_46 , n2253 );
buf ( RI1754aae0_60 , n2254 );
buf ( RI1754acc0_56 , n2255 );
buf ( RI1754a978_63 , n2256 );
buf ( RI19ad1588_2202 , n2257 );
buf ( RI1754b620_36 , n2258 );
buf ( RI1754bd28_21 , n2259 );
buf ( RI1754b9e0_28 , n2260 );
buf ( RI1754bb48_25 , n2261 );
buf ( RI1754ab58_59 , n2262 );
buf ( RI1754abd0_58 , n2263 );
buf ( RI1754b2d8_43 , n2264 );
buf ( RI1754c598_3 , n2265 );
buf ( RI19ad1858_2201 , n2266 );
buf ( RI1754b4b8_39 , n2267 );
buf ( RI1754b0f8_47 , n2268 );
buf ( RI1754c0e8_13 , n2269 );
buf ( RI1754bff8_15 , n2270 );
buf ( RI1754b698_35 , n2271 );
buf ( RI19ad1c18_2200 , n2272 );
buf ( RI1754c520_4 , n2273 );
buf ( RI1754b968_29 , n2274 );
buf ( RI19ad1ee8_2199 , n2275 );
buf ( RI1754b008_49 , n2276 );
buf ( RI1754c4a8_5 , n2277 );
buf ( RI1754b710_34 , n2278 );
buf ( RI1754a9f0_62 , n2279 );
buf ( RI1754b8f0_30 , n2280 );
buf ( RI19ad0958_2207 , n2281 );
buf ( n2282 , R_147ef_11ce6748 );
buf ( n2283 , R_5f38_10569f58 );
buf ( n2284 , R_13287_11ce6b08 );
buf ( n2285 , R_c94b_102f7608 );
buf ( n2286 , R_20a_1204ce78 );
buf ( n2287 , R_12f29_10571bb8 );
buf ( n2288 , R_13a43_13a1dec8 );
buf ( n2289 , R_1474d_1056fbd8 );
buf ( n2290 , R_14493_12657988 );
buf ( n2291 , R_11fd1_11ce17e8 );
buf ( n2292 , R_14705_1264d248 );
buf ( n2293 , R_105_f8cc2b8 );
buf ( n2294 , R_13cb9_11ce3c28 );
buf ( n2295 , R_138ee_13309fa8 );
buf ( n2296 , R_129dc_11543018 );
buf ( n2297 , R_10bcf_11ce1ba8 );
buf ( n2298 , R_13b6e_13a1e648 );
buf ( n2299 , R_14840_13a13ec8 );
buf ( n2300 , R_13482_10563838 );
buf ( n2301 , R_12d08_12650088 );
buf ( n2302 , R_10303_12b42dd8 );
buf ( n2303 , R_1437c_1056ac78 );
buf ( n2304 , R_87e9_1056cd98 );
buf ( n2305 , R_a30d_13320588 );
buf ( n2306 , R_144a2_133222e8 );
buf ( n2307 , R_1236b_13a1c8e8 );
buf ( n2308 , R_1396e_105627f8 );
buf ( n2309 , R_9ba7_10567258 );
buf ( n2310 , R_1f3_13797a68 );
buf ( n2311 , R_11c_13796528 );
buf ( n2312 , R_7a_1331e148 );
buf ( n2313 , R_117c9_1264ba88 );
buf ( n2314 , R_13b3f_1153ed38 );
buf ( n2315 , R_11abc_1264c2a8 );
buf ( n2316 , R_20d_137962a8 );
buf ( n2317 , R_207_1265a548 );
buf ( n2318 , R_14828_1207a118 );
buf ( n2319 , R_148eb_105aa7d8 );
buf ( n2320 , R_f3a4_10568bf8 );
buf ( n2321 , R_1b6_13799d68 );
buf ( n2322 , R_13429_1207f4d8 );
buf ( n2323 , R_14506_1056e878 );
buf ( n2324 , R_159_12b3d158 );
buf ( n2325 , R_108_105aaeb8 );
buf ( n2326 , R_102_13794cc8 );
buf ( n2327 , R_b1_12053638 );
buf ( n2328 , R_54_13309d28 );
buf ( n2329 , R_145d8_12b3ae58 );
buf ( n2330 , R_1278a_12083718 );
buf ( n2331 , R_13640_11cdeae8 );
buf ( n2332 , R_f706_11542578 );
buf ( n2333 , R_dc82_1153ebf8 );
buf ( n2334 , R_1491b_1265ef08 );
buf ( n2335 , R_14a05_10569738 );
buf ( n2336 , R_13fc5_102eac28 );
buf ( n2337 , R_1405a_115415d8 );
buf ( n2338 , R_136b3_126461c8 );
buf ( n2339 , R_1a0_132f9c88 );
buf ( n2340 , R_16f_1265bee8 );
buf ( n2341 , R_1480d_105a9dd8 );
buf ( n2342 , R_61_13304288 );
buf ( n2343 , R_e082_13798fa8 );
buf ( n2344 , R_10c7d_12082bd8 );
buf ( n2345 , R_14793_1379e188 );
buf ( n2346 , R_11ee1_102f4688 );
buf ( n2347 , R_128ba_12b27758 );
buf ( n2348 , R_70_120513d8 );
buf ( n2349 , R_129f0_12049bd8 );
buf ( n2350 , R_117e7_102f5588 );
buf ( n2351 , R_fee6_13309e68 );
buf ( n2352 , R_148f7_132f3ce8 );
buf ( n2353 , R_1362d_11ce39a8 );
buf ( n2354 , R_10693_126510c8 );
buf ( n2355 , R_11998_12656808 );
buf ( n2356 , R_143ec_11537df8 );
buf ( n2357 , R_138e8_1264afe8 );
buf ( n2358 , R_12650_12649b48 );
buf ( n2359 , R_137a1_105b63f8 );
buf ( n2360 , R_13afd_120772d8 );
buf ( n2361 , R_1490c_1264a7c8 );
buf ( n2362 , R_105e5_13306f88 );
buf ( n2363 , R_12e2b_132fa868 );
buf ( n2364 , R_144e7_12b38e78 );
buf ( n2365 , R_143e4_11cddf08 );
buf ( n2366 , R_1324a_1264c348 );
buf ( n2367 , R_1215a_11542ed8 );
buf ( n2368 , R_f685_11541678 );
buf ( n2369 , R_149ba_102ecb68 );
buf ( n2370 , R_135dc_12646088 );
buf ( n2371 , R_1476c_11cd7928 );
buf ( n2372 , R_146bd_11537998 );
buf ( n2373 , R_1df_12b39378 );
buf ( n2374 , R_13ee8_133069e8 );
buf ( n2375 , R_130_1265ac28 );
buf ( n2376 , R_65_12047c98 );
buf ( n2377 , R_13d75_1330d6a8 );
buf ( n2378 , R_13933_12081198 );
buf ( n2379 , R_133b5_12648388 );
buf ( n2380 , R_125a0_13311488 );
buf ( n2381 , R_8c_1379a808 );
buf ( n2382 , R_eadc_1207ead8 );
buf ( n2383 , R_134c7_126487e8 );
buf ( n2384 , R_11df5_1056e9b8 );
buf ( n2385 , R_144d5_102f8aa8 );
buf ( n2386 , R_12b2a_102eed28 );
buf ( n2387 , R_143d2_11538898 );
buf ( n2388 , R_1462c_102f8508 );
buf ( n2389 , R_13269_11543658 );
buf ( n2390 , R_f4_1331e0a8 );
buf ( n2391 , R_d7_132fde28 );
buf ( n2392 , R_238_1204ec78 );
buf ( n2393 , R_21b_1265e508 );
buf ( n2394 , R_12f3d_12b38b58 );
buf ( n2395 , R_112f1_1153c858 );
buf ( n2396 , R_f09_f8c93d8 );
buf ( n2397 , R_1487c_11cd99a8 );
buf ( n2398 , R_c08f_1207cb98 );
buf ( n2399 , R_923a_13a1ab88 );
buf ( n2400 , R_14042_102f2108 );
buf ( n2401 , R_143e8_102f3b48 );
buf ( n2402 , R_c2e7_13a19e68 );
buf ( n2403 , R_c175_12045118 );
buf ( n2404 , R_1450f_102f8b48 );
buf ( n2405 , R_12b14_12077238 );
buf ( n2406 , R_149e4_13a1c528 );
buf ( n2407 , R_12a04_11ce2968 );
buf ( n2408 , R_145ed_13a14e68 );
buf ( n2409 , R_13884_13796488 );
buf ( n2410 , R_13b0b_1330a688 );
buf ( n2411 , R_b5a4_102f4868 );
buf ( n2412 , R_14584_1056ec38 );
buf ( n2413 , R_13cee_12653148 );
buf ( n2414 , R_10bed_12080ab8 );
buf ( n2415 , R_117f0_102ef4a8 );
buf ( n2416 , R_10a2a_133048c8 );
buf ( n2417 , R_1be_137995e8 );
buf ( n2418 , R_151_12b448b8 );
buf ( n2419 , R_ef06_10563c98 );
buf ( n2420 , R_f9d4_1056b178 );
buf ( n2421 , R_e88a_13a13a68 );
buf ( n2422 , R_13c67_102f38c8 );
buf ( n2423 , R_128eb_10568dd8 );
buf ( n2424 , R_12eaf_f8c3118 );
buf ( n2425 , R_204_12039778 );
buf ( n2426 , R_14951_1265ebe8 );
buf ( n2427 , R_149c3_11ce5348 );
buf ( n2428 , R_1ad_12b28e78 );
buf ( n2429 , R_13f99_102f0da8 );
buf ( n2430 , R_162_12b25e58 );
buf ( n2431 , R_12003_11cdf628 );
buf ( n2432 , R_10b_11539478 );
buf ( n2433 , R_ff_1203c6f8 );
buf ( n2434 , R_1484f_1153ea18 );
buf ( n2435 , R_a8_12b425b8 );
buf ( n2436 , R_5d_13312068 );
buf ( n2437 , R_210_12043bd8 );
buf ( n2438 , R_13d84_102f4188 );
buf ( n2439 , R_142e1_10568658 );
buf ( n2440 , R_10f30_11cd9ae8 );
buf ( n2441 , R_1293d_12b43d78 );
buf ( n2442 , R_10b34_1056da18 );
buf ( n2443 , R_11a07_102eb4e8 );
buf ( n2444 , R_145b1_12082db8 );
buf ( n2445 , R_12c96_13a190a8 );
buf ( n2446 , R_d3b0_10565958 );
buf ( n2447 , R_13f2c_102f4b88 );
buf ( n2448 , R_fb8a_13a18608 );
buf ( n2449 , R_130d5_13319c88 );
buf ( n2450 , R_13f89_102f36e8 );
buf ( n2451 , R_146ff_13a1a4a8 );
buf ( n2452 , R_10ccb_1264f868 );
buf ( n2453 , R_124c3_1056f138 );
buf ( n2454 , R_10786_102f2568 );
buf ( n2455 , R_12a16_10568e78 );
buf ( n2456 , R_10726_102ef408 );
buf ( n2457 , R_137d3_12656da8 );
buf ( n2458 , R_13863_11cddb48 );
buf ( n2459 , R_14993_102f27e8 );
buf ( n2460 , R_bab1_1264a2c8 );
buf ( n2461 , R_1451e_10565818 );
buf ( n2462 , R_12a46_126515c8 );
buf ( n2463 , R_e7da_102f3508 );
buf ( n2464 , R_12756_13a1f0e8 );
buf ( n2465 , R_c4_13797ba8 );
buf ( n2466 , R_128da_1207ec18 );
buf ( n2467 , R_c282_12076838 );
buf ( n2468 , R_1272e_1056cbb8 );
buf ( n2469 , R_14a5f_120797b8 );
buf ( n2470 , R_14448_12663648 );
buf ( n2471 , R_c2_12048058 );
buf ( n2472 , R_1372d_11ce2aa8 );
buf ( n2473 , R_f878_1207c7d8 );
buf ( n2474 , R_13a76_13797888 );
buf ( n2475 , R_13a17_13796b68 );
buf ( n2476 , R_1cb_12044ad8 );
buf ( n2477 , R_14462_12b3f8b8 );
buf ( n2478 , R_6021_1379bd48 );
buf ( n2479 , R_144_13795128 );
buf ( n2480 , R_1383e_105671b8 );
buf ( n2481 , R_147ab_1056a6d8 );
buf ( n2482 , R_c6_1330e0a8 );
buf ( n2483 , R_249_12654368 );
buf ( n2484 , R_1305a_13796ca8 );
buf ( n2485 , R_12e4b_13307348 );
buf ( n2486 , R_14a38_137a1e28 );
buf ( n2487 , R_d1de_11cd9ea8 );
buf ( n2488 , R_138e2_11cd83c8 );
buf ( n2489 , R_13e62_1056dab8 );
buf ( n2490 , R_114a7_1331d748 );
buf ( n2491 , R_12f53_13319648 );
buf ( n2492 , R_f8a4_11543a18 );
buf ( n2493 , R_11ec3_13a157c8 );
buf ( n2494 , R_12c06_11cdac68 );
buf ( n2495 , R_12be8_12649788 );
buf ( n2496 , R_136c6_11cdc6a8 );
buf ( n2497 , R_1482e_13a1a228 );
buf ( n2498 , R_10ba7_115431f8 );
buf ( n2499 , R_89f2_11545098 );
buf ( n2500 , R_11953_1153c538 );
buf ( n2501 , R_9e64_11ce48a8 );
buf ( n2502 , R_e77d_11ce3ea8 );
buf ( n2503 , R_1091c_13a1a2c8 );
buf ( n2504 , R_114ec_12650628 );
buf ( n2505 , R_1286a_11cdcd88 );
buf ( n2506 , R_10d6d_1265db08 );
buf ( n2507 , R_1228f_1331f0e8 );
buf ( n2508 , R_1c5_126590a8 );
buf ( n2509 , R_14490_132f7d48 );
buf ( n2510 , R_1a1_1264a408 );
buf ( n2511 , R_976e_12056398 );
buf ( n2512 , R_6845_12648ec8 );
buf ( n2513 , R_16e_1379a3a8 );
buf ( n2514 , R_14a_12657528 );
buf ( n2515 , R_12718_10566fd8 );
buf ( n2516 , R_145c9_12075438 );
buf ( n2517 , R_c0_132fa5e8 );
buf ( n2518 , R_9c_12655f48 );
buf ( n2519 , R_d230_102edec8 );
buf ( n2520 , R_69_12658888 );
buf ( n2521 , R_13097_11ce5b68 );
buf ( n2522 , R_11051_1264a5e8 );
buf ( n2523 , R_145f0_11536818 );
buf ( n2524 , R_13ccd_132f9288 );
buf ( n2525 , R_e0_12661ac8 );
buf ( n2526 , R_22f_1331df68 );
buf ( n2527 , R_12a2a_11cd9f48 );
buf ( n2528 , R_10a54_11540458 );
buf ( n2529 , R_d027_13795628 );
buf ( n2530 , R_144d2_105677f8 );
buf ( n2531 , R_14638_11cd9228 );
buf ( n2532 , R_1454b_10568338 );
buf ( n2533 , R_147fe_1265bb28 );
buf ( n2534 , R_e861_12650448 );
buf ( n2535 , R_c03c_137931e8 );
buf ( n2536 , R_13574_102f97c8 );
buf ( n2537 , R_10e6d_102ec0c8 );
buf ( n2538 , R_c8_1331c348 );
buf ( n2539 , R_247_12b3bad8 );
buf ( n2540 , R_77_126636e8 );
buf ( n2541 , R_13a50_1056bb78 );
buf ( n2542 , R_129a5_11543798 );
buf ( n2543 , R_ef35_102f6d48 );
buf ( n2544 , R_1028c_137951c8 );
buf ( n2545 , R_1348b_12051838 );
buf ( n2546 , R_11f8b_11cdc428 );
buf ( n2547 , R_1452d_f8c5878 );
buf ( n2548 , R_12a3b_12650308 );
buf ( n2549 , R_13fd5_12079d58 );
buf ( n2550 , R_dd89_13302de8 );
buf ( n2551 , R_13dcc_102f7ec8 );
buf ( n2552 , R_14822_102f5768 );
buf ( n2553 , R_baf1_12084e38 );
buf ( n2554 , R_1315c_11ce75a8 );
buf ( n2555 , R_df0e_12654d68 );
buf ( n2556 , R_efea_11cdc248 );
buf ( n2557 , R_fe90_13a14a08 );
buf ( n2558 , R_1453c_102ec208 );
buf ( n2559 , R_aaa7_102edba8 );
buf ( n2560 , R_13c4e_13a1c988 );
buf ( n2561 , R_f758_13a13d88 );
buf ( n2562 , R_1485e_12b38f18 );
buf ( n2563 , R_ece9_1264c488 );
buf ( n2564 , R_14a35_12037f18 );
buf ( n2565 , R_1190c_102ecfc8 );
buf ( n2566 , R_12810_12650d08 );
buf ( n2567 , R_f016_12044df8 );
buf ( n2568 , R_1494e_13a14f08 );
buf ( n2569 , R_14344_1264eaa8 );
buf ( n2570 , R_10e_1265af48 );
buf ( n2571 , R_13f62_12075758 );
buf ( n2572 , R_fc_133201c8 );
buf ( n2573 , R_1378e_11cdd8c8 );
buf ( n2574 , R_147eb_120847f8 );
buf ( n2575 , R_13331_13308ec8 );
buf ( n2576 , R_213_12654f48 );
buf ( n2577 , R_146ae_1265dc48 );
buf ( n2578 , R_201_1153b138 );
buf ( n2579 , R_11d47_f8cc0d8 );
buf ( n2580 , R_c820_13a19328 );
buf ( n2581 , R_edbe_132fbd08 );
buf ( n2582 , R_be_132f4148 );
buf ( n2583 , R_a1_12043c78 );
buf ( n2584 , R_131b9_102f29c8 );
buf ( n2585 , R_12eb9_1153f738 );
buf ( n2586 , R_146e1_1153fb98 );
buf ( n2587 , R_1487f_13a173e8 );
buf ( n2588 , R_13fb4_11544af8 );
buf ( n2589 , R_1446b_10568798 );
buf ( n2590 , R_ef60_1264cf28 );
buf ( n2591 , R_1463b_1207bd38 );
buf ( n2592 , R_13166_1153aff8 );
buf ( n2593 , R_10a4b_10565bd8 );
buf ( n2594 , R_14599_12080c98 );
buf ( n2595 , R_10b18_12080018 );
buf ( n2596 , R_7254_12055078 );
buf ( n2597 , R_db04_1207b3d8 );
buf ( n2598 , R_149f9_10570cb8 );
buf ( n2599 , R_14a4a_1265d608 );
buf ( n2600 , R_14796_1264b808 );
buf ( n2601 , R_120d3_1379f3a8 );
buf ( n2602 , R_119cb_102f2068 );
buf ( n2603 , R_12acb_10565458 );
buf ( n2604 , R_145b4_12083358 );
buf ( n2605 , R_11ae9_12651528 );
buf ( n2606 , R_13af6_f8ce6f8 );
buf ( n2607 , R_13451_102f0128 );
buf ( n2608 , R_ef8c_1204e098 );
buf ( n2609 , R_ca_12b3e058 );
buf ( n2610 , R_245_f8c5ff8 );
buf ( n2611 , R_af_12b2a8b8 );
buf ( n2612 , R_10e57_11544eb8 );
buf ( n2613 , R_b243_f8c5698 );
buf ( n2614 , R_13633_13a13248 );
buf ( n2615 , R_11c97_10562078 );
buf ( n2616 , R_13838_102f5e48 );
buf ( n2617 , R_efb7_13a1bc68 );
buf ( n2618 , R_d4db_10566038 );
buf ( n2619 , R_10bc8_11ce66a8 );
buf ( n2620 , R_c9c0_102eee68 );
buf ( n2621 , R_13608_10563798 );
buf ( n2622 , R_8f_12b299b8 );
buf ( n2623 , R_59_133089c8 );
buf ( n2624 , R_134f1_102ebf88 );
buf ( n2625 , R_10499_1331e828 );
buf ( n2626 , R_14424_102f8f08 );
buf ( n2627 , R_1d6_133209e8 );
buf ( n2628 , R_ebe2_13a18568 );
buf ( n2629 , R_139_12b44ef8 );
buf ( n2630 , R_97_13792c48 );
buf ( n2631 , R_144ed_105660d8 );
buf ( n2632 , R_120c8_11541d58 );
buf ( n2633 , R_11736_11cde408 );
buf ( n2634 , R_149a8_13317528 );
buf ( n2635 , R_1450c_1056eff8 );
buf ( n2636 , R_147d9_120828b8 );
buf ( n2637 , R_11ea5_1264a9a8 );
buf ( n2638 , R_11425_1207c918 );
buf ( n2639 , R_d53e_1207c2d8 );
buf ( n2640 , R_14787_12b352b8 );
buf ( n2641 , R_13cf3_10571078 );
buf ( n2642 , R_13f36_1330ebe8 );
buf ( n2643 , R_d00d_102ee968 );
buf ( n2644 , R_a1e6_11cde368 );
buf ( n2645 , R_13f77_13a19648 );
buf ( n2646 , R_118_132f5f48 );
buf ( n2647 , R_13688_120832b8 );
buf ( n2648 , R_1f7_105a9978 );
buf ( n2649 , R_f630_1056b858 );
buf ( n2650 , R_136a1_1153fa58 );
buf ( n2651 , R_1b7_126577a8 );
buf ( n2652 , R_158_12b27938 );
buf ( n2653 , R_ec_1330a868 );
buf ( n2654 , R_223_f8c32f8 );
buf ( n2655 , R_133bf_11543338 );
buf ( n2656 , R_f2a8_102f47c8 );
buf ( n2657 , R_e112_12076e78 );
buf ( n2658 , R_12b72_1056c6b8 );
buf ( n2659 , R_2f00_102f3d28 );
buf ( n2660 , R_14819_1331de28 );
buf ( n2661 , R_e809_13313c48 );
buf ( n2662 , R_14358_11cd8788 );
buf ( n2663 , R_1473e_11543b58 );
buf ( n2664 , R_139c7_102ed1a8 );
buf ( n2665 , R_13d65_12036a78 );
buf ( n2666 , R_12c10_102ea548 );
buf ( n2667 , R_13870_11ce5e88 );
buf ( n2668 , R_dede_13a16448 );
buf ( n2669 , R_12c49_12b27438 );
buf ( n2670 , R_1192b_12645e08 );
buf ( n2671 , R_bd66_126533c8 );
buf ( n2672 , R_13fa2_1379f6c8 );
buf ( n2673 , R_13407_1056df18 );
buf ( n2674 , R_118b0_1204acb8 );
buf ( n2675 , R_13c3e_126496e8 );
buf ( n2676 , R_1438a_11cda268 );
buf ( n2677 , R_11e51_102fa268 );
buf ( n2678 , R_102b9_132f6588 );
buf ( n2679 , R_d9_1330dec8 );
buf ( n2680 , R_bc_13799c28 );
buf ( n2681 , R_236_13795f88 );
buf ( n2682 , R_ffee_1264d568 );
buf ( n2683 , R_10ea9_102f8788 );
buf ( n2684 , R_14852_13a154a8 );
buf ( n2685 , R_e696_11cdce28 );
buf ( n2686 , R_1ae_1203c3d8 );
buf ( n2687 , R_1457e_133027e8 );
buf ( n2688 , R_161_12656c68 );
buf ( n2689 , R_127_12b3cc58 );
buf ( n2690 , R_ea26_1265a4a8 );
buf ( n2691 , R_1e8_11539298 );
buf ( n2692 , R_139e4_102f59e8 );
buf ( n2693 , R_1477b_1204f218 );
buf ( n2694 , R_1459c_12056a78 );
buf ( n2695 , R_1336e_11545138 );
buf ( n2696 , R_108cd_102f7ce8 );
buf ( n2697 , R_13b4f_13305c28 );
buf ( n2698 , R_1a2_12b423d8 );
buf ( n2699 , R_16d_12664c28 );
buf ( n2700 , R_14656_11ce6ce8 );
buf ( n2701 , R_827e_1207e998 );
buf ( n2702 , R_11ab0_1204a358 );
buf ( n2703 , R_144ab_12b39af8 );
buf ( n2704 , R_144c3_12080338 );
buf ( n2705 , R_12794_102f5b28 );
buf ( n2706 , R_13149_102f7888 );
buf ( n2707 , R_144e4_12b28838 );
buf ( n2708 , R_13e_12660da8 );
buf ( n2709 , R_123_1330d888 );
buf ( n2710 , R_e7_137956c8 );
buf ( n2711 , R_cc_12038918 );
buf ( n2712 , R_137c7_102f79c8 );
buf ( n2713 , R_243_13796d48 );
buf ( n2714 , R_13795_13795588 );
buf ( n2715 , R_228_10570c18 );
buf ( n2716 , R_13f01_1056e2d8 );
buf ( n2717 , R_13d8e_11cd77e8 );
buf ( n2718 , R_1ec_12039ef8 );
buf ( n2719 , R_f175_13a17ca8 );
buf ( n2720 , R_1d1_126540e8 );
buf ( n2721 , R_14409_12b434b8 );
buf ( n2722 , R_138b2_102f06c8 );
buf ( n2723 , R_14653_1207e0d8 );
buf ( n2724 , R_13044_102f7a68 );
buf ( n2725 , R_13133_13a1ae08 );
buf ( n2726 , R_10b8f_1265ad68 );
buf ( n2727 , R_12e35_12b3b858 );
buf ( n2728 , R_12df0_12050bb8 );
buf ( n2729 , R_fc88_1207be78 );
buf ( n2730 , R_13804_102ef548 );
buf ( n2731 , R_13b68_137a1ba8 );
buf ( n2732 , R_134_13312b68 );
buf ( n2733 , R_14990_1331ae08 );
buf ( n2734 , R_1db_12043db8 );
buf ( n2735 , R_ccdc_102f6488 );
buf ( n2736 , R_1494b_11ce61a8 );
buf ( n2737 , R_12c39_10562ed8 );
buf ( n2738 , R_131c2_11ce4b28 );
buf ( n2739 , R_12d97_126626a8 );
buf ( n2740 , R_12d59_12b26b78 );
buf ( n2741 , R_1352d_13315188 );
buf ( n2742 , R_12c4f_13321d48 );
buf ( n2743 , R_1343e_10562d98 );
buf ( n2744 , R_1345b_102fa088 );
buf ( n2745 , R_1167d_115410d8 );
buf ( n2746 , R_14008_1264dec8 );
buf ( n2747 , R_11bc8_11544e18 );
buf ( n2748 , R_13c9a_1207e178 );
buf ( n2749 , R_148be_12b27f78 );
buf ( n2750 , R_14360_105ad078 );
buf ( n2751 , R_13aa3_12078138 );
buf ( n2752 , R_116da_13a1a7c8 );
buf ( n2753 , R_14732_102f5448 );
buf ( n2754 , R_cec6_132f3608 );
buf ( n2755 , R_133dc_13a1ea08 );
buf ( n2756 , R_14942_f8c5058 );
buf ( n2757 , R_13a0f_10563018 );
buf ( n2758 , R_bd10_f8ce978 );
buf ( n2759 , R_12da1_12647528 );
buf ( n2760 , R_12af5_12052418 );
buf ( n2761 , R_13cf9_13a1c0c8 );
buf ( n2762 , R_13658_12646628 );
buf ( n2763 , R_149bd_1204adf8 );
buf ( n2764 , R_13233_11cde908 );
buf ( n2765 , R_12585_1207a898 );
buf ( n2766 , R_118e9_10564a58 );
buf ( n2767 , R_1359a_13a18928 );
buf ( n2768 , R_12451_13a1d568 );
buf ( n2769 , R_dcbb_1265bf88 );
buf ( n2770 , R_f424_13a1b948 );
buf ( n2771 , R_1226a_11cdef48 );
buf ( n2772 , R_14641_13a12d48 );
buf ( n2773 , R_1257c_11ce4448 );
buf ( n2774 , R_e309_120806f8 );
buf ( n2775 , R_11ccc_13314be8 );
buf ( n2776 , R_146c0_13a15908 );
buf ( n2777 , R_14843_13a196e8 );
buf ( n2778 , R_11d00_1207f9d8 );
buf ( n2779 , R_14a1d_13a14c88 );
buf ( n2780 , R_13d54_11ce00c8 );
buf ( n2781 , R_135b5_132fdd88 );
buf ( n2782 , R_d40b_10569058 );
buf ( n2783 , R_145f9_102ee148 );
buf ( n2784 , R_14882_1056d838 );
buf ( n2785 , R_101a4_f8c2ad8 );
buf ( n2786 , R_13abf_13a15188 );
buf ( n2787 , R_eab3_126509e8 );
buf ( n2788 , R_8296_13322608 );
buf ( n2789 , R_6d_12036618 );
buf ( n2790 , R_50_12b3c118 );
buf ( n2791 , R_11b19_102ee508 );
buf ( n2792 , R_de1d_13a193c8 );
buf ( n2793 , R_14477_11cdcc48 );
buf ( n2794 , R_1195d_12038198 );
buf ( n2795 , R_14527_102eb6c8 );
buf ( n2796 , R_be8c_126504e8 );
buf ( n2797 , R_11e87_12b3c398 );
buf ( n2798 , R_14a02_13309aa8 );
buf ( n2799 , R_12b_1203e6d8 );
buf ( n2800 , R_f1_13799ea8 );
buf ( n2801 , R_21e_126608a8 );
buf ( n2802 , R_1e4_12b28338 );
buf ( n2803 , R_115ff_13304148 );
buf ( n2804 , R_10d8e_1264cfc8 );
buf ( n2805 , R_11500_12083c18 );
buf ( n2806 , R_c4bc_137945e8 );
buf ( n2807 , R_1465c_10568f18 );
buf ( n2808 , R_133e6_11cd9048 );
buf ( n2809 , R_7c4f_11ce4a88 );
buf ( n2810 , R_11f78_12b2c118 );
buf ( n2811 , R_1013a_132f59a8 );
buf ( n2812 , R_149e1_105b62b8 );
buf ( n2813 , R_150_1330cac8 );
buf ( n2814 , R_111_12b3e238 );
buf ( n2815 , R_f9_1204ba78 );
buf ( n2816 , R_ba_1331bc68 );
buf ( n2817 , R_4b_1264c028 );
buf ( n2818 , R_216_1204a038 );
buf ( n2819 , R_13733_f8d0098 );
buf ( n2820 , R_1fe_120539f8 );
buf ( n2821 , R_146de_12648748 );
buf ( n2822 , R_1bf_1265cd48 );
buf ( n2823 , R_74_1331da68 );
buf ( n2824 , R_f5c3_1264d108 );
buf ( n2825 , R_f1f7_120367f8 );
buf ( n2826 , R_e338_13301ac8 );
buf ( n2827 , R_1486d_1056e558 );
buf ( n2828 , R_13e2d_12047fb8 );
buf ( n2829 , R_12344_137a0de8 );
buf ( n2830 , R_14729_10570178 );
buf ( n2831 , R_13364_105717f8 );
buf ( n2832 , R_11160_1153e298 );
buf ( n2833 , R_10a01_11cde228 );
buf ( n2834 , R_13c6f_12041658 );
buf ( n2835 , R_148c4_10568978 );
buf ( n2836 , R_11c81_132f7348 );
buf ( n2837 , R_10ec5_11cdb028 );
buf ( n2838 , R_14441_12659008 );
buf ( n2839 , R_cbab_105a9a18 );
buf ( n2840 , R_1238a_126482e8 );
buf ( n2841 , R_a6_12660448 );
buf ( n2842 , R_12b36_11ce6428 );
buf ( n2843 , R_dc46_10566498 );
buf ( n2844 , R_11f_137936e8 );
buf ( n2845 , R_ce_12055fd8 );
buf ( n2846 , R_241_132fd748 );
buf ( n2847 , R_147f8_1207ccd8 );
buf ( n2848 , R_1f0_13798a08 );
buf ( n2849 , R_1467d_1056bcb8 );
buf ( n2850 , R_14668_11546178 );
buf ( n2851 , R_132cc_1153edd8 );
buf ( n2852 , R_136ba_11ce37c8 );
buf ( n2853 , R_12c23_102f1d48 );
buf ( n2854 , R_106be_1264edc8 );
buf ( n2855 , R_11bde_10564878 );
buf ( n2856 , R_11a1a_11cd9a48 );
buf ( n2857 , R_9548_11ce6ba8 );
buf ( n2858 , R_f451_11542438 );
buf ( n2859 , R_119b7_105663f8 );
buf ( n2860 , R_142e5_102f2388 );
buf ( n2861 , R_147e4_13a19dc8 );
buf ( n2862 , R_d862_12661348 );
buf ( n2863 , R_d940_13a19d28 );
buf ( n2864 , R_eb8c_13a19288 );
buf ( n2865 , R_1175e_11cda088 );
buf ( n2866 , R_146f9_11ce4768 );
buf ( n2867 , R_14551_102eae08 );
buf ( n2868 , R_14578_12b3a6d8 );
buf ( n2869 , R_1467a_13a13568 );
buf ( n2870 , R_1130e_1056bfd8 );
buf ( n2871 , R_1493f_1056d3d8 );
buf ( n2872 , R_14948_102f76a8 );
buf ( n2873 , R_10230_1153d1b8 );
buf ( n2874 , R_f4d1_13a17848 );
buf ( n2875 , R_14772_11cda8a8 );
buf ( n2876 , R_1466e_1203e138 );
buf ( n2877 , R_14999_120382d8 );
buf ( n2878 , R_9d72_102f18e8 );
buf ( n2879 , R_eeaf_10566f38 );
buf ( n2880 , R_13083_12b3ff98 );
buf ( n2881 , R_e288_11541fd8 );
buf ( n2882 , R_13969_102ea408 );
buf ( n2883 , R_13825_1264d928 );
buf ( n2884 , R_134a8_13a13c48 );
buf ( n2885 , R_fcde_115390b8 );
buf ( n2886 , R_14566_102f6988 );
buf ( n2887 , R_f5eb_11544558 );
buf ( n2888 , R_12318_102ec348 );
buf ( n2889 , R_d2c9_11cd9408 );
buf ( n2890 , R_16c_132f7ca8 );
buf ( n2891 , R_d894_1056f778 );
buf ( n2892 , R_12323_102ec8e8 );
buf ( n2893 , R_1a3_13303108 );
buf ( n2894 , R_118ba_13307ac8 );
buf ( n2895 , R_12704_10562938 );
buf ( n2896 , R_148c7_1264d888 );
buf ( n2897 , R_148bb_12661d48 );
buf ( n2898 , R_1221a_13a1d248 );
buf ( n2899 , R_135b0_12651348 );
buf ( n2900 , R_1470e_10562898 );
buf ( n2901 , R_efa_1207d1d8 );
buf ( n2902 , R_ce1e_102f95e8 );
buf ( n2903 , R_126e3_105b5c78 );
buf ( n2904 , R_14026_102ecd48 );
buf ( n2905 , R_11e36_102ed608 );
buf ( n2906 , R_11515_12039318 );
buf ( n2907 , R_108e3_1056dd38 );
buf ( n2908 , R_128f4_1207aa78 );
buf ( n2909 , R_147ae_1207ce18 );
buf ( n2910 , R_12235_12650e48 );
buf ( n2911 , R_12183_12052eb8 );
buf ( n2912 , R_14647_102f04e8 );
buf ( n2913 , R_13aef_11cdd968 );
buf ( n2914 , R_1249f_102f9368 );
buf ( n2915 , R_f34d_13a18ec8 );
buf ( n2916 , R_12c3f_f8cfd78 );
buf ( n2917 , R_13d5d_1153d4d8 );
buf ( n2918 , R_12126_102ef228 );
buf ( n2919 , R_ad_12b3b358 );
buf ( n2920 , R_92_13312d48 );
buf ( n2921 , R_113db_f8cb4f8 );
buf ( n2922 , R_10d98_f8c6318 );
buf ( n2923 , R_1481f_1264dce8 );
buf ( n2924 , R_ad98_102f3aa8 );
buf ( n2925 , R_55_132f50e8 );
buf ( n2926 , R_102d5_f8ced38 );
buf ( n2927 , R_144ae_11545ef8 );
buf ( n2928 , R_a3e0_12655308 );
buf ( n2929 , R_5dbf_13a15f48 );
buf ( n2930 , R_e2_1203f858 );
buf ( n2931 , R_22d_1379de68 );
buf ( n2932 , R_135c4_105b5bd8 );
buf ( n2933 , R_13cff_13a16308 );
buf ( n2934 , R_12692_102eb8a8 );
buf ( n2935 , R_13375_13794a48 );
buf ( n2936 , R_12f6a_10562438 );
buf ( n2937 , R_128c4_102ea5e8 );
buf ( n2938 , R_122f0_12650f88 );
buf ( n2939 , R_14855_12056f78 );
buf ( n2940 , R_14885_13795a88 );
buf ( n2941 , R_bb92_11ce0ca8 );
buf ( n2942 , R_8b04_1265cf28 );
buf ( n2943 , R_e71c_115426b8 );
buf ( n2944 , R_14a23_120545d8 );
buf ( n2945 , R_149_1330f408 );
buf ( n2946 , R_b8_13305048 );
buf ( n2947 , R_1c6_1379cce8 );
buf ( n2948 , R_e13d_102eb448 );
buf ( n2949 , R_14617_11ce2f08 );
buf ( n2950 , R_13557_11545778 );
buf ( n2951 , R_148cd_12082c78 );
buf ( n2952 , R_11768_1264ffe8 );
buf ( n2953 , R_12503_11cdd008 );
buf ( n2954 , R_1239d_1330d1a8 );
buf ( n2955 , R_1448c_105662b8 );
buf ( n2956 , R_160_f8c0d78 );
buf ( n2957 , R_143_13795e48 );
buf ( n2958 , R_1252c_102f1208 );
buf ( n2959 , R_1cc_f8cc858 );
buf ( n2960 , R_149de_11cde7c8 );
buf ( n2961 , R_1af_12b40678 );
buf ( n2962 , R_a28f_11ce5708 );
buf ( n2963 , R_f7ae_11ce57a8 );
buf ( n2964 , R_1243d_10571118 );
buf ( n2965 , R_d0df_126478e8 );
buf ( n2966 , R_1498d_1153fe18 );
buf ( n2967 , R_10350_11cda6c8 );
buf ( n2968 , R_103a6_10569878 );
buf ( n2969 , R_128b0_1056c118 );
buf ( n2970 , R_14936_10561e98 );
buf ( n2971 , R_10d1b_11cd7748 );
buf ( n2972 , R_ed92_102eea08 );
buf ( n2973 , R_145d2_11cdb208 );
buf ( n2974 , R_109f6_1153ca38 );
buf ( n2975 , R_cc46_1207b298 );
buf ( n2976 , R_11006_126501c8 );
buf ( n2977 , R_188_1265c348 );
buf ( n2978 , R_187_12b25d18 );
buf ( n2979 , R_12f_1379dbe8 );
buf ( n2980 , R_db_12663f08 );
buf ( n2981 , R_84_12652ce8 );
buf ( n2982 , R_81_12042a58 );
buf ( n2983 , R_234_12b43af8 );
buf ( n2984 , R_1e0_133037e8 );
buf ( n2985 , R_13ed7_1207ad98 );
buf ( n2986 , R_189_f8c6458 );
buf ( n2987 , R_186_126553a8 );
buf ( n2988 , R_157_132f7a28 );
buf ( n2989 , R_d0_105aa238 );
buf ( n2990 , R_23f_13307848 );
buf ( n2991 , R_11399_12b3c1b8 );
buf ( n2992 , R_1b8_11537358 );
buf ( n2993 , R_f82c_f8cdc58 );
buf ( n2994 , R_d9ca_10562bb8 );
buf ( n2995 , R_145f6_f8c3398 );
buf ( n2996 , R_1449c_11ce71e8 );
buf ( n2997 , R_13850_13a1fe08 );
buf ( n2998 , R_135e3_13306da8 );
buf ( n2999 , R_ec0b_132fa368 );
buf ( n3000 , R_147e0_13a12fc8 );
buf ( n3001 , R_13add_132ff728 );
buf ( n3002 , R_f65b_12084578 );
buf ( n3003 , R_10cb4_11cdf9e8 );
buf ( n3004 , R_18a_133173e8 );
buf ( n3005 , R_185_12042cd8 );
buf ( n3006 , R_134d0_12651028 );
buf ( n3007 , R_144f3_102f3fa8 );
buf ( n3008 , R_12dd1_f8c52d8 );
buf ( n3009 , R_135a9_10567938 );
buf ( n3010 , R_11b39_102ec988 );
buf ( n3011 , R_1386a_102ebda8 );
buf ( n3012 , R_14747_12042b98 );
buf ( n3013 , R_148d0_137a0a28 );
buf ( n3014 , R_11f4d_137986e8 );
buf ( n3015 , R_13d05_12081378 );
buf ( n3016 , R_f56e_102f2608 );
buf ( n3017 , R_62_12b26498 );
buf ( n3018 , R_10e0b_1056abd8 );
buf ( n3019 , R_ba73_1264c8e8 );
buf ( n3020 , R_14888_12653288 );
buf ( n3021 , R_fc34_1379c428 );
buf ( n3022 , R_18b_12663fa8 );
buf ( n3023 , R_184_1153acd8 );
buf ( n3024 , R_119d5_1331dc48 );
buf ( n3025 , R_122b5_13305688 );
buf ( n3026 , R_e051_12649f08 );
buf ( n3027 , R_ca0a_10567438 );
buf ( n3028 , R_10a84_115427f8 );
buf ( n3029 , R_668e_10563f18 );
buf ( n3030 , R_14539_102f7108 );
buf ( n3031 , R_c3d6_11cdb7a8 );
buf ( n3032 , R_11703_132fa728 );
buf ( n3033 , R_1472f_105708f8 );
buf ( n3034 , R_1307a_11cdc1a8 );
buf ( n3035 , R_fdae_1153d258 );
buf ( n3036 , R_13ac5_102ee3c8 );
buf ( n3037 , R_120bd_1153ff58 );
buf ( n3038 , R_13f6e_12649dc8 );
buf ( n3039 , R_1177b_1207fbb8 );
buf ( n3040 , R_f804_1379efe8 );
buf ( n3041 , R_111d5_13a17c08 );
buf ( n3042 , R_14750_13304008 );
buf ( n3043 , R_137d9_12055e98 );
buf ( n3044 , R_87_132ffa48 );
buf ( n3045 , R_7e_137949a8 );
buf ( n3046 , R_f140_1056f598 );
buf ( n3047 , R_d43f_12079678 );
buf ( n3048 , R_11900_1056f6d8 );
buf ( n3049 , R_18c_12660e48 );
buf ( n3050 , R_c969_1330f9a8 );
buf ( n3051 , R_183_126587e8 );
buf ( n3052 , R_11093_102f60c8 );
buf ( n3053 , R_f31e_120770f8 );
buf ( n3054 , R_f06_1265f728 );
buf ( n3055 , R_d5cf_102f5128 );
buf ( n3056 , R_10874_12037838 );
buf ( n3057 , R_11324_13a1f228 );
buf ( n3058 , R_13621_120823b8 );
buf ( n3059 , R_120dd_f8cdcf8 );
buf ( n3060 , R_148d3_12049a98 );
buf ( n3061 , R_13e42_12648888 );
buf ( n3062 , R_144c0_12078db8 );
buf ( n3063 , R_12978_13316d08 );
buf ( n3064 , R_11b5e_13a1b088 );
buf ( n3065 , R_13025_13a1ef08 );
buf ( n3066 , R_e615_12084bb8 );
buf ( n3067 , R_149b7_102ea4a8 );
buf ( n3068 , R_1497e_1207ef38 );
buf ( n3069 , R_11fee_12b2a3b8 );
buf ( n3070 , R_11b_12b43198 );
buf ( n3071 , R_5e_126647c8 );
buf ( n3072 , R_1f4_1265d108 );
buf ( n3073 , R_1445f_13792888 );
buf ( n3074 , R_13981_13798aa8 );
buf ( n3075 , R_14569_11cdbfc8 );
buf ( n3076 , R_114_12b3e4b8 );
buf ( n3077 , R_f6_12664188 );
buf ( n3078 , R_9f_12054d58 );
buf ( n3079 , R_66_13308068 );
buf ( n3080 , R_219_1203c338 );
buf ( n3081 , R_132a5_12654868 );
buf ( n3082 , R_f9aa_11cdd5a8 );
buf ( n3083 , R_1fb_126610c8 );
buf ( n3084 , R_1a4_13798648 );
buf ( n3085 , R_16b_1331a2c8 );
buf ( n3086 , R_9a_12658568 );
buf ( n3087 , R_13c54_102f6e88 );
buf ( n3088 , R_14933_1207e5d8 );
buf ( n3089 , R_a6b7_1264b588 );
buf ( n3090 , R_10fad_13a15548 );
buf ( n3091 , R_18d_13321a28 );
buf ( n3092 , R_182_13315cc8 );
buf ( n3093 , R_14a58_102f65c8 );
buf ( n3094 , R_c8f6_132f4a08 );
buf ( n3095 , R_1458d_13a17ac8 );
buf ( n3096 , R_126d9_11545598 );
buf ( n3097 , R_10942_102f85a8 );
buf ( n3098 , R_14a32_12654ea8 );
buf ( n3099 , R_b7bc_12b28798 );
buf ( n3100 , R_1389f_11cda3a8 );
buf ( n3101 , R_14602_102ed7e8 );
buf ( n3102 , R_100bf_1330b9e8 );
buf ( n3103 , R_112eb_115386b8 );
buf ( n3104 , R_146d5_105b59f8 );
buf ( n3105 , R_1206a_1207c878 );
buf ( n3106 , R_e2de_1264ce88 );
buf ( n3107 , R_13b3a_11cddaa8 );
buf ( n3108 , R_13739_10563bf8 );
buf ( n3109 , R_148d6_11cd86e8 );
buf ( n3110 , R_1319d_11544918 );
buf ( n3111 , R_12f7f_12077eb8 );
buf ( n3112 , R_1242c_f8cda78 );
buf ( n3113 , R_14483_12054fd8 );
buf ( n3114 , R_14456_102ea728 );
buf ( n3115 , R_6b42_120790d8 );
buf ( n3116 , R_1186d_f8cbb38 );
buf ( n3117 , R_147d3_12648e28 );
buf ( n3118 , R_11add_1056c4d8 );
buf ( n3119 , R_13c18_1264df68 );
buf ( n3120 , R_13e19_132f7c08 );
buf ( n3121 , R_b6_1265e148 );
buf ( n3122 , R_13bb8_1265edc8 );
buf ( n3123 , R_146a8_12050118 );
buf ( n3124 , R_18e_12043ef8 );
buf ( n3125 , R_181_12647a28 );
buf ( n3126 , R_b677_12083178 );
buf ( n3127 , R_1176f_1379f8a8 );
buf ( n3128 , R_11d7b_102f2d88 );
buf ( n3129 , R_145bd_1207cff8 );
buf ( n3130 , R_13bae_105700d8 );
buf ( n3131 , R_10fed_1330ad68 );
buf ( n3132 , R_1479f_11cde4a8 );
buf ( n3133 , R_71_1265e8c8 );
buf ( n3134 , R_3ca5_102eebe8 );
buf ( n3135 , R_14769_1056b718 );
buf ( n3136 , R_139ba_11ce35e8 );
buf ( n3137 , R_ccf5_13a128e8 );
buf ( n3138 , R_13964_1207def8 );
buf ( n3139 , R_13920_133128e8 );
buf ( n3140 , R_13b74_11cd8dc8 );
buf ( n3141 , R_13e6d_11cd90e8 );
buf ( n3142 , R_13ae8_11545db8 );
buf ( n3143 , R_e946_13796668 );
buf ( n3144 , R_12db3_10562b18 );
buf ( n3145 , R_7b5f_1264bc68 );
buf ( n3146 , R_139f5_132fc348 );
buf ( n3147 , R_cd6e_10562a78 );
buf ( n3148 , R_13626_12077cd8 );
buf ( n3149 , R_148dc_102f3c88 );
buf ( n3150 , R_11db0_13302748 );
buf ( n3151 , R_1470b_115413f8 );
buf ( n3152 , R_fd8e_120835d8 );
buf ( n3153 , R_142aa_102f2a68 );
buf ( n3154 , R_1267b_1056b538 );
buf ( n3155 , R_10df7_1264ae08 );
buf ( n3156 , R_b753_102ebe48 );
buf ( n3157 , R_14a47_102eeb48 );
buf ( n3158 , R_12f94_1379c068 );
buf ( n3159 , R_f3d0_1264e3c8 );
buf ( n3160 , R_13cd6_10565638 );
buf ( n3161 , R_123b1_12b3e378 );
buf ( n3162 , R_144cf_f8c96f8 );
buf ( n3163 , R_13d0c_102f6168 );
buf ( n3164 , R_13c61_12081d78 );
buf ( n3165 , R_134f6_11ce6608 );
buf ( n3166 , R_112c2_12b294b8 );
buf ( n3167 , R_11922_1056c898 );
buf ( n3168 , R_11971_1207dbd8 );
buf ( n3169 , R_138_1265b308 );
buf ( n3170 , R_d2_12654c28 );
buf ( n3171 , R_23d_12656088 );
buf ( n3172 , R_8a_1379cba8 );
buf ( n3173 , R_38ad_12048418 );
buf ( n3174 , R_7b_12651de8 );
buf ( n3175 , R_13889_10564918 );
buf ( n3176 , R_13188_12079c18 );
buf ( n3177 , R_13b8c_13a15728 );
buf ( n3178 , R_947f_1056eaf8 );
buf ( n3179 , R_1d7_12649648 );
buf ( n3180 , R_149db_102f1668 );
buf ( n3181 , R_ac1d_120826d8 );
buf ( n3182 , R_13a06_105668f8 );
buf ( n3183 , R_18f_132fc988 );
buf ( n3184 , R_180_1265fea8 );
buf ( n3185 , R_10e36_11ce6d88 );
buf ( n3186 , R_136a7_12035cb8 );
buf ( n3187 , R_148df_13a1d608 );
buf ( n3188 , R_1380f_12080838 );
buf ( n3189 , R_1485b_1265a688 );
buf ( n3190 , R_14930_102f1a28 );
buf ( n3191 , R_10044_102f1c08 );
buf ( n3192 , R_d2a3_1207bbf8 );
buf ( n3193 , R_1c0_1203c0b8 );
buf ( n3194 , R_14f_12b25778 );
buf ( n3195 , R_8472_126654e8 );
buf ( n3196 , R_1483d_11ce0d48 );
buf ( n3197 , R_12b67_11cdf3a8 );
buf ( n3198 , R_11346_12655448 );
buf ( n3199 , R_13893_12084d98 );
buf ( n3200 , R_103f0_1207ecb8 );
buf ( n3201 , R_1308d_1379eea8 );
buf ( n3202 , R_f8ce_102f10c8 );
buf ( n3203 , R_13f82_11543978 );
buf ( n3204 , R_12359_133022e8 );
buf ( n3205 , R_12cd3_13a1f728 );
buf ( n3206 , R_13546_1153efb8 );
buf ( n3207 , R_143b6_115408b8 );
buf ( n3208 , R_148e5_10568518 );
buf ( n3209 , R_10a79_11545278 );
buf ( n3210 , R_1368d_102f3be8 );
buf ( n3211 , R_14002_12047518 );
buf ( n3212 , R_febc_1207caf8 );
buf ( n3213 , R_14987_10571d98 );
buf ( n3214 , R_14894_126569e8 );
buf ( n3215 , R_13e23_102f1708 );
buf ( n3216 , R_12304_10569e18 );
buf ( n3217 , R_12daa_f8cc218 );
buf ( n3218 , R_1289e_13316128 );
buf ( n3219 , R_146ea_132fd6a8 );
buf ( n3220 , R_104_12b414d8 );
buf ( n3221 , R_e9_12055a78 );
buf ( n3222 , R_226_12652568 );
buf ( n3223 , R_20b_12656bc8 );
buf ( n3224 , R_1484c_1056c078 );
buf ( n3225 , R_149fc_12077a58 );
buf ( n3226 , R_143f0_120442b8 );
buf ( n3227 , R_107_1203f538 );
buf ( n3228 , R_208_12b260d8 );
buf ( n3229 , R_1d2_1203ce78 );
buf ( n3230 , R_1442a_102f6668 );
buf ( n3231 , R_13d_1379c568 );
buf ( n3232 , R_134be_13a19148 );
buf ( n3233 , R_145cf_13304328 );
buf ( n3234 , R_12fa4_1153e0b8 );
buf ( n3235 , R_1053d_12079858 );
buf ( n3236 , R_ee_f8c86b8 );
buf ( n3237 , R_221_12652888 );
buf ( n3238 , R_13eb5_132f7ac8 );
buf ( n3239 , R_190_133178e8 );
buf ( n3240 , R_17f_115396f8 );
buf ( n3241 , R_137af_11ce6e28 );
buf ( n3242 , R_1455a_102ed748 );
buf ( n3243 , R_10db8_102f74c8 );
buf ( n3244 , R_ab_1264cde8 );
buf ( n3245 , R_1187e_12077698 );
buf ( n3246 , R_5a_126653a8 );
buf ( n3247 , R_7e57_13a1a188 );
buf ( n3248 , R_146ed_1153a238 );
buf ( n3249 , R_1b0_12b29918 );
buf ( n3250 , R_15f_1265f188 );
buf ( n3251 , R_138b8_1264a368 );
buf ( n3252 , R_13bd6_102f9188 );
buf ( n3253 , R_14a17_102f0ee8 );
buf ( n3254 , R_143a6_133121a8 );
buf ( n3255 , R_11f57_12649328 );
buf ( n3256 , R_14972_13302608 );
buf ( n3257 , R_10701_1207f1b8 );
buf ( n3258 , R_14503_1203e3b8 );
buf ( n3259 , R_a4_12b36e98 );
buf ( n3260 , R_6a_12b40178 );
buf ( n3261 , R_aeba_105624d8 );
buf ( n3262 , R_1379b_11ce6ec8 );
buf ( n3263 , R_134e2_13a1e3c8 );
buf ( n3264 , R_10973_12663008 );
buf ( n3265 , R_11c66_102f7ba8 );
buf ( n3266 , R_1325f_126468a8 );
buf ( n3267 , R_1327d_10570d58 );
buf ( n3268 , R_13417_102f3968 );
buf ( n3269 , R_101_1264f048 );
buf ( n3270 , R_95_133017a8 );
buf ( n3271 , R_20e_1265e788 );
buf ( n3272 , R_13c59_105b5638 );
buf ( n3273 , R_13ca1_12652f68 );
buf ( n3274 , R_1481c_11cdb988 );
buf ( n3275 , R_14611_11545458 );
buf ( n3276 , R_12fae_102f7388 );
buf ( n3277 , R_1469f_1207d138 );
buf ( n3278 , R_142dd_13314828 );
buf ( n3279 , R_1279d_12079fd8 );
buf ( n3280 , R_12646_1056b2b8 );
buf ( n3281 , R_11486_102ee788 );
buf ( n3282 , R_13389_1207fb18 );
buf ( n3283 , R_1492d_11ce64c8 );
buf ( n3284 , R_12d46_12648928 );
buf ( n3285 , R_145b7_12b3d5b8 );
buf ( n3286 , R_b211_12048c38 );
buf ( n3287 , R_143aa_13795c68 );
buf ( n3288 , R_1110c_11cdc928 );
buf ( n3289 , R_1a5_12b3c618 );
buf ( n3290 , R_16a_137a1248 );
buf ( n3291 , R_df67_1207b8d8 );
buf ( n3292 , R_124f6_1264f2c8 );
buf ( n3293 , R_12b54_102f2248 );
buf ( n3294 , R_d7dc_13a17de8 );
buf ( n3295 , R_1247b_11ce4808 );
buf ( n3296 , R_149ea_11540598 );
buf ( n3297 , R_10a_12b30678 );
buf ( n3298 , R_13c77_13a1cc08 );
buf ( n3299 , R_205_12653dc8 );
buf ( n3300 , R_14753_1264efa8 );
buf ( n3301 , R_191_12043d18 );
buf ( n3302 , R_17e_132f8568 );
buf ( n3303 , R_11c4b_13a15c28 );
buf ( n3304 , R_13208_11542758 );
buf ( n3305 , R_e0ad_133021a8 );
buf ( n3306 , R_11a3f_12b3e9b8 );
buf ( n3307 , R_1230e_f8cb598 );
buf ( n3308 , R_eee_1056adb8 );
buf ( n3309 , R_14444_12648108 );
buf ( n3310 , R_1dc_11538d98 );
buf ( n3311 , R_12b7a_1264f188 );
buf ( n3312 , R_133_13313888 );
buf ( n3313 , R_147b1_105b5a98 );
buf ( n3314 , R_f116_11ce1068 );
buf ( n3315 , R_13a5c_1379a268 );
buf ( n3316 , R_14340_12078458 );
buf ( n3317 , R_e522_1330ed28 );
buf ( n3318 , R_146f0_1153da78 );
buf ( n3319 , R_136f4_12649148 );
buf ( n3320 , R_119e8_1153e798 );
buf ( n3321 , R_1391b_12b277f8 );
buf ( n3322 , R_fd37_120394f8 );
buf ( n3323 , R_1461d_11539dd8 );
buf ( n3324 , R_ee50_102eb9e8 );
buf ( n3325 , R_dd_132f61c8 );
buf ( n3326 , R_232_105afa58 );
buf ( n3327 , R_4c_12652b08 );
buf ( n3328 , R_135a0_1153f0f8 );
buf ( n3329 , R_125d0_12b3f6d8 );
buf ( n3330 , R_b4_13302988 );
buf ( n3331 , R_51_13309648 );
buf ( n3332 , R_f925_12048b98 );
buf ( n3333 , R_14034_f8cf198 );
buf ( n3334 , R_123e9_f8c0eb8 );
buf ( n3335 , R_14726_1203bc58 );
buf ( n3336 , R_10894_1153ad78 );
buf ( n3337 , R_1b9_1379b7a8 );
buf ( n3338 , R_156_137927e8 );
buf ( n3339 , R_1471a_1379da08 );
buf ( n3340 , R_13d4e_11544f58 );
buf ( n3341 , R_112ae_115429d8 );
buf ( n3342 , R_dcb0_10564e18 );
buf ( n3343 , R_13ae3_12083498 );
buf ( n3344 , R_11a90_13a1ba88 );
buf ( n3345 , R_13f1a_10566998 );
buf ( n3346 , R_fdd5_1264d068 );
buf ( n3347 , R_13acb_13a17988 );
buf ( n3348 , R_ef1_13a16ee8 );
buf ( n3349 , R_145e1_12b40d58 );
buf ( n3350 , R_14915_102f7748 );
buf ( n3351 , R_ed3c_120760b8 );
buf ( n3352 , R_13cdc_11542398 );
buf ( n3353 , R_f544_102f5d08 );
buf ( n3354 , R_147e7_13793fa8 );
buf ( n3355 , R_e4_133095a8 );
buf ( n3356 , R_8d_1153d078 );
buf ( n3357 , R_78_12044178 );
buf ( n3358 , R_22b_12b3b538 );
buf ( n3359 , R_128ff_105b6178 );
buf ( n3360 , R_148ac_102f0f88 );
buf ( n3361 , R_1e9_133208a8 );
buf ( n3362 , R_192_12b44a98 );
buf ( n3363 , R_17d_12661f28 );
buf ( n3364 , R_12b83_13305e08 );
buf ( n3365 , R_fbb3_10567078 );
buf ( n3366 , R_126_12660588 );
buf ( n3367 , R_cfc6_1264a868 );
buf ( n3368 , R_1492a_13a1e1e8 );
buf ( n3369 , R_116bb_1207d6d8 );
buf ( n3370 , R_144d8_1330d9c8 );
buf ( n3371 , R_e6f2_102ecc08 );
buf ( n3372 , R_14a14_1207bdd8 );
buf ( n3373 , R_10f70_11544a58 );
buf ( n3374 , R_119fa_1207f2f8 );
buf ( n3375 , R_cef5_1265b6c8 );
buf ( n3376 , R_115b3_12082458 );
buf ( n3377 , R_211_1265c028 );
buf ( n3378 , R_146cc_11542618 );
buf ( n3379 , R_fe_120448f8 );
buf ( n3380 , R_119df_1056bad8 );
buf ( n3381 , R_13787_11ce21e8 );
buf ( n3382 , R_147dd_11ce6068 );
buf ( n3383 , R_14695_11cdf8a8 );
buf ( n3384 , R_149b1_102fa128 );
buf ( n3385 , R_110af_1379aee8 );
buf ( n3386 , R_14560_1330b3a8 );
buf ( n3387 , R_143ff_11cdca68 );
buf ( n3388 , R_d4_12654a48 );
buf ( n3389 , R_23b_13799408 );
buf ( n3390 , R_1c7_132fc0c8 );
buf ( n3391 , R_148_105aacd8 );
buf ( n3392 , R_13d6d_13a17668 );
buf ( n3393 , R_ce64_1056f9f8 );
buf ( n3394 , R_14474_13307a28 );
buf ( n3395 , R_12bde_102f62a8 );
buf ( n3396 , R_1436a_102eefa8 );
buf ( n3397 , R_14957_11540db8 );
buf ( n3398 , R_b634_11cdc068 );
buf ( n3399 , R_1460e_11ce2dc8 );
buf ( n3400 , R_f24f_11ce2fa8 );
buf ( n3401 , R_13763_105679d8 );
buf ( n3402 , R_f0b2_102f7f68 );
buf ( n3403 , R_14620_11ce6108 );
buf ( n3404 , R_131f5_12084618 );
buf ( n3405 , R_1490f_12651e88 );
buf ( n3406 , R_136cc_1264fcc8 );
buf ( n3407 , R_f227_1207a398 );
buf ( n3408 , R_13959_1153f918 );
buf ( n3409 , R_142cf_12659aa8 );
buf ( n3410 , R_f6b2_11cdfb28 );
buf ( n3411 , R_1ed_1203f5d8 );
buf ( n3412 , R_a2f6_11cdb3e8 );
buf ( n3413 , R_fc5e_13a18888 );
buf ( n3414 , R_122_12663d28 );
buf ( n3415 , R_13f67_12083b78 );
buf ( n3416 , R_13740_11cdb348 );
buf ( n3417 , R_146c9_1153fd78 );
buf ( n3418 , R_145db_13a12b68 );
buf ( n3419 , R_101ae_13a1fae8 );
buf ( n3420 , R_bb03_12b29ff8 );
buf ( n3421 , R_1101b_12045f38 );
buf ( n3422 , R_12bfd_10564b98 );
buf ( n3423 , R_121a5_1056a138 );
buf ( n3424 , R_127df_1330a728 );
buf ( n3425 , R_11617_105656d8 );
buf ( n3426 , R_13f90_12080518 );
buf ( n3427 , R_13be9_12662388 );
buf ( n3428 , R_12760_1331ab88 );
buf ( n3429 , R_126bb_10563b58 );
buf ( n3430 , R_147c6_12081cd8 );
buf ( n3431 , R_21c_12b41398 );
buf ( n3432 , R_13b33_102f0588 );
buf ( n3433 , R_1f8_132f5fe8 );
buf ( n3434 , R_11d2f_105665d8 );
buf ( n3435 , R_1227d_1265f2c8 );
buf ( n3436 , R_11a35_102f44a8 );
buf ( n3437 , R_1479c_1056c758 );
buf ( n3438 , R_116e4_12659828 );
buf ( n3439 , R_14662_1207ceb8 );
buf ( n3440 , R_14515_12079ad8 );
buf ( n3441 , R_117_12650c68 );
buf ( n3442 , R_115ca_11ce5fc8 );
buf ( n3443 , R_f3_1379bde8 );
buf ( n3444 , R_e229_102ecca8 );
buf ( n3445 , R_202_12b3f098 );
buf ( n3446 , R_1e5_1203a218 );
buf ( n3447 , R_12a_1331fea8 );
buf ( n3448 , R_10d_1330bda8 );
buf ( n3449 , R_135d6_1056fef8 );
buf ( n3450 , R_14918_13a1d888 );
buf ( n3451 , R_1452a_10564378 );
buf ( n3452 , R_14984_1056bc18 );
buf ( n3453 , R_1cd_1265c8e8 );
buf ( n3454 , R_eb34_11cda628 );
buf ( n3455 , R_125ac_11ce4308 );
buf ( n3456 , R_193_f8c7cb8 );
buf ( n3457 , R_1216d_1264d7e8 );
buf ( n3458 , R_17c_132fe648 );
buf ( n3459 , R_142_13792ce8 );
buf ( n3460 , R_cdb8_102f4f48 );
buf ( n3461 , R_144bd_11cdeb88 );
buf ( n3462 , R_131ae_1056bd58 );
buf ( n3463 , R_14909_1379f768 );
buf ( n3464 , R_14924_12b3adb8 );
buf ( n3465 , R_102a2_12b41e38 );
buf ( n3466 , R_13aa8_120525f8 );
buf ( n3467 , R_d3ca_102ef7c8 );
buf ( n3468 , R_1459f_120792b8 );
buf ( n3469 , R_120b3_12b407b8 );
buf ( n3470 , R_127a7_105683d8 );
buf ( n3471 , R_14545_1056b218 );
buf ( n3472 , R_12056_1204f178 );
buf ( n3473 , R_11f2a_10563ab8 );
buf ( n3474 , R_e021_12b26718 );
buf ( n3475 , R_f377_1056d1f8 );
buf ( n3476 , R_127ca_13a16da8 );
buf ( n3477 , R_14689_120838f8 );
buf ( n3478 , R_11be7_1207a6b8 );
buf ( n3479 , R_139a1_1264c668 );
buf ( n3480 , R_14536_12b42978 );
buf ( n3481 , R_13c2d_11cdd828 );
buf ( n3482 , R_14906_11544ff8 );
buf ( n3483 , R_11a5d_132f52c8 );
buf ( n3484 , R_ca63_1331c8e8 );
buf ( n3485 , R_14714_102f77e8 );
buf ( n3486 , R_14799_137933c8 );
buf ( n3487 , R_1390f_13a14828 );
buf ( n3488 , R_1234f_12083858 );
buf ( n3489 , R_142c6_12081738 );
buf ( n3490 , R_127ae_12b3ccf8 );
buf ( n3491 , R_13590_12079a38 );
buf ( n3492 , R_148b8_102eaa48 );
buf ( n3493 , R_5735_137a0988 );
buf ( n3494 , R_1a6_12038698 );
buf ( n3495 , R_169_1203e458 );
buf ( n3496 , R_127c1_12082638 );
buf ( n3497 , R_1288a_137a1ec8 );
buf ( n3498 , R_1488e_102f6708 );
buf ( n3499 , R_113b9_1264ea08 );
buf ( n3500 , R_1430f_11cd8fa8 );
buf ( n3501 , R_f97f_13304dc8 );
buf ( n3502 , R_104fa_120761f8 );
buf ( n3503 , R_119ae_11cdfa88 );
buf ( n3504 , R_12c78_1207ca58 );
buf ( n3505 , R_d606_11ce46c8 );
buf ( n3506 , R_146a5_102f90e8 );
buf ( n3507 , R_14900_120781d8 );
buf ( n3508 , R_1374f_13a16808 );
buf ( n3509 , R_ff3c_11ce1f68 );
buf ( n3510 , R_e834_10564238 );
buf ( n3511 , R_14a5e_105aa4b8 );
buf ( n3512 , R_13465_13316bc8 );
buf ( n3513 , R_13d25_11540b38 );
buf ( n3514 , R_56_13308248 );
buf ( n3515 , R_ef7_1153e838 );
buf ( n3516 , R_13193_102ec7a8 );
buf ( n3517 , R_132f1_13a145a8 );
buf ( n3518 , R_1291e_1056ee18 );
buf ( n3519 , R_14921_105640f8 );
buf ( n3520 , R_1371a_12083fd8 );
buf ( n3521 , R_14837_132f32e8 );
buf ( n3522 , R_13a37_12b3d338 );
buf ( n3523 , R_dad2_1379c6a8 );
buf ( n3524 , R_1495d_12b43878 );
buf ( n3525 , R_149f3_12b27c58 );
buf ( n3526 , R_107c6_1203f998 );
buf ( n3527 , R_1456c_12b437d8 );
buf ( n3528 , R_11888_13794868 );
buf ( n3529 , R_13b62_13a13428 );
buf ( n3530 , R_1360f_10563158 );
buf ( n3531 , R_1b1_12657ac8 );
buf ( n3532 , R_10844_1153e1f8 );
buf ( n3533 , R_194_1331d4c8 );
buf ( n3534 , R_17b_1265ea08 );
buf ( n3535 , R_15e_126544a8 );
buf ( n3536 , R_be25_102ec028 );
buf ( n3537 , R_148fd_102eb768 );
buf ( n3538 , R_14683_13a1d9c8 );
buf ( n3539 , R_a069_12080298 );
buf ( n3540 , R_1233a_13a143c8 );
buf ( n3541 , R_6e_13304b48 );
buf ( n3542 , R_1334f_1204e598 );
buf ( n3543 , R_121e7_1207ff78 );
buf ( n3544 , R_12bb7_102f3e68 );
buf ( n3545 , R_12bcc_12652608 );
buf ( n3546 , R_f783_13797b08 );
buf ( n3547 , R_14680_12076fb8 );
buf ( n3548 , R_13d2b_12085338 );
buf ( n3549 , R_11bbe_1153de38 );
buf ( n3550 , R_148e8_1264bda8 );
buf ( n3551 , R_148fa_102f5948 );
buf ( n3552 , R_149d8_132fc168 );
buf ( n3553 , R_148ee_120808d8 );
buf ( n3554 , R_148f4_11cd8468 );
buf ( n3555 , R_ff98_12b41618 );
buf ( n3556 , R_13bc3_102f8d28 );
buf ( n3557 , R_12b1f_120564d8 );
buf ( n3558 , R_c961_12080f18 );
buf ( n3559 , R_214_12655588 );
buf ( n3560 , R_dff5_102ed9c8 );
buf ( n3561 , R_13d49_13a16bc8 );
buf ( n3562 , R_fb_1379f808 );
buf ( n3563 , R_12958_102f1848 );
buf ( n3564 , R_12220_1379e908 );
buf ( n3565 , R_144de_12076798 );
buf ( n3566 , R_c6d1_10566178 );
buf ( n3567 , R_11547_1264cc08 );
buf ( n3568 , R_138ac_102eb128 );
buf ( n3569 , R_12853_105b58b8 );
buf ( n3570 , R_1f1_12655268 );
buf ( n3571 , R_11e_12b29b98 );
buf ( n3572 , R_13d30_1207b658 );
buf ( n3573 , R_b2_105aa0f8 );
buf ( n3574 , R_d5a1_105690f8 );
buf ( n3575 , R_c700_13304788 );
buf ( n3576 , R_a359_12662888 );
buf ( n3577 , R_1449f_12055898 );
buf ( n3578 , R_14587_10565ef8 );
buf ( n3579 , R_14759_1056e378 );
buf ( n3580 , R_1385d_1056ab38 );
buf ( n3581 , R_1401f_132fb588 );
buf ( n3582 , R_1245b_12658f68 );
buf ( n3583 , R_fe3a_11cdb168 );
buf ( n3584 , R_a47d_13a18f68 );
buf ( n3585 , R_145ea_1056c438 );
buf ( n3586 , R_99a4_102f5bc8 );
buf ( n3587 , R_1491e_12661528 );
buf ( n3588 , R_1c1_126618e8 );
buf ( n3589 , R_b180_12039a98 );
buf ( n3590 , R_14e_12b29e18 );
buf ( n3591 , R_13b1f_12052c38 );
buf ( n3592 , R_146e4_f8cb638 );
buf ( n3593 , R_14581_10571b18 );
buf ( n3594 , R_1354d_12040078 );
buf ( n3595 , R_13508_120842f8 );
buf ( n3596 , R_148d9_13a14d28 );
buf ( n3597 , R_149c0_102ed068 );
buf ( n3598 , R_1477e_10568fb8 );
buf ( n3599 , R_14735_105680b8 );
buf ( n3600 , R_13d35_11ce1108 );
buf ( n3601 , R_4d49_102f8dc8 );
buf ( n3602 , R_133aa_11545b38 );
buf ( n3603 , R_14518_102f67a8 );
buf ( n3604 , R_bf1d_1153d618 );
buf ( n3605 , R_a9_1204d4b8 );
buf ( n3606 , R_14702_12b3d0b8 );
buf ( n3607 , R_1431c_11cde188 );
buf ( n3608 , R_9323_1331d068 );
buf ( n3609 , R_14a2f_12075ed8 );
buf ( n3610 , R_1e1_13321ca8 );
buf ( n3611 , R_12e_105af9b8 );
buf ( n3612 , R_9d_1379c9c8 );
buf ( n3613 , R_12caa_126508a8 );
buf ( n3614 , R_115df_10566c18 );
buf ( n3615 , R_144fd_102f1b68 );
buf ( n3616 , R_127f1_12b2a098 );
buf ( n3617 , R_137eb_12082138 );
buf ( n3618 , R_11b9a_12b3f278 );
buf ( n3619 , R_1483a_12081f58 );
buf ( n3620 , R_7d2b_11ce4948 );
buf ( n3621 , R_13a49_102f8e68 );
buf ( n3622 , R_1493c_11cdc568 );
buf ( n3623 , R_14a3e_102ed428 );
buf ( n3624 , R_195_12045cb8 );
buf ( n3625 , R_14489_12b3fe58 );
buf ( n3626 , R_17a_1330dc48 );
buf ( n3627 , R_1066b_1264a228 );
buf ( n3628 , R_139b5_11536318 );
buf ( n3629 , R_12775_126513e8 );
buf ( n3630 , R_13d43_13a1c168 );
buf ( n3631 , R_13e78_1056a598 );
buf ( n3632 , R_90_f8cccb8 );
buf ( n3633 , R_75_12b443b8 );
buf ( n3634 , R_14816_10565db8 );
buf ( n3635 , R_e4c7_10571398 );
buf ( n3636 , R_14354_13317348 );
buf ( n3637 , R_146c3_12b3bfd8 );
buf ( n3638 , R_db95_12b2ff98 );
buf ( n3639 , R_b45b_11ce7508 );
buf ( n3640 , R_145de_1056b5d8 );
buf ( n3641 , R_13c7d_1056d798 );
buf ( n3642 , R_c7c0_102ed4c8 );
buf ( n3643 , R_1ff_13315c28 );
buf ( n3644 , R_1361a_102f01c8 );
buf ( n3645 , R_110_1204b938 );
buf ( n3646 , R_10c17_13a13888 );
buf ( n3647 , R_d6_1264b1c8 );
buf ( n3648 , R_239_12b2a958 );
buf ( n3649 , R_144a8_115369f8 );
buf ( n3650 , R_12516_13305188 );
buf ( n3651 , R_14699_10567e38 );
buf ( n3652 , R_12de4_12045b18 );
buf ( n3653 , R_10fd9_11ce1928 );
buf ( n3654 , R_145c6_13a1cb68 );
buf ( n3655 , R_147c3_13a177a8 );
buf ( n3656 , R_1313e_1207a1b8 );
buf ( n3657 , R_e9a6_1153dcf8 );
buf ( n3658 , R_123a6_12077418 );
buf ( n3659 , R_e669_1056eb98 );
buf ( n3660 , R_eea5_13793c88 );
buf ( n3661 , R_8e12_f8c7538 );
buf ( n3662 , R_11a2c_12b3f1d8 );
buf ( n3663 , R_bc89_12664548 );
buf ( n3664 , R_b132_13300a88 );
buf ( n3665 , R_14626_102f4ae8 );
buf ( n3666 , R_125c9_11ce5c08 );
buf ( n3667 , R_14891_1265e0a8 );
buf ( n3668 , R_13ba9_1056f4f8 );
buf ( n3669 , R_11299_1056a4f8 );
buf ( n3670 , R_1395f_1207ba18 );
buf ( n3671 , R_1085f_13312a28 );
buf ( n3672 , R_c642_12b41b18 );
buf ( n3673 , R_1445c_f8ce478 );
buf ( n3674 , R_14981_12b3f598 );
buf ( n3675 , R_148e2_12650b28 );
buf ( n3676 , R_988f_13a1e968 );
buf ( n3677 , R_962b_105647d8 );
buf ( n3678 , R_124a7_12079498 );
buf ( n3679 , R_fe64_1153f378 );
buf ( n3680 , R_11f16_102eb088 );
buf ( n3681 , R_13e03_1379bf28 );
buf ( n3682 , R_14927_11cdf808 );
buf ( n3683 , R_1ba_1330eb48 );
buf ( n3684 , R_14471_13793be8 );
buf ( n3685 , R_121fd_11ce3048 );
buf ( n3686 , R_14499_1207a9d8 );
buf ( n3687 , R_155_12b43f58 );
buf ( n3688 , R_98_12048af8 );
buf ( n3689 , R_e916_105699b8 );
buf ( n3690 , R_e1ea_1056b998 );
buf ( n3691 , R_11af3_13793788 );
buf ( n3692 , R_13bcf_12650948 );
buf ( n3693 , R_10070_12077e18 );
buf ( n3694 , R_f2f6_126613e8 );
buf ( n3695 , R_104a3_11542d98 );
buf ( n3696 , R_149ae_10565138 );
buf ( n3697 , R_1430b_1204c8d8 );
buf ( n3698 , R_ede8_1056dfb8 );
buf ( n3699 , R_13495_13a1e008 );
buf ( n3700 , R_df_132f6808 );
buf ( n3701 , R_230_12664a48 );
buf ( n3702 , R_136ac_102eacc8 );
buf ( n3703 , R_dd20_137974c8 );
buf ( n3704 , R_14741_132f2c08 );
buf ( n3705 , R_137c1_11543dd8 );
buf ( n3706 , R_14364_11ce6568 );
buf ( n3707 , R_11d60_132fc8e8 );
buf ( n3708 , R_14a44_105b60d8 );
buf ( n3709 , R_13749_11543518 );
buf ( n3710 , R_854a_1207fed8 );
buf ( n3711 , R_14a11_12045a78 );
buf ( n3712 , R_1a7_12659b48 );
buf ( n3713 , R_168_105b3158 );
buf ( n3714 , R_f03_13a17208 );
buf ( n3715 , R_1274c_12653fa8 );
buf ( n3716 , R_147b7_12079df8 );
buf ( n3717 , R_a2_1379e228 );
buf ( n3718 , R_63_f8c7b78 );
buf ( n3719 , R_13c49_102ecac8 );
buf ( n3720 , R_d68f_12078a98 );
buf ( n3721 , R_148f1_11cde688 );
buf ( n3722 , R_196_11536778 );
buf ( n3723 , R_179_13301c08 );
buf ( n3724 , R_11c1b_120757f8 );
buf ( n3725 , R_1181a_10565098 );
buf ( n3726 , R_14912_13300628 );
buf ( n3727 , R_10c93_13310768 );
buf ( n3728 , R_147f2_10571618 );
buf ( n3729 , R_c832_12075f78 );
buf ( n3730 , R_14530_11540778 );
buf ( n3731 , R_e8ba_11ce3b88 );
buf ( n3732 , R_14903_11ce50c8 );
buf ( n3733 , R_14629_115412b8 );
buf ( n3734 , R_11966_10562118 );
buf ( n3735 , R_f8fa_105b4d78 );
buf ( n3736 , R_1d8_1331f5e8 );
buf ( n3737 , R_1281b_1207f6b8 );
buf ( n3738 , R_137_1331a7c8 );
buf ( n3739 , R_5f_12b428d8 );
buf ( n3740 , R_12288_126495a8 );
buf ( n3741 , R_a469_13a14648 );
buf ( n3742 , R_130cc_13a17348 );
buf ( n3743 , R_136e6_11cdcb08 );
buf ( n3744 , R_d806_102f5a88 );
buf ( n3745 , R_fd98_12052d78 );
buf ( n3746 , R_144b4_1153eab8 );
buf ( n3747 , R_1482b_12b3b3f8 );
buf ( n3748 , R_13858_12081e18 );
buf ( n3749 , R_1d3_1265ae08 );
buf ( n3750 , R_13c_1265b1c8 );
buf ( n3751 , R_14596_12048558 );
buf ( n3752 , R_eb_1153bf98 );
buf ( n3753 , R_224_12b29698 );
buf ( n3754 , R_13d3c_132f70c8 );
buf ( n3755 , R_c353_102f31e8 );
buf ( n3756 , R_1092e_13a140a8 );
buf ( n3757 , R_1018e_10563478 );
buf ( n3758 , R_12875_1153eb58 );
buf ( n3759 , R_13693_13795448 );
buf ( n3760 , R_123bb_11ce7008 );
buf ( n3761 , R_dfc9_12647208 );
buf ( n3762 , R_da6d_12082098 );
buf ( n3763 , R_1198e_1153d758 );
buf ( n3764 , R_149ff_1264c848 );
buf ( n3765 , R_1180e_12648248 );
buf ( n3766 , R_12535_126604e8 );
buf ( n3767 , R_12780_10568b58 );
buf ( n3768 , R_9dc0_102f6f28 );
buf ( n3769 , R_c4a7_1330a908 );
buf ( n3770 , R_11bfb_12649968 );
buf ( n3771 , R_13fe4_105622f8 );
buf ( n3772 , R_12e0c_13797388 );
buf ( n3773 , R_1454e_11ce1c48 );
buf ( n3774 , R_14069_1153db18 );
buf ( n3775 , R_10c0e_120464d8 );
buf ( n3776 , R_13c1f_f8c8938 );
buf ( n3777 , R_d910_1056e418 );
buf ( n3778 , R_cfae_13a15368 );
buf ( n3779 , R_10806_1264d608 );
buf ( n3780 , R_13706_13319b48 );
buf ( n3781 , R_12e21_1330cb68 );
buf ( n3782 , R_f8_12665808 );
buf ( n3783 , R_67_105aac38 );
buf ( n3784 , R_217_105b3fb8 );
buf ( n3785 , R_12a8e_1264ef08 );
buf ( n3786 , R_e5ea_115436f8 );
buf ( n3787 , R_14858_10571c58 );
buf ( n3788 , R_111b8_102ebbc8 );
buf ( n3789 , R_12ba4_12b28ab8 );
buf ( n3790 , R_108f1_102f35a8 );
buf ( n3791 , R_138a5_1264e468 );
buf ( n3792 , R_131ff_13a1eaa8 );
buf ( n3793 , R_11448_11ce41c8 );
buf ( n3794 , R_11534_13a13ce8 );
buf ( n3795 , R_12d1d_1207c238 );
buf ( n3796 , R_134e8_13a1e8c8 );
buf ( n3797 , R_b82e_1153c2b8 );
buf ( n3798 , R_11572_11ce43a8 );
buf ( n3799 , R_14897_1265c988 );
buf ( n3800 , R_125fa_1265b128 );
buf ( n3801 , R_b95d_102f8008 );
buf ( n3802 , R_14436_10570718 );
buf ( n3803 , R_f951_132fcde8 );
buf ( n3804 , R_10246_1056ae58 );
buf ( n3805 , R_12041_11ce0ac8 );
buf ( n3806 , R_138cd_1153e018 );
buf ( n3807 , R_1b2_12660f88 );
buf ( n3808 , R_197_1379a768 );
buf ( n3809 , R_121dd_12659328 );
buf ( n3810 , R_178_12658d88 );
buf ( n3811 , R_15d_133195a8 );
buf ( n3812 , R_13f24_13318428 );
buf ( n3813 , R_146f6_132fbc68 );
buf ( n3814 , R_b880_12083d58 );
buf ( n3815 , R_12ab4_132f57c8 );
buf ( n3816 , R_ed14_133110c8 );
buf ( n3817 , R_144f0_132ff0e8 );
buf ( n3818 , R_10aa5_12053f98 );
buf ( n3819 , R_1290a_11ce1388 );
buf ( n3820 , R_9d4e_11cddbe8 );
buf ( n3821 , R_e6_12b344f8 );
buf ( n3822 , R_b0_12b3f458 );
buf ( n3823 , R_229_126659e8 );
buf ( n3824 , R_12b3f_105b6538 );
buf ( n3825 , R_1f5_1203e958 );
buf ( n3826 , R_f624_1265b808 );
buf ( n3827 , R_14711_11ce2828 );
buf ( n3828 , R_fe05_102f9548 );
buf ( n3829 , R_1118b_11cdb8e8 );
buf ( n3830 , R_1c8_f8c6b38 );
buf ( n3831 , R_147_12b38c98 );
buf ( n3832 , R_11a_1204b438 );
buf ( n3833 , R_14778_13a1f688 );
buf ( n3834 , R_137fd_11544418 );
buf ( n3835 , R_f0_13795d08 );
buf ( n3836 , R_c3_132ff188 );
buf ( n3837 , R_21f_1265a2c8 );
buf ( n3838 , R_12e60_132f3a68 );
buf ( n3839 , R_4a02_12646e48 );
buf ( n3840 , R_c5_12657e88 );
buf ( n3841 , R_132ae_1056ef58 );
buf ( n3842 , R_d400_133126a8 );
buf ( n3843 , R_128a8_f8c9978 );
buf ( n3844 , R_ecbd_12040a78 );
buf ( n3845 , R_146ba_11cd8c88 );
buf ( n3846 , R_ea59_102f5088 );
buf ( n3847 , R_1183a_1204a498 );
buf ( n3848 , R_13d1f_1207ddb8 );
buf ( n3849 , R_136e0_11ce7148 );
buf ( n3850 , R_ddb7_12078b38 );
buf ( n3851 , R_14575_13307c08 );
buf ( n3852 , R_14864_13a1b768 );
buf ( n3853 , R_1471d_12040bb8 );
buf ( n3854 , R_11237_1056f958 );
buf ( n3855 , R_13fee_12663288 );
buf ( n3856 , R_c1_1204fd58 );
buf ( n3857 , R_14632_11cd85a8 );
buf ( n3858 , R_4d_12662d88 );
buf ( n3859 , R_b895_1264a4a8 );
buf ( n3860 , R_11b87_12648b08 );
buf ( n3861 , R_111c4_12076658 );
buf ( n3862 , R_a534_12b3d018 );
buf ( n3863 , R_11805_12b41578 );
buf ( n3864 , R_c901_126603a8 );
buf ( n3865 , R_13bde_13a1bbc8 );
buf ( n3866 , R_149b4_10564d78 );
buf ( n3867 , R_c7_126589c8 );
buf ( n3868 , R_248_1331ef08 );
buf ( n3869 , R_5b_12655088 );
buf ( n3870 , R_13720_102f3f08 );
buf ( n3871 , R_b9b1_1056c9d8 );
buf ( n3872 , R_f1cc_10567ed8 );
buf ( n3873 , R_cd0b_11542f78 );
buf ( n3874 , R_1497b_11cdfda8 );
buf ( n3875 , R_12d6f_13799b88 );
buf ( n3876 , R_14305_120844d8 );
buf ( n3877 , R_145ae_102efe08 );
buf ( n3878 , R_147d6_12b27b18 );
buf ( n3879 , R_13dc3_11cdbf28 );
buf ( n3880 , R_dc22_1153d438 );
buf ( n3881 , R_5970_11cdbe88 );
buf ( n3882 , R_113_1265c528 );
buf ( n3883 , R_82_f8cbc78 );
buf ( n3884 , R_1fc_12050078 );
buf ( n3885 , R_b00a_1153e658 );
buf ( n3886 , R_1346e_10567bb8 );
buf ( n3887 , R_1dd_12b395f8 );
buf ( n3888 , R_10390_1207ed58 );
buf ( n3889 , R_12cf4_13310ee8 );
buf ( n3890 , R_10675_1203cab8 );
buf ( n3891 , R_1399b_1264c3e8 );
buf ( n3892 , R_132_120518d8 );
buf ( n3893 , R_d8_12b3c938 );
buf ( n3894 , R_237_105a9fb8 );
buf ( n3895 , R_d4b2_1265bda8 );
buf ( n3896 , R_14453_12649d28 );
buf ( n3897 , R_10e2c_102ecde8 );
buf ( n3898 , R_52_13799868 );
buf ( n3899 , R_143dc_120824f8 );
buf ( n3900 , R_13ebe_11ce4128 );
buf ( n3901 , R_14053_102f21a8 );
buf ( n3902 , R_10960_133050e8 );
buf ( n3903 , R_1037b_1264a048 );
buf ( n3904 , R_7fe6_12b3f638 );
buf ( n3905 , R_12685_11cdf088 );
buf ( n3906 , R_135e9_11ce0de8 );
buf ( n3907 , R_bf_1379fa88 );
buf ( n3908 , R_85_12b41898 );
buf ( n3909 , R_149d5_11541358 );
buf ( n3910 , R_13f4d_10561fd8 );
buf ( n3911 , R_d0f1_1056a1d8 );
buf ( n3912 , R_a3f3_12646da8 );
buf ( n3913 , R_1311d_13a131a8 );
buf ( n3914 , R_1026e_11541ad8 );
buf ( n3915 , R_139de_13310588 );
buf ( n3916 , R_144cc_11ce23c8 );
buf ( n3917 , R_1403a_1331cc08 );
buf ( n3918 , R_1ce_12656628 );
buf ( n3919 , R_198_12b3fdb8 );
buf ( n3920 , R_d37f_1379a1c8 );
buf ( n3921 , R_177_1330de28 );
buf ( n3922 , R_141_12b3cf78 );
buf ( n3923 , R_14500_102f92c8 );
buf ( n3924 , R_c9_12b28fb8 );
buf ( n3925 , R_246_1203df58 );
buf ( n3926 , R_93_12659be8 );
buf ( n3927 , R_72_132fe788 );
buf ( n3928 , R_125bf_105685b8 );
buf ( n3929 , R_1a8_137a0d48 );
buf ( n3930 , R_147a5_1264a728 );
buf ( n3931 , R_167_1204f678 );
buf ( n3932 , R_7f_105ac998 );
buf ( n3933 , R_149f0_13a1fea8 );
buf ( n3934 , R_12210_13793aa8 );
buf ( n3935 , R_13db7_11ce11a8 );
buf ( n3936 , R_100e9_132f3ec8 );
buf ( n3937 , R_5362_13a18108 );
buf ( n3938 , R_124d7_13a18e28 );
buf ( n3939 , R_14a55_133001c8 );
buf ( n3940 , R_12419_1153d398 );
buf ( n3941 , R_108b6_1264e0a8 );
buf ( n3942 , R_10d4d_11cded68 );
buf ( n3943 , R_1464a_13a15b88 );
buf ( n3944 , R_c7f2_11cdc748 );
buf ( n3945 , R_13c83_11544698 );
buf ( n3946 , R_1489a_f8c6c78 );
buf ( n3947 , R_125b6_12040b18 );
buf ( n3948 , R_c00b_12079718 );
buf ( n3949 , R_eeb_13a13608 );
buf ( n3950 , R_f088_1330ba88 );
buf ( n3951 , R_1365e_1207b838 );
buf ( n3952 , R_fa81_12052198 );
buf ( n3953 , R_145f3_13a14788 );
buf ( n3954 , R_10995_102f3148 );
buf ( n3955 , R_123f8_13a13388 );
buf ( n3956 , R_6358_1204fe98 );
buf ( n3957 , R_14763_11ce4c68 );
buf ( n3958 , R_1433c_12077c38 );
buf ( n3959 , R_dde7_13a141e8 );
buf ( n3960 , R_13ef9_1204a858 );
buf ( n3961 , R_14810_1056db58 );
buf ( n3962 , R_13fdc_102f15c8 );
buf ( n3963 , R_d995_11ce0fc8 );
buf ( n3964 , R_117fc_12056078 );
buf ( n3965 , R_8d57_11ce53e8 );
buf ( n3966 , R_11bb4_12b39cd8 );
buf ( n3967 , R_13b97_1207a438 );
buf ( n3968 , R_14068_11cdc108 );
buf ( n3969 , R_1335a_105b5ef8 );
buf ( n3970 , R_1043d_13a1c5c8 );
buf ( n3971 , R_128cf_11cdabc8 );
buf ( n3972 , R_1219b_1207a938 );
buf ( n3973 , R_10dce_105631f8 );
buf ( n3974 , R_bbfa_10564418 );
buf ( n3975 , R_11864_12b44318 );
buf ( n3976 , R_12435_11ce4088 );
buf ( n3977 , R_a7_1265a5e8 );
buf ( n3978 , R_111f4_11cdf6c8 );
buf ( n3979 , R_135cf_1207eb78 );
buf ( n3980 , R_102ef_1153c218 );
buf ( n3981 , R_12ca0_11ce0668 );
buf ( n3982 , R_1c2_1330f228 );
buf ( n3983 , R_c6f4_12056438 );
buf ( n3984 , R_1404f_12b3e738 );
buf ( n3985 , R_ee7b_1379a628 );
buf ( n3986 , R_127e9_f8c8078 );
buf ( n3987 , R_14d_1203cbf8 );
buf ( n3988 , R_bd_1203f3f8 );
buf ( n3989 , R_48_13301848 );
buf ( n3990 , R_10afa_13a15d68 );
buf ( n3991 , R_ed66_11ce3368 );
buf ( n3992 , R_13a92_102f0bc8 );
buf ( n3993 , R_e9fb_12646268 );
buf ( n3994 , R_10d30_12084078 );
buf ( n3995 , R_149ab_1153d7f8 );
buf ( n3996 , R_88_13300d08 );
buf ( n3997 , R_6b_105aaff8 );
buf ( n3998 , R_11c31_115418f8 );
buf ( n3999 , R_13677_102f9868 );
buf ( n4000 , R_133f2_1379f088 );
buf ( n4001 , R_13edf_120837b8 );
buf ( n4002 , R_d399_137980a8 );
buf ( n4003 , R_1446e_1207d958 );
buf ( n4004 , R_1382d_1207d9f8 );
buf ( n4005 , R_cb_1331fa48 );
buf ( n4006 , R_244_1264c708 );
buf ( n4007 , R_12dc8_13a1f548 );
buf ( n4008 , R_12299_1265d1a8 );
buf ( n4009 , R_1474a_12076dd8 );
buf ( n4010 , R_13844_12663aa8 );
buf ( n4011 , R_13c11_1153d578 );
buf ( n4012 , R_14650_1056f278 );
buf ( n4013 , R_146fc_12647848 );
buf ( n4014 , R_10f84_1207bab8 );
buf ( n4015 , R_131cc_12b272f8 );
buf ( n4016 , R_1451b_10567cf8 );
buf ( n4017 , R_14390_10567c58 );
buf ( n4018 , R_13754_12082318 );
buf ( n4019 , R_1bb_12664868 );
buf ( n4020 , R_154_1204e1d8 );
buf ( n4021 , R_14831_1264f408 );
buf ( n4022 , R_7c_105b1cb8 );
buf ( n4023 , R_f1a0_12075938 );
buf ( n4024 , R_e9d0_1153f558 );
buf ( n4025 , R_f0eb_102f7568 );
buf ( n4026 , R_fb0c_1331a368 );
buf ( n4027 , R_1397b_1331b268 );
buf ( n4028 , R_e589_1379bb68 );
buf ( n4029 , R_1381a_120547b8 );
buf ( n4030 , R_1463e_105703f8 );
buf ( n4031 , R_12e76_11cd9908 );
buf ( n4032 , R_199_132fb3a8 );
buf ( n4033 , R_176_12b265d8 );
buf ( n4034 , R_125_13798008 );
buf ( n4035 , R_11ad2_102ed108 );
buf ( n4036 , R_1ea_1265a868 );
buf ( n4037 , R_10764_11cd9548 );
buf ( n4038 , R_14563_1264d6a8 );
buf ( n4039 , R_12c1a_102f0268 );
buf ( n4040 , R_146d2_1203a998 );
buf ( n4041 , R_147bd_102f9048 );
buf ( n4042 , R_fa57_1207f398 );
buf ( n4043 , R_c5a3_120849d8 );
buf ( n4044 , R_11dc9_f8c9b58 );
buf ( n4045 , R_11d95_1153f198 );
buf ( n4046 , R_1329b_11cd95e8 );
buf ( n4047 , R_14861_f8c41f8 );
buf ( n4048 , R_1064a_10561f38 );
buf ( n4049 , R_ce07_f8c8f78 );
buf ( n4050 , R_14720_11ce07a8 );
buf ( n4051 , R_13ca7_12078098 );
buf ( n4052 , R_147f5_1207a078 );
buf ( n4053 , R_142d3_12036758 );
buf ( n4054 , R_13dee_12083a38 );
buf ( n4055 , R_ec91_126490a8 );
buf ( n4056 , R_13421_11544c38 );
buf ( n4057 , R_cf92_11cdfee8 );
buf ( n4058 , R_4c49_13a1d748 );
buf ( n4059 , R_114d1_13307de8 );
buf ( n4060 , R_cff7_12076bf8 );
buf ( n4061 , R_142ff_11ce1b08 );
buf ( n4062 , R_139c0_13a1e5a8 );
buf ( n4063 , R_143cc_1056e738 );
buf ( n4064 , R_ba4e_13a1d388 );
buf ( n4065 , R_12485_105b6358 );
buf ( n4066 , R_11f0c_13a1aea8 );
buf ( n4067 , R_14867_12054b78 );
buf ( n4068 , R_137b5_10569cd8 );
buf ( n4069 , R_11d1b_12649288 );
buf ( n4070 , R_13d7b_102f56c8 );
buf ( n4071 , R_14a2c_102f12a8 );
buf ( n4072 , R_14608_13a155e8 );
buf ( n4073 , R_144c9_10571578 );
buf ( n4074 , R_fc0a_11541858 );
buf ( n4075 , R_144fa_120775f8 );
buf ( n4076 , R_129_1331c988 );
buf ( n4077 , R_13561_1330d068 );
buf ( n4078 , R_e1_12661708 );
buf ( n4079 , R_1299a_1207b158 );
buf ( n4080 , R_1489d_105686f8 );
buf ( n4081 , R_22e_132f2ac8 );
buf ( n4082 , R_6d01_102f72e8 );
buf ( n4083 , R_ffc3_12656e48 );
buf ( n4084 , R_1496f_102f9908 );
buf ( n4085 , R_1e6_13792a68 );
buf ( n4086 , R_14760_11ce3868 );
buf ( n4087 , R_d2d1_13793468 );
buf ( n4088 , R_12145_1207b978 );
buf ( n4089 , R_f5_11537038 );
buf ( n4090 , R_bb_13799cc8 );
buf ( n4091 , R_21a_1265b088 );
buf ( n4092 , R_14975_11541998 );
buf ( n4093 , R_147c0_11ce20a8 );
buf ( n4094 , R_13b7f_1153a198 );
buf ( n4095 , R_13615_12084c58 );
buf ( n4096 , R_14a29_10571438 );
buf ( n4097 , R_13526_102f49a8 );
buf ( n4098 , R_11215_12075b18 );
buf ( n4099 , R_10e4c_13a169e8 );
buf ( n4100 , R_13d97_105651d8 );
buf ( n4101 , R_1b3_1379b348 );
buf ( n4102 , R_13fab_11538758 );
buf ( n4103 , R_10ff9_105aad78 );
buf ( n4104 , R_145c0_11cd7f68 );
buf ( n4105 , R_145fc_120476f8 );
buf ( n4106 , R_15c_137992c8 );
buf ( n4107 , R_67bc_13311028 );
buf ( n4108 , R_efc2_11cdefe8 );
buf ( n4109 , R_145cc_132f8388 );
buf ( n4110 , R_ae_1379c1a8 );
buf ( n4111 , R_1263c_11cdf768 );
buf ( n4112 , R_57_126522e8 );
buf ( n4113 , R_14659_1264e1e8 );
buf ( n4114 , R_13899_133075c8 );
buf ( n4115 , R_125e5_13311348 );
buf ( n4116 , R_113fb_11ce7288 );
buf ( n4117 , R_11e0e_102f4908 );
buf ( n4118 , R_11270_12b29a58 );
buf ( n4119 , R_f61a_13305cc8 );
buf ( n4120 , R_1499f_133198c8 );
buf ( n4121 , R_121_13795808 );
buf ( n4122 , R_106_12b25a98 );
buf ( n4123 , R_1458a_102eb268 );
buf ( n4124 , R_126cf_13a19788 );
buf ( n4125 , R_209_1379cb08 );
buf ( n4126 , R_1ee_12656268 );
buf ( n4127 , R_12c5a_102ef688 );
buf ( n4128 , R_1270e_11cdb708 );
buf ( n4129 , R_e437_102f2c48 );
buf ( n4130 , R_147cf_11ce5168 );
buf ( n4131 , R_e233_1056d338 );
buf ( n4132 , R_13bbe_11ce55c8 );
buf ( n4133 , R_11e6b_1207d458 );
buf ( n4134 , R_13f0b_12b42f18 );
buf ( n4135 , R_103_12b41c58 );
buf ( n4136 , R_cd_12b39a58 );
buf ( n4137 , R_242_12654688 );
buf ( n4138 , R_20c_12b43c38 );
buf ( n4139 , R_11ce5_1379e048 );
buf ( n4140 , R_ef4_1056dc98 );
buf ( n4141 , R_11823_13a15fe8 );
buf ( n4142 , R_130b8_13a12988 );
buf ( n4143 , R_12baf_12648ba8 );
buf ( n4144 , R_119a4_102f3288 );
buf ( n4145 , R_f4e5_1264b308 );
buf ( n4146 , R_12c6f_11cdea48 );
buf ( n4147 , R_1473b_102fa308 );
buf ( n4148 , R_8b_132f8608 );
buf ( n4149 , R_11467_105659f8 );
buf ( n4150 , R_11b4a_11ce1568 );
buf ( n4151 , R_137f7_12077878 );
buf ( n4152 , R_e5b5_1153d938 );
buf ( n4153 , R_14775_13a1bda8 );
buf ( n4154 , R_14671_1264ab88 );
buf ( n4155 , R_14066_12084258 );
buf ( n4156 , R_13954_12076518 );
buf ( n4157 , R_de4d_12b26538 );
buf ( n4158 , R_149f6_11cda308 );
buf ( n4159 , R_aff6_102f4a48 );
buf ( n4160 , R_d75d_1207c0f8 );
buf ( n4161 , R_10f46_12081ff8 );
buf ( n4162 , R_c50b_11cdd3c8 );
buf ( n4163 , R_136ed_12082ef8 );
buf ( n4164 , R_101d1_1056e198 );
buf ( n4165 , R_1a9_12037658 );
buf ( n4166 , R_166_120507f8 );
buf ( n4167 , R_9b_12b3b178 );
buf ( n4168 , R_bb16_12650268 );
buf ( n4169 , R_1265a_105635b8 );
buf ( n4170 , R_b802_1265dba8 );
buf ( n4171 , R_131ea_102f4cc8 );
buf ( n4172 , R_14a0e_10570e98 );
buf ( n4173 , R_19a_12662068 );
buf ( n4174 , R_175_12b3fc78 );
buf ( n4175 , R_109_12b2c7f8 );
buf ( n4176 , R_206_105b5b38 );
buf ( n4177 , R_146b4_1153fcd8 );
buf ( n4178 , R_11e21_11cd9e08 );
buf ( n4179 , R_104ba_f8c7218 );
buf ( n4180 , R_13fbc_11541218 );
buf ( n4181 , R_144ba_102f8c88 );
buf ( n4182 , R_11622_102ed388 );
buf ( n4183 , R_13c02_12b29198 );
buf ( n4184 , R_13ba3_105626b8 );
buf ( n4185 , R_ff0f_12081918 );
buf ( n4186 , R_123d6_11541e98 );
buf ( n4187 , R_fd64_102f3328 );
buf ( n4188 , R_14486_102ef728 );
buf ( n4189 , R_13776_1379fd08 );
buf ( n4190 , R_14665_132f5ae8 );
buf ( n4191 , R_10098_13793968 );
buf ( n4192 , R_11072_13a1ed28 );
buf ( n4193 , R_14554_10565778 );
buf ( n4194 , R_137a8_1056b678 );
buf ( n4195 , R_11b55_12649a08 );
buf ( n4196 , R_14411_12663508 );
buf ( n4197 , R_84a7_12b40fd8 );
buf ( n4198 , R_133fc_1153ee78 );
buf ( n4199 , R_da_1331b088 );
buf ( n4200 , R_a0_1379b2a8 );
buf ( n4201 , R_235_1264d4c8 );
buf ( n4202 , R_1333b_11542c58 );
buf ( n4203 , R_132e7_11ce28c8 );
buf ( n4204 , R_1357d_1153feb8 );
buf ( n4205 , R_14644_1056d978 );
buf ( n4206 , R_100_1265f0e8 );
buf ( n4207 , R_79_137a1388 );
buf ( n4208 , R_e0d7_126556c8 );
buf ( n4209 , R_11b42_1264b6c8 );
buf ( n4210 , R_20f_12b28018 );
buf ( n4211 , R_f4db_1207bfb8 );
buf ( n4212 , R_1193e_13a19968 );
buf ( n4213 , R_138d5_1379b848 );
buf ( n4214 , R_13e4c_1207f118 );
buf ( n4215 , R_13a7e_102f6ac8 );
buf ( n4216 , R_12d79_102ee468 );
buf ( n4217 , R_116a8_12084398 );
buf ( n4218 , R_116_1265f868 );
buf ( n4219 , R_148a3_11cdecc8 );
buf ( n4220 , R_13273_13a1a688 );
buf ( n4221 , R_1f9_1379ddc8 );
buf ( n4222 , R_1025b_1330bee8 );
buf ( n4223 , R_122e8_12b39878 );
buf ( n4224 , R_11ba2_11544738 );
buf ( n4225 , R_12521_1056c258 );
buf ( n4226 , R_e8e6_f8cf4b8 );
buf ( n4227 , R_8cd2_1264ac28 );
buf ( n4228 , R_11a11_126477a8 );
buf ( n4229 , R_143c6_120850b8 );
buf ( n4230 , R_13e99_12039e58 );
buf ( n4231 , R_1466b_13306808 );
buf ( n4232 , R_14465_1207a758 );
buf ( n4233 , R_134b3_102f3468 );
buf ( n4234 , R_11fe7_1330c3e8 );
buf ( n4235 , R_1258d_13a14dc8 );
buf ( n4236 , R_14677_105712f8 );
buf ( n4237 , R_1367d_102eb628 );
buf ( n4238 , R_1e2_12663c88 );
buf ( n4239 , R_b9_12661848 );
buf ( n4240 , R_12d_12660268 );
buf ( n4241 , R_f47c_1153ded8 );
buf ( n4242 , R_1468c_13a1aae8 );
buf ( n4243 , R_145ba_120815f8 );
buf ( n4244 , R_14790_11cd9cc8 );
buf ( n4245 , R_14419_12048f58 );
buf ( n4246 , R_13bb3_1207b6f8 );
buf ( n4247 , R_1046b_105688d8 );
buf ( n4248 , R_1232e_13314008 );
buf ( n4249 , R_1170d_1264c528 );
buf ( n4250 , R_14a41_1056fa98 );
buf ( n4251 , R_14459_11cd92c8 );
buf ( n4252 , R_14480_11cdcf68 );
buf ( n4253 , R_13a88_11ce3f48 );
buf ( n4254 , R_c8f0_102f0d08 );
buf ( n4255 , R_134ff_1056bf38 );
buf ( n4256 , R_aac5_13a18748 );
buf ( n4257 , R_14509_13a1e148 );
buf ( n4258 , R_cebc_12039d18 );
buf ( n4259 , R_135bd_12081058 );
buf ( n4260 , R_147ba_12078ef8 );
buf ( n4261 , R_f4a6_105654f8 );
buf ( n4262 , R_1182e_13a19aa8 );
buf ( n4263 , R_142eb_11cdec28 );
buf ( n4264 , R_13bf5_10568ab8 );
buf ( n4265 , R_12093_12077058 );
buf ( n4266 , R_13dac_13a15688 );
buf ( n4267 , R_dc51_13304f08 );
buf ( n4268 , R_13e8f_1264a0e8 );
buf ( n4269 , R_13c89_12b39f58 );
buf ( n4270 , R_f0be_102f1de8 );
buf ( n4271 , R_9373_10563e78 );
buf ( n4272 , R_11a48_13a195a8 );
buf ( n4273 , R_f3f9_1153f9b8 );
buf ( n4274 , R_1d4_12b42fb8 );
buf ( n4275 , R_e3f1_12b25bd8 );
buf ( n4276 , R_13c27_13309b48 );
buf ( n4277 , R_240_105ab4f8 );
buf ( n4278 , R_cf_13311a28 );
buf ( n4279 , R_13c38_1204a3f8 );
buf ( n4280 , R_13b_13300f88 );
buf ( n4281 , R_11ef6_11cd7888 );
buf ( n4282 , R_135c9_11ce6888 );
buf ( n4283 , R_116d1_1153d898 );
buf ( n4284 , R_149d2_12080158 );
buf ( n4285 , R_ba5b_12b403f8 );
buf ( n4286 , R_ea84_1330ca28 );
buf ( n4287 , R_f59a_11ce3908 );
buf ( n4288 , R_1496c_1331e968 );
buf ( n4289 , R_12bd5_11ce3fe8 );
buf ( n4290 , R_1253e_105b6678 );
buf ( n4291 , R_14873_11cd79c8 );
buf ( n4292 , R_149a5_132ff868 );
buf ( n4293 , R_14512_11540bd8 );
buf ( n4294 , R_14756_10565318 );
buf ( n4295 , R_1c9_13313a68 );
buf ( n4296 , R_d09b_12660948 );
buf ( n4297 , R_203_12050cf8 );
buf ( n4298 , R_10c_12038058 );
buf ( n4299 , R_146_12b42298 );
buf ( n4300 , R_136c1_12b276b8 );
buf ( n4301 , R_1480a_12649e68 );
buf ( n4302 , R_1d9_1379e7c8 );
buf ( n4303 , R_13e84_1056ad18 );
buf ( n4304 , R_1021c_1056fc78 );
buf ( n4305 , R_136_132fe6e8 );
buf ( n4306 , R_145ff_102ef2c8 );
buf ( n4307 , R_19b_12b28dd8 );
buf ( n4308 , R_1031a_11540e58 );
buf ( n4309 , R_1f2_11538438 );
buf ( n4310 , R_13114_102f3648 );
buf ( n4311 , R_ec36_12042af8 );
buf ( n4312 , R_222_133189c8 );
buf ( n4313 , R_6f_12b3a458 );
buf ( n4314 , R_96_1203c838 );
buf ( n4315 , R_ed_1203deb8 );
buf ( n4316 , R_11d_1204c838 );
buf ( n4317 , R_174_13318928 );
buf ( n4318 , R_119f1_13316588 );
buf ( n4319 , R_1486a_13a1d428 );
buf ( n4320 , R_11717_1207d778 );
buf ( n4321 , R_14781_115447d8 );
buf ( n4322 , R_13995_12038738 );
buf ( n4323 , R_e4f5_12049598 );
buf ( n4324 , R_74a9_12645d68 );
buf ( n4325 , R_10208_12038558 );
buf ( n4326 , R_145ab_12b3f9f8 );
buf ( n4327 , R_227_1331e508 );
buf ( n4328 , R_e8_133028e8 );
buf ( n4329 , R_13809_1153faf8 );
buf ( n4330 , R_f732_12649008 );
buf ( n4331 , R_14524_137968e8 );
buf ( n4332 , R_146d8_11cd94a8 );
buf ( n4333 , R_14064_1264d2e8 );
buf ( n4334 , R_12dfa_11cd88c8 );
buf ( n4335 , R_135ef_102f0a88 );
buf ( n4336 , R_10ee5_12047798 );
buf ( n4337 , R_14548_120493b8 );
buf ( n4338 , R_11030_11cdbca8 );
buf ( n4339 , R_1400f_13a1a368 );
buf ( n4340 , R_f051_1264e6e8 );
buf ( n4341 , R_de7c_102eafe8 );
buf ( n4342 , R_13538_120754d8 );
buf ( n4343 , R_13e56_12b297d8 );
buf ( n4344 , R_84eb_1331c2a8 );
buf ( n4345 , R_1498a_1207e3f8 );
buf ( n4346 , R_148a6_115459f8 );
buf ( n4347 , R_212_1330bd08 );
buf ( n4348 , R_fd_13307d48 );
buf ( n4349 , R_144a5_13a1c028 );
buf ( n4350 , R_10110_120369d8 );
buf ( n4351 , R_12b5e_12651208 );
buf ( n4352 , R_149ed_13303428 );
buf ( n4353 , R_144db_12078598 );
buf ( n4354 , R_bf9f_11cd9b88 );
buf ( n4355 , R_14017_f8c20d8 );
buf ( n4356 , R_13a3d_f8ca918 );
buf ( n4357 , R_13b2d_120830d8 );
buf ( n4358 , R_8e_132f37e8 );
buf ( n4359 , R_12aeb_120810f8 );
buf ( n4360 , R_a23e_11ce5ca8 );
buf ( n4361 , R_12ce9_12081c38 );
buf ( n4362 , R_f00_1207c058 );
buf ( n4363 , R_c1fe_1264be48 );
buf ( n4364 , R_f2d2_11cdf948 );
buf ( n4365 , R_14385_12044c18 );
buf ( n4366 , R_143c0_1265fb88 );
buf ( n4367 , R_14496_13a1c668 );
buf ( n4368 , R_14738_12b28bf8 );
buf ( n4369 , R_cab9_102f99a8 );
buf ( n4370 , R_1255c_f8c61d8 );
buf ( n4371 , R_143ba_11cde868 );
buf ( n4372 , R_147c9_13a18ce8 );
buf ( n4373 , R_13311_13a198c8 );
buf ( n4374 , R_147a2_102f2ce8 );
buf ( n4375 , R_fbe0_13a1b628 );
buf ( n4376 , R_dcc6_12664ae8 );
buf ( n4377 , R_103cf_12085158 );
buf ( n4378 , R_13909_1204f5d8 );
buf ( n4379 , R_1197b_115433d8 );
buf ( n4380 , R_144e1_13a1f4a8 );
buf ( n4381 , R_145a2_11cd7ce8 );
buf ( n4382 , R_12d50_120851f8 );
buf ( n4383 , R_12380_10563338 );
buf ( n4384 , R_107a7_1379f9e8 );
buf ( n4385 , R_10e8a_102ea688 );
buf ( n4386 , R_122fb_13a17708 );
buf ( n4387 , R_12aa7_12037798 );
buf ( n4388 , R_12107_1264d428 );
buf ( n4389 , R_14533_1330c8e8 );
buf ( n4390 , R_14542_120759d8 );
buf ( n4391 , R_4276_102effe8 );
buf ( n4392 , R_1478d_115453b8 );
buf ( n4393 , R_130c1_11542258 );
buf ( n4394 , R_13ff8_102f9fe8 );
buf ( n4395 , R_1aa_13795268 );
buf ( n4396 , R_116b1_13a159a8 );
buf ( n4397 , R_1bc_126536e8 );
buf ( n4398 , R_b76e_1153c8f8 );
buf ( n4399 , R_4e_13792e28 );
buf ( n4400 , R_60_12b44bd8 );
buf ( n4401 , R_a5_13311668 );
buf ( n4402 , R_b7_1379f948 );
buf ( n4403 , R_153_13793288 );
buf ( n4404 , R_165_13306948 );
buf ( n4405 , R_f9fe_102f9408 );
buf ( n4406 , R_14431_12080478 );
buf ( n4407 , R_1c3_12047158 );
buf ( n4408 , R_64_f8c1bd8 );
buf ( n4409 , R_14c_120387d8 );
buf ( n4410 , R_12471_102f7068 );
buf ( n4411 , R_148c1_13316f88 );
buf ( n4412 , R_11433_1265f048 );
buf ( n4413 , R_13ce2_1264aa48 );
buf ( n4414 , R_121bd_115449b8 );
buf ( n4415 , R_14813_10566d58 );
buf ( n4416 , R_147fb_102f83c8 );
buf ( n4417 , R_146ab_12051658 );
buf ( n4418 , R_12c65_1264cb68 );
buf ( n4419 , R_e2b4_f8c0f58 );
buf ( n4420 , R_10c61_120805b8 );
buf ( n4421 , R_10f1d_10566df8 );
buf ( n4422 , R_10de4_1379b5c8 );
buf ( n4423 , R_ae51_105ab098 );
buf ( n4424 , R_146f3_12659d28 );
buf ( n4425 , R_d03f_126484c8 );
buf ( n4426 , R_9fe2_11543fb8 );
buf ( n4427 , R_10b79_12657028 );
buf ( n4428 , R_64c2_12662748 );
buf ( n4429 , R_139d0_102f1fc8 );
buf ( n4430 , R_13639_1207f578 );
buf ( n4431 , R_1b4_12654728 );
buf ( n4432 , R_1cf_133184c8 );
buf ( n4433 , R_e214_1207ae38 );
buf ( n4434 , R_140_12665448 );
buf ( n4435 , R_15b_f8c0378 );
buf ( n4436 , R_1435c_13304d28 );
buf ( n4437 , R_10745_12056898 );
buf ( n4438 , R_1044f_120557f8 );
buf ( n4439 , R_10824_11ce3188 );
buf ( n4440 , R_13820_12b41438 );
buf ( n4441 , R_69b8_11cdc888 );
buf ( n4442 , R_124b9_1056d658 );
buf ( n4443 , R_143f4_102edd88 );
buf ( n4444 , R_142f5_1264a908 );
buf ( n4445 , R_76_f8ca198 );
buf ( n4446 , R_ac_12660a88 );
buf ( n4447 , R_1269b_11cd9368 );
buf ( n4448 , R_147b4_120766f8 );
buf ( n4449 , R_14834_13a16a88 );
buf ( n4450 , R_12e88_102f8a08 );
buf ( n4451 , R_f021_102ec168 );
buf ( n4452 , R_f6dd_13a163a8 );
buf ( n4453 , R_145e4_126463a8 );
buf ( n4454 , R_14723_1264db08 );
buf ( n4455 , R_173_f8c3438 );
buf ( n4456 , R_19c_12b40218 );
buf ( n4457 , R_11142_10562f78 );
buf ( n4458 , R_23e_1265bc68 );
buf ( n4459 , R_d1_13311f28 );
buf ( n4460 , R_13512_12080dd8 );
buf ( n4461 , R_7859_11cdaee8 );
buf ( n4462 , R_14593_115458b8 );
buf ( n4463 , R_148a9_12647ac8 );
buf ( n4464 , R_10577_11545318 );
buf ( n4465 , R_133ca_1203e098 );
buf ( n4466 , R_13b92_13a14be8 );
buf ( n4467 , R_10efd_102ec3e8 );
buf ( n4468 , R_f0b_1153f4b8 );
buf ( n4469 , R_12e15_10568018 );
buf ( n4470 , R_200_12b29eb8 );
buf ( n4471 , R_21d_137a03e8 );
buf ( n4472 , R_f2_12652ec8 );
buf ( n4473 , R_10f_12b3e5f8 );
buf ( n4474 , R_ca13_11ce4628 );
buf ( n4475 , R_14966_11546218 );
buf ( n4476 , R_13ad8_1203a358 );
buf ( n4477 , R_12d8d_105b5db8 );
buf ( n4478 , R_10165_1264cac8 );
buf ( n4479 , R_1337f_13a12c08 );
buf ( n4480 , R_53_f8c2a38 );
buf ( n4481 , R_149c9_132f4fa8 );
buf ( n4482 , R_10aae_1207c558 );
buf ( n4483 , R_13aad_11541a38 );
buf ( n4484 , R_12362_10563dd8 );
buf ( n4485 , R_5c4e_1056ced8 );
buf ( n4486 , R_130f5_1056a098 );
buf ( n4487 , R_12a7c_11cdde68 );
buf ( n4488 , R_14415_12b2a318 );
buf ( n4489 , R_1488b_13a189c8 );
buf ( n4490 , R_14062_1204cf18 );
buf ( n4491 , R_14784_11cd8508 );
buf ( n4492 , R_1032f_10570f38 );
buf ( n4493 , R_9bdf_102ee5a8 );
buf ( n4494 , R_13bf0_1331c528 );
buf ( n4495 , R_11b90_11ce0208 );
buf ( n4496 , R_149cf_13a17b68 );
buf ( n4497 , R_12021_11ce25a8 );
buf ( n4498 , R_1de_12056d98 );
buf ( n4499 , R_49_1331f4a8 );
buf ( n4500 , R_131_105ab3b8 );
buf ( n4501 , R_1462f_13794688 );
buf ( n4502 , R_10628_1203d2d8 );
buf ( n4503 , R_122bf_10570038 );
buf ( n4504 , R_11387_11540d18 );
buf ( n4505 , R_11fa6_13306308 );
buf ( n4506 , R_85b5_120819b8 );
buf ( n4507 , R_142ef_102eec88 );
buf ( n4508 , R_1434c_102f13e8 );
buf ( n4509 , R_22c_1379b708 );
buf ( n4510 , R_5c_137944a8 );
buf ( n4511 , R_e3_1203e778 );
buf ( n4512 , R_b948_1153a5f8 );
buf ( n4513 , R_e169_11cd7a68 );
buf ( n4514 , R_d051_11536ef8 );
buf ( n4515 , R_10e01_120551b8 );
buf ( n4516 , R_233_12b392d8 );
buf ( n4517 , R_68_12b283d8 );
buf ( n4518 , R_dc_13300768 );
buf ( n4519 , R_13bfb_13316a88 );
buf ( n4520 , R_10ad6_10565598 );
buf ( n4521 , R_14870_10570538 );
buf ( n4522 , R_12260_13a1b268 );
buf ( n4523 , R_d661_1265cfc8 );
buf ( n4524 , R_14572_11cd9d68 );
buf ( n4525 , R_130ff_12078318 );
buf ( n4526 , R_a98a_11cdaf88 );
buf ( n4527 , R_14978_12b321f8 );
buf ( n4528 , R_14a1a_115445f8 );
buf ( n4529 , R_14a26_13792568 );
buf ( n4530 , R_b327_12648568 );
buf ( n4531 , R_108fb_105b5e58 );
buf ( n4532 , R_1440d_11544238 );
buf ( n4533 , R_10cff_13a1dc48 );
buf ( n4534 , R_139ae_11cd8b48 );
buf ( n4535 , R_14338_11cda808 );
buf ( n4536 , R_106b3_13a16088 );
buf ( n4537 , R_c4f8_11ce12e8 );
buf ( n4538 , R_215_1265b948 );
buf ( n4539 , R_fa_133070c8 );
buf ( n4540 , R_11b68_1264ec88 );
buf ( n4541 , R_129b1_1056f098 );
buf ( n4542 , R_13670_10564558 );
buf ( n4543 , R_1439c_11cdd148 );
buf ( n4544 , R_107e6_11cdbc08 );
buf ( n4545 , R_f279_13a1acc8 );
buf ( n4546 , R_12ed9_102edf68 );
buf ( n4547 , R_12bc1_13a1f048 );
buf ( n4548 , R_13b19_12b2ba38 );
buf ( n4549 , R_e361_120812d8 );
buf ( n4550 , R_bef9_11ce0528 );
buf ( n4551 , R_13ce8_120793f8 );
buf ( n4552 , R_a235_12084a78 );
buf ( n4553 , R_14521_1264f228 );
buf ( n4554 , R_13cad_13a1edc8 );
buf ( n4555 , R_148af_11540098 );
buf ( n4556 , R_10968_13304968 );
buf ( n4557 , R_13fcb_102f0c68 );
buf ( n4558 , R_11645_13304e68 );
buf ( n4559 , R_bf09_1056b498 );
buf ( n4560 , R_12553_13310308 );
buf ( n4561 , R_145d5_132fa228 );
buf ( n4562 , R_146a2_1207bf18 );
buf ( n4563 , R_136fc_12076018 );
buf ( n4564 , R_149a2_1264d1a8 );
buf ( n4565 , R_12b9a_13a14968 );
buf ( n4566 , R_137cc_10569af8 );
buf ( n4567 , R_c5ef_12081238 );
buf ( n4568 , R_1184d_11cd9188 );
buf ( n4569 , R_13c8f_102ed568 );
buf ( n4570 , R_109bf_1379c248 );
buf ( n4571 , R_14326_13301528 );
buf ( n4572 , R_11123_12045258 );
buf ( n4573 , R_e197_11ce3228 );
buf ( n4574 , R_172_126656c8 );
buf ( n4575 , R_19d_132ffb88 );
buf ( n4576 , R_c306_f8c5418 );
buf ( n4577 , R_b5_133157c8 );
buf ( n4578 , R_13902_13799ae8 );
buf ( n4579 , R_14348_1056c398 );
buf ( n4580 , R_1457b_102f5628 );
buf ( n4581 , R_14766_105674d8 );
buf ( n4582 , R_d2c1_12036e38 );
buf ( n4583 , R_1f6_1330dce8 );
buf ( n4584 , R_10c28_12080e78 );
buf ( n4585 , R_119_133166c8 );
buf ( n4586 , R_1300e_12646bc8 );
buf ( n4587 , R_13129_10567b18 );
buf ( n4588 , R_1394d_1056f318 );
buf ( n4589 , R_14846_13798b48 );
buf ( n4590 , R_146cf_1379e868 );
buf ( n4591 , R_10019_11542118 );
buf ( n4592 , R_fb35_132fb4e8 );
buf ( n4593 , R_11a23_126506c8 );
buf ( n4594 , R_9aae_1056dbf8 );
buf ( n4595 , R_14468_1264aea8 );
buf ( n4596 , R_7aaf_f8c22b8 );
buf ( n4597 , R_b5af_1264e508 );
buf ( n4598 , R_13f11_11cd7b08 );
buf ( n4599 , R_e6c6_12075cf8 );
buf ( n4600 , R_14374_102f0768 );
buf ( n4601 , R_14605_13a182e8 );
buf ( n4602 , R_13de4_102f94a8 );
buf ( n4603 , R_102c2_1264ed28 );
buf ( n4604 , R_91_13799548 );
buf ( n4605 , R_135f5_11cda4e8 );
buf ( n4606 , R_14807_1331e288 );
buf ( n4607 , R_14a08_11cdc388 );
buf ( n4608 , R_cb44_12b3ee18 );
buf ( n4609 , R_13a63_11544198 );
buf ( n4610 , R_109ca_1264cd48 );
buf ( n4611 , R_12e41_10569198 );
buf ( n4612 , R_e46a_13a181a8 );
buf ( n4613 , R_12963_13a1afe8 );
buf ( n4614 , R_14a5a_12b42158 );
buf ( n4615 , R_13e38_1207efd8 );
buf ( n4616 , R_144ea_1264f5e8 );
buf ( n4617 , R_11668_137a1d88 );
buf ( n4618 , R_13ec7_11540318 );
buf ( n4619 , R_ff67_13799688 );
buf ( n4620 , R_13b27_102eb588 );
buf ( n4621 , R_fa2a_1056e0f8 );
buf ( n4622 , R_145a5_132f4dc8 );
buf ( n4623 , R_14060_13a15ae8 );
buf ( n4624 , R_164_12b27118 );
buf ( n4625 , R_104d9_120779b8 );
buf ( n4626 , R_1ab_f8c2998 );
buf ( n4627 , R_23c_13319328 );
buf ( n4628 , R_bbdf_133063a8 );
buf ( n4629 , R_d3_12659968 );
buf ( n4630 , R_cc7b_13a1b128 );
buf ( n4631 , R_12ffe_1331cd48 );
buf ( n4632 , R_1323e_126561c8 );
buf ( n4633 , R_1207f_133190a8 );
buf ( n4634 , R_10f99_126549a8 );
buf ( n4635 , R_913d_12646b28 );
buf ( n4636 , R_c3ee_102f6848 );
buf ( n4637 , R_13b12_13a1a728 );
buf ( n4638 , R_10a0c_11cdf1c8 );
buf ( n4639 , R_13974_13a19008 );
buf ( n4640 , R_13602_126635a8 );
buf ( n4641 , R_124e1_11cdb668 );
buf ( n4642 , R_142d7_12b30d58 );
buf ( n4643 , R_14960_105b5598 );
buf ( n4644 , R_f86d_120385f8 );
buf ( n4645 , R_148a0_12b38ab8 );
buf ( n4646 , R_e63f_f8cb9f8 );
buf ( n4647 , R_12741_105642d8 );
buf ( n4648 , R_684e_1056aa98 );
buf ( n4649 , R_13b04_12081558 );
buf ( n4650 , R_1453f_11ce2328 );
buf ( n4651 , R_148b5_1207f898 );
buf ( n4652 , R_1499c_12080658 );
buf ( n4653 , R_128e2_12647668 );
buf ( n4654 , R_13345_11ce0988 );
buf ( n4655 , R_cd4f_102f2f68 );
buf ( n4656 , R_13dd3_1204cd38 );
buf ( n4657 , R_13ea4_11ce0708 );
buf ( n4658 , R_f16b_11cda448 );
buf ( n4659 , R_139fe_1153e5b8 );
buf ( n4660 , R_12eed_102ee1e8 );
buf ( n4661 , R_13479_13306b28 );
buf ( n4662 , R_1135b_1056d158 );
buf ( n4663 , R_131a5_1153dc58 );
buf ( n4664 , R_14744_1264b3a8 );
buf ( n4665 , R_144c6_1056d5b8 );
buf ( n4666 , R_13109_f8c4798 );
buf ( n4667 , R_137bb_10564058 );
buf ( n4668 , R_146db_1056a818 );
buf ( n4669 , R_119c2_13a1a548 );
buf ( n4670 , R_eb5e_1056d018 );
buf ( n4671 , R_b0d7_1153e3d8 );
buf ( n4672 , R_13b9e_12083038 );
buf ( n4673 , R_1116a_13a15868 );
buf ( n4674 , R_12a65_10564c38 );
buf ( n4675 , R_14969_11cdb2a8 );
buf ( n4676 , R_1464d_12075618 );
buf ( n4677 , R_e3c5_12080a18 );
buf ( n4678 , R_1469c_120511f8 );
buf ( n4679 , R_d50f_12663828 );
buf ( n4680 , R_137f0_12079358 );
buf ( n4681 , R_11593_1207a258 );
buf ( n4682 , R_14350_1207d8b8 );
buf ( n4683 , R_cbe2_11536a98 );
buf ( n4684 , R_110ed_10563d38 );
buf ( n4685 , R_1125d_102f86e8 );
buf ( n4686 , R_13c09_11ce4268 );
buf ( n4687 , R_135fc_13795948 );
buf ( n4688 , R_14557_11cdcec8 );
buf ( n4689 , R_112_13312248 );
buf ( n4690 , R_1fd_133221a8 );
buf ( n4691 , R_9e_11539838 );
buf ( n4692 , R_143b2_11cddd28 );
buf ( n4693 , R_12fec_102efea8 );
buf ( n4694 , R_c4d7_13a1f408 );
buf ( n4695 , R_1398e_13320bc8 );
buf ( n4696 , R_12894_11ce1428 );
buf ( n4697 , R_b6f4_102f9ea8 );
buf ( n4698 , R_fcb3_12649be8 );
buf ( n4699 , R_12375_1207edf8 );
buf ( n4700 , R_146b1_102ed248 );
buf ( n4701 , R_11b11_11545818 );
buf ( n4702 , R_58_13317a28 );
buf ( n4703 , R_73_12b3e0f8 );
buf ( n4704 , R_bd7c_11ce2be8 );
buf ( n4705 , R_12fd8_10565278 );
buf ( n4706 , R_14876_12054678 );
buf ( n4707 , R_138da_1153dbb8 );
buf ( n4708 , R_14825_12647168 );
buf ( n4709 , R_14a4d_12646ee8 );
buf ( n4710 , R_124_1203edb8 );
buf ( n4711 , R_15a_f8c6958 );
buf ( n4712 , R_1b5_1331afe8 );
buf ( n4713 , R_1eb_12038d78 );
buf ( n4714 , R_1475d_11546038 );
buf ( n4715 , R_171_105aa5f8 );
buf ( n4716 , R_106ea_102f6528 );
buf ( n4717 , R_19e_1331e788 );
buf ( n4718 , R_11a86_1204ffd8 );
buf ( n4719 , R_fad7_102f5ee8 );
buf ( n4720 , R_e21e_1056b7b8 );
buf ( n4721 , R_12933_11cd7c48 );
buf ( n4722 , R_6c_12040938 );
buf ( n4723 , R_99_12b27618 );
buf ( n4724 , R_1353d_1153d9d8 );
buf ( n4725 , R_b283_1330acc8 );
buf ( n4726 , R_143ae_13a1cca8 );
buf ( n4727 , R_14801_11540c78 );
buf ( n4728 , R_149e7_10568298 );
buf ( n4729 , R_14708_1203c018 );
buf ( n4730 , R_14450_13a17028 );
buf ( n4731 , R_128_12b43b98 );
buf ( n4732 , R_145_1265aa48 );
buf ( n4733 , R_1ca_1265ff48 );
buf ( n4734 , R_1e7_12b3d798 );
buf ( n4735 , R_7741_13a16128 );
buf ( n4736 , R_da39_12b40718 );
buf ( n4737 , R_e38d_12651168 );
buf ( n4738 , R_12fc4_11544878 );
buf ( n4739 , R_145e7_11544058 );
buf ( n4740 , R_1465f_105676b8 );
buf ( n4741 , R_10fc1_12078638 );
buf ( n4742 , R_704f_11ce4da8 );
buf ( n4743 , R_13a8d_13318108 );
buf ( n4744 , R_145c3_1264da68 );
buf ( n4745 , R_faad_13a1fd68 );
buf ( n4746 , R_12738_10570678 );
buf ( n4747 , R_11935_13a1ff48 );
buf ( n4748 , R_11720_1330eaa8 );
buf ( n4749 , R_d16a_11ce5de8 );
buf ( n4750 , R_13e0d_13a1b4e8 );
buf ( n4751 , R_1447d_11ce3a48 );
buf ( n4752 , R_152_12b3c4d8 );
buf ( n4753 , R_105ba_13306bc8 );
buf ( n4754 , R_b1aa_12649468 );
buf ( n4755 , R_1bd_12653be8 );
buf ( n4756 , R_14a50_13a161c8 );
buf ( n4757 , R_13a83_10567a78 );
buf ( n4758 , R_123c2_13797108 );
buf ( n4759 , R_144b7_13305d68 );
buf ( n4760 , R_13814_137926a8 );
buf ( n4761 , R_12cbd_13a14328 );
buf ( n4762 , R_11bab_120768d8 );
buf ( n4763 , R_c07e_13a18b08 );
buf ( n4764 , R_142f9_11545e58 );
buf ( n4765 , R_1478a_12652928 );
buf ( n4766 , R_14a3b_11ce2d28 );
buf ( n4767 , R_c3a2_13a19508 );
buf ( n4768 , R_aa_126535a8 );
buf ( n4769 , R_146e7_10566538 );
buf ( n4770 , R_138fb_12082778 );
buf ( n4771 , R_13988_133186a8 );
buf ( n4772 , R_13c43_1264cca8 );
buf ( n4773 , R_14590_132f3b08 );
buf ( n4774 , R_110cf_137940e8 );
buf ( n4775 , R_13326_12648d88 );
buf ( n4776 , R_13153_10567118 );
buf ( n4777 , R_1405e_f8c95b8 );
buf ( n4778 , R_1051f_13793b48 );
buf ( n4779 , R_f518_12075bb8 );
buf ( n4780 , R_143a2_12079038 );
buf ( n4781 , R_147a8_12657de8 );
buf ( n4782 , R_13cb3_102f6fc8 );
buf ( n4783 , R_10c3d_f8c5b98 );
buf ( n4784 , R_e7ab_1264f7c8 );
buf ( n4785 , R_13449_12077378 );
buf ( n4786 , R_14403_12b29418 );
buf ( n4787 , R_148b2_132fc708 );
buf ( n4788 , R_1468f_10562cf8 );
buf ( n4789 , R_f7_13309828 );
buf ( n4790 , R_13f54_102f4e08 );
buf ( n4791 , R_218_12050258 );
buf ( n4792 , R_83_1379cd88 );
buf ( n4793 , R_12f16_137a0b68 );
buf ( n4794 , R_10598_102ead68 );
buf ( n4795 , R_10365_12051478 );
buf ( n4796 , R_13ab4_13a12ca8 );
buf ( n4797 , R_13393_10568a18 );
buf ( n4798 , R_13683_1207cf58 );
buf ( n4799 , R_13a_105ac2b8 );
buf ( n4800 , R_127d5_11cdf268 );
buf ( n4801 , R_11917_11ce1248 );
buf ( n4802 , R_1d5_1265e468 );
buf ( n4803 , R_12e98_1204e778 );
buf ( n4804 , R_b3_12655ea8 );
buf ( n4805 , R_149cc_10564cd8 );
buf ( n4806 , R_134d9_10565f98 );
buf ( n4807 , R_fd0b_102ec488 );
buf ( n4808 , R_af25_133136a8 );
buf ( n4809 , R_11948_12b288d8 );
buf ( n4810 , R_149c6_1207b018 );
buf ( n4811 , R_14b_12b28a18 );
buf ( n4812 , R_1c4_12652e28 );
buf ( n4813 , R_10199_13a1f368 );
buf ( n4814 , R_80_12055438 );
buf ( n4815 , R_10b70_f8cd438 );
buf ( n4816 , R_10cdf_115401d8 );
buf ( n4817 , R_11a66_1207dc78 );
buf ( n4818 , R_132fc_13307708 );
buf ( n4819 , R_8c7b_12076b58 );
buf ( n4820 , R_1495a_1207a2f8 );
buf ( n4821 , R_1201a_10570218 );
buf ( n4822 , R_132d6_11ce0348 );
buf ( n4823 , R_14963_13304be8 );
buf ( n4824 , R_1285e_11545c78 );
buf ( n4825 , R_130de_102f58a8 );
buf ( n4826 , R_fb5f_13a1e288 );
buf ( n4827 , R_13ecf_1207c5f8 );
buf ( n4828 , R_1456f_13a1f5e8 );
buf ( n4829 , R_ea_1331a9a8 );
buf ( n4830 , R_120_12b400d8 );
buf ( n4831 , R_13eac_11ce2a08 );
buf ( n4832 , R_12568_1056b0d8 );
buf ( n4833 , R_e3ba_1207df98 );
buf ( n4834 , R_dcf2_12085298 );
buf ( n4835 , R_1ef_f8c2cb8 );
buf ( n4836 , R_225_12b3a318 );
buf ( n4837 , R_f7da_1204e9f8 );
buf ( n4838 , R_f857_13a13748 );
buf ( n4839 , R_1461a_13301988 );
buf ( n4840 , R_146b7_13a15228 );
buf ( n4841 , R_1384a_126503a8 );
buf ( n4842 , R_c8e7_105b6498 );
buf ( n4843 , R_86_137a1a68 );
buf ( n4844 , R_a3_126621a8 );
buf ( n4845 , R_f862_13a1a908 );
buf ( n4846 , R_10ab7_102f7b08 );
buf ( n4847 , R_11890_102eb308 );
buf ( n4848 , R_df3c_120774b8 );
buf ( n4849 , R_1369b_1330c2a8 );
buf ( n4850 , R_12e03_132ff368 );
buf ( n4851 , R_1356b_102f5da8 );
buf ( n4852 , R_10e42_1207e718 );
buf ( n4853 , R_10f59_f8c2c18 );
buf ( n4854 , R_127b6_12b412f8 );
buf ( n4855 , R_120e7_12b44818 );
buf ( n4856 , R_12492_1265b9e8 );
buf ( n4857 , R_10d12_13792b08 );
buf ( n4858 , R_130ae_12044b78 );
buf ( n4859 , R_13652_11ce1ce8 );
buf ( n4860 , R_117a7_12080fb8 );
buf ( n4861 , R_14674_13a13ba8 );
buf ( n4862 , R_11306_11540638 );
buf ( n4863 , R_d5_126617a8 );
buf ( n4864 , R_de_1265ce88 );
buf ( n4865 , R_12c_1379b488 );
buf ( n4866 , R_135_f8c6f98 );
buf ( n4867 , R_1da_12664b88 );
buf ( n4868 , R_1e3_1153c498 );
buf ( n4869 , R_122dd_13a1b6c8 );
buf ( n4870 , R_231_1379a6c8 );
buf ( n4871 , R_23a_12660b28 );
buf ( n4872 , R_1240e_13a150e8 );
buf ( n4873 , R_14686_13a137e8 );
buf ( n4874 , R_146c6_f8cf918 );
buf ( n4875 , R_13f5b_1207c738 );
buf ( n4876 , R_ebb7_102efd68 );
buf ( n4877 , R_1447a_105697d8 );
buf ( n4878 , R_13c95_12650ee8 );
buf ( n4879 , R_11de0_12083cb8 );
buf ( n4880 , R_11552_12648c48 );
buf ( n4881 , R_11cb2_1207ab18 );
buf ( n4882 , R_14849_11ce0028 );
buf ( n4883 , R_13f45_13a134c8 );
buf ( n4884 , R_13726_12084f78 );
buf ( n4885 , R_121f2_102f30a8 );
buf ( n4886 , R_ef_1379b0c8 );
buf ( n4887 , R_163_12b38a18 );
buf ( n4888 , R_1ac_12b29558 );
buf ( n4889 , R_220_12b25638 );
buf ( n4890 , R_14623_13a12a28 );
buf ( n4891 , R_1393a_11ce3408 );
buf ( n4892 , R_139ea_11cd8828 );
buf ( n4893 , R_cf49_11541718 );
buf ( n4894 , R_b889_1056a458 );
buf ( n4895 , R_1349f_1204fdf8 );
buf ( n4896 , R_170_120440d8 );
buf ( n4897 , R_19f_133087e8 );
buf ( n4898 , R_a9d8_102f22e8 );
buf ( n4899 , R_7d_12660308 );
buf ( n4900 , R_1460b_10569a58 );
buf ( n4901 , R_11983_13318568 );
buf ( n4902 , R_a6e4_13314648 );
buf ( n4903 , R_144b1_1207b478 );
buf ( n4904 , R_14614_12664f48 );
buf ( n4905 , R_139d7_132fda68 );
buf ( n4906 , R_ec64_11ce6248 );
buf ( n4907 , R_12d32_115454f8 );
buf ( n4908 , R_82bb_1204a678 );
buf ( n4909 , R_1472c_13a139c8 );
buf ( n4910 , R_144f7_10565e58 );
buf ( n4911 , R_10dad_12082f98 );
buf ( n4912 , R_b05c_1330b4e8 );
buf ( n4913 , R_13ef1_105714d8 );
buf ( n4914 , R_14635_12b3b038 );
buf ( n4915 , R_117b5_1056fdb8 );
buf ( n4916 , R_14692_11cdf128 );
buf ( n4917 , R_13f_1203dd78 );
buf ( n4918 , R_1055c_105672f8 );
buf ( n4919 , R_1d0_12040258 );
buf ( n4920 , R_13aba_1265cde8 );
buf ( n4921 , R_131e1_102f2ec8 );
buf ( n4922 , R_eb07_1153ef18 );
buf ( n4923 , R_9c9a_1056c578 );
buf ( n4924 , R_10605_11545d18 );
buf ( n4925 , R_13a97_12079218 );
buf ( n4926 , R_1331b_102efc28 );
buf ( n4927 , R_14879_11ce58e8 );
buf ( n4928 , R_14996_102eb3a8 );
buf ( n4929 , R_1405c_11ce34a8 );
buf ( n4930 , R_14945_1056e238 );
buf ( n4931 , R_b65f_11cdba28 );
buf ( n4932 , R_13f3e_13a1e508 );
buf ( n4933 , R_dbc0_132fb9e8 );
buf ( n4934 , R_1351c_13797068 );
buf ( n4935 , R_14804_120788b8 );
buf ( n4936 , R_14a0b_133206c8 );
buf ( n4937 , R_89_126595a8 );
buf ( n4938 , R_13c33_11ce3688 );
buf ( n4939 , R_4f_12b44d18 );
buf ( n4940 , R_cb5a_12b256d8 );
buf ( n4941 , R_13b85_10571258 );
buf ( n4942 , R_138f4_1330a9a8 );
buf ( n4943 , R_ee1a_1264fae8 );
buf ( n4944 , R_10411_102f8828 );
buf ( n4945 , R_14331_1056be98 );
buf ( n4946 , R_14717_1153a378 );
buf ( n4947 , R_94_1330ee68 );
buf ( n4948 , R_e5_1153cfd8 );
buf ( n4949 , R_22a_12b43698 );
buf ( n4950 , R_cba1_13a16e48 );
buf ( n4951 , R_129d1_12047978 );
buf ( n4952 , R_143d8_11cdc2e8 );
buf ( n4953 , R_13070_1264b268 );
buf ( n4954 , R_12915_1056d518 );
buf ( n4955 , R_12942_11cdd0a8 );
buf ( n4956 , R_145a8_12662608 );
buf ( n4957 , R_fda2_1264e328 );
buf ( n4958 , R_ee25_13a16588 );
buf ( n4959 , R_13a1f_11cde2c8 );
buf ( n4960 , R_1432d_11cdddc8 );
buf ( n4961 , R_13be3_12036bb8 );
buf ( n4962 , R_fe10_13a14468 );
buf ( n4963 , R_12610_1204bcf8 );
buf ( n4964 , R_13701_11cdc608 );
buf ( n4965 , R_12597_105711b8 );
buf ( n4966 , R_1441d_12035d58 );
buf ( n4967 , R_1443c_137979c8 );
buf ( n4968 , R_139a7_11ce70a8 );
buf ( n4969 , R_13ad3_1056bdf8 );
buf ( n4970 , R_143e0_102efcc8 );
buf ( n4971 , R_147cc_13315ae8 );
buf ( n4972 , R_1444b_11cdad08 );
buf ( n4973 , R_12631_12036c58 );
buf ( n4974 , R_13dda_102f4fe8 );
buf ( n4975 , R_efd_13a14fa8 );
buf ( n4976 , R_14954_12054358 );
buf ( n4977 , R_1287f_115422f8 );
buf ( n4978 , R_1169f_102f8968 );
buf ( n4979 , R_13a2b_1264b628 );
buf ( n4980 , R_11285_102f9e08 );
buf ( n4981 , R_12548_1056ce38 );
buf ( n4982 , R_1173e_12649fa8 );
buf ( n4983 , R_10b51_13a18a68 );
buf ( n4984 , R_148ca_13a18c48 );
buf ( n4985 , R_12c82_102f0448 );
buf ( n4986 , R_13b79_11543d38 );
buf ( n4987 , R_14057_f8cd618 );
buf ( n4988 , R_a2e4_1056c618 );
buf ( n4989 , R_101e6_1330c7a8 );
buf ( n4990 , R_13a56_f8c0a58 );
buf ( n4991 , R_d6bc_13a1ca28 );
buf ( n4992 , R_4a_1265e648 );
buf ( n4993 , R_115_13316c68 );
buf ( n4994 , R_1224c_12b3d478 );
buf ( n4995 , R_1fa_1265d388 );
buf ( n4996 , R_eeda_11cd81e8 );
buf ( n4997 , R_1455d_11cd9fe8 );
buf ( n4998 , R_1402e_1264dc48 );
buf ( n4999 , R_c753_12039098 );
buf ( n5000 , R_1283c_13a1da68 );
buf ( n5001 , R_aeda_13a1d6a8 );
buf ( n5002 , R_14939_1379f448 );
buf ( n5003 , R_14a20_13a13e28 );
buf ( n5004 , R_13a9d_12081698 );
buf ( n5005 , R_117c0_11ce3e08 );
buf ( n5006 , R_114e1_132f28e8 );
buf ( n5007 , R_1476f_132fb768 );
buf ( R_147ef_11ce6748 , n27686 );
buf ( R_5f38_10569f58 , n29617 );
buf ( R_13287_11ce6b08 , n30747 );
buf ( R_c94b_102f7608 , n31386 );
buf ( R_20a_1204ce78 , n31387 );
buf ( R_12f29_10571bb8 , n31931 );
buf ( R_13a43_13a1dec8 , n32487 );
buf ( R_1474d_1056fbd8 , n32490 );
buf ( R_14493_12657988 , n32493 );
buf ( R_11fd1_11ce17e8 , n32869 );
buf ( R_14705_1264d248 , n32872 );
buf ( R_105_f8cc2b8 , n32873 );
buf ( R_13cb9_11ce3c28 , n33181 );
buf ( R_138ee_13309fa8 , n33511 );
buf ( R_129dc_11543018 , n33784 );
buf ( R_10bcf_11ce1ba8 , n34047 );
buf ( R_13b6e_13a1e648 , n34257 );
buf ( R_14840_13a13ec8 , n34260 );
buf ( R_13482_10563838 , n34481 );
buf ( R_12d08_12650088 , n34650 );
buf ( R_10303_12b42dd8 , n34843 );
buf ( R_1437c_1056ac78 , n34864 );
buf ( R_87e9_1056cd98 , n35075 );
buf ( R_a30d_13320588 , n35279 );
buf ( R_144a2_133222e8 , n35282 );
buf ( R_1236b_13a1c8e8 , n35464 );
buf ( R_1396e_105627f8 , n35603 );
buf ( R_9ba7_10567258 , n35646 );
buf ( R_1f3_13797a68 , n35647 );
buf ( R_11c_13796528 , n35648 );
buf ( R_7a_1331e148 , n35649 );
buf ( R_117c9_1264ba88 , n35848 );
buf ( R_13b3f_1153ed38 , n35861 );
buf ( R_11abc_1264c2a8 , n36009 );
buf ( R_20d_137962a8 , n36010 );
buf ( R_207_1265a548 , n36011 );
buf ( R_14828_1207a118 , n36014 );
buf ( R_148eb_105aa7d8 , n36017 );
buf ( R_f3a4_10568bf8 , n36108 );
buf ( R_1b6_13799d68 , n36109 );
buf ( R_13429_1207f4d8 , n36165 );
buf ( R_14506_1056e878 , n36168 );
buf ( R_159_12b3d158 , n36169 );
buf ( R_108_105aaeb8 , n36170 );
buf ( R_102_13794cc8 , n36171 );
buf ( R_b1_12053638 , n36172 );
buf ( R_54_13309d28 , n36173 );
buf ( R_145d8_12b3ae58 , n36176 );
buf ( R_1278a_12083718 , n36258 );
buf ( R_13640_11cdeae8 , n36299 );
buf ( R_f706_11542578 , n36407 );
buf ( R_dc82_1153ebf8 , n36470 );
buf ( R_1491b_1265ef08 , n36473 );
buf ( R_14a05_10569738 , n36476 );
buf ( R_13fc5_102eac28 , n36660 );
buf ( R_1405a_115415d8 , n36662 );
buf ( R_136b3_126461c8 , n36708 );
buf ( R_1a0_132f9c88 , n36709 );
buf ( R_16f_1265bee8 , n36710 );
buf ( R_1480d_105a9dd8 , n36713 );
buf ( R_61_13304288 , n36714 );
buf ( R_e082_13798fa8 , n36880 );
buf ( R_10c7d_12082bd8 , n36953 );
buf ( R_14793_1379e188 , n36956 );
buf ( R_11ee1_102f4688 , n37110 );
buf ( R_128ba_12b27758 , n37215 );
buf ( R_70_120513d8 , n37216 );
buf ( R_129f0_12049bd8 , n37272 );
buf ( R_117e7_102f5588 , n37346 );
buf ( R_fee6_13309e68 , n37380 );
buf ( R_148f7_132f3ce8 , n37383 );
buf ( R_1362d_11ce39a8 , n37496 );
buf ( R_10693_126510c8 , n37657 );
buf ( R_11998_12656808 , n37820 );
buf ( R_143ec_11537df8 , n37830 );
buf ( R_138e8_1264afe8 , n37921 );
buf ( R_12650_12649b48 , n38043 );
buf ( R_137a1_105b63f8 , n38195 );
buf ( R_13afd_120772d8 , n38290 );
buf ( R_1490c_1264a7c8 , n38293 );
buf ( R_105e5_13306f88 , n38378 );
buf ( R_12e2b_132fa868 , n38454 );
buf ( R_144e7_12b38e78 , n38457 );
buf ( R_143e4_11cddf08 , n38467 );
buf ( R_1324a_1264c348 , n38502 );
buf ( R_1215a_11542ed8 , n38600 );
buf ( R_f685_11541678 , n38654 );
buf ( R_149ba_102ecb68 , n38657 );
buf ( R_135dc_12646088 , n38731 );
buf ( R_1476c_11cd7928 , n38734 );
buf ( R_146bd_11537998 , n38737 );
buf ( R_1df_12b39378 , n38738 );
buf ( R_13ee8_133069e8 , n38826 );
buf ( R_130_1265ac28 , n38827 );
buf ( R_65_12047c98 , n38828 );
buf ( R_13d75_1330d6a8 , n38843 );
buf ( R_13933_12081198 , n38895 );
buf ( R_133b5_12648388 , n38957 );
buf ( R_125a0_13311488 , n39071 );
buf ( R_8c_1379a808 , n39072 );
buf ( R_eadc_1207ead8 , n39108 );
buf ( R_134c7_126487e8 , n39160 );
buf ( R_11df5_1056e9b8 , n39189 );
buf ( R_144d5_102f8aa8 , n39192 );
buf ( R_12b2a_102eed28 , n39226 );
buf ( R_143d2_11538898 , n39240 );
buf ( R_1462c_102f8508 , n39243 );
buf ( R_13269_11543658 , n39296 );
buf ( R_f4_1331e0a8 , n39297 );
buf ( R_d7_132fde28 , n39298 );
buf ( R_238_1204ec78 , n39299 );
buf ( R_21b_1265e508 , n39300 );
buf ( R_12f3d_12b38b58 , n39312 );
buf ( R_112f1_1153c858 , n39353 );
buf ( R_f09_f8c93d8 , n39355 );
buf ( R_1487c_11cd99a8 , n39358 );
buf ( R_c08f_1207cb98 , n39431 );
buf ( R_923a_13a1ab88 , n39484 );
buf ( R_14042_102f2108 , n39569 );
buf ( R_143e8_102f3b48 , n39579 );
buf ( R_c2e7_13a19e68 , n39662 );
buf ( R_c175_12045118 , n39715 );
buf ( R_1450f_102f8b48 , n39718 );
buf ( R_12b14_12077238 , n39752 );
buf ( R_149e4_13a1c528 , n39755 );
buf ( R_12a04_11ce2968 , n39826 );
buf ( R_145ed_13a14e68 , n39829 );
buf ( R_13884_13796488 , n39892 );
buf ( R_13b0b_1330a688 , n39958 );
buf ( R_b5a4_102f4868 , n40057 );
buf ( R_14584_1056ec38 , n40060 );
buf ( R_13cee_12653148 , n40075 );
buf ( R_10bed_12080ab8 , n40125 );
buf ( R_117f0_102ef4a8 , n40175 );
buf ( R_10a2a_133048c8 , n40222 );
buf ( R_1be_137995e8 , n40223 );
buf ( R_151_12b448b8 , n40224 );
buf ( R_ef06_10563c98 , n40265 );
buf ( R_f9d4_1056b178 , n40325 );
buf ( R_e88a_13a13a68 , n40388 );
buf ( R_13c67_102f38c8 , n40443 );
buf ( R_128eb_10568dd8 , n40522 );
buf ( R_12eaf_f8c3118 , n40534 );
buf ( R_204_12039778 , n40535 );
buf ( R_14951_1265ebe8 , n40538 );
buf ( R_149c3_11ce5348 , n40541 );
buf ( R_1ad_12b28e78 , n40542 );
buf ( R_13f99_102f0da8 , n40592 );
buf ( R_162_12b25e58 , n40593 );
buf ( R_12003_11cdf628 , n40606 );
buf ( R_10b_11539478 , n40607 );
buf ( R_ff_1203c6f8 , n40608 );
buf ( R_1484f_1153ea18 , n40611 );
buf ( R_a8_12b425b8 , n40612 );
buf ( R_5d_13312068 , n40613 );
buf ( R_210_12043bd8 , n40614 );
buf ( R_13d84_102f4188 , n40637 );
buf ( R_142e1_10568658 , n40646 );
buf ( R_10f30_11cd9ae8 , n40672 );
buf ( R_1293d_12b43d78 , n40724 );
buf ( R_10b34_1056da18 , n40752 );
buf ( R_11a07_102eb4e8 , n40783 );
buf ( R_145b1_12082db8 , n40786 );
buf ( R_12c96_13a190a8 , n40837 );
buf ( R_d3b0_10565958 , n40865 );
buf ( R_13f2c_102f4b88 , n40896 );
buf ( R_fb8a_13a18608 , n40921 );
buf ( R_130d5_13319c88 , n40973 );
buf ( R_13f89_102f36e8 , n40986 );
buf ( R_146ff_13a1a4a8 , n40989 );
buf ( R_10ccb_1264f868 , n41015 );
buf ( R_124c3_1056f138 , n41027 );
buf ( R_10786_102f2568 , n41074 );
buf ( R_12a16_10568e78 , n41105 );
buf ( R_10726_102ef408 , n41136 );
buf ( R_137d3_12656da8 , n41158 );
buf ( R_13863_11cddb48 , n41176 );
buf ( R_14993_102f27e8 , n41179 );
buf ( R_bab1_1264a2c8 , n41222 );
buf ( R_1451e_10565818 , n41225 );
buf ( R_12a46_126515c8 , n41250 );
buf ( R_e7da_102f3508 , n41262 );
buf ( R_12756_13a1f0e8 , n41293 );
buf ( R_c4_13797ba8 , n41294 );
buf ( R_128da_1207ec18 , n41325 );
buf ( R_c282_12076838 , n41335 );
buf ( R_1272e_1056cbb8 , n41350 );
buf ( R_14a5f_120797b8 , n41353 );
buf ( R_14448_12663648 , n41356 );
buf ( R_c2_12048058 , n41357 );
buf ( R_1372d_11ce2aa8 , n41398 );
buf ( R_f878_1207c7d8 , n41410 );
buf ( R_13a76_13797888 , n41441 );
buf ( R_13a17_13796b68 , n41456 );
buf ( R_1cb_12044ad8 , n41457 );
buf ( R_14462_12b3f8b8 , n41460 );
buf ( R_6021_1379bd48 , n41510 );
buf ( R_144_13795128 , n41511 );
buf ( R_1383e_105671b8 , n41552 );
buf ( R_147ab_1056a6d8 , n41555 );
buf ( R_c6_1330e0a8 , n41556 );
buf ( R_249_12654368 , n41557 );
buf ( R_1305a_13796ca8 , n41569 );
buf ( R_12e4b_13307348 , n41597 );
buf ( R_14a38_137a1e28 , n41600 );
buf ( R_d1de_11cd9ea8 , n41637 );
buf ( R_138e2_11cd83c8 , n41671 );
buf ( R_13e62_1056dab8 , n41698 );
buf ( R_114a7_1331d748 , n41710 );
buf ( R_12f53_13319648 , n41722 );
buf ( R_f8a4_11543a18 , n41750 );
buf ( R_11ec3_13a157c8 , n41778 );
buf ( R_12c06_11cdac68 , n41825 );
buf ( R_12be8_12649788 , n41835 );
buf ( R_136c6_11cdc6a8 , n41863 );
buf ( R_1482e_13a1a228 , n41866 );
buf ( R_10ba7_115431f8 , n41891 );
buf ( R_89f2_11545098 , n41903 );
buf ( R_11953_1153c538 , n41915 );
buf ( R_9e64_11ce48a8 , n41942 );
buf ( R_e77d_11ce3ea8 , n41957 );
buf ( R_1091c_13a1a2c8 , n41969 );
buf ( R_114ec_12650628 , n42000 );
buf ( R_1286a_11cdcd88 , n42015 );
buf ( R_10d6d_1265db08 , n42056 );
buf ( R_1228f_1331f0e8 , n42064 );
buf ( R_1c5_126590a8 , n42065 );
buf ( R_14490_132f7d48 , n42068 );
buf ( R_1a1_1264a408 , n42069 );
buf ( R_976e_12056398 , n42081 );
buf ( R_6845_12648ec8 , n42091 );
buf ( R_16e_1379a3a8 , n42092 );
buf ( R_14a_12657528 , n42093 );
buf ( R_12718_10566fd8 , n42105 );
buf ( R_145c9_12075438 , n42108 );
buf ( R_c0_132fa5e8 , n42109 );
buf ( R_9c_12655f48 , n42110 );
buf ( R_d230_102edec8 , n42122 );
buf ( R_69_12658888 , n42123 );
buf ( R_13097_11ce5b68 , n42131 );
buf ( R_11051_1264a5e8 , n42143 );
buf ( R_145f0_11536818 , n42146 );
buf ( R_13ccd_132f9288 , n42154 );
buf ( R_e0_12661ac8 , n42155 );
buf ( R_22f_1331df68 , n42156 );
buf ( R_12a2a_11cd9f48 , n42168 );
buf ( R_10a54_11540458 , n42199 );
buf ( R_d027_13795628 , n42211 );
buf ( R_144d2_105677f8 , n42214 );
buf ( R_14638_11cd9228 , n42217 );
buf ( R_1454b_10568338 , n42220 );
buf ( R_147fe_1265bb28 , n42223 );
buf ( R_e861_12650448 , n42233 );
buf ( R_c03c_137931e8 , n42245 );
buf ( R_13574_102f97c8 , n42276 );
buf ( R_10e6d_102ec0c8 , n42288 );
buf ( R_c8_1331c348 , n42289 );
buf ( R_247_12b3bad8 , n42290 );
buf ( R_77_126636e8 , n42291 );
buf ( R_13a50_1056bb78 , n42315 );
buf ( R_129a5_11543798 , n42330 );
buf ( R_ef35_102f6d48 , n42355 );
buf ( R_1028c_137951c8 , n42367 );
buf ( R_1348b_12051838 , n42386 );
buf ( R_11f8b_11cdc428 , n42394 );
buf ( R_1452d_f8c5878 , n42397 );
buf ( R_12a3b_12650308 , n42407 );
buf ( R_13fd5_12079d58 , n42419 );
buf ( R_dd89_13302de8 , n42427 );
buf ( R_13dcc_102f7ec8 , n42439 );
buf ( R_14822_102f5768 , n42442 );
buf ( R_baf1_12084e38 , n42454 );
buf ( R_1315c_11ce75a8 , n42466 );
buf ( R_df0e_12654d68 , n42478 );
buf ( R_efea_11cdc248 , n42490 );
buf ( R_fe90_13a14a08 , n42515 );
buf ( R_1453c_102ec208 , n42518 );
buf ( R_aaa7_102edba8 , n42530 );
buf ( R_13c4e_13a1c988 , n42561 );
buf ( R_f758_13a13d88 , n42569 );
buf ( R_1485e_12b38f18 , n42572 );
buf ( R_ece9_1264c488 , n42584 );
buf ( R_14a35_12037f18 , n42587 );
buf ( R_1190c_102ecfc8 , n42641 );
buf ( R_12810_12650d08 , n42653 );
buf ( R_f016_12044df8 , n42661 );
buf ( R_1494e_13a14f08 , n42664 );
buf ( R_14344_1264eaa8 , n42675 );
buf ( R_10e_1265af48 , n42676 );
buf ( R_13f62_12075758 , n42688 );
buf ( R_fc_133201c8 , n42689 );
buf ( R_1378e_11cdd8c8 , n42697 );
buf ( R_147eb_120847f8 , n42700 );
buf ( R_13331_13308ec8 , n42708 );
buf ( R_213_12654f48 , n42709 );
buf ( R_146ae_1265dc48 , n42712 );
buf ( R_201_1153b138 , n42713 );
buf ( R_11d47_f8cc0d8 , n42721 );
buf ( R_c820_13a19328 , n42733 );
buf ( R_edbe_132fbd08 , n42745 );
buf ( R_be_132f4148 , n42746 );
buf ( R_a1_12043c78 , n42747 );
buf ( R_131b9_102f29c8 , n42759 );
buf ( R_12eb9_1153f738 , n42769 );
buf ( R_146e1_1153fb98 , n42772 );
buf ( R_1487f_13a173e8 , n42775 );
buf ( R_13fb4_11544af8 , n42783 );
buf ( R_1446b_10568798 , n42786 );
buf ( R_ef60_1264cf28 , n42798 );
buf ( R_1463b_1207bd38 , n42801 );
buf ( R_13166_1153aff8 , n42809 );
buf ( R_10a4b_10565bd8 , n42815 );
buf ( R_14599_12080c98 , n42818 );
buf ( R_10b18_12080018 , n42830 );
buf ( R_7254_12055078 , n42842 );
buf ( R_db04_1207b3d8 , n42854 );
buf ( R_149f9_10570cb8 , n42857 );
buf ( R_14a4a_1265d608 , n42860 );
buf ( R_14796_1264b808 , n42863 );
buf ( R_120d3_1379f3a8 , n42871 );
buf ( R_119cb_102f2068 , n42883 );
buf ( R_12acb_10565458 , n42893 );
buf ( R_145b4_12083358 , n42896 );
buf ( R_11ae9_12651528 , n42908 );
buf ( R_13af6_f8ce6f8 , n42920 );
buf ( R_13451_102f0128 , n42930 );
buf ( R_ef8c_1204e098 , n42955 );
buf ( R_ca_12b3e058 , n42956 );
buf ( R_245_f8c5ff8 , n42957 );
buf ( R_af_12b2a8b8 , n42958 );
buf ( R_10e57_11544eb8 , n42966 );
buf ( R_b243_f8c5698 , n42978 );
buf ( R_13633_13a13248 , n42990 );
buf ( R_11c97_10562078 , n43002 );
buf ( R_13838_102f5e48 , n43010 );
buf ( R_efb7_13a1bc68 , n43020 );
buf ( R_d4db_10566038 , n43033 );
buf ( R_10bc8_11ce66a8 , n43045 );
buf ( R_c9c0_102eee68 , n43055 );
buf ( R_13608_10563798 , n43067 );
buf ( R_8f_12b299b8 , n43068 );
buf ( R_59_133089c8 , n43069 );
buf ( R_134f1_102ebf88 , n43077 );
buf ( R_10499_1331e828 , n43085 );
buf ( R_14424_102f8f08 , n43091 );
buf ( R_1d6_133209e8 , n43092 );
buf ( R_ebe2_13a18568 , n43104 );
buf ( R_139_12b44ef8 , n43105 );
buf ( R_97_13792c48 , n43106 );
buf ( R_144ed_105660d8 , n43109 );
buf ( R_120c8_11541d58 , n43119 );
buf ( R_11736_11cde408 , n43127 );
buf ( R_149a8_13317528 , n43130 );
buf ( R_1450c_1056eff8 , n43133 );
buf ( R_147d9_120828b8 , n43136 );
buf ( R_11ea5_1264a9a8 , n43146 );
buf ( R_11425_1207c918 , n43158 );
buf ( R_d53e_1207c2d8 , n43170 );
buf ( R_14787_12b352b8 , n43173 );
buf ( R_13cf3_10571078 , n43185 );
buf ( R_13f36_1330ebe8 , n43193 );
buf ( R_d00d_102ee968 , n43205 );
buf ( R_a1e6_11cde368 , n43217 );
buf ( R_13f77_13a19648 , n43225 );
buf ( R_118_132f5f48 , n43226 );
buf ( R_13688_120832b8 , n43234 );
buf ( R_1f7_105a9978 , n43235 );
buf ( R_f630_1056b858 , n43247 );
buf ( R_136a1_1153fa58 , n43255 );
buf ( R_1b7_126577a8 , n43256 );
buf ( R_158_12b27938 , n43257 );
buf ( R_ec_1330a868 , n43258 );
buf ( R_223_f8c32f8 , n43259 );
buf ( R_133bf_11543338 , n43290 );
buf ( R_f2a8_102f47c8 , n43302 );
buf ( R_e112_12076e78 , n43310 );
buf ( R_12b72_1056c6b8 , n43322 );
buf ( R_2f00_102f3d28 , n43332 );
buf ( R_14819_1331de28 , n43335 );
buf ( R_e809_13313c48 , n43347 );
buf ( R_14358_11cd8788 , n43358 );
buf ( R_1473e_11543b58 , n43361 );
buf ( R_139c7_102ed1a8 , n43369 );
buf ( R_13d65_12036a78 , n43379 );
buf ( R_12c10_102ea548 , n43389 );
buf ( R_13870_11ce5e88 , n43395 );
buf ( R_dede_13a16448 , n43407 );
buf ( R_12c49_12b27438 , n43419 );
buf ( R_1192b_12645e08 , n43431 );
buf ( R_bd66_126533c8 , n43437 );
buf ( R_13fa2_1379f6c8 , n43445 );
buf ( R_13407_1056df18 , n43473 );
buf ( R_118b0_1204acb8 , n43504 );
buf ( R_13c3e_126496e8 , n43512 );
buf ( R_1438a_11cda268 , n43522 );
buf ( R_11e51_102fa268 , n43532 );
buf ( R_102b9_132f6588 , n43544 );
buf ( R_d9_1330dec8 , n43545 );
buf ( R_bc_13799c28 , n43546 );
buf ( R_236_13795f88 , n43547 );
buf ( R_ffee_1264d568 , n43553 );
buf ( R_10ea9_102f8788 , n43561 );
buf ( R_14852_13a154a8 , n43564 );
buf ( R_e696_11cdce28 , n43576 );
buf ( R_1ae_1203c3d8 , n43577 );
buf ( R_1457e_133027e8 , n43580 );
buf ( R_161_12656c68 , n43581 );
buf ( R_127_12b3cc58 , n43582 );
buf ( R_ea26_1265a4a8 , n43594 );
buf ( R_1e8_11539298 , n43595 );
buf ( R_139e4_102f59e8 , n43603 );
buf ( R_1477b_1204f218 , n43606 );
buf ( R_1459c_12056a78 , n43609 );
buf ( R_1336e_11545138 , n43619 );
buf ( R_108cd_102f7ce8 , n43631 );
buf ( R_13b4f_13305c28 , n43643 );
buf ( R_1a2_12b423d8 , n43644 );
buf ( R_16d_12664c28 , n43645 );
buf ( R_14656_11ce6ce8 , n43648 );
buf ( R_827e_1207e998 , n43660 );
buf ( R_11ab0_1204a358 , n43672 );
buf ( R_144ab_12b39af8 , n43675 );
buf ( R_144c3_12080338 , n43678 );
buf ( R_12794_102f5b28 , n43688 );
buf ( R_13149_102f7888 , n43700 );
buf ( R_144e4_12b28838 , n43703 );
buf ( R_13e_12660da8 , n43704 );
buf ( R_123_1330d888 , n43705 );
buf ( R_e7_137956c8 , n43706 );
buf ( R_cc_12038918 , n43707 );
buf ( R_137c7_102f79c8 , n43719 );
buf ( R_243_13796d48 , n43720 );
buf ( R_13795_13795588 , n43732 );
buf ( R_228_10570c18 , n43733 );
buf ( R_13f01_1056e2d8 , n43743 );
buf ( R_13d8e_11cd77e8 , n43755 );
buf ( R_1ec_12039ef8 , n43756 );
buf ( R_f175_13a17ca8 , n43762 );
buf ( R_1d1_126540e8 , n43763 );
buf ( R_14409_12b434b8 , n43778 );
buf ( R_138b2_102f06c8 , n43784 );
buf ( R_14653_1207e0d8 , n43787 );
buf ( R_13044_102f7a68 , n43795 );
buf ( R_13133_13a1ae08 , n43807 );
buf ( R_10b8f_1265ad68 , n43819 );
buf ( R_12e35_12b3b858 , n43831 );
buf ( R_12df0_12050bb8 , n43837 );
buf ( R_fc88_1207be78 , n43845 );
buf ( R_13804_102ef548 , n43855 );
buf ( R_13b68_137a1ba8 , n43865 );
buf ( R_134_13312b68 , n43866 );
buf ( R_14990_1331ae08 , n43869 );
buf ( R_1db_12043db8 , n43870 );
buf ( R_ccdc_102f6488 , n43882 );
buf ( R_1494b_11ce61a8 , n43885 );
buf ( R_12c39_10562ed8 , n43893 );
buf ( R_131c2_11ce4b28 , n43899 );
buf ( R_12d97_126626a8 , n43909 );
buf ( R_12d59_12b26b78 , n43921 );
buf ( R_1352d_13315188 , n43933 );
buf ( R_12c4f_13321d48 , n43943 );
buf ( R_1343e_10562d98 , n43955 );
buf ( R_1345b_102fa088 , n43967 );
buf ( R_1167d_115410d8 , n43979 );
buf ( R_14008_1264dec8 , n44002 );
buf ( R_11bc8_11544e18 , n44010 );
buf ( R_13c9a_1207e178 , n44016 );
buf ( R_148be_12b27f78 , n44019 );
buf ( R_14360_105ad078 , n44027 );
buf ( R_13aa3_12078138 , n44035 );
buf ( R_116da_13a1a7c8 , n44045 );
buf ( R_14732_102f5448 , n44048 );
buf ( R_cec6_132f3608 , n44056 );
buf ( R_133dc_13a1ea08 , n44064 );
buf ( R_14942_f8c5058 , n44067 );
buf ( R_13a0f_10563018 , n44077 );
buf ( R_bd10_f8ce978 , n44083 );
buf ( R_12da1_12647528 , n44093 );
buf ( R_12af5_12052418 , n44105 );
buf ( R_13cf9_13a1c0c8 , n44113 );
buf ( R_13658_12646628 , n44121 );
buf ( R_149bd_1204adf8 , n44124 );
buf ( R_13233_11cde908 , n44132 );
buf ( R_12585_1207a898 , n44157 );
buf ( R_118e9_10564a58 , n44169 );
buf ( R_1359a_13a18928 , n44181 );
buf ( R_12451_13a1d568 , n44191 );
buf ( R_dcbb_1265bf88 , n44199 );
buf ( R_f424_13a1b948 , n44211 );
buf ( R_1226a_11cdef48 , n44219 );
buf ( R_14641_13a12d48 , n44222 );
buf ( R_1257c_11ce4448 , n44234 );
buf ( R_e309_120806f8 , n44242 );
buf ( R_11ccc_13314be8 , n44252 );
buf ( R_146c0_13a15908 , n44255 );
buf ( R_14843_13a196e8 , n44258 );
buf ( R_11d00_1207f9d8 , n44264 );
buf ( R_14a1d_13a14c88 , n44267 );
buf ( R_13d54_11ce00c8 , n44273 );
buf ( R_135b5_132fdd88 , n44285 );
buf ( R_d40b_10569058 , n44295 );
buf ( R_145f9_102ee148 , n44298 );
buf ( R_14882_1056d838 , n44301 );
buf ( R_101a4_f8c2ad8 , n44313 );
buf ( R_13abf_13a15188 , n44321 );
buf ( R_eab3_126509e8 , n44331 );
buf ( R_8296_13322608 , n44343 );
buf ( R_6d_12036618 , n44344 );
buf ( R_50_12b3c118 , n44345 );
buf ( R_11b19_102ee508 , n44357 );
buf ( R_de1d_13a193c8 , n44363 );
buf ( R_14477_11cdcc48 , n44366 );
buf ( R_1195d_12038198 , n44374 );
buf ( R_14527_102eb6c8 , n44377 );
buf ( R_be8c_126504e8 , n44387 );
buf ( R_11e87_12b3c398 , n44399 );
buf ( R_14a02_13309aa8 , n44402 );
buf ( R_12b_1203e6d8 , n44403 );
buf ( R_f1_13799ea8 , n44404 );
buf ( R_21e_126608a8 , n44405 );
buf ( R_1e4_12b28338 , n44406 );
buf ( R_115ff_13304148 , n44416 );
buf ( R_10d8e_1264cfc8 , n44424 );
buf ( R_11500_12083c18 , n44430 );
buf ( R_c4bc_137945e8 , n44442 );
buf ( R_1465c_10568f18 , n44445 );
buf ( R_133e6_11cd9048 , n44457 );
buf ( R_7c4f_11ce4a88 , n44469 );
buf ( R_11f78_12b2c118 , n44481 );
buf ( R_1013a_132f59a8 , n44489 );
buf ( R_149e1_105b62b8 , n44492 );
buf ( R_150_1330cac8 , n44493 );
buf ( R_111_12b3e238 , n44494 );
buf ( R_f9_1204ba78 , n44495 );
buf ( R_ba_1331bc68 , n44496 );
buf ( R_4b_1264c028 , n44497 );
buf ( R_216_1204a038 , n44498 );
buf ( R_13733_f8d0098 , n44506 );
buf ( R_1fe_120539f8 , n44507 );
buf ( R_146de_12648748 , n44510 );
buf ( R_1bf_1265cd48 , n44511 );
buf ( R_74_1331da68 , n44512 );
buf ( R_f5c3_1264d108 , n44522 );
buf ( R_f1f7_120367f8 , n44534 );
buf ( R_e338_13301ac8 , n44542 );
buf ( R_1486d_1056e558 , n44545 );
buf ( R_13e2d_12047fb8 , n44555 );
buf ( R_12344_137a0de8 , n44565 );
buf ( R_14729_10570178 , n44568 );
buf ( R_13364_105717f8 , n44580 );
buf ( R_11160_1153e298 , n44590 );
buf ( R_10a01_11cde228 , n44598 );
buf ( R_13c6f_12041658 , n44608 );
buf ( R_148c4_10568978 , n44611 );
buf ( R_11c81_132f7348 , n44623 );
buf ( R_10ec5_11cdb028 , n44633 );
buf ( R_14441_12659008 , n44637 );
buf ( R_cbab_105a9a18 , n44643 );
buf ( R_1238a_126482e8 , n44653 );
buf ( R_a6_12660448 , n44654 );
buf ( R_12b36_11ce6428 , n44660 );
buf ( R_dc46_10566498 , n44670 );
buf ( R_11f_137936e8 , n44671 );
buf ( R_ce_12055fd8 , n44672 );
buf ( R_241_132fd748 , n44673 );
buf ( R_147f8_1207ccd8 , n44676 );
buf ( R_1f0_13798a08 , n44677 );
buf ( R_1467d_1056bcb8 , n44680 );
buf ( R_14668_11546178 , n44683 );
buf ( R_132cc_1153edd8 , n44695 );
buf ( R_136ba_11ce37c8 , n44703 );
buf ( R_12c23_102f1d48 , n44711 );
buf ( R_106be_1264edc8 , n44719 );
buf ( R_11bde_10564878 , n44727 );
buf ( R_11a1a_11cd9a48 , n44737 );
buf ( R_9548_11ce6ba8 , n44745 );
buf ( R_f451_11542438 , n44753 );
buf ( R_119b7_105663f8 , n44765 );
buf ( R_142e5_102f2388 , n44774 );
buf ( R_147e4_13a19dc8 , n44777 );
buf ( R_d862_12661348 , n44789 );
buf ( R_d940_13a19d28 , n44797 );
buf ( R_eb8c_13a19288 , n44807 );
buf ( R_1175e_11cda088 , n44817 );
buf ( R_146f9_11ce4768 , n44820 );
buf ( R_14551_102eae08 , n44823 );
buf ( R_14578_12b3a6d8 , n44826 );
buf ( R_1467a_13a13568 , n44829 );
buf ( R_1130e_1056bfd8 , n44837 );
buf ( R_1493f_1056d3d8 , n44840 );
buf ( R_14948_102f76a8 , n44843 );
buf ( R_10230_1153d1b8 , n44855 );
buf ( R_f4d1_13a17848 , n44863 );
buf ( R_14772_11cda8a8 , n44866 );
buf ( R_1466e_1203e138 , n44869 );
buf ( R_14999_120382d8 , n44872 );
buf ( R_9d72_102f18e8 , n44884 );
buf ( R_eeaf_10566f38 , n44896 );
buf ( R_13083_12b3ff98 , n44908 );
buf ( R_e288_11541fd8 , n44920 );
buf ( R_13969_102ea408 , n44928 );
buf ( R_13825_1264d928 , n44940 );
buf ( R_134a8_13a13c48 , n44950 );
buf ( R_fcde_115390b8 , n44958 );
buf ( R_14566_102f6988 , n44961 );
buf ( R_f5eb_11544558 , n44969 );
buf ( R_12318_102ec348 , n44981 );
buf ( R_d2c9_11cd9408 , n44993 );
buf ( R_16c_132f7ca8 , n44994 );
buf ( R_d894_1056f778 , n45002 );
buf ( R_12323_102ec8e8 , n45014 );
buf ( R_1a3_13303108 , n45015 );
buf ( R_118ba_13307ac8 , n45023 );
buf ( R_12704_10562938 , n45031 );
buf ( R_148c7_1264d888 , n45034 );
buf ( R_148bb_12661d48 , n45037 );
buf ( R_1221a_13a1d248 , n45049 );
buf ( R_135b0_12651348 , n45055 );
buf ( R_1470e_10562898 , n45058 );
buf ( R_efa_1207d1d8 , n45060 );
buf ( R_ce1e_102f95e8 , n45068 );
buf ( R_126e3_105b5c78 , n45080 );
buf ( R_14026_102ecd48 , n45092 );
buf ( R_11e36_102ed608 , n45100 );
buf ( R_11515_12039318 , n45106 );
buf ( R_108e3_1056dd38 , n45118 );
buf ( R_128f4_1207aa78 , n45124 );
buf ( R_147ae_1207ce18 , n45127 );
buf ( R_12235_12650e48 , n45139 );
buf ( R_12183_12052eb8 , n45149 );
buf ( R_14647_102f04e8 , n45152 );
buf ( R_13aef_11cdd968 , n45162 );
buf ( R_1249f_102f9368 , n45170 );
buf ( R_f34d_13a18ec8 , n45180 );
buf ( R_12c3f_f8cfd78 , n45190 );
buf ( R_13d5d_1153d4d8 , n45202 );
buf ( R_12126_102ef228 , n45210 );
buf ( R_ad_12b3b358 , n45211 );
buf ( R_92_13312d48 , n45212 );
buf ( R_113db_f8cb4f8 , n45222 );
buf ( R_10d98_f8c6318 , n45234 );
buf ( R_1481f_1264dce8 , n45237 );
buf ( R_ad98_102f3aa8 , n45245 );
buf ( R_55_132f50e8 , n45246 );
buf ( R_102d5_f8ced38 , n45256 );
buf ( R_144ae_11545ef8 , n45259 );
buf ( R_a3e0_12655308 , n45267 );
buf ( R_5dbf_13a15f48 , n45275 );
buf ( R_e2_1203f858 , n45276 );
buf ( R_22d_1379de68 , n45277 );
buf ( R_135c4_105b5bd8 , n45289 );
buf ( R_13cff_13a16308 , n45297 );
buf ( R_12692_102eb8a8 , n45305 );
buf ( R_13375_13794a48 , n45317 );
buf ( R_12f6a_10562438 , n45329 );
buf ( R_128c4_102ea5e8 , n45339 );
buf ( R_122f0_12650f88 , n45345 );
buf ( R_14855_12056f78 , n45348 );
buf ( R_14885_13795a88 , n45351 );
buf ( R_bb92_11ce0ca8 , n45357 );
buf ( R_8b04_1265cf28 , n45365 );
buf ( R_e71c_115426b8 , n45377 );
buf ( R_14a23_120545d8 , n45380 );
buf ( R_149_1330f408 , n45381 );
buf ( R_b8_13305048 , n45382 );
buf ( R_1c6_1379cce8 , n45383 );
buf ( R_e13d_102eb448 , n45393 );
buf ( R_14617_11ce2f08 , n45396 );
buf ( R_13557_11545778 , n45404 );
buf ( R_148cd_12082c78 , n45407 );
buf ( R_11768_1264ffe8 , n45413 );
buf ( R_12503_11cdd008 , n45425 );
buf ( R_1239d_1330d1a8 , n45431 );
buf ( R_1448c_105662b8 , n45434 );
buf ( R_160_f8c0d78 , n45435 );
buf ( R_143_13795e48 , n45436 );
buf ( R_1252c_102f1208 , n45446 );
buf ( R_1cc_f8cc858 , n45447 );
buf ( R_149de_11cde7c8 , n45450 );
buf ( R_1af_12b40678 , n45451 );
buf ( R_a28f_11ce5708 , n45461 );
buf ( R_f7ae_11ce57a8 , n45471 );
buf ( R_1243d_10571118 , n45481 );
buf ( R_d0df_126478e8 , n45493 );
buf ( R_1498d_1153fe18 , n45496 );
buf ( R_10350_11cda6c8 , n45506 );
buf ( R_103a6_10569878 , n45512 );
buf ( R_128b0_1056c118 , n45524 );
buf ( R_14936_10561e98 , n45527 );
buf ( R_10d1b_11cd7748 , n45539 );
buf ( R_ed92_102eea08 , n45551 );
buf ( R_145d2_11cdb208 , n45554 );
buf ( R_109f6_1153ca38 , n45562 );
buf ( R_cc46_1207b298 , n45570 );
buf ( R_11006_126501c8 , n45578 );
buf ( R_188_1265c348 , n45579 );
buf ( R_187_12b25d18 , n45580 );
buf ( R_12f_1379dbe8 , n45581 );
buf ( R_db_12663f08 , n45582 );
buf ( R_84_12652ce8 , n45583 );
buf ( R_81_12042a58 , n45584 );
buf ( R_234_12b43af8 , n45585 );
buf ( R_1e0_133037e8 , n45586 );
buf ( R_13ed7_1207ad98 , n45596 );
buf ( R_189_f8c6458 , n45597 );
buf ( R_186_126553a8 , n45598 );
buf ( R_157_132f7a28 , n45599 );
buf ( R_d0_105aa238 , n45600 );
buf ( R_23f_13307848 , n45601 );
buf ( R_11399_12b3c1b8 , n45609 );
buf ( R_1b8_11537358 , n45610 );
buf ( R_f82c_f8cdc58 , n45622 );
buf ( R_d9ca_10562bb8 , n45634 );
buf ( R_145f6_f8c3398 , n45637 );
buf ( R_1449c_11ce71e8 , n45640 );
buf ( R_13850_13a1fe08 , n45648 );
buf ( R_135e3_13306da8 , n45656 );
buf ( R_ec0b_132fa368 , n45662 );
buf ( R_147e0_13a12fc8 , n45665 );
buf ( R_13add_132ff728 , n45677 );
buf ( R_f65b_12084578 , n45685 );
buf ( R_10cb4_11cdf9e8 , n45695 );
buf ( R_18a_133173e8 , n45696 );
buf ( R_185_12042cd8 , n45697 );
buf ( R_134d0_12651028 , n45705 );
buf ( R_144f3_102f3fa8 , n45708 );
buf ( R_12dd1_f8c52d8 , n45714 );
buf ( R_135a9_10567938 , n45726 );
buf ( R_11b39_102ec988 , n45738 );
buf ( R_1386a_102ebda8 , n45744 );
buf ( R_14747_12042b98 , n45747 );
buf ( R_148d0_137a0a28 , n45750 );
buf ( R_11f4d_137986e8 , n45760 );
buf ( R_13d05_12081378 , n45770 );
buf ( R_f56e_102f2608 , n45776 );
buf ( R_62_12b26498 , n45777 );
buf ( R_10e0b_1056abd8 , n45787 );
buf ( R_ba73_1264c8e8 , n45799 );
buf ( R_14888_12653288 , n45802 );
buf ( R_fc34_1379c428 , n45814 );
buf ( R_18b_12663fa8 , n45815 );
buf ( R_184_1153acd8 , n45816 );
buf ( R_119d5_1331dc48 , n45824 );
buf ( R_122b5_13305688 , n45836 );
buf ( R_e051_12649f08 , n45844 );
buf ( R_ca0a_10567438 , n45854 );
buf ( R_10a84_115427f8 , n45862 );
buf ( R_668e_10563f18 , n45868 );
buf ( R_14539_102f7108 , n45871 );
buf ( R_c3d6_11cdb7a8 , n45883 );
buf ( R_11703_132fa728 , n45891 );
buf ( R_1472f_105708f8 , n45894 );
buf ( R_1307a_11cdc1a8 , n45902 );
buf ( R_fdae_1153d258 , n45910 );
buf ( R_13ac5_102ee3c8 , n45920 );
buf ( R_120bd_1153ff58 , n45932 );
buf ( R_13f6e_12649dc8 , n45940 );
buf ( R_1177b_1207fbb8 , n45952 );
buf ( R_f804_1379efe8 , n45960 );
buf ( R_111d5_13a17c08 , n45968 );
buf ( R_14750_13304008 , n45971 );
buf ( R_137d9_12055e98 , n45977 );
buf ( R_87_132ffa48 , n45978 );
buf ( R_7e_137949a8 , n45979 );
buf ( R_f140_1056f598 , n45987 );
buf ( R_d43f_12079678 , n45993 );
buf ( R_11900_1056f6d8 , n46005 );
buf ( R_18c_12660e48 , n46006 );
buf ( R_c969_1330f9a8 , n46016 );
buf ( R_183_126587e8 , n46017 );
buf ( R_11093_102f60c8 , n46025 );
buf ( R_f31e_120770f8 , n46031 );
buf ( R_f06_1265f728 , n46033 );
buf ( R_d5cf_102f5128 , n46045 );
buf ( R_10874_12037838 , n46051 );
buf ( R_11324_13a1f228 , n46057 );
buf ( R_13621_120823b8 , n46067 );
buf ( R_120dd_f8cdcf8 , n46077 );
buf ( R_148d3_12049a98 , n46080 );
buf ( R_13e42_12648888 , n46088 );
buf ( R_144c0_12078db8 , n46091 );
buf ( R_12978_13316d08 , n46099 );
buf ( R_11b5e_13a1b088 , n46109 );
buf ( R_13025_13a1ef08 , n46121 );
buf ( R_e615_12084bb8 , n46127 );
buf ( R_149b7_102ea4a8 , n46130 );
buf ( R_1497e_1207ef38 , n46133 );
buf ( R_11fee_12b2a3b8 , n46145 );
buf ( R_11b_12b43198 , n46146 );
buf ( R_5e_126647c8 , n46147 );
buf ( R_1f4_1265d108 , n46148 );
buf ( R_1445f_13792888 , n46151 );
buf ( R_13981_13798aa8 , n46161 );
buf ( R_14569_11cdbfc8 , n46164 );
buf ( R_114_12b3e4b8 , n46165 );
buf ( R_f6_12664188 , n46166 );
buf ( R_9f_12054d58 , n46167 );
buf ( R_66_13308068 , n46168 );
buf ( R_219_1203c338 , n46169 );
buf ( R_132a5_12654868 , n46179 );
buf ( R_f9aa_11cdd5a8 , n46191 );
buf ( R_1fb_126610c8 , n46192 );
buf ( R_1a4_13798648 , n46193 );
buf ( R_16b_1331a2c8 , n46194 );
buf ( R_9a_12658568 , n46195 );
buf ( R_13c54_102f6e88 , n46207 );
buf ( R_14933_1207e5d8 , n46210 );
buf ( R_a6b7_1264b588 , n46218 );
buf ( R_10fad_13a15548 , n46226 );
buf ( R_18d_13321a28 , n46227 );
buf ( R_182_13315cc8 , n46228 );
buf ( R_14a58_102f65c8 , n46233 );
buf ( R_c8f6_132f4a08 , n46241 );
buf ( R_1458d_13a17ac8 , n46244 );
buf ( R_126d9_11545598 , n46252 );
buf ( R_10942_102f85a8 , n46262 );
buf ( R_14a32_12654ea8 , n46265 );
buf ( R_b7bc_12b28798 , n46275 );
buf ( R_1389f_11cda3a8 , n46283 );
buf ( R_14602_102ed7e8 , n46286 );
buf ( R_100bf_1330b9e8 , n46294 );
buf ( R_112eb_115386b8 , n46300 );
buf ( R_146d5_105b59f8 , n46303 );
buf ( R_1206a_1207c878 , n46309 );
buf ( R_e2de_1264ce88 , n46317 );
buf ( R_13b3a_11cddaa8 , n46325 );
buf ( R_13739_10563bf8 , n46331 );
buf ( R_148d6_11cd86e8 , n46334 );
buf ( R_1319d_11544918 , n46340 );
buf ( R_12f7f_12077eb8 , n46348 );
buf ( R_1242c_f8cda78 , n46356 );
buf ( R_14483_12054fd8 , n46359 );
buf ( R_14456_102ea728 , n46362 );
buf ( R_6b42_120790d8 , n46370 );
buf ( R_1186d_f8cbb38 , n46378 );
buf ( R_147d3_12648e28 , n46381 );
buf ( R_11add_1056c4d8 , n46389 );
buf ( R_13c18_1264df68 , n46401 );
buf ( R_13e19_132f7c08 , n46411 );
buf ( R_b6_1265e148 , n46412 );
buf ( R_13bb8_1265edc8 , n46420 );
buf ( R_146a8_12050118 , n46423 );
buf ( R_18e_12043ef8 , n46424 );
buf ( R_181_12647a28 , n46425 );
buf ( R_b677_12083178 , n46437 );
buf ( R_1176f_1379f8a8 , n46447 );
buf ( R_11d7b_102f2d88 , n46455 );
buf ( R_145bd_1207cff8 , n46458 );
buf ( R_13bae_105700d8 , n46466 );
buf ( R_10fed_1330ad68 , n46474 );
buf ( R_1479f_11cde4a8 , n46477 );
buf ( R_71_1265e8c8 , n46478 );
buf ( R_3ca5_102eebe8 , n46486 );
buf ( R_14769_1056b718 , n46489 );
buf ( R_139ba_11ce35e8 , n46495 );
buf ( R_ccf5_13a128e8 , n46505 );
buf ( R_13964_1207def8 , n46513 );
buf ( R_13920_133128e8 , n46521 );
buf ( R_13b74_11cd8dc8 , n46533 );
buf ( R_13e6d_11cd90e8 , n46539 );
buf ( R_13ae8_11545db8 , n46547 );
buf ( R_e946_13796668 , n46555 );
buf ( R_12db3_10562b18 , n46563 );
buf ( R_7b5f_1264bc68 , n46571 );
buf ( R_139f5_132fc348 , n46583 );
buf ( R_cd6e_10562a78 , n46591 );
buf ( R_13626_12077cd8 , n46601 );
buf ( R_148dc_102f3c88 , n46604 );
buf ( R_11db0_13302748 , n46610 );
buf ( R_1470b_115413f8 , n46613 );
buf ( R_fd8e_120835d8 , n46621 );
buf ( R_142aa_102f2a68 , n46625 );
buf ( R_1267b_1056b538 , n46637 );
buf ( R_10df7_1264ae08 , n46643 );
buf ( R_b753_102ebe48 , n46653 );
buf ( R_14a47_102eeb48 , n46656 );
buf ( R_12f94_1379c068 , n46668 );
buf ( R_f3d0_1264e3c8 , n46676 );
buf ( R_13cd6_10565638 , n46684 );
buf ( R_123b1_12b3e378 , n46690 );
buf ( R_144cf_f8c96f8 , n46693 );
buf ( R_13d0c_102f6168 , n46703 );
buf ( R_13c61_12081d78 , n46713 );
buf ( R_134f6_11ce6608 , n46719 );
buf ( R_112c2_12b294b8 , n46731 );
buf ( R_11922_1056c898 , n46743 );
buf ( R_11971_1207dbd8 , n46751 );
buf ( R_138_1265b308 , n46752 );
buf ( R_d2_12654c28 , n46753 );
buf ( R_23d_12656088 , n46754 );
buf ( R_8a_1379cba8 , n46755 );
buf ( R_38ad_12048418 , n46761 );
buf ( R_7b_12651de8 , n46762 );
buf ( R_13889_10564918 , n46770 );
buf ( R_13188_12079c18 , n46776 );
buf ( R_13b8c_13a15728 , n46788 );
buf ( R_947f_1056eaf8 , n46796 );
buf ( R_1d7_12649648 , n46797 );
buf ( R_149db_102f1668 , n46800 );
buf ( R_ac1d_120826d8 , n46810 );
buf ( R_13a06_105668f8 , n46822 );
buf ( R_18f_132fc988 , n46823 );
buf ( R_180_1265fea8 , n46824 );
buf ( R_10e36_11ce6d88 , n46836 );
buf ( R_136a7_12035cb8 , n46846 );
buf ( R_148df_13a1d608 , n46849 );
buf ( R_1380f_12080838 , n46861 );
buf ( R_1485b_1265a688 , n46864 );
buf ( R_14930_102f1a28 , n46867 );
buf ( R_10044_102f1c08 , n46875 );
buf ( R_d2a3_1207bbf8 , n46883 );
buf ( R_1c0_1203c0b8 , n46884 );
buf ( R_14f_12b25778 , n46885 );
buf ( R_8472_126654e8 , n46897 );
buf ( R_1483d_11ce0d48 , n46900 );
buf ( R_12b67_11cdf3a8 , n46908 );
buf ( R_11346_12655448 , n46914 );
buf ( R_13893_12084d98 , n46926 );
buf ( R_103f0_1207ecb8 , n46932 );
buf ( R_1308d_1379eea8 , n46940 );
buf ( R_f8ce_102f10c8 , n46948 );
buf ( R_13f82_11543978 , n46956 );
buf ( R_12359_133022e8 , n46964 );
buf ( R_12cd3_13a1f728 , n46976 );
buf ( R_13546_1153efb8 , n46988 );
buf ( R_143b6_115408b8 , n47000 );
buf ( R_148e5_10568518 , n47003 );
buf ( R_10a79_11545278 , n47009 );
buf ( R_1368d_102f3be8 , n47017 );
buf ( R_14002_12047518 , n47029 );
buf ( R_febc_1207caf8 , n47041 );
buf ( R_14987_10571d98 , n47044 );
buf ( R_14894_126569e8 , n47047 );
buf ( R_13e23_102f1708 , n47055 );
buf ( R_12304_10569e18 , n47061 );
buf ( R_12daa_f8cc218 , n47073 );
buf ( R_1289e_13316128 , n47081 );
buf ( R_146ea_132fd6a8 , n47084 );
buf ( R_104_12b414d8 , n47085 );
buf ( R_e9_12055a78 , n47086 );
buf ( R_226_12652568 , n47087 );
buf ( R_20b_12656bc8 , n47088 );
buf ( R_1484c_1056c078 , n47091 );
buf ( R_149fc_12077a58 , n47094 );
buf ( R_143f0_120442b8 , n47099 );
buf ( R_107_1203f538 , n47100 );
buf ( R_208_12b260d8 , n47101 );
buf ( R_1d2_1203ce78 , n47102 );
buf ( R_1442a_102f6668 , n47106 );
buf ( R_13d_1379c568 , n47107 );
buf ( R_134be_13a19148 , n47115 );
buf ( R_145cf_13304328 , n47118 );
buf ( R_12fa4_1153e0b8 , n47124 );
buf ( R_1053d_12079858 , n47134 );
buf ( R_ee_f8c86b8 , n47135 );
buf ( R_221_12652888 , n47136 );
buf ( R_13eb5_132f7ac8 , n47144 );
buf ( R_190_133178e8 , n47145 );
buf ( R_17f_115396f8 , n47146 );
buf ( R_137af_11ce6e28 , n47152 );
buf ( R_1455a_102ed748 , n47155 );
buf ( R_10db8_102f74c8 , n47165 );
buf ( R_ab_1264cde8 , n47166 );
buf ( R_1187e_12077698 , n47178 );
buf ( R_5a_126653a8 , n47179 );
buf ( R_7e57_13a1a188 , n47187 );
buf ( R_146ed_1153a238 , n47190 );
buf ( R_1b0_12b29918 , n47191 );
buf ( R_15f_1265f188 , n47192 );
buf ( R_138b8_1264a368 , n47200 );
buf ( R_13bd6_102f9188 , n47208 );
buf ( R_14a17_102f0ee8 , n47211 );
buf ( R_143a6_133121a8 , n47223 );
buf ( R_11f57_12649328 , n47231 );
buf ( R_14972_13302608 , n47234 );
buf ( R_10701_1207f1b8 , n47240 );
buf ( R_14503_1203e3b8 , n47243 );
buf ( R_a4_12b36e98 , n47244 );
buf ( R_6a_12b40178 , n47245 );
buf ( R_aeba_105624d8 , n47253 );
buf ( R_1379b_11ce6ec8 , n47261 );
buf ( R_134e2_13a1e3c8 , n47267 );
buf ( R_10973_12663008 , n47273 );
buf ( R_11c66_102f7ba8 , n47279 );
buf ( R_1325f_126468a8 , n47285 );
buf ( R_1327d_10570d58 , n47293 );
buf ( R_13417_102f3968 , n47301 );
buf ( R_101_1264f048 , n47302 );
buf ( R_95_133017a8 , n47303 );
buf ( R_20e_1265e788 , n47304 );
buf ( R_13c59_105b5638 , n47316 );
buf ( R_13ca1_12652f68 , n47324 );
buf ( R_1481c_11cdb988 , n47327 );
buf ( R_14611_11545458 , n47330 );
buf ( R_12fae_102f7388 , n47342 );
buf ( R_1469f_1207d138 , n47345 );
buf ( R_142dd_13314828 , n47352 );
buf ( R_1279d_12079fd8 , n47360 );
buf ( R_12646_1056b2b8 , n47368 );
buf ( R_11486_102ee788 , n47378 );
buf ( R_13389_1207fb18 , n47384 );
buf ( R_1492d_11ce64c8 , n47387 );
buf ( R_12d46_12648928 , n47395 );
buf ( R_145b7_12b3d5b8 , n47398 );
buf ( R_b211_12048c38 , n47406 );
buf ( R_143aa_13795c68 , n47418 );
buf ( R_1110c_11cdc928 , n47426 );
buf ( R_1a5_12b3c618 , n47427 );
buf ( R_16a_137a1248 , n47428 );
buf ( R_df67_1207b8d8 , n47440 );
buf ( R_124f6_1264f2c8 , n47450 );
buf ( R_12b54_102f2248 , n47458 );
buf ( R_d7dc_13a17de8 , n47464 );
buf ( R_1247b_11ce4808 , n47470 );
buf ( R_149ea_11540598 , n47473 );
buf ( R_10a_12b30678 , n47474 );
buf ( R_13c77_13a1cc08 , n47480 );
buf ( R_205_12653dc8 , n47481 );
buf ( R_14753_1264efa8 , n47484 );
buf ( R_191_12043d18 , n47485 );
buf ( R_17e_132f8568 , n47486 );
buf ( R_11c4b_13a15c28 , n47492 );
buf ( R_13208_11542758 , n47498 );
buf ( R_e0ad_133021a8 , n47504 );
buf ( R_11a3f_12b3e9b8 , n47510 );
buf ( R_1230e_f8cb598 , n47520 );
buf ( R_eee_1056adb8 , n47522 );
buf ( R_14444_12648108 , n47525 );
buf ( R_1dc_11538d98 , n47526 );
buf ( R_12b7a_1264f188 , n47538 );
buf ( R_133_13313888 , n47539 );
buf ( R_147b1_105b5a98 , n47542 );
buf ( R_f116_11ce1068 , n47550 );
buf ( R_13a5c_1379a268 , n47560 );
buf ( R_14340_12078458 , n47571 );
buf ( R_e522_1330ed28 , n47581 );
buf ( R_146f0_1153da78 , n47584 );
buf ( R_136f4_12649148 , n47592 );
buf ( R_119e8_1153e798 , n47600 );
buf ( R_1391b_12b277f8 , n47612 );
buf ( R_fd37_120394f8 , n47620 );
buf ( R_1461d_11539dd8 , n47623 );
buf ( R_ee50_102eb9e8 , n47629 );
buf ( R_dd_132f61c8 , n47630 );
buf ( R_232_105afa58 , n47631 );
buf ( R_4c_12652b08 , n47632 );
buf ( R_135a0_1153f0f8 , n47644 );
buf ( R_125d0_12b3f6d8 , n47654 );
buf ( R_b4_13302988 , n47655 );
buf ( R_51_13309648 , n47656 );
buf ( R_f925_12048b98 , n47664 );
buf ( R_14034_f8cf198 , n47670 );
buf ( R_123e9_f8c0eb8 , n47676 );
buf ( R_14726_1203bc58 , n47679 );
buf ( R_10894_1153ad78 , n47687 );
buf ( R_1b9_1379b7a8 , n47688 );
buf ( R_156_137927e8 , n47689 );
buf ( R_1471a_1379da08 , n47692 );
buf ( R_13d4e_11544f58 , n47700 );
buf ( R_112ae_115429d8 , n47708 );
buf ( R_dcb0_10564e18 , n47714 );
buf ( R_13ae3_12083498 , n47722 );
buf ( R_11a90_13a1ba88 , n47728 );
buf ( R_13f1a_10566998 , n47736 );
buf ( R_fdd5_1264d068 , n47742 );
buf ( R_13acb_13a17988 , n47750 );
buf ( R_ef1_13a16ee8 , n47752 );
buf ( R_145e1_12b40d58 , n47755 );
buf ( R_14915_102f7748 , n47758 );
buf ( R_ed3c_120760b8 , n47766 );
buf ( R_13cdc_11542398 , n47776 );
buf ( R_f544_102f5d08 , n47788 );
buf ( R_147e7_13793fa8 , n47791 );
buf ( R_e4_133095a8 , n47792 );
buf ( R_8d_1153d078 , n47793 );
buf ( R_78_12044178 , n47794 );
buf ( R_22b_12b3b538 , n47795 );
buf ( R_128ff_105b6178 , n47801 );
buf ( R_148ac_102f0f88 , n47804 );
buf ( R_1e9_133208a8 , n47805 );
buf ( R_192_12b44a98 , n47806 );
buf ( R_17d_12661f28 , n47807 );
buf ( R_12b83_13305e08 , n47813 );
buf ( R_fbb3_10567078 , n47821 );
buf ( R_126_12660588 , n47822 );
buf ( R_cfc6_1264a868 , n47834 );
buf ( R_1492a_13a1e1e8 , n47837 );
buf ( R_116bb_1207d6d8 , n47845 );
buf ( R_144d8_1330d9c8 , n47848 );
buf ( R_e6f2_102ecc08 , n47860 );
buf ( R_14a14_1207bdd8 , n47863 );
buf ( R_10f70_11544a58 , n47871 );
buf ( R_119fa_1207f2f8 , n47879 );
buf ( R_cef5_1265b6c8 , n47885 );
buf ( R_115b3_12082458 , n47893 );
buf ( R_211_1265c028 , n47894 );
buf ( R_146cc_11542618 , n47897 );
buf ( R_fe_120448f8 , n47898 );
buf ( R_119df_1056bad8 , n47904 );
buf ( R_13787_11ce21e8 , n47914 );
buf ( R_147dd_11ce6068 , n47917 );
buf ( R_14695_11cdf8a8 , n47920 );
buf ( R_149b1_102fa128 , n47923 );
buf ( R_110af_1379aee8 , n47929 );
buf ( R_14560_1330b3a8 , n47932 );
buf ( R_143ff_11cdca68 , n47936 );
buf ( R_d4_12654a48 , n47937 );
buf ( R_23b_13799408 , n47938 );
buf ( R_1c7_132fc0c8 , n47939 );
buf ( R_148_105aacd8 , n47940 );
buf ( R_13d6d_13a17668 , n47946 );
buf ( R_ce64_1056f9f8 , n47954 );
buf ( R_14474_13307a28 , n47957 );
buf ( R_12bde_102f62a8 , n47967 );
buf ( R_1436a_102eefa8 , n47979 );
buf ( R_14957_11540db8 , n47982 );
buf ( R_b634_11cdc068 , n47994 );
buf ( R_1460e_11ce2dc8 , n47997 );
buf ( R_f24f_11ce2fa8 , n48003 );
buf ( R_13763_105679d8 , n48011 );
buf ( R_f0b2_102f7f68 , n48019 );
buf ( R_14620_11ce6108 , n48022 );
buf ( R_131f5_12084618 , n48034 );
buf ( R_1490f_12651e88 , n48037 );
buf ( R_136cc_1264fcc8 , n48045 );
buf ( R_f227_1207a398 , n48053 );
buf ( R_13959_1153f918 , n48061 );
buf ( R_142cf_12659aa8 , n48070 );
buf ( R_f6b2_11cdfb28 , n48076 );
buf ( R_1ed_1203f5d8 , n48077 );
buf ( R_a2f6_11cdb3e8 , n48083 );
buf ( R_fc5e_13a18888 , n48089 );
buf ( R_122_12663d28 , n48090 );
buf ( R_13f67_12083b78 , n48098 );
buf ( R_13740_11cdb348 , n48104 );
buf ( R_146c9_1153fd78 , n48107 );
buf ( R_145db_13a12b68 , n48110 );
buf ( R_101ae_13a1fae8 , n48122 );
buf ( R_bb03_12b29ff8 , n48128 );
buf ( R_1101b_12045f38 , n48136 );
buf ( R_12bfd_10564b98 , n48142 );
buf ( R_121a5_1056a138 , n48148 );
buf ( R_127df_1330a728 , n48154 );
buf ( R_11617_105656d8 , n48160 );
buf ( R_13f90_12080518 , n48166 );
buf ( R_13be9_12662388 , n48178 );
buf ( R_12760_1331ab88 , n48188 );
buf ( R_126bb_10563b58 , n48194 );
buf ( R_147c6_12081cd8 , n48197 );
buf ( R_21c_12b41398 , n48198 );
buf ( R_13b33_102f0588 , n48206 );
buf ( R_1f8_132f5fe8 , n48207 );
buf ( R_11d2f_105665d8 , n48215 );
buf ( R_1227d_1265f2c8 , n48221 );
buf ( R_11a35_102f44a8 , n48227 );
buf ( R_1479c_1056c758 , n48230 );
buf ( R_116e4_12659828 , n48238 );
buf ( R_14662_1207ceb8 , n48241 );
buf ( R_14515_12079ad8 , n48244 );
buf ( R_117_12650c68 , n48245 );
buf ( R_115ca_11ce5fc8 , n48251 );
buf ( R_f3_1379bde8 , n48252 );
buf ( R_e229_102ecca8 , n48260 );
buf ( R_202_12b3f098 , n48261 );
buf ( R_1e5_1203a218 , n48262 );
buf ( R_12a_1331fea8 , n48263 );
buf ( R_10d_1330bda8 , n48264 );
buf ( R_135d6_1056fef8 , n48272 );
buf ( R_14918_13a1d888 , n48275 );
buf ( R_1452a_10564378 , n48278 );
buf ( R_14984_1056bc18 , n48281 );
buf ( R_1cd_1265c8e8 , n48282 );
buf ( R_eb34_11cda628 , n48294 );
buf ( R_125ac_11ce4308 , n48302 );
buf ( R_193_f8c7cb8 , n48303 );
buf ( R_1216d_1264d7e8 , n48315 );
buf ( R_17c_132fe648 , n48316 );
buf ( R_142_13792ce8 , n48317 );
buf ( R_cdb8_102f4f48 , n48325 );
buf ( R_144bd_11cdeb88 , n48328 );
buf ( R_131ae_1056bd58 , n48334 );
buf ( R_14909_1379f768 , n48337 );
buf ( R_14924_12b3adb8 , n48340 );
buf ( R_102a2_12b41e38 , n48350 );
buf ( R_13aa8_120525f8 , n48358 );
buf ( R_d3ca_102ef7c8 , n48364 );
buf ( R_1459f_120792b8 , n48367 );
buf ( R_120b3_12b407b8 , n48373 );
buf ( R_127a7_105683d8 , n48385 );
buf ( R_14545_1056b218 , n48388 );
buf ( R_12056_1204f178 , n48396 );
buf ( R_11f2a_10563ab8 , n48404 );
buf ( R_e021_12b26718 , n48410 );
buf ( R_f377_1056d1f8 , n48418 );
buf ( R_127ca_13a16da8 , n48424 );
buf ( R_14689_120838f8 , n48427 );
buf ( R_11be7_1207a6b8 , n48435 );
buf ( R_139a1_1264c668 , n48441 );
buf ( R_14536_12b42978 , n48444 );
buf ( R_13c2d_11cdd828 , n48456 );
buf ( R_14906_11544ff8 , n48459 );
buf ( R_11a5d_132f52c8 , n48465 );
buf ( R_ca63_1331c8e8 , n48473 );
buf ( R_14714_102f77e8 , n48476 );
buf ( R_14799_137933c8 , n48479 );
buf ( R_1390f_13a14828 , n48487 );
buf ( R_1234f_12083858 , n48495 );
buf ( R_142c6_12081738 , n48502 );
buf ( R_127ae_12b3ccf8 , n48510 );
buf ( R_13590_12079a38 , n48516 );
buf ( R_148b8_102eaa48 , n48519 );
buf ( R_5735_137a0988 , n48525 );
buf ( R_1a6_12038698 , n48526 );
buf ( R_169_1203e458 , n48527 );
buf ( R_127c1_12082638 , n48533 );
buf ( R_1288a_137a1ec8 , n48541 );
buf ( R_1488e_102f6708 , n48544 );
buf ( R_113b9_1264ea08 , n48554 );
buf ( R_1430f_11cd8fa8 , n48562 );
buf ( R_f97f_13304dc8 , n48568 );
buf ( R_104fa_120761f8 , n48574 );
buf ( R_119ae_11cdfa88 , n48580 );
buf ( R_12c78_1207ca58 , n48590 );
buf ( R_d606_11ce46c8 , n48598 );
buf ( R_146a5_102f90e8 , n48601 );
buf ( R_14900_120781d8 , n48604 );
buf ( R_1374f_13a16808 , n48610 );
buf ( R_ff3c_11ce1f68 , n48618 );
buf ( R_e834_10564238 , n48624 );
buf ( R_14a5e_105aa4b8 , n48628 );
buf ( R_13465_13316bc8 , n48638 );
buf ( R_13d25_11540b38 , n48648 );
buf ( R_56_13308248 , n48649 );
buf ( R_ef7_1153e838 , n48651 );
buf ( R_13193_102ec7a8 , n48657 );
buf ( R_132f1_13a145a8 , n48665 );
buf ( R_1291e_1056ee18 , n48671 );
buf ( R_14921_105640f8 , n48674 );
buf ( R_1371a_12083fd8 , n48680 );
buf ( R_14837_132f32e8 , n48683 );
buf ( R_13a37_12b3d338 , n48695 );
buf ( R_dad2_1379c6a8 , n48701 );
buf ( R_1495d_12b43878 , n48704 );
buf ( R_149f3_12b27c58 , n48707 );
buf ( R_107c6_1203f998 , n48713 );
buf ( R_1456c_12b437d8 , n48716 );
buf ( R_11888_13794868 , n48724 );
buf ( R_13b62_13a13428 , n48730 );
buf ( R_1360f_10563158 , n48742 );
buf ( R_1b1_12657ac8 , n48743 );
buf ( R_10844_1153e1f8 , n48753 );
buf ( R_194_1331d4c8 , n48754 );
buf ( R_17b_1265ea08 , n48755 );
buf ( R_15e_126544a8 , n48756 );
buf ( R_be25_102ec028 , n48762 );
buf ( R_148fd_102eb768 , n48765 );
buf ( R_14683_13a1d9c8 , n48768 );
buf ( R_a069_12080298 , n48776 );
buf ( R_1233a_13a143c8 , n48784 );
buf ( R_6e_13304b48 , n48785 );
buf ( R_1334f_1204e598 , n48791 );
buf ( R_121e7_1207ff78 , n48797 );
buf ( R_12bb7_102f3e68 , n48809 );
buf ( R_12bcc_12652608 , n48815 );
buf ( R_f783_13797b08 , n48823 );
buf ( R_14680_12076fb8 , n48826 );
buf ( R_13d2b_12085338 , n48836 );
buf ( R_11bbe_1153de38 , n48844 );
buf ( R_148e8_1264bda8 , n48847 );
buf ( R_148fa_102f5948 , n48850 );
buf ( R_149d8_132fc168 , n48853 );
buf ( R_148ee_120808d8 , n48856 );
buf ( R_148f4_11cd8468 , n48859 );
buf ( R_ff98_12b41618 , n48865 );
buf ( R_13bc3_102f8d28 , n48873 );
buf ( R_12b1f_120564d8 , n48881 );
buf ( R_c961_12080f18 , n48889 );
buf ( R_214_12655588 , n48890 );
buf ( R_dff5_102ed9c8 , n48900 );
buf ( R_13d49_13a16bc8 , n48908 );
buf ( R_fb_1379f808 , n48909 );
buf ( R_12958_102f1848 , n48921 );
buf ( R_12220_1379e908 , n48927 );
buf ( R_144de_12076798 , n48930 );
buf ( R_c6d1_10566178 , n48942 );
buf ( R_11547_1264cc08 , n48948 );
buf ( R_138ac_102eb128 , n48960 );
buf ( R_12853_105b58b8 , n48970 );
buf ( R_1f1_12655268 , n48971 );
buf ( R_11e_12b29b98 , n48972 );
buf ( R_13d30_1207b658 , n48982 );
buf ( R_b2_105aa0f8 , n48983 );
buf ( R_d5a1_105690f8 , n48991 );
buf ( R_c700_13304788 , n48997 );
buf ( R_a359_12662888 , n49003 );
buf ( R_1449f_12055898 , n49006 );
buf ( R_14587_10565ef8 , n49009 );
buf ( R_14759_1056e378 , n49012 );
buf ( R_1385d_1056ab38 , n49018 );
buf ( R_1401f_132fb588 , n49026 );
buf ( R_1245b_12658f68 , n49034 );
buf ( R_fe3a_11cdb168 , n49042 );
buf ( R_a47d_13a18f68 , n49048 );
buf ( R_145ea_1056c438 , n49051 );
buf ( R_99a4_102f5bc8 , n49059 );
buf ( R_1491e_12661528 , n49062 );
buf ( R_1c1_126618e8 , n49063 );
buf ( R_b180_12039a98 , n49075 );
buf ( R_14e_12b29e18 , n49076 );
buf ( R_13b1f_12052c38 , n49086 );
buf ( R_146e4_f8cb638 , n49089 );
buf ( R_14581_10571b18 , n49092 );
buf ( R_1354d_12040078 , n49100 );
buf ( R_13508_120842f8 , n49106 );
buf ( R_148d9_13a14d28 , n49109 );
buf ( R_149c0_102ed068 , n49112 );
buf ( R_1477e_10568fb8 , n49115 );
buf ( R_14735_105680b8 , n49118 );
buf ( R_13d35_11ce1108 , n49126 );
buf ( R_4d49_102f8dc8 , n49132 );
buf ( R_133aa_11545b38 , n49140 );
buf ( R_14518_102f67a8 , n49143 );
buf ( R_bf1d_1153d618 , n49155 );
buf ( R_a9_1204d4b8 , n49156 );
buf ( R_14702_12b3d0b8 , n49159 );
buf ( R_1431c_11cde188 , n49168 );
buf ( R_9323_1331d068 , n49174 );
buf ( R_14a2f_12075ed8 , n49177 );
buf ( R_1e1_13321ca8 , n49178 );
buf ( R_12e_105af9b8 , n49179 );
buf ( R_9d_1379c9c8 , n49180 );
buf ( R_12caa_126508a8 , n49188 );
buf ( R_115df_10566c18 , n49196 );
buf ( R_144fd_102f1b68 , n49199 );
buf ( R_127f1_12b2a098 , n49207 );
buf ( R_137eb_12082138 , n49215 );
buf ( R_11b9a_12b3f278 , n49223 );
buf ( R_1483a_12081f58 , n49226 );
buf ( R_7d2b_11ce4948 , n49232 );
buf ( R_13a49_102f8e68 , n49242 );
buf ( R_1493c_11cdc568 , n49245 );
buf ( R_14a3e_102ed428 , n49248 );
buf ( R_195_12045cb8 , n49249 );
buf ( R_14489_12b3fe58 , n49252 );
buf ( R_17a_1330dc48 , n49253 );
buf ( R_1066b_1264a228 , n49259 );
buf ( R_139b5_11536318 , n49265 );
buf ( R_12775_126513e8 , n49271 );
buf ( R_13d43_13a1c168 , n49279 );
buf ( R_13e78_1056a598 , n49285 );
buf ( R_90_f8cccb8 , n49286 );
buf ( R_75_12b443b8 , n49287 );
buf ( R_14816_10565db8 , n49290 );
buf ( R_e4c7_10571398 , n49302 );
buf ( R_14354_13317348 , n49313 );
buf ( R_146c3_12b3bfd8 , n49316 );
buf ( R_db95_12b2ff98 , n49322 );
buf ( R_b45b_11ce7508 , n49328 );
buf ( R_145de_1056b5d8 , n49331 );
buf ( R_13c7d_1056d798 , n49337 );
buf ( R_c7c0_102ed4c8 , n49352 );
buf ( R_1ff_13315c28 , n49353 );
buf ( R_1361a_102f01c8 , n49359 );
buf ( R_110_1204b938 , n49360 );
buf ( R_10c17_13a13888 , n49370 );
buf ( R_d6_1264b1c8 , n49371 );
buf ( R_239_12b2a958 , n49372 );
buf ( R_144a8_115369f8 , n49375 );
buf ( R_12516_13305188 , n49383 );
buf ( R_14699_10567e38 , n49386 );
buf ( R_12de4_12045b18 , n49392 );
buf ( R_10fd9_11ce1928 , n49400 );
buf ( R_145c6_13a1cb68 , n49403 );
buf ( R_147c3_13a177a8 , n49406 );
buf ( R_1313e_1207a1b8 , n49414 );
buf ( R_e9a6_1153dcf8 , n49420 );
buf ( R_123a6_12077418 , n49432 );
buf ( R_e669_1056eb98 , n49438 );
buf ( R_eea5_13793c88 , n49444 );
buf ( R_8e12_f8c7538 , n49452 );
buf ( R_11a2c_12b3f1d8 , n49462 );
buf ( R_bc89_12664548 , n49470 );
buf ( R_b132_13300a88 , n49478 );
buf ( R_14626_102f4ae8 , n49481 );
buf ( R_125c9_11ce5c08 , n49487 );
buf ( R_14891_1265e0a8 , n49490 );
buf ( R_13ba9_1056f4f8 , n49502 );
buf ( R_11299_1056a4f8 , n49510 );
buf ( R_1395f_1207ba18 , n49522 );
buf ( R_1085f_13312a28 , n49532 );
buf ( R_c642_12b41b18 , n49538 );
buf ( R_1445c_f8ce478 , n49541 );
buf ( R_14981_12b3f598 , n49544 );
buf ( R_148e2_12650b28 , n49547 );
buf ( R_988f_13a1e968 , n49559 );
buf ( R_962b_105647d8 , n49571 );
buf ( R_124a7_12079498 , n49583 );
buf ( R_fe64_1153f378 , n49593 );
buf ( R_11f16_102eb088 , n49601 );
buf ( R_13e03_1379bf28 , n49609 );
buf ( R_14927_11cdf808 , n49612 );
buf ( R_1ba_1330eb48 , n49613 );
buf ( R_14471_13793be8 , n49616 );
buf ( R_121fd_11ce3048 , n49622 );
buf ( R_14499_1207a9d8 , n49625 );
buf ( R_155_12b43f58 , n49626 );
buf ( R_98_12048af8 , n49627 );
buf ( R_e916_105699b8 , n49635 );
buf ( R_e1ea_1056b998 , n49645 );
buf ( R_11af3_13793788 , n49651 );
buf ( R_13bcf_12650948 , n49657 );
buf ( R_10070_12077e18 , n49663 );
buf ( R_f2f6_126613e8 , n49671 );
buf ( R_104a3_11542d98 , n49677 );
buf ( R_149ae_10565138 , n49680 );
buf ( R_1430b_1204c8d8 , n49687 );
buf ( R_ede8_1056dfb8 , n49693 );
buf ( R_13495_13a1e008 , n49701 );
buf ( R_df_132f6808 , n49702 );
buf ( R_230_12664a48 , n49703 );
buf ( R_136ac_102eacc8 , n49713 );
buf ( R_dd20_137974c8 , n49721 );
buf ( R_14741_132f2c08 , n49724 );
buf ( R_137c1_11543dd8 , n49730 );
buf ( R_14364_11ce6568 , n49738 );
buf ( R_11d60_132fc8e8 , n49744 );
buf ( R_14a44_105b60d8 , n49747 );
buf ( R_13749_11543518 , n49755 );
buf ( R_854a_1207fed8 , n49761 );
buf ( R_14a11_12045a78 , n49764 );
buf ( R_1a7_12659b48 , n49765 );
buf ( R_168_105b3158 , n49766 );
buf ( R_f03_13a17208 , n49768 );
buf ( R_1274c_12653fa8 , n49778 );
buf ( R_147b7_12079df8 , n49781 );
buf ( R_a2_1379e228 , n49782 );
buf ( R_63_f8c7b78 , n49783 );
buf ( R_13c49_102ecac8 , n49789 );
buf ( R_d68f_12078a98 , n49797 );
buf ( R_148f1_11cde688 , n49800 );
buf ( R_196_11536778 , n49801 );
buf ( R_179_13301c08 , n49802 );
buf ( R_11c1b_120757f8 , n49808 );
buf ( R_1181a_10565098 , n49814 );
buf ( R_14912_13300628 , n49817 );
buf ( R_10c93_13310768 , n49827 );
buf ( R_147f2_10571618 , n49830 );
buf ( R_c832_12075f78 , n49836 );
buf ( R_14530_11540778 , n49839 );
buf ( R_e8ba_11ce3b88 , n49845 );
buf ( R_14903_11ce50c8 , n49848 );
buf ( R_14629_115412b8 , n49851 );
buf ( R_11966_10562118 , n49859 );
buf ( R_f8fa_105b4d78 , n49865 );
buf ( R_1d8_1331f5e8 , n49866 );
buf ( R_1281b_1207f6b8 , n49872 );
buf ( R_137_1331a7c8 , n49873 );
buf ( R_5f_12b428d8 , n49874 );
buf ( R_12288_126495a8 , n49880 );
buf ( R_a469_13a14648 , n49888 );
buf ( R_130cc_13a17348 , n49896 );
buf ( R_136e6_11cdcb08 , n49906 );
buf ( R_d806_102f5a88 , n49914 );
buf ( R_fd98_12052d78 , n49922 );
buf ( R_144b4_1153eab8 , n49925 );
buf ( R_1482b_12b3b3f8 , n49928 );
buf ( R_13858_12081e18 , n49934 );
buf ( R_1d3_1265ae08 , n49935 );
buf ( R_13c_1265b1c8 , n49936 );
buf ( R_14596_12048558 , n49939 );
buf ( R_eb_1153bf98 , n49940 );
buf ( R_224_12b29698 , n49941 );
buf ( R_13d3c_132f70c8 , n49947 );
buf ( R_c353_102f31e8 , n49953 );
buf ( R_1092e_13a140a8 , n49959 );
buf ( R_1018e_10563478 , n49971 );
buf ( R_12875_1153eb58 , n49979 );
buf ( R_13693_13795448 , n49985 );
buf ( R_123bb_11ce7008 , n49991 );
buf ( R_dfc9_12647208 , n49997 );
buf ( R_da6d_12082098 , n50003 );
buf ( R_1198e_1153d758 , n50013 );
buf ( R_149ff_1264c848 , n50016 );
buf ( R_1180e_12648248 , n50026 );
buf ( R_12535_126604e8 , n50036 );
buf ( R_12780_10568b58 , n50042 );
buf ( R_9dc0_102f6f28 , n50050 );
buf ( R_c4a7_1330a908 , n50062 );
buf ( R_11bfb_12649968 , n50070 );
buf ( R_13fe4_105622f8 , n50078 );
buf ( R_12e0c_13797388 , n50086 );
buf ( R_1454e_11ce1c48 , n50089 );
buf ( R_14069_1153db18 , n50091 );
buf ( R_10c0e_120464d8 , n50097 );
buf ( R_13c1f_f8c8938 , n50103 );
buf ( R_d910_1056e418 , n50109 );
buf ( R_cfae_13a15368 , n50115 );
buf ( R_10806_1264d608 , n50121 );
buf ( R_13706_13319b48 , n50133 );
buf ( R_12e21_1330cb68 , n50143 );
buf ( R_f8_12665808 , n50144 );
buf ( R_67_105aac38 , n50145 );
buf ( R_217_105b3fb8 , n50146 );
buf ( R_12a8e_1264ef08 , n50152 );
buf ( R_e5ea_115436f8 , n50158 );
buf ( R_14858_10571c58 , n50161 );
buf ( R_111b8_102ebbc8 , n50169 );
buf ( R_12ba4_12b28ab8 , n50177 );
buf ( R_108f1_102f35a8 , n50185 );
buf ( R_138a5_1264e468 , n50195 );
buf ( R_131ff_13a1eaa8 , n50201 );
buf ( R_11448_11ce41c8 , n50207 );
buf ( R_11534_13a13ce8 , n50213 );
buf ( R_12d1d_1207c238 , n50221 );
buf ( R_134e8_13a1e8c8 , n50227 );
buf ( R_b82e_1153c2b8 , n50237 );
buf ( R_11572_11ce43a8 , n50245 );
buf ( R_14897_1265c988 , n50248 );
buf ( R_125fa_1265b128 , n50256 );
buf ( R_b95d_102f8008 , n50264 );
buf ( R_14436_10570718 , n50268 );
buf ( R_f951_132fcde8 , n50274 );
buf ( R_10246_1056ae58 , n50282 );
buf ( R_12041_11ce0ac8 , n50288 );
buf ( R_138cd_1153e018 , n50294 );
buf ( R_1b2_12660f88 , n50295 );
buf ( R_197_1379a768 , n50296 );
buf ( R_121dd_12659328 , n50302 );
buf ( R_178_12658d88 , n50303 );
buf ( R_15d_133195a8 , n50304 );
buf ( R_13f24_13318428 , n50310 );
buf ( R_146f6_132fbc68 , n50313 );
buf ( R_b880_12083d58 , n50319 );
buf ( R_12ab4_132f57c8 , n50325 );
buf ( R_ed14_133110c8 , n50331 );
buf ( R_144f0_132ff0e8 , n50334 );
buf ( R_10aa5_12053f98 , n50340 );
buf ( R_1290a_11ce1388 , n50346 );
buf ( R_9d4e_11cddbe8 , n50352 );
buf ( R_e6_12b344f8 , n50353 );
buf ( R_b0_12b3f458 , n50354 );
buf ( R_229_126659e8 , n50355 );
buf ( R_12b3f_105b6538 , n50361 );
buf ( R_1f5_1203e958 , n50362 );
buf ( R_f624_1265b808 , n50370 );
buf ( R_14711_11ce2828 , n50373 );
buf ( R_fe05_102f9548 , n50379 );
buf ( R_1118b_11cdb8e8 , n50385 );
buf ( R_1c8_f8c6b38 , n50386 );
buf ( R_147_12b38c98 , n50387 );
buf ( R_11a_1204b438 , n50388 );
buf ( R_14778_13a1f688 , n50391 );
buf ( R_137fd_11544418 , n50397 );
buf ( R_f0_13795d08 , n50398 );
buf ( R_c3_132ff188 , n50399 );
buf ( R_21f_1265a2c8 , n50400 );
buf ( R_12e60_132f3a68 , n50410 );
buf ( R_4a02_12646e48 , n50416 );
buf ( R_c5_12657e88 , n50417 );
buf ( R_132ae_1056ef58 , n50423 );
buf ( R_d400_133126a8 , n50435 );
buf ( R_128a8_f8c9978 , n50441 );
buf ( R_ecbd_12040a78 , n50449 );
buf ( R_146ba_11cd8c88 , n50452 );
buf ( R_ea59_102f5088 , n50462 );
buf ( R_1183a_1204a498 , n50472 );
buf ( R_13d1f_1207ddb8 , n50478 );
buf ( R_136e0_11ce7148 , n50490 );
buf ( R_ddb7_12078b38 , n50496 );
buf ( R_14575_13307c08 , n50499 );
buf ( R_14864_13a1b768 , n50502 );
buf ( R_1471d_12040bb8 , n50505 );
buf ( R_11237_1056f958 , n50511 );
buf ( R_13fee_12663288 , n50517 );
buf ( R_c1_1204fd58 , n50518 );
buf ( R_14632_11cd85a8 , n50521 );
buf ( R_4d_12662d88 , n50522 );
buf ( R_b895_1264a4a8 , n50528 );
buf ( R_11b87_12648b08 , n50538 );
buf ( R_111c4_12076658 , n50546 );
buf ( R_a534_12b3d018 , n50552 );
buf ( R_11805_12b41578 , n50558 );
buf ( R_c901_126603a8 , n50566 );
buf ( R_13bde_13a1bbc8 , n50572 );
buf ( R_149b4_10564d78 , n50575 );
buf ( R_c7_126589c8 , n50576 );
buf ( R_248_1331ef08 , n50577 );
buf ( R_5b_12655088 , n50578 );
buf ( R_13720_102f3f08 , n50586 );
buf ( R_b9b1_1056c9d8 , n50592 );
buf ( R_f1cc_10567ed8 , n50598 );
buf ( R_cd0b_11542f78 , n50604 );
buf ( R_1497b_11cdfda8 , n50607 );
buf ( R_12d6f_13799b88 , n50613 );
buf ( R_14305_120844d8 , n50620 );
buf ( R_145ae_102efe08 , n50623 );
buf ( R_147d6_12b27b18 , n50626 );
buf ( R_13dc3_11cdbf28 , n50632 );
buf ( R_dc22_1153d438 , n50638 );
buf ( R_5970_11cdbe88 , n50644 );
buf ( R_113_1265c528 , n50645 );
buf ( R_82_f8cbc78 , n50646 );
buf ( R_1fc_12050078 , n50647 );
buf ( R_b00a_1153e658 , n50653 );
buf ( R_1346e_10567bb8 , n50661 );
buf ( R_1dd_12b395f8 , n50662 );
buf ( R_10390_1207ed58 , n50668 );
buf ( R_12cf4_13310ee8 , n50674 );
buf ( R_10675_1203cab8 , n50680 );
buf ( R_1399b_1264c3e8 , n50686 );
buf ( R_132_120518d8 , n50687 );
buf ( R_d8_12b3c938 , n50688 );
buf ( R_237_105a9fb8 , n50689 );
buf ( R_d4b2_1265bda8 , n50697 );
buf ( R_14453_12649d28 , n50700 );
buf ( R_10e2c_102ecde8 , n50706 );
buf ( R_52_13799868 , n50707 );
buf ( R_143dc_120824f8 , n50712 );
buf ( R_13ebe_11ce4128 , n50720 );
buf ( R_14053_102f21a8 , n50726 );
buf ( R_10960_133050e8 , n50734 );
buf ( R_1037b_1264a048 , n50740 );
buf ( R_7fe6_12b3f638 , n50748 );
buf ( R_12685_11cdf088 , n50754 );
buf ( R_135e9_11ce0de8 , n50762 );
buf ( R_bf_1379fa88 , n50763 );
buf ( R_85_12b41898 , n50764 );
buf ( R_149d5_11541358 , n50767 );
buf ( R_13f4d_10561fd8 , n50773 );
buf ( R_d0f1_1056a1d8 , n50779 );
buf ( R_a3f3_12646da8 , n50787 );
buf ( R_1311d_13a131a8 , n50795 );
buf ( R_1026e_11541ad8 , n50801 );
buf ( R_139de_13310588 , n50807 );
buf ( R_144cc_11ce23c8 , n50810 );
buf ( R_1403a_1331cc08 , n50818 );
buf ( R_1ce_12656628 , n50819 );
buf ( R_198_12b3fdb8 , n50820 );
buf ( R_d37f_1379a1c8 , n50828 );
buf ( R_177_1330de28 , n50829 );
buf ( R_141_12b3cf78 , n50830 );
buf ( R_14500_102f92c8 , n50833 );
buf ( R_c9_12b28fb8 , n50834 );
buf ( R_246_1203df58 , n50835 );
buf ( R_93_12659be8 , n50836 );
buf ( R_72_132fe788 , n50837 );
buf ( R_125bf_105685b8 , n50843 );
buf ( R_1a8_137a0d48 , n50844 );
buf ( R_147a5_1264a728 , n50847 );
buf ( R_167_1204f678 , n50848 );
buf ( R_7f_105ac998 , n50849 );
buf ( R_149f0_13a1fea8 , n50852 );
buf ( R_12210_13793aa8 , n50860 );
buf ( R_13db7_11ce11a8 , n50866 );
buf ( R_100e9_132f3ec8 , n50872 );
buf ( R_5362_13a18108 , n50878 );
buf ( R_124d7_13a18e28 , n50884 );
buf ( R_14a55_133001c8 , n50888 );
buf ( R_12419_1153d398 , n50894 );
buf ( R_108b6_1264e0a8 , n50900 );
buf ( R_10d4d_11cded68 , n50906 );
buf ( R_1464a_13a15b88 , n50909 );
buf ( R_c7f2_11cdc748 , n50915 );
buf ( R_13c83_11544698 , n50921 );
buf ( R_1489a_f8c6c78 , n50924 );
buf ( R_125b6_12040b18 , n50930 );
buf ( R_c00b_12079718 , n50936 );
buf ( R_eeb_13a13608 , n50942 );
buf ( R_f088_1330ba88 , n50948 );
buf ( R_1365e_1207b838 , n50956 );
buf ( R_fa81_12052198 , n50962 );
buf ( R_145f3_13a14788 , n50965 );
buf ( R_10995_102f3148 , n50973 );
buf ( R_123f8_13a13388 , n50979 );
buf ( R_6358_1204fe98 , n50987 );
buf ( R_14763_11ce4c68 , n50990 );
buf ( R_1433c_12077c38 , n51001 );
buf ( R_dde7_13a141e8 , n51007 );
buf ( R_13ef9_1204a858 , n51013 );
buf ( R_14810_1056db58 , n51016 );
buf ( R_13fdc_102f15c8 , n51024 );
buf ( R_d995_11ce0fc8 , n51030 );
buf ( R_117fc_12056078 , n51036 );
buf ( R_8d57_11ce53e8 , n51042 );
buf ( R_11bb4_12b39cd8 , n51048 );
buf ( R_13b97_1207a438 , n51058 );
buf ( R_14068_11cdc108 , n51060 );
buf ( R_1335a_105b5ef8 , n51068 );
buf ( R_1043d_13a1c5c8 , n51074 );
buf ( R_128cf_11cdabc8 , n51084 );
buf ( R_1219b_1207a938 , n51092 );
buf ( R_10dce_105631f8 , n51098 );
buf ( R_bbfa_10564418 , n51104 );
buf ( R_11864_12b44318 , n51110 );
buf ( R_12435_11ce4088 , n51118 );
buf ( R_a7_1265a5e8 , n51119 );
buf ( R_111f4_11cdf6c8 , n51129 );
buf ( R_135cf_1207eb78 , n51135 );
buf ( R_102ef_1153c218 , n51141 );
buf ( R_12ca0_11ce0668 , n51149 );
buf ( R_1c2_1330f228 , n51150 );
buf ( R_c6f4_12056438 , n51158 );
buf ( R_1404f_12b3e738 , n51164 );
buf ( R_ee7b_1379a628 , n51170 );
buf ( R_127e9_f8c8078 , n51176 );
buf ( R_14d_1203cbf8 , n51177 );
buf ( R_bd_1203f3f8 , n51178 );
buf ( R_48_13301848 , n51179 );
buf ( R_10afa_13a15d68 , n51185 );
buf ( R_ed66_11ce3368 , n51191 );
buf ( R_13a92_102f0bc8 , n51197 );
buf ( R_e9fb_12646268 , n51205 );
buf ( R_10d30_12084078 , n51211 );
buf ( R_149ab_1153d7f8 , n51214 );
buf ( R_88_13300d08 , n51215 );
buf ( R_6b_105aaff8 , n51216 );
buf ( R_11c31_115418f8 , n51222 );
buf ( R_13677_102f9868 , n51228 );
buf ( R_133f2_1379f088 , n51236 );
buf ( R_13edf_120837b8 , n51244 );
buf ( R_d399_137980a8 , n51252 );
buf ( R_1446e_1207d958 , n51255 );
buf ( R_1382d_1207d9f8 , n51261 );
buf ( R_cb_1331fa48 , n51262 );
buf ( R_244_1264c708 , n51263 );
buf ( R_12dc8_13a1f548 , n51269 );
buf ( R_12299_1265d1a8 , n51277 );
buf ( R_1474a_12076dd8 , n51280 );
buf ( R_13844_12663aa8 , n51290 );
buf ( R_13c11_1153d578 , n51298 );
buf ( R_14650_1056f278 , n51301 );
buf ( R_146fc_12647848 , n51304 );
buf ( R_10f84_1207bab8 , n51310 );
buf ( R_131cc_12b272f8 , n51318 );
buf ( R_1451b_10567cf8 , n51321 );
buf ( R_14390_10567c58 , n51328 );
buf ( R_13754_12082318 , n51334 );
buf ( R_1bb_12664868 , n51335 );
buf ( R_154_1204e1d8 , n51336 );
buf ( R_14831_1264f408 , n51339 );
buf ( R_7c_105b1cb8 , n51340 );
buf ( R_f1a0_12075938 , n51346 );
buf ( R_e9d0_1153f558 , n51352 );
buf ( R_f0eb_102f7568 , n51362 );
buf ( R_fb0c_1331a368 , n51368 );
buf ( R_1397b_1331b268 , n51374 );
buf ( R_e589_1379bb68 , n51380 );
buf ( R_1381a_120547b8 , n51386 );
buf ( R_1463e_105703f8 , n51389 );
buf ( R_12e76_11cd9908 , n51395 );
buf ( R_199_132fb3a8 , n51396 );
buf ( R_176_12b265d8 , n51397 );
buf ( R_125_13798008 , n51398 );
buf ( R_11ad2_102ed108 , n51406 );
buf ( R_1ea_1265a868 , n51407 );
buf ( R_10764_11cd9548 , n51415 );
buf ( R_14563_1264d6a8 , n51418 );
buf ( R_12c1a_102f0268 , n51428 );
buf ( R_146d2_1203a998 , n51431 );
buf ( R_147bd_102f9048 , n51434 );
buf ( R_fa57_1207f398 , n51440 );
buf ( R_c5a3_120849d8 , n51450 );
buf ( R_11dc9_f8c9b58 , n51458 );
buf ( R_11d95_1153f198 , n51466 );
buf ( R_1329b_11cd95e8 , n51472 );
buf ( R_14861_f8c41f8 , n51475 );
buf ( R_1064a_10561f38 , n51481 );
buf ( R_ce07_f8c8f78 , n51487 );
buf ( R_14720_11ce07a8 , n51490 );
buf ( R_13ca7_12078098 , n51496 );
buf ( R_147f5_1207a078 , n51499 );
buf ( R_142d3_12036758 , n51508 );
buf ( R_13dee_12083a38 , n51516 );
buf ( R_ec91_126490a8 , n51522 );
buf ( R_13421_11544c38 , n51528 );
buf ( R_cf92_11cdfee8 , n51534 );
buf ( R_4c49_13a1d748 , n51540 );
buf ( R_114d1_13307de8 , n51546 );
buf ( R_cff7_12076bf8 , n51552 );
buf ( R_142ff_11ce1b08 , n51559 );
buf ( R_139c0_13a1e5a8 , n51567 );
buf ( R_143cc_1056e738 , n51580 );
buf ( R_ba4e_13a1d388 , n51588 );
buf ( R_12485_105b6358 , n51596 );
buf ( R_11f0c_13a1aea8 , n51602 );
buf ( R_14867_12054b78 , n51605 );
buf ( R_137b5_10569cd8 , n51611 );
buf ( R_11d1b_12649288 , n51617 );
buf ( R_13d7b_102f56c8 , n51625 );
buf ( R_14a2c_102f12a8 , n51628 );
buf ( R_14608_13a155e8 , n51631 );
buf ( R_144c9_10571578 , n51634 );
buf ( R_fc0a_11541858 , n51642 );
buf ( R_144fa_120775f8 , n51645 );
buf ( R_129_1331c988 , n51646 );
buf ( R_13561_1330d068 , n51652 );
buf ( R_e1_12661708 , n51653 );
buf ( R_1299a_1207b158 , n51659 );
buf ( R_1489d_105686f8 , n51662 );
buf ( R_22e_132f2ac8 , n51663 );
buf ( R_6d01_102f72e8 , n51669 );
buf ( R_ffc3_12656e48 , n51675 );
buf ( R_1496f_102f9908 , n51678 );
buf ( R_1e6_13792a68 , n51679 );
buf ( R_14760_11ce3868 , n51682 );
buf ( R_d2d1_13793468 , n51692 );
buf ( R_12145_1207b978 , n51698 );
buf ( R_f5_11537038 , n51699 );
buf ( R_bb_13799cc8 , n51700 );
buf ( R_21a_1265b088 , n51701 );
buf ( R_14975_11541998 , n51704 );
buf ( R_147c0_11ce20a8 , n51707 );
buf ( R_13b7f_1153a198 , n51713 );
buf ( R_13615_12084c58 , n51719 );
buf ( R_14a29_10571438 , n51722 );
buf ( R_13526_102f49a8 , n51728 );
buf ( R_11215_12075b18 , n51734 );
buf ( R_10e4c_13a169e8 , n51740 );
buf ( R_13d97_105651d8 , n51746 );
buf ( R_1b3_1379b348 , n51747 );
buf ( R_13fab_11538758 , n51753 );
buf ( R_10ff9_105aad78 , n51759 );
buf ( R_145c0_11cd7f68 , n51762 );
buf ( R_145fc_120476f8 , n51765 );
buf ( R_15c_137992c8 , n51766 );
buf ( R_67bc_13311028 , n51772 );
buf ( R_efc2_11cdefe8 , n51778 );
buf ( R_145cc_132f8388 , n51781 );
buf ( R_ae_1379c1a8 , n51782 );
buf ( R_1263c_11cdf768 , n51788 );
buf ( R_57_126522e8 , n51789 );
buf ( R_14659_1264e1e8 , n51792 );
buf ( R_13899_133075c8 , n51800 );
buf ( R_125e5_13311348 , n51810 );
buf ( R_113fb_11ce7288 , n51818 );
buf ( R_11e0e_102f4908 , n51824 );
buf ( R_11270_12b29a58 , n51830 );
buf ( R_f61a_13305cc8 , n51836 );
buf ( R_1499f_133198c8 , n51839 );
buf ( R_121_13795808 , n51840 );
buf ( R_106_12b25a98 , n51841 );
buf ( R_1458a_102eb268 , n51844 );
buf ( R_126cf_13a19788 , n51850 );
buf ( R_209_1379cb08 , n51851 );
buf ( R_1ee_12656268 , n51852 );
buf ( R_12c5a_102ef688 , n51858 );
buf ( R_1270e_11cdb708 , n51864 );
buf ( R_e437_102f2c48 , n51870 );
buf ( R_147cf_11ce5168 , n51873 );
buf ( R_e233_1056d338 , n51879 );
buf ( R_13bbe_11ce55c8 , n51889 );
buf ( R_11e6b_1207d458 , n51895 );
buf ( R_13f0b_12b42f18 , n51901 );
buf ( R_103_12b41c58 , n51902 );
buf ( R_cd_12b39a58 , n51903 );
buf ( R_242_12654688 , n51904 );
buf ( R_20c_12b43c38 , n51905 );
buf ( R_11ce5_1379e048 , n51911 );
buf ( R_ef4_1056dc98 , n51913 );
buf ( R_11823_13a15fe8 , n51919 );
buf ( R_130b8_13a12988 , n51925 );
buf ( R_12baf_12648ba8 , n51933 );
buf ( R_119a4_102f3288 , n51939 );
buf ( R_f4e5_1264b308 , n51945 );
buf ( R_12c6f_11cdea48 , n51951 );
buf ( R_1473b_102fa308 , n51954 );
buf ( R_8b_132f8608 , n51955 );
buf ( R_11467_105659f8 , n51961 );
buf ( R_11b4a_11ce1568 , n51967 );
buf ( R_137f7_12077878 , n51975 );
buf ( R_e5b5_1153d938 , n51981 );
buf ( R_14775_13a1bda8 , n51984 );
buf ( R_14671_1264ab88 , n51987 );
buf ( R_14066_12084258 , n51989 );
buf ( R_13954_12076518 , n51995 );
buf ( R_de4d_12b26538 , n52003 );
buf ( R_149f6_11cda308 , n52006 );
buf ( R_aff6_102f4a48 , n52012 );
buf ( R_d75d_1207c0f8 , n52018 );
buf ( R_10f46_12081ff8 , n52024 );
buf ( R_c50b_11cdd3c8 , n52032 );
buf ( R_136ed_12082ef8 , n52038 );
buf ( R_101d1_1056e198 , n52046 );
buf ( R_1a9_12037658 , n52047 );
buf ( R_166_120507f8 , n52048 );
buf ( R_9b_12b3b178 , n52049 );
buf ( R_bb16_12650268 , n52057 );
buf ( R_1265a_105635b8 , n52063 );
buf ( R_b802_1265dba8 , n52069 );
buf ( R_131ea_102f4cc8 , n52077 );
buf ( R_14a0e_10570e98 , n52080 );
buf ( R_19a_12662068 , n52081 );
buf ( R_175_12b3fc78 , n52082 );
buf ( R_109_12b2c7f8 , n52083 );
buf ( R_206_105b5b38 , n52084 );
buf ( R_146b4_1153fcd8 , n52087 );
buf ( R_11e21_11cd9e08 , n52093 );
buf ( R_104ba_f8c7218 , n52101 );
buf ( R_13fbc_11541218 , n52107 );
buf ( R_144ba_102f8c88 , n52110 );
buf ( R_11622_102ed388 , n52118 );
buf ( R_13c02_12b29198 , n52124 );
buf ( R_13ba3_105626b8 , n52132 );
buf ( R_ff0f_12081918 , n52140 );
buf ( R_123d6_11541e98 , n52146 );
buf ( R_fd64_102f3328 , n52152 );
buf ( R_14486_102ef728 , n52155 );
buf ( R_13776_1379fd08 , n52161 );
buf ( R_14665_132f5ae8 , n52164 );
buf ( R_10098_13793968 , n52170 );
buf ( R_11072_13a1ed28 , n52176 );
buf ( R_14554_10565778 , n52179 );
buf ( R_137a8_1056b678 , n52191 );
buf ( R_11b55_12649a08 , n52197 );
buf ( R_14411_12663508 , n52207 );
buf ( R_84a7_12b40fd8 , n52215 );
buf ( R_133fc_1153ee78 , n52221 );
buf ( R_da_1331b088 , n52222 );
buf ( R_a0_1379b2a8 , n52223 );
buf ( R_235_1264d4c8 , n52224 );
buf ( R_1333b_11542c58 , n52232 );
buf ( R_132e7_11ce28c8 , n52238 );
buf ( R_1357d_1153feb8 , n52244 );
buf ( R_14644_1056d978 , n52247 );
buf ( R_100_1265f0e8 , n52248 );
buf ( R_79_137a1388 , n52249 );
buf ( R_e0d7_126556c8 , n52259 );
buf ( R_11b42_1264b6c8 , n52265 );
buf ( R_20f_12b28018 , n52266 );
buf ( R_f4db_1207bfb8 , n52272 );
buf ( R_1193e_13a19968 , n52278 );
buf ( R_138d5_1379b848 , n52284 );
buf ( R_13e4c_1207f118 , n52292 );
buf ( R_13a7e_102f6ac8 , n52298 );
buf ( R_12d79_102ee468 , n52304 );
buf ( R_116a8_12084398 , n52310 );
buf ( R_116_1265f868 , n52311 );
buf ( R_148a3_11cdecc8 , n52314 );
buf ( R_13273_13a1a688 , n52322 );
buf ( R_1f9_1379ddc8 , n52323 );
buf ( R_1025b_1330bee8 , n52329 );
buf ( R_122e8_12b39878 , n52335 );
buf ( R_11ba2_11544738 , n52343 );
buf ( R_12521_1056c258 , n52353 );
buf ( R_e8e6_f8cf4b8 , n52359 );
buf ( R_8cd2_1264ac28 , n52365 );
buf ( R_11a11_126477a8 , n52371 );
buf ( R_143c6_120850b8 , n52384 );
buf ( R_13e99_12039e58 , n52390 );
buf ( R_1466b_13306808 , n52393 );
buf ( R_14465_1207a758 , n52396 );
buf ( R_134b3_102f3468 , n52402 );
buf ( R_11fe7_1330c3e8 , n52408 );
buf ( R_1258d_13a14dc8 , n52416 );
buf ( R_14677_105712f8 , n52419 );
buf ( R_1367d_102eb628 , n52425 );
buf ( R_1e2_12663c88 , n52426 );
buf ( R_b9_12661848 , n52427 );
buf ( R_12d_12660268 , n52428 );
buf ( R_f47c_1153ded8 , n52436 );
buf ( R_1468c_13a1aae8 , n52439 );
buf ( R_145ba_120815f8 , n52442 );
buf ( R_14790_11cd9cc8 , n52445 );
buf ( R_14419_12048f58 , n52450 );
buf ( R_13bb3_1207b6f8 , n52456 );
buf ( R_1046b_105688d8 , n52462 );
buf ( R_1232e_13314008 , n52468 );
buf ( R_1170d_1264c528 , n52474 );
buf ( R_14a41_1056fa98 , n52477 );
buf ( R_14459_11cd92c8 , n52480 );
buf ( R_14480_11cdcf68 , n52483 );
buf ( R_13a88_11ce3f48 , n52489 );
buf ( R_c8f0_102f0d08 , n52495 );
buf ( R_134ff_1056bf38 , n52501 );
buf ( R_aac5_13a18748 , n52509 );
buf ( R_14509_13a1e148 , n52512 );
buf ( R_cebc_12039d18 , n52520 );
buf ( R_135bd_12081058 , n52526 );
buf ( R_147ba_12078ef8 , n52529 );
buf ( R_f4a6_105654f8 , n52535 );
buf ( R_1182e_13a19aa8 , n52541 );
buf ( R_142eb_11cdec28 , n52548 );
buf ( R_13bf5_10568ab8 , n52554 );
buf ( R_12093_12077058 , n52560 );
buf ( R_13dac_13a15688 , n52566 );
buf ( R_dc51_13304f08 , n52574 );
buf ( R_13e8f_1264a0e8 , n52580 );
buf ( R_13c89_12b39f58 , n52588 );
buf ( R_f0be_102f1de8 , n52594 );
buf ( R_9373_10563e78 , n52602 );
buf ( R_11a48_13a195a8 , n52608 );
buf ( R_f3f9_1153f9b8 , n52614 );
buf ( R_1d4_12b42fb8 , n52615 );
buf ( R_e3f1_12b25bd8 , n52621 );
buf ( R_13c27_13309b48 , n52627 );
buf ( R_240_105ab4f8 , n52628 );
buf ( R_cf_13311a28 , n52629 );
buf ( R_13c38_1204a3f8 , n52635 );
buf ( R_13b_13300f88 , n52636 );
buf ( R_11ef6_11cd7888 , n52642 );
buf ( R_135c9_11ce6888 , n52648 );
buf ( R_116d1_1153d898 , n52654 );
buf ( R_149d2_12080158 , n52657 );
buf ( R_ba5b_12b403f8 , n52663 );
buf ( R_ea84_1330ca28 , n52669 );
buf ( R_f59a_11ce3908 , n52675 );
buf ( R_1496c_1331e968 , n52678 );
buf ( R_12bd5_11ce3fe8 , n52684 );
buf ( R_1253e_105b6678 , n52690 );
buf ( R_14873_11cd79c8 , n52693 );
buf ( R_149a5_132ff868 , n52696 );
buf ( R_14512_11540bd8 , n52699 );
buf ( R_14756_10565318 , n52702 );
buf ( R_1c9_13313a68 , n52703 );
buf ( R_d09b_12660948 , n52709 );
buf ( R_203_12050cf8 , n52710 );
buf ( R_10c_12038058 , n52711 );
buf ( R_146_12b42298 , n52712 );
buf ( R_136c1_12b276b8 , n52718 );
buf ( R_1480a_12649e68 , n52721 );
buf ( R_1d9_1379e7c8 , n52722 );
buf ( R_13e84_1056ad18 , n52728 );
buf ( R_1021c_1056fc78 , n52734 );
buf ( R_136_132fe6e8 , n52735 );
buf ( R_145ff_102ef2c8 , n52738 );
buf ( R_19b_12b28dd8 , n52739 );
buf ( R_1031a_11540e58 , n52745 );
buf ( R_1f2_11538438 , n52746 );
buf ( R_13114_102f3648 , n52752 );
buf ( R_ec36_12042af8 , n52760 );
buf ( R_222_133189c8 , n52761 );
buf ( R_6f_12b3a458 , n52762 );
buf ( R_96_1203c838 , n52763 );
buf ( R_ed_1203deb8 , n52764 );
buf ( R_11d_1204c838 , n52765 );
buf ( R_174_13318928 , n52766 );
buf ( R_119f1_13316588 , n52774 );
buf ( R_1486a_13a1d428 , n52777 );
buf ( R_11717_1207d778 , n52783 );
buf ( R_14781_115447d8 , n52786 );
buf ( R_13995_12038738 , n52792 );
buf ( R_e4f5_12049598 , n52798 );
buf ( R_74a9_12645d68 , n52804 );
buf ( R_10208_12038558 , n52812 );
buf ( R_145ab_12b3f9f8 , n52815 );
buf ( R_227_1331e508 , n52816 );
buf ( R_e8_133028e8 , n52817 );
buf ( R_13809_1153faf8 , n52823 );
buf ( R_f732_12649008 , n52829 );
buf ( R_14524_137968e8 , n52832 );
buf ( R_146d8_11cd94a8 , n52835 );
buf ( R_14064_1264d2e8 , n52837 );
buf ( R_12dfa_11cd88c8 , n52843 );
buf ( R_135ef_102f0a88 , n52849 );
buf ( R_10ee5_12047798 , n52855 );
buf ( R_14548_120493b8 , n52858 );
buf ( R_11030_11cdbca8 , n52864 );
buf ( R_1400f_13a1a368 , n52870 );
buf ( R_f051_1264e6e8 , n52876 );
buf ( R_de7c_102eafe8 , n52884 );
buf ( R_13538_120754d8 , n52890 );
buf ( R_13e56_12b297d8 , n52898 );
buf ( R_84eb_1331c2a8 , n52904 );
buf ( R_1498a_1207e3f8 , n52907 );
buf ( R_148a6_115459f8 , n52910 );
buf ( R_212_1330bd08 , n52911 );
buf ( R_fd_13307d48 , n52912 );
buf ( R_144a5_13a1c028 , n52915 );
buf ( R_10110_120369d8 , n52921 );
buf ( R_12b5e_12651208 , n52927 );
buf ( R_149ed_13303428 , n52930 );
buf ( R_144db_12078598 , n52933 );
buf ( R_bf9f_11cd9b88 , n52941 );
buf ( R_14017_f8c20d8 , n52947 );
buf ( R_13a3d_f8ca918 , n52953 );
buf ( R_13b2d_120830d8 , n52959 );
buf ( R_8e_132f37e8 , n52960 );
buf ( R_12aeb_120810f8 , n52966 );
buf ( R_a23e_11ce5ca8 , n52972 );
buf ( R_12ce9_12081c38 , n52978 );
buf ( R_f00_1207c058 , n52980 );
buf ( R_c1fe_1264be48 , n52986 );
buf ( R_f2d2_11cdf948 , n52994 );
buf ( R_14385_12044c18 , n53007 );
buf ( R_143c0_1265fb88 , n53020 );
buf ( R_14496_13a1c668 , n53023 );
buf ( R_14738_12b28bf8 , n53026 );
buf ( R_cab9_102f99a8 , n53032 );
buf ( R_1255c_f8c61d8 , n53038 );
buf ( R_143ba_11cde868 , n53050 );
buf ( R_147c9_13a18ce8 , n53053 );
buf ( R_13311_13a198c8 , n53059 );
buf ( R_147a2_102f2ce8 , n53062 );
buf ( R_fbe0_13a1b628 , n53068 );
buf ( R_dcc6_12664ae8 , n53074 );
buf ( R_103cf_12085158 , n53080 );
buf ( R_13909_1204f5d8 , n53086 );
buf ( R_1197b_115433d8 , n53092 );
buf ( R_144e1_13a1f4a8 , n53095 );
buf ( R_145a2_11cd7ce8 , n53098 );
buf ( R_12d50_120851f8 , n53104 );
buf ( R_12380_10563338 , n53110 );
buf ( R_107a7_1379f9e8 , n53116 );
buf ( R_10e8a_102ea688 , n53122 );
buf ( R_122fb_13a17708 , n53128 );
buf ( R_12aa7_12037798 , n53134 );
buf ( R_12107_1264d428 , n53140 );
buf ( R_14533_1330c8e8 , n53143 );
buf ( R_14542_120759d8 , n53146 );
buf ( R_4276_102effe8 , n53152 );
buf ( R_1478d_115453b8 , n53155 );
buf ( R_130c1_11542258 , n53161 );
buf ( R_13ff8_102f9fe8 , n53167 );
buf ( R_1aa_13795268 , n53168 );
buf ( R_116b1_13a159a8 , n53174 );
buf ( R_1bc_126536e8 , n53175 );
buf ( R_b76e_1153c8f8 , n53181 );
buf ( R_4e_13792e28 , n53182 );
buf ( R_60_12b44bd8 , n53183 );
buf ( R_a5_13311668 , n53184 );
buf ( R_b7_1379f948 , n53185 );
buf ( R_153_13793288 , n53186 );
buf ( R_165_13306948 , n53187 );
buf ( R_f9fe_102f9408 , n53193 );
buf ( R_14431_12080478 , n53197 );
buf ( R_1c3_12047158 , n53198 );
buf ( R_64_f8c1bd8 , n53199 );
buf ( R_14c_120387d8 , n53200 );
buf ( R_12471_102f7068 , n53206 );
buf ( R_148c1_13316f88 , n53209 );
buf ( R_11433_1265f048 , n53221 );
buf ( R_13ce2_1264aa48 , n53227 );
buf ( R_121bd_115449b8 , n53233 );
buf ( R_14813_10566d58 , n53236 );
buf ( R_147fb_102f83c8 , n53239 );
buf ( R_146ab_12051658 , n53242 );
buf ( R_12c65_1264cb68 , n53248 );
buf ( R_e2b4_f8c0f58 , n53254 );
buf ( R_10c61_120805b8 , n53260 );
buf ( R_10f1d_10566df8 , n53266 );
buf ( R_10de4_1379b5c8 , n53272 );
buf ( R_ae51_105ab098 , n53278 );
buf ( R_146f3_12659d28 , n53281 );
buf ( R_d03f_126484c8 , n53287 );
buf ( R_9fe2_11543fb8 , n53293 );
buf ( R_10b79_12657028 , n53301 );
buf ( R_64c2_12662748 , n53307 );
buf ( R_139d0_102f1fc8 , n53313 );
buf ( R_13639_1207f578 , n53319 );
buf ( R_1b4_12654728 , n53320 );
buf ( R_1cf_133184c8 , n53321 );
buf ( R_e214_1207ae38 , n53327 );
buf ( R_140_12665448 , n53328 );
buf ( R_15b_f8c0378 , n53329 );
buf ( R_1435c_13304d28 , n53337 );
buf ( R_10745_12056898 , n53343 );
buf ( R_1044f_120557f8 , n53349 );
buf ( R_10824_11ce3188 , n53355 );
buf ( R_13820_12b41438 , n53361 );
buf ( R_69b8_11cdc888 , n53367 );
buf ( R_124b9_1056d658 , n53373 );
buf ( R_143f4_102edd88 , n53378 );
buf ( R_142f5_1264a908 , n53385 );
buf ( R_76_f8ca198 , n53386 );
buf ( R_ac_12660a88 , n53387 );
buf ( R_1269b_11cd9368 , n53393 );
buf ( R_147b4_120766f8 , n53396 );
buf ( R_14834_13a16a88 , n53399 );
buf ( R_12e88_102f8a08 , n53405 );
buf ( R_f021_102ec168 , n53411 );
buf ( R_f6dd_13a163a8 , n53417 );
buf ( R_145e4_126463a8 , n53420 );
buf ( R_14723_1264db08 , n53423 );
buf ( R_173_f8c3438 , n53424 );
buf ( R_19c_12b40218 , n53425 );
buf ( R_11142_10562f78 , n53431 );
buf ( R_23e_1265bc68 , n53432 );
buf ( R_d1_13311f28 , n53433 );
buf ( R_13512_12080dd8 , n53439 );
buf ( R_7859_11cdaee8 , n53445 );
buf ( R_14593_115458b8 , n53448 );
buf ( R_148a9_12647ac8 , n53451 );
buf ( R_10577_11545318 , n53457 );
buf ( R_133ca_1203e098 , n53463 );
buf ( R_13b92_13a14be8 , n53471 );
buf ( R_10efd_102ec3e8 , n53477 );
buf ( R_f0b_1153f4b8 , n53479 );
buf ( R_12e15_10568018 , n53485 );
buf ( R_200_12b29eb8 , n53486 );
buf ( R_21d_137a03e8 , n53487 );
buf ( R_f2_12652ec8 , n53488 );
buf ( R_10f_12b3e5f8 , n53489 );
buf ( R_ca13_11ce4628 , n53495 );
buf ( R_14966_11546218 , n53498 );
buf ( R_13ad8_1203a358 , n53504 );
buf ( R_12d8d_105b5db8 , n53510 );
buf ( R_10165_1264cac8 , n53516 );
buf ( R_1337f_13a12c08 , n53522 );
buf ( R_53_f8c2a38 , n53523 );
buf ( R_149c9_132f4fa8 , n53526 );
buf ( R_10aae_1207c558 , n53532 );
buf ( R_13aad_11541a38 , n53538 );
buf ( R_12362_10563dd8 , n53544 );
buf ( R_5c4e_1056ced8 , n53550 );
buf ( R_130f5_1056a098 , n53556 );
buf ( R_12a7c_11cdde68 , n53562 );
buf ( R_14415_12b2a318 , n53567 );
buf ( R_1488b_13a189c8 , n53570 );
buf ( R_14062_1204cf18 , n53572 );
buf ( R_14784_11cd8508 , n53575 );
buf ( R_1032f_10570f38 , n53581 );
buf ( R_9bdf_102ee5a8 , n53587 );
buf ( R_13bf0_1331c528 , n53593 );
buf ( R_11b90_11ce0208 , n53599 );
buf ( R_149cf_13a17b68 , n53602 );
buf ( R_12021_11ce25a8 , n53608 );
buf ( R_1de_12056d98 , n53609 );
buf ( R_49_1331f4a8 , n53610 );
buf ( R_131_105ab3b8 , n53611 );
buf ( R_1462f_13794688 , n53614 );
buf ( R_10628_1203d2d8 , n53620 );
buf ( R_122bf_10570038 , n53626 );
buf ( R_11387_11540d18 , n53632 );
buf ( R_11fa6_13306308 , n53638 );
buf ( R_85b5_120819b8 , n53644 );
buf ( R_142ef_102eec88 , n53653 );
buf ( R_1434c_102f13e8 , n53664 );
buf ( R_22c_1379b708 , n53665 );
buf ( R_5c_137944a8 , n53666 );
buf ( R_e3_1203e778 , n53667 );
buf ( R_b948_1153a5f8 , n53673 );
buf ( R_e169_11cd7a68 , n53679 );
buf ( R_d051_11536ef8 , n53685 );
buf ( R_10e01_120551b8 , n53691 );
buf ( R_233_12b392d8 , n53692 );
buf ( R_68_12b283d8 , n53693 );
buf ( R_dc_13300768 , n53694 );
buf ( R_13bfb_13316a88 , n53700 );
buf ( R_10ad6_10565598 , n53706 );
buf ( R_14870_10570538 , n53709 );
buf ( R_12260_13a1b268 , n53715 );
buf ( R_d661_1265cfc8 , n53721 );
buf ( R_14572_11cd9d68 , n53724 );
buf ( R_130ff_12078318 , n53730 );
buf ( R_a98a_11cdaf88 , n53740 );
buf ( R_14978_12b321f8 , n53743 );
buf ( R_14a1a_115445f8 , n53746 );
buf ( R_14a26_13792568 , n53749 );
buf ( R_b327_12648568 , n53755 );
buf ( R_108fb_105b5e58 , n53761 );
buf ( R_1440d_11544238 , n53771 );
buf ( R_10cff_13a1dc48 , n53777 );
buf ( R_139ae_11cd8b48 , n53783 );
buf ( R_14338_11cda808 , n53794 );
buf ( R_106b3_13a16088 , n53800 );
buf ( R_c4f8_11ce12e8 , n53806 );
buf ( R_215_1265b948 , n53807 );
buf ( R_fa_133070c8 , n53808 );
buf ( R_11b68_1264ec88 , n53814 );
buf ( R_129b1_1056f098 , n53820 );
buf ( R_13670_10564558 , n53826 );
buf ( R_1439c_11cdd148 , n53832 );
buf ( R_107e6_11cdbc08 , n53838 );
buf ( R_f279_13a1acc8 , n53844 );
buf ( R_12ed9_102edf68 , n53850 );
buf ( R_12bc1_13a1f048 , n53856 );
buf ( R_13b19_12b2ba38 , n53862 );
buf ( R_e361_120812d8 , n53868 );
buf ( R_bef9_11ce0528 , n53874 );
buf ( R_13ce8_120793f8 , n53880 );
buf ( R_a235_12084a78 , n53886 );
buf ( R_14521_1264f228 , n53889 );
buf ( R_13cad_13a1edc8 , n53895 );
buf ( R_148af_11540098 , n53898 );
buf ( R_10968_13304968 , n53904 );
buf ( R_13fcb_102f0c68 , n53910 );
buf ( R_11645_13304e68 , n53916 );
buf ( R_bf09_1056b498 , n53922 );
buf ( R_12553_13310308 , n53928 );
buf ( R_145d5_132fa228 , n53931 );
buf ( R_146a2_1207bf18 , n53934 );
buf ( R_136fc_12076018 , n53940 );
buf ( R_149a2_1264d1a8 , n53943 );
buf ( R_12b9a_13a14968 , n53949 );
buf ( R_137cc_10569af8 , n53955 );
buf ( R_c5ef_12081238 , n53963 );
buf ( R_1184d_11cd9188 , n53969 );
buf ( R_13c8f_102ed568 , n53975 );
buf ( R_109bf_1379c248 , n53981 );
buf ( R_14326_13301528 , n53989 );
buf ( R_11123_12045258 , n53995 );
buf ( R_e197_11ce3228 , n54001 );
buf ( R_172_126656c8 , n54002 );
buf ( R_19d_132ffb88 , n54003 );
buf ( R_c306_f8c5418 , n54009 );
buf ( R_b5_133157c8 , n54010 );
buf ( R_13902_13799ae8 , n54016 );
buf ( R_14348_1056c398 , n54024 );
buf ( R_1457b_102f5628 , n54027 );
buf ( R_14766_105674d8 , n54030 );
buf ( R_d2c1_12036e38 , n54036 );
buf ( R_1f6_1330dce8 , n54037 );
buf ( R_10c28_12080e78 , n54043 );
buf ( R_119_133166c8 , n54044 );
buf ( R_1300e_12646bc8 , n54050 );
buf ( R_13129_10567b18 , n54056 );
buf ( R_1394d_1056f318 , n54062 );
buf ( R_14846_13798b48 , n54065 );
buf ( R_146cf_1379e868 , n54068 );
buf ( R_10019_11542118 , n54074 );
buf ( R_fb35_132fb4e8 , n54080 );
buf ( R_11a23_126506c8 , n54086 );
buf ( R_9aae_1056dbf8 , n54092 );
buf ( R_14468_1264aea8 , n54095 );
buf ( R_7aaf_f8c22b8 , n54101 );
buf ( R_b5af_1264e508 , n54109 );
buf ( R_13f11_11cd7b08 , n54115 );
buf ( R_e6c6_12075cf8 , n54121 );
buf ( R_14374_102f0768 , n54134 );
buf ( R_14605_13a182e8 , n54137 );
buf ( R_13de4_102f94a8 , n54143 );
buf ( R_102c2_1264ed28 , n54151 );
buf ( R_91_13799548 , n54152 );
buf ( R_135f5_11cda4e8 , n54158 );
buf ( R_14807_1331e288 , n54161 );
buf ( R_14a08_11cdc388 , n54164 );
buf ( R_cb44_12b3ee18 , n54170 );
buf ( R_13a63_11544198 , n54180 );
buf ( R_109ca_1264cd48 , n54186 );
buf ( R_12e41_10569198 , n54192 );
buf ( R_e46a_13a181a8 , n54198 );
buf ( R_12963_13a1afe8 , n54204 );
buf ( R_14a5a_12b42158 , n54208 );
buf ( R_13e38_1207efd8 , n54214 );
buf ( R_144ea_1264f5e8 , n54217 );
buf ( R_11668_137a1d88 , n54225 );
buf ( R_13ec7_11540318 , n54231 );
buf ( R_ff67_13799688 , n54237 );
buf ( R_13b27_102eb588 , n54243 );
buf ( R_fa2a_1056e0f8 , n54249 );
buf ( R_145a5_132f4dc8 , n54252 );
buf ( R_14060_13a15ae8 , n54254 );
buf ( R_164_12b27118 , n54255 );
buf ( R_104d9_120779b8 , n54261 );
buf ( R_1ab_f8c2998 , n54262 );
buf ( R_23c_13319328 , n54263 );
buf ( R_bbdf_133063a8 , n54269 );
buf ( R_d3_12659968 , n54270 );
buf ( R_cc7b_13a1b128 , n54276 );
buf ( R_12ffe_1331cd48 , n54282 );
buf ( R_1323e_126561c8 , n54288 );
buf ( R_1207f_133190a8 , n54294 );
buf ( R_10f99_126549a8 , n54300 );
buf ( R_913d_12646b28 , n54306 );
buf ( R_c3ee_102f6848 , n54312 );
buf ( R_13b12_13a1a728 , n54318 );
buf ( R_10a0c_11cdf1c8 , n54324 );
buf ( R_13974_13a19008 , n54330 );
buf ( R_13602_126635a8 , n54336 );
buf ( R_124e1_11cdb668 , n54342 );
buf ( R_142d7_12b30d58 , n54351 );
buf ( R_14960_105b5598 , n54354 );
buf ( R_f86d_120385f8 , n54360 );
buf ( R_148a0_12b38ab8 , n54363 );
buf ( R_e63f_f8cb9f8 , n54369 );
buf ( R_12741_105642d8 , n54375 );
buf ( R_684e_1056aa98 , n54381 );
buf ( R_13b04_12081558 , n54387 );
buf ( R_1453f_11ce2328 , n54390 );
buf ( R_148b5_1207f898 , n54393 );
buf ( R_1499c_12080658 , n54396 );
buf ( R_128e2_12647668 , n54402 );
buf ( R_13345_11ce0988 , n54408 );
buf ( R_cd4f_102f2f68 , n54414 );
buf ( R_13dd3_1204cd38 , n54420 );
buf ( R_13ea4_11ce0708 , n54426 );
buf ( R_f16b_11cda448 , n54432 );
buf ( R_139fe_1153e5b8 , n54438 );
buf ( R_12eed_102ee1e8 , n54444 );
buf ( R_13479_13306b28 , n54450 );
buf ( R_1135b_1056d158 , n54456 );
buf ( R_131a5_1153dc58 , n54462 );
buf ( R_14744_1264b3a8 , n54465 );
buf ( R_144c6_1056d5b8 , n54468 );
buf ( R_13109_f8c4798 , n54474 );
buf ( R_137bb_10564058 , n54480 );
buf ( R_146db_1056a818 , n54483 );
buf ( R_119c2_13a1a548 , n54489 );
buf ( R_eb5e_1056d018 , n54495 );
buf ( R_b0d7_1153e3d8 , n54501 );
buf ( R_13b9e_12083038 , n54507 );
buf ( R_1116a_13a15868 , n54513 );
buf ( R_12a65_10564c38 , n54519 );
buf ( R_14969_11cdb2a8 , n54522 );
buf ( R_1464d_12075618 , n54525 );
buf ( R_e3c5_12080a18 , n54531 );
buf ( R_1469c_120511f8 , n54534 );
buf ( R_d50f_12663828 , n54540 );
buf ( R_137f0_12079358 , n54546 );
buf ( R_11593_1207a258 , n54552 );
buf ( R_14350_1207d8b8 , n54560 );
buf ( R_cbe2_11536a98 , n54566 );
buf ( R_110ed_10563d38 , n54572 );
buf ( R_1125d_102f86e8 , n54578 );
buf ( R_13c09_11ce4268 , n54584 );
buf ( R_135fc_13795948 , n54590 );
buf ( R_14557_11cdcec8 , n54593 );
buf ( R_112_13312248 , n54594 );
buf ( R_1fd_133221a8 , n54595 );
buf ( R_9e_11539838 , n54596 );
buf ( R_143b2_11cddd28 , n54608 );
buf ( R_12fec_102efea8 , n54614 );
buf ( R_c4d7_13a1f408 , n54620 );
buf ( R_1398e_13320bc8 , n54626 );
buf ( R_12894_11ce1428 , n54632 );
buf ( R_b6f4_102f9ea8 , n54638 );
buf ( R_fcb3_12649be8 , n54644 );
buf ( R_12375_1207edf8 , n54650 );
buf ( R_146b1_102ed248 , n54653 );
buf ( R_11b11_11545818 , n54659 );
buf ( R_58_13317a28 , n54660 );
buf ( R_73_12b3e0f8 , n54661 );
buf ( R_bd7c_11ce2be8 , n54667 );
buf ( R_12fd8_10565278 , n54673 );
buf ( R_14876_12054678 , n54676 );
buf ( R_138da_1153dbb8 , n54682 );
buf ( R_14825_12647168 , n54685 );
buf ( R_14a4d_12646ee8 , n54688 );
buf ( R_124_1203edb8 , n54689 );
buf ( R_15a_f8c6958 , n54690 );
buf ( R_1b5_1331afe8 , n54691 );
buf ( R_1eb_12038d78 , n54692 );
buf ( R_1475d_11546038 , n54695 );
buf ( R_171_105aa5f8 , n54696 );
buf ( R_106ea_102f6528 , n54702 );
buf ( R_19e_1331e788 , n54703 );
buf ( R_11a86_1204ffd8 , n54711 );
buf ( R_fad7_102f5ee8 , n54717 );
buf ( R_e21e_1056b7b8 , n54723 );
buf ( R_12933_11cd7c48 , n54729 );
buf ( R_6c_12040938 , n54730 );
buf ( R_99_12b27618 , n54731 );
buf ( R_1353d_1153d9d8 , n54737 );
buf ( R_b283_1330acc8 , n54743 );
buf ( R_143ae_13a1cca8 , n54755 );
buf ( R_14801_11540c78 , n54758 );
buf ( R_149e7_10568298 , n54761 );
buf ( R_14708_1203c018 , n54764 );
buf ( R_14450_13a17028 , n54768 );
buf ( R_128_12b43b98 , n54769 );
buf ( R_145_1265aa48 , n54770 );
buf ( R_1ca_1265ff48 , n54771 );
buf ( R_1e7_12b3d798 , n54772 );
buf ( R_7741_13a16128 , n54778 );
buf ( R_da39_12b40718 , n54784 );
buf ( R_e38d_12651168 , n54790 );
buf ( R_12fc4_11544878 , n54796 );
buf ( R_145e7_11544058 , n54799 );
buf ( R_1465f_105676b8 , n54802 );
buf ( R_10fc1_12078638 , n54808 );
buf ( R_704f_11ce4da8 , n54814 );
buf ( R_13a8d_13318108 , n54820 );
buf ( R_145c3_1264da68 , n54823 );
buf ( R_faad_13a1fd68 , n54829 );
buf ( R_12738_10570678 , n54835 );
buf ( R_11935_13a1ff48 , n54841 );
buf ( R_11720_1330eaa8 , n54847 );
buf ( R_d16a_11ce5de8 , n54858 );
buf ( R_13e0d_13a1b4e8 , n54864 );
buf ( R_1447d_11ce3a48 , n54867 );
buf ( R_152_12b3c4d8 , n54868 );
buf ( R_105ba_13306bc8 , n54874 );
buf ( R_b1aa_12649468 , n54880 );
buf ( R_1bd_12653be8 , n54881 );
buf ( R_14a50_13a161c8 , n54884 );
buf ( R_13a83_10567a78 , n54890 );
buf ( R_123c2_13797108 , n54896 );
buf ( R_144b7_13305d68 , n54899 );
buf ( R_13814_137926a8 , n54905 );
buf ( R_12cbd_13a14328 , n54911 );
buf ( R_11bab_120768d8 , n54917 );
buf ( R_c07e_13a18b08 , n54923 );
buf ( R_142f9_11545e58 , n54932 );
buf ( R_1478a_12652928 , n54935 );
buf ( R_14a3b_11ce2d28 , n54938 );
buf ( R_c3a2_13a19508 , n54944 );
buf ( R_aa_126535a8 , n54945 );
buf ( R_146e7_10566538 , n54948 );
buf ( R_138fb_12082778 , n54954 );
buf ( R_13988_133186a8 , n54960 );
buf ( R_13c43_1264cca8 , n54966 );
buf ( R_14590_132f3b08 , n54969 );
buf ( R_110cf_137940e8 , n54975 );
buf ( R_13326_12648d88 , n54981 );
buf ( R_13153_10567118 , n54987 );
buf ( R_1405e_f8c95b8 , n54989 );
buf ( R_1051f_13793b48 , n54997 );
buf ( R_f518_12075bb8 , n55003 );
buf ( R_143a2_12079038 , n55016 );
buf ( R_147a8_12657de8 , n55019 );
buf ( R_13cb3_102f6fc8 , n55025 );
buf ( R_10c3d_f8c5b98 , n55031 );
buf ( R_e7ab_1264f7c8 , n55037 );
buf ( R_13449_12077378 , n55043 );
buf ( R_14403_12b29418 , n55053 );
buf ( R_148b2_132fc708 , n55056 );
buf ( R_1468f_10562cf8 , n55059 );
buf ( R_f7_13309828 , n55060 );
buf ( R_13f54_102f4e08 , n55066 );
buf ( R_218_12050258 , n55067 );
buf ( R_83_1379cd88 , n55068 );
buf ( R_12f16_137a0b68 , n55074 );
buf ( R_10598_102ead68 , n55080 );
buf ( R_10365_12051478 , n55086 );
buf ( R_13ab4_13a12ca8 , n55092 );
buf ( R_13393_10568a18 , n55098 );
buf ( R_13683_1207cf58 , n55104 );
buf ( R_13a_105ac2b8 , n55105 );
buf ( R_127d5_11cdf268 , n55111 );
buf ( R_11917_11ce1248 , n55117 );
buf ( R_1d5_1265e468 , n55118 );
buf ( R_12e98_1204e778 , n55124 );
buf ( R_b3_12655ea8 , n55125 );
buf ( R_149cc_10564cd8 , n55128 );
buf ( R_134d9_10565f98 , n55134 );
buf ( R_fd0b_102ec488 , n55140 );
buf ( R_af25_133136a8 , n55146 );
buf ( R_11948_12b288d8 , n55152 );
buf ( R_149c6_1207b018 , n55155 );
buf ( R_14b_12b28a18 , n55156 );
buf ( R_1c4_12652e28 , n55157 );
buf ( R_10199_13a1f368 , n55163 );
buf ( R_80_12055438 , n55164 );
buf ( R_10b70_f8cd438 , n55170 );
buf ( R_10cdf_115401d8 , n55176 );
buf ( R_11a66_1207dc78 , n55182 );
buf ( R_132fc_13307708 , n55188 );
buf ( R_8c7b_12076b58 , n55194 );
buf ( R_1495a_1207a2f8 , n55197 );
buf ( R_1201a_10570218 , n55203 );
buf ( R_132d6_11ce0348 , n55209 );
buf ( R_14963_13304be8 , n55212 );
buf ( R_1285e_11545c78 , n55218 );
buf ( R_130de_102f58a8 , n55224 );
buf ( R_fb5f_13a1e288 , n55230 );
buf ( R_13ecf_1207c5f8 , n55236 );
buf ( R_1456f_13a1f5e8 , n55239 );
buf ( R_ea_1331a9a8 , n55240 );
buf ( R_120_12b400d8 , n55241 );
buf ( R_13eac_11ce2a08 , n55249 );
buf ( R_12568_1056b0d8 , n55255 );
buf ( R_e3ba_1207df98 , n55261 );
buf ( R_dcf2_12085298 , n55267 );
buf ( R_1ef_f8c2cb8 , n55268 );
buf ( R_225_12b3a318 , n55269 );
buf ( R_f7da_1204e9f8 , n55275 );
buf ( R_f857_13a13748 , n55281 );
buf ( R_1461a_13301988 , n55284 );
buf ( R_146b7_13a15228 , n55287 );
buf ( R_1384a_126503a8 , n55293 );
buf ( R_c8e7_105b6498 , n55299 );
buf ( R_86_137a1a68 , n55300 );
buf ( R_a3_126621a8 , n55301 );
buf ( R_f862_13a1a908 , n55307 );
buf ( R_10ab7_102f7b08 , n55313 );
buf ( R_11890_102eb308 , n55319 );
buf ( R_df3c_120774b8 , n55325 );
buf ( R_1369b_1330c2a8 , n55331 );
buf ( R_12e03_132ff368 , n55337 );
buf ( R_1356b_102f5da8 , n55343 );
buf ( R_10e42_1207e718 , n55349 );
buf ( R_10f59_f8c2c18 , n55355 );
buf ( R_127b6_12b412f8 , n55361 );
buf ( R_120e7_12b44818 , n55367 );
buf ( R_12492_1265b9e8 , n55373 );
buf ( R_10d12_13792b08 , n55379 );
buf ( R_130ae_12044b78 , n55385 );
buf ( R_13652_11ce1ce8 , n55391 );
buf ( R_117a7_12080fb8 , n55397 );
buf ( R_14674_13a13ba8 , n55400 );
buf ( R_11306_11540638 , n55406 );
buf ( R_d5_126617a8 , n55407 );
buf ( R_de_1265ce88 , n55408 );
buf ( R_12c_1379b488 , n55409 );
buf ( R_135_f8c6f98 , n55410 );
buf ( R_1da_12664b88 , n55411 );
buf ( R_1e3_1153c498 , n55412 );
buf ( R_122dd_13a1b6c8 , n55418 );
buf ( R_231_1379a6c8 , n55419 );
buf ( R_23a_12660b28 , n55420 );
buf ( R_1240e_13a150e8 , n55426 );
buf ( R_14686_13a137e8 , n55429 );
buf ( R_146c6_f8cf918 , n55432 );
buf ( R_13f5b_1207c738 , n55438 );
buf ( R_ebb7_102efd68 , n55444 );
buf ( R_1447a_105697d8 , n55447 );
buf ( R_13c95_12650ee8 , n55453 );
buf ( R_11de0_12083cb8 , n55459 );
buf ( R_11552_12648c48 , n55465 );
buf ( R_11cb2_1207ab18 , n55471 );
buf ( R_14849_11ce0028 , n55474 );
buf ( R_13f45_13a134c8 , n55480 );
buf ( R_13726_12084f78 , n55486 );
buf ( R_121f2_102f30a8 , n55492 );
buf ( R_ef_1379b0c8 , n55493 );
buf ( R_163_12b38a18 , n55494 );
buf ( R_1ac_12b29558 , n55495 );
buf ( R_220_12b25638 , n55496 );
buf ( R_14623_13a12a28 , n55499 );
buf ( R_1393a_11ce3408 , n55505 );
buf ( R_139ea_11cd8828 , n55511 );
buf ( R_cf49_11541718 , n55517 );
buf ( R_b889_1056a458 , n55523 );
buf ( R_1349f_1204fdf8 , n55529 );
buf ( R_170_120440d8 , n55530 );
buf ( R_19f_133087e8 , n55531 );
buf ( R_a9d8_102f22e8 , n55537 );
buf ( R_7d_12660308 , n55538 );
buf ( R_1460b_10569a58 , n55541 );
buf ( R_11983_13318568 , n55547 );
buf ( R_a6e4_13314648 , n55553 );
buf ( R_144b1_1207b478 , n55556 );
buf ( R_14614_12664f48 , n55559 );
buf ( R_139d7_132fda68 , n55565 );
buf ( R_ec64_11ce6248 , n55571 );
buf ( R_12d32_115454f8 , n55577 );
buf ( R_82bb_1204a678 , n55583 );
buf ( R_1472c_13a139c8 , n55586 );
buf ( R_144f7_10565e58 , n55589 );
buf ( R_10dad_12082f98 , n55595 );
buf ( R_b05c_1330b4e8 , n55601 );
buf ( R_13ef1_105714d8 , n55607 );
buf ( R_14635_12b3b038 , n55610 );
buf ( R_117b5_1056fdb8 , n55616 );
buf ( R_14692_11cdf128 , n55619 );
buf ( R_13f_1203dd78 , n55620 );
buf ( R_1055c_105672f8 , n55626 );
buf ( R_1d0_12040258 , n55627 );
buf ( R_13aba_1265cde8 , n55633 );
buf ( R_131e1_102f2ec8 , n55639 );
buf ( R_eb07_1153ef18 , n55645 );
buf ( R_9c9a_1056c578 , n55651 );
buf ( R_10605_11545d18 , n55657 );
buf ( R_13a97_12079218 , n55663 );
buf ( R_1331b_102efc28 , n55669 );
buf ( R_14879_11ce58e8 , n55672 );
buf ( R_14996_102eb3a8 , n55675 );
buf ( R_1405c_11ce34a8 , n55677 );
buf ( R_14945_1056e238 , n55680 );
buf ( R_b65f_11cdba28 , n55686 );
buf ( R_13f3e_13a1e508 , n55692 );
buf ( R_dbc0_132fb9e8 , n55698 );
buf ( R_1351c_13797068 , n55704 );
buf ( R_14804_120788b8 , n55707 );
buf ( R_14a0b_133206c8 , n55710 );
buf ( R_89_126595a8 , n55711 );
buf ( R_13c33_11ce3688 , n55717 );
buf ( R_4f_12b44d18 , n55718 );
buf ( R_cb5a_12b256d8 , n55724 );
buf ( R_13b85_10571258 , n55730 );
buf ( R_138f4_1330a9a8 , n55736 );
buf ( R_ee1a_1264fae8 , n55742 );
buf ( R_10411_102f8828 , n55748 );
buf ( R_14331_1056be98 , n55756 );
buf ( R_14717_1153a378 , n55759 );
buf ( R_94_1330ee68 , n55760 );
buf ( R_e5_1153cfd8 , n55761 );
buf ( R_22a_12b43698 , n55762 );
buf ( R_cba1_13a16e48 , n55773 );
buf ( R_129d1_12047978 , n55779 );
buf ( R_143d8_11cdc2e8 , n55792 );
buf ( R_13070_1264b268 , n55798 );
buf ( R_12915_1056d518 , n55804 );
buf ( R_12942_11cdd0a8 , n55810 );
buf ( R_145a8_12662608 , n55813 );
buf ( R_fda2_1264e328 , n55819 );
buf ( R_ee25_13a16588 , n55825 );
buf ( R_13a1f_11cde2c8 , n55831 );
buf ( R_1432d_11cdddc8 , n55842 );
buf ( R_13be3_12036bb8 , n55848 );
buf ( R_fe10_13a14468 , n55854 );
buf ( R_12610_1204bcf8 , n55860 );
buf ( R_13701_11cdc608 , n55866 );
buf ( R_12597_105711b8 , n55872 );
buf ( R_1441d_12035d58 , n55877 );
buf ( R_1443c_137979c8 , n55881 );
buf ( R_139a7_11ce70a8 , n55887 );
buf ( R_13ad3_1056bdf8 , n55893 );
buf ( R_143e0_102efcc8 , n55903 );
buf ( R_147cc_13315ae8 , n55906 );
buf ( R_1444b_11cdad08 , n55909 );
buf ( R_12631_12036c58 , n55915 );
buf ( R_13dda_102f4fe8 , n55921 );
buf ( R_efd_13a14fa8 , n55923 );
buf ( R_14954_12054358 , n55926 );
buf ( R_1287f_115422f8 , n55932 );
buf ( R_1169f_102f8968 , n55938 );
buf ( R_13a2b_1264b628 , n55944 );
buf ( R_11285_102f9e08 , n55950 );
buf ( R_12548_1056ce38 , n55956 );
buf ( R_1173e_12649fa8 , n55962 );
buf ( R_10b51_13a18a68 , n55968 );
buf ( R_148ca_13a18c48 , n55971 );
buf ( R_12c82_102f0448 , n55977 );
buf ( R_13b79_11543d38 , n55983 );
buf ( R_14057_f8cd618 , n55985 );
buf ( R_a2e4_1056c618 , n55991 );
buf ( R_101e6_1330c7a8 , n55997 );
buf ( R_13a56_f8c0a58 , n56003 );
buf ( R_d6bc_13a1ca28 , n56009 );
buf ( R_4a_1265e648 , n56010 );
buf ( R_115_13316c68 , n56011 );
buf ( R_1224c_12b3d478 , n56017 );
buf ( R_1fa_1265d388 , n56018 );
buf ( R_eeda_11cd81e8 , n56024 );
buf ( R_1455d_11cd9fe8 , n56027 );
buf ( R_1402e_1264dc48 , n56033 );
buf ( R_c753_12039098 , n56039 );
buf ( R_1283c_13a1da68 , n56045 );
buf ( R_aeda_13a1d6a8 , n56051 );
buf ( R_14939_1379f448 , n56054 );
buf ( R_14a20_13a13e28 , n56057 );
buf ( R_13a9d_12081698 , n56063 );
buf ( R_117c0_11ce3e08 , n56069 );
buf ( R_114e1_132f28e8 , n56075 );
buf ( R_1476f_132fb768 , n56078 );
not ( n27676 , RI19a22f70_2797);
and ( n27677 , n27676 , RI1754a798_67);
not ( n27678 , RI19a23e70_2789);
and ( n27679 , n27677 , n27678 );
and ( n27680 , RI19a22f70_2797 , n27678 );
or ( n27681 , n27679 , n27680 );
not ( n27682 , RI19ad04a8_2209);
and ( n27683 , n27681 , n27682 );
not ( n10016 , n27683 );
and ( n10017 , n10016 , RI19a859b8_2755);
and ( n10018 , RI19a23510_2794 , n27683 );
or ( n27684 , n10017 , n10018 );
not ( n10019 , RI1754c610_2);
and ( n10020 , n10019 , n27684 );
and ( n10021 , C0 , RI1754c610_2);
or ( n27685 , n10020 , n10021 );
buf ( n27686 , n27685 );
xor ( n27687 , RI19a8fd50_2684 , RI17465568_1242);
not ( n27688 , RI1753aa78_586);
and ( n27689 , RI19a23e70_2789 , n27688 );
not ( n10022 , n27689 );
and ( n10023 , n10022 , RI17465568_1242);
and ( n10024 , n27687 , n27689 );
or ( n27690 , n10023 , n10024 );
xor ( n27691 , RI19ab7530_2399 , RI1749f948_958);
not ( n10025 , n27689 );
and ( n10026 , n10025 , RI1749f948_958);
and ( n10027 , n27691 , n27689 );
or ( n27692 , n10026 , n10027 );
buf ( n27693 , RI17534808_603);
xor ( n27694 , n27692 , n27693 );
buf ( n27695 , RI173ba970_1846);
xor ( n27696 , n27694 , n27695 );
buf ( n27697 , RI17403660_1491);
xor ( n27698 , n27696 , n27697 );
buf ( n27699 , RI173efea8_1586);
xor ( n27700 , n27698 , n27699 );
xor ( n27701 , n27690 , n27700 );
xor ( n27702 , RI19a9a160_2611 , RI174741a8_1170);
not ( n10028 , n27689 );
and ( n10029 , n10028 , RI174741a8_1170);
and ( n10030 , n27702 , n27689 );
or ( n27703 , n10029 , n10030 );
xor ( n27704 , RI19ac9938_2258 , RI174bfb80_814);
not ( n10031 , n27689 );
and ( n10032 , n10031 , RI174bfb80_814);
and ( n10033 , n27704 , n27689 );
or ( n27705 , n10032 , n10033 );
xor ( n27706 , n27703 , n27705 );
buf ( n27707 , RI1738f1d0_2058);
xor ( n27708 , n27706 , n27707 );
buf ( n27709 , RI173d7ec0_1703);
xor ( n27710 , n27708 , n27709 );
buf ( n27711 , RI1744f998_1348);
xor ( n27712 , n27710 , n27711 );
xor ( n27713 , n27701 , n27712 );
xor ( n27714 , RI19ac4460_2297 , RI174cedd8_767);
not ( n10034 , n27689 );
and ( n10035 , n10034 , RI174cedd8_767);
and ( n10036 , n27714 , n27689 );
or ( n27715 , n10035 , n10036 );
xor ( n27716 , RI19a8a2d8_2723 , RI1746f630_1193);
not ( n10037 , n27689 );
and ( n10038 , n10037 , RI1746f630_1193);
and ( n10039 , n27716 , n27689 );
or ( n27717 , n10038 , n10039 );
xor ( n27718 , RI19abbe50_2368 , RI174b8308_838);
not ( n10040 , n27689 );
and ( n10041 , n10040 , RI174b8308_838);
and ( n10042 , n27718 , n27689 );
or ( n27719 , n10041 , n10042 );
xor ( n27720 , n27717 , n27719 );
buf ( n27721 , RI1738a658_2081);
xor ( n27722 , n27720 , n27721 );
buf ( n27723 , RI173d3348_1726);
xor ( n27724 , n27722 , n27723 );
buf ( n27725 , RI1744ae20_1371);
xor ( n27726 , n27724 , n27725 );
xor ( n27727 , n27715 , n27726 );
xor ( n27728 , RI19aa5560_2527 , RI1747e270_1121);
not ( n10043 , n27689 );
and ( n10044 , n10043 , RI1747e270_1121);
and ( n10045 , n27728 , n27689 );
or ( n27729 , n10044 , n10045 );
xor ( n27730 , RI19a869a8_2748 , RI174cf300_766);
not ( n10046 , n27689 );
and ( n10047 , n10046 , RI174cf300_766);
and ( n10048 , n27730 , n27689 );
or ( n27731 , n10047 , n10048 );
xor ( n27732 , n27729 , n27731 );
buf ( n27733 , RI17398f50_2010);
xor ( n27734 , n27732 , n27733 );
buf ( n27735 , RI173e1c40_1655);
xor ( n27736 , n27734 , n27735 );
buf ( n27737 , RI17459a60_1299);
xor ( n27738 , n27736 , n27737 );
xor ( n27739 , n27727 , n27738 );
not ( n27740 , n27739 );
buf ( n27741 , RI173a7500_1940);
xor ( n27742 , RI19a93fe0_2654 , RI1747dbe0_1123);
not ( n10049 , n27689 );
and ( n10050 , n10049 , RI1747dbe0_1123);
and ( n10051 , n27742 , n27689 );
or ( n27743 , n10050 , n10051 );
xor ( n27744 , RI19ac4280_2298 , RI174ce8b0_768);
not ( n10052 , n27689 );
and ( n10053 , n10052 , RI174ce8b0_768);
and ( n10054 , n27744 , n27689 );
or ( n27745 , n10053 , n10054 );
xor ( n27746 , n27743 , n27745 );
buf ( n27747 , RI173988c0_2012);
xor ( n27748 , n27746 , n27747 );
buf ( n27749 , RI173e15b0_1657);
xor ( n27750 , n27748 , n27749 );
buf ( n27751 , RI174593d0_1301);
xor ( n27752 , n27750 , n27751 );
xor ( n27753 , n27741 , n27752 );
xor ( n27754 , RI19aa7e28_2510 , RI1749b118_980);
not ( n10055 , n27689 );
and ( n10056 , n10055 , RI1749b118_980);
and ( n10057 , n27754 , n27689 );
or ( n27755 , n10056 , n10057 );
xor ( n27756 , RI19a89e28_2725 , RI1752d698_625);
not ( n10058 , n27689 );
and ( n10059 , n10058 , RI1752d698_625);
and ( n10060 , n27756 , n27689 );
or ( n27757 , n10059 , n10060 );
xor ( n27758 , n27755 , n27757 );
buf ( n27759 , RI173b5df8_1869);
xor ( n27760 , n27758 , n27759 );
buf ( n27761 , RI173fee30_1513);
xor ( n27762 , n27760 , n27761 );
buf ( n27763 , RI173c2620_1808);
xor ( n27764 , n27762 , n27763 );
xor ( n27765 , n27753 , n27764 );
and ( n27766 , n27740 , n27765 );
xor ( n27767 , n27713 , n27766 );
buf ( n27768 , RI1740fb40_1431);
xor ( n27769 , RI19aaac18_2490 , RI174944d0_1013);
not ( n10061 , n27689 );
and ( n10062 , n10061 , RI174944d0_1013);
and ( n10063 , n27769 , n27689 );
or ( n27770 , n10062 , n10063 );
xor ( n27771 , RI19aa5a88_2525 , RI17522c70_658);
not ( n10064 , n27689 );
and ( n10065 , n10064 , RI17522c70_658);
and ( n10066 , n27771 , n27689 );
or ( n27772 , n10065 , n10066 );
xor ( n27773 , n27770 , n27772 );
buf ( n27774 , RI173af1b0_1902);
xor ( n27775 , n27773 , n27774 );
buf ( n27776 , RI173f7ea0_1547);
xor ( n27777 , n27775 , n27776 );
buf ( n27778 , RI1733d8d0_2141);
xor ( n27779 , n27777 , n27778 );
xor ( n27780 , n27768 , n27779 );
xor ( n27781 , RI19a8d410_2702 , RI17468d30_1225);
not ( n10067 , n27689 );
and ( n10068 , n10067 , RI17468d30_1225);
and ( n10069 , n27781 , n27689 );
or ( n27782 , n10068 , n10069 );
xor ( n27783 , RI19abe4c0_2347 , RI174b1a08_870);
not ( n10070 , n27689 );
and ( n10071 , n10070 , RI174b1a08_870);
and ( n10072 , n27783 , n27689 );
or ( n27784 , n10071 , n10072 );
xor ( n27785 , n27782 , n27784 );
buf ( n27786 , RI17343168_2114);
xor ( n27787 , n27785 , n27786 );
buf ( n27788 , RI173cc6e8_1759);
xor ( n27789 , n27787 , n27788 );
buf ( n27790 , RI17415720_1403);
xor ( n27791 , n27789 , n27790 );
xor ( n27792 , n27780 , n27791 );
not ( n27793 , n27713 );
and ( n27794 , n27793 , n27739 );
xor ( n27795 , n27792 , n27794 );
buf ( n27796 , RI1745d570_1281);
xor ( n27797 , RI19a99698_2616 , RI17473488_1174);
not ( n10073 , n27689 );
and ( n10074 , n10073 , RI17473488_1174);
and ( n10075 , n27797 , n27689 );
or ( n27798 , n10074 , n10075 );
xor ( n27799 , RI19ac90c8_2262 , RI174be6e0_818);
not ( n10076 , n27689 );
and ( n10077 , n10076 , RI174be6e0_818);
and ( n10078 , n27799 , n27689 );
or ( n27800 , n10077 , n10078 );
xor ( n27801 , n27798 , n27800 );
buf ( n27802 , RI1738e4b0_2062);
xor ( n27803 , n27801 , n27802 );
buf ( n27804 , RI173d71a0_1707);
xor ( n27805 , n27803 , n27804 );
buf ( n27806 , RI1744ec78_1352);
xor ( n27807 , n27805 , n27806 );
xor ( n27808 , n27796 , n27807 );
xor ( n27809 , RI19aad468_2473 , RI174909c0_1031);
not ( n10079 , n27689 );
and ( n10080 , n10079 , RI174909c0_1031);
and ( n10081 , n27809 , n27689 );
or ( n27810 , n10080 , n10081 );
xor ( n27811 , RI19abe2e0_2348 , RI1751cfa0_676);
not ( n10082 , n27689 );
and ( n10083 , n10082 , RI1751cfa0_676);
and ( n10084 , n27811 , n27689 );
or ( n27812 , n10083 , n10084 );
xor ( n27813 , n27810 , n27812 );
buf ( n27814 , RI173ab6a0_1920);
xor ( n27815 , n27813 , n27814 );
buf ( n27816 , RI173f4390_1565);
xor ( n27817 , n27815 , n27816 );
buf ( n27818 , RI1750ecc0_720);
xor ( n27819 , n27817 , n27818 );
xor ( n27820 , n27808 , n27819 );
xor ( n27821 , RI19aaa510_2493 , RI17497608_998);
not ( n10085 , n27689 );
and ( n10086 , n10085 , RI17497608_998);
and ( n10087 , n27821 , n27689 );
or ( n27822 , n10086 , n10087 );
xor ( n27823 , RI19aa0970_2564 , RI17488d10_1069);
not ( n10088 , n27689 );
and ( n10089 , n10088 , RI17488d10_1069);
and ( n10090 , n27823 , n27689 );
or ( n27824 , n10089 , n10090 );
xor ( n27825 , RI19acf680_2215 , RI17510bb0_714);
not ( n10091 , n27689 );
and ( n10092 , n10091 , RI17510bb0_714);
and ( n10093 , n27825 , n27689 );
or ( n27826 , n10092 , n10093 );
xor ( n27827 , n27824 , n27826 );
buf ( n27828 , RI173a3d38_1957);
xor ( n27829 , n27827 , n27828 );
buf ( n27830 , RI173eca28_1602);
xor ( n27831 , n27829 , n27830 );
buf ( n27832 , RI17483130_1097);
xor ( n27833 , n27831 , n27832 );
xor ( n27834 , n27822 , n27833 );
xor ( n27835 , RI19ab2148_2439 , RI174a6590_925);
not ( n10094 , n27689 );
and ( n10095 , n10094 , RI174a6590_925);
and ( n10096 , n27835 , n27689 );
or ( n27836 , n10095 , n10096 );
buf ( n27837 , RI17337cf0_2169);
xor ( n27838 , n27836 , n27837 );
buf ( n27839 , RI173c1270_1814);
xor ( n27840 , n27838 , n27839 );
buf ( n27841 , RI17409f60_1459);
xor ( n27842 , n27840 , n27841 );
buf ( n27843 , RI17460d38_1264);
xor ( n27844 , n27842 , n27843 );
xor ( n27845 , n27834 , n27844 );
not ( n27846 , n27845 );
buf ( n27847 , RI17335c20_2179);
xor ( n27848 , RI19aabb90_2484 , RI17495bc8_1006);
not ( n10097 , n27689 );
and ( n10098 , n10097 , RI17495bc8_1006);
and ( n10099 , n27848 , n27689 );
or ( n27849 , n10098 , n10099 );
xor ( n27850 , RI19aaf448_2459 , RI17525088_651);
not ( n10100 , n27689 );
and ( n10101 , n10100 , RI17525088_651);
and ( n10102 , n27850 , n27689 );
or ( n27851 , n10101 , n10102 );
xor ( n27852 , n27849 , n27851 );
buf ( n27853 , RI173b08a8_1895);
xor ( n27854 , n27852 , n27853 );
buf ( n27855 , RI173f9598_1540);
xor ( n27856 , n27854 , n27855 );
buf ( n27857 , RI1738bd50_2074);
xor ( n27858 , n27856 , n27857 );
xor ( n27859 , n27847 , n27858 );
xor ( n27860 , RI19a8bbb0_2713 , RI1746a428_1218);
not ( n10103 , n27689 );
and ( n10104 , n10103 , RI1746a428_1218);
and ( n10105 , n27860 , n27689 );
or ( n27861 , n10104 , n10105 );
xor ( n27862 , RI19abd188_2358 , RI174b3100_863);
not ( n10106 , n27689 );
and ( n10107 , n10106 , RI174b3100_863);
and ( n10108 , n27862 , n27689 );
or ( n27863 , n10107 , n10108 );
xor ( n27864 , n27861 , n27863 );
buf ( n27865 , RI17344860_2107);
xor ( n27866 , n27864 , n27865 );
buf ( n27867 , RI173ce128_1751);
xor ( n27868 , n27866 , n27867 );
buf ( n27869 , RI17445c18_1396);
xor ( n27870 , n27868 , n27869 );
xor ( n27871 , n27859 , n27870 );
and ( n27872 , n27846 , n27871 );
xor ( n27873 , n27820 , n27872 );
xor ( n27874 , n27795 , n27873 );
buf ( n27875 , RI17444ef8_1400);
xor ( n27876 , RI19ab52f8_2415 , RI174a3ae8_938);
not ( n10109 , n27689 );
and ( n10110 , n10109 , RI174a3ae8_938);
and ( n10111 , n27876 , n27689 );
or ( n27877 , n10110 , n10111 );
buf ( n27878 , RI17335590_2181);
xor ( n27879 , n27877 , n27878 );
buf ( n27880 , RI173beb10_1826);
xor ( n27881 , n27879 , n27880 );
buf ( n27882 , RI17407800_1471);
xor ( n27883 , n27881 , n27882 );
buf ( n27884 , RI17447ce8_1386);
xor ( n27885 , n27883 , n27884 );
xor ( n27886 , n27875 , n27885 );
xor ( n27887 , RI19a97dc0_2627 , RI17478690_1149);
not ( n10112 , n27689 );
and ( n10113 , n10112 , RI17478690_1149);
and ( n10114 , n27887 , n27689 );
or ( n27888 , n10113 , n10114 );
xor ( n27889 , RI19ac7b38_2272 , RI174c62a0_794);
not ( n10115 , n27689 );
and ( n10116 , n10115 , RI174c62a0_794);
and ( n10117 , n27889 , n27689 );
or ( n27890 , n10116 , n10117 );
xor ( n27891 , n27888 , n27890 );
buf ( n27892 , RI17393370_2038);
xor ( n27893 , n27891 , n27892 );
buf ( n27894 , RI173dc060_1683);
xor ( n27895 , n27893 , n27894 );
buf ( n27896 , RI17453b38_1328);
xor ( n27897 , n27895 , n27896 );
xor ( n27898 , n27886 , n27897 );
xor ( n27899 , RI19a8ffa8_2683 , RI17465bf8_1240);
not ( n10118 , n27689 );
and ( n10119 , n10118 , RI17465bf8_1240);
and ( n10120 , n27899 , n27689 );
or ( n27900 , n10119 , n10120 );
xor ( n27901 , RI19ac0680_2328 , RI174ae8d0_885);
not ( n10121 , n27689 );
and ( n10122 , n10121 , RI174ae8d0_885);
and ( n10123 , n27901 , n27689 );
or ( n27902 , n10122 , n10123 );
xor ( n27903 , n27900 , n27902 );
buf ( n27904 , RI17340030_2129);
xor ( n27905 , n27903 , n27904 );
buf ( n27906 , RI173c95b0_1774);
xor ( n27907 , n27905 , n27906 );
buf ( n27908 , RI174125e8_1418);
xor ( n27909 , n27907 , n27908 );
xor ( n27910 , n27703 , n27909 );
xor ( n27911 , RI19aa3aa8_2540 , RI17482de8_1098);
not ( n10124 , n27689 );
and ( n10125 , n10124 , RI17482de8_1098);
and ( n10126 , n27911 , n27689 );
or ( n27912 , n10125 , n10126 );
xor ( n27913 , RI19a84e00_2760 , RI17507628_743);
not ( n10127 , n27689 );
and ( n10128 , n10127 , RI17507628_743);
and ( n10129 , n27913 , n27689 );
or ( n27914 , n10128 , n10129 );
xor ( n27915 , n27912 , n27914 );
buf ( n27916 , RI1739dac8_1987);
xor ( n27917 , n27915 , n27916 );
buf ( n27918 , RI173e6b00_1631);
xor ( n27919 , n27917 , n27918 );
buf ( n27920 , RI1745e5d8_1276);
xor ( n27921 , n27919 , n27920 );
xor ( n27922 , n27910 , n27921 );
not ( n27923 , n27922 );
xor ( n27924 , RI19a82f88_2773 , RI17508ff0_738);
not ( n10130 , n27689 );
and ( n10131 , n10130 , RI17508ff0_738);
and ( n10132 , n27924 , n27689 );
or ( n27925 , n10131 , n10132 );
xor ( n27926 , RI19a98630_2623 , RI17475210_1165);
not ( n10133 , n27689 );
and ( n10134 , n10133 , RI17475210_1165);
and ( n10135 , n27926 , n27689 );
or ( n27927 , n10134 , n10135 );
xor ( n27928 , RI19ac81c8_2269 , RI174c1548_809);
not ( n10136 , n27689 );
and ( n10137 , n10136 , RI174c1548_809);
and ( n10138 , n27928 , n27689 );
or ( n27929 , n10137 , n10138 );
xor ( n27930 , n27927 , n27929 );
buf ( n27931 , RI17390238_2053);
xor ( n27932 , n27930 , n27931 );
buf ( n27933 , RI173d8f28_1698);
xor ( n27934 , n27932 , n27933 );
buf ( n27935 , RI17450a00_1343);
xor ( n27936 , n27934 , n27935 );
xor ( n27937 , n27925 , n27936 );
xor ( n27938 , RI19aac6d0_2480 , RI17492a90_1021);
not ( n10139 , n27689 );
and ( n10140 , n10139 , RI17492a90_1021);
and ( n10141 , n27938 , n27689 );
or ( n27939 , n10140 , n10141 );
xor ( n27940 , RI19ab3c00_2425 , RI17520330_666);
not ( n10142 , n27689 );
and ( n10143 , n10142 , RI17520330_666);
and ( n10144 , n27940 , n27689 );
or ( n27941 , n10143 , n10144 );
xor ( n27942 , n27939 , n27941 );
buf ( n27943 , RI173ad770_1910);
xor ( n27944 , n27942 , n27943 );
buf ( n27945 , RI173f6460_1555);
xor ( n27946 , n27944 , n27945 );
buf ( n27947 , RI1752f060_620);
xor ( n27948 , n27946 , n27947 );
xor ( n27949 , n27937 , n27948 );
and ( n27950 , n27923 , n27949 );
xor ( n27951 , n27898 , n27950 );
xor ( n27952 , n27874 , n27951 );
buf ( n27953 , RI174c8be0_786);
xor ( n27954 , RI19aa4a98_2532 , RI174809d0_1109);
not ( n10145 , n27689 );
and ( n10146 , n10145 , RI174809d0_1109);
and ( n10147 , n27954 , n27689 );
or ( n27955 , n10146 , n10147 );
xor ( n27956 , RI19a85e68_2753 , RI17501ef8_754);
not ( n10148 , n27689 );
and ( n10149 , n10148 , RI17501ef8_754);
and ( n10150 , n27956 , n27689 );
or ( n27957 , n10149 , n10150 );
xor ( n27958 , n27955 , n27957 );
buf ( n27959 , RI1739b6b0_1998);
xor ( n27960 , n27958 , n27959 );
buf ( n27961 , RI173e43a0_1643);
xor ( n27962 , n27960 , n27961 );
buf ( n27963 , RI1745c1c0_1287);
xor ( n27964 , n27962 , n27963 );
xor ( n27965 , n27953 , n27964 );
xor ( n27966 , RI19ab8d90_2389 , RI1749df08_966);
not ( n10151 , n27689 );
and ( n10152 , n10151 , RI1749df08_966);
and ( n10153 , n27966 , n27689 );
or ( n27967 , n10152 , n10153 );
buf ( n27968 , RI17531ec8_611);
xor ( n27969 , n27967 , n27968 );
buf ( n27970 , RI173b8f30_1854);
xor ( n27971 , n27969 , n27970 );
buf ( n27972 , RI17401c20_1499);
xor ( n27973 , n27971 , n27972 );
buf ( n27974 , RI173dfeb8_1664);
xor ( n27975 , n27973 , n27974 );
xor ( n27976 , n27965 , n27975 );
xor ( n27977 , RI19ab4380_2422 , RI174a5f00_927);
not ( n10154 , n27689 );
and ( n10155 , n10154 , RI174a5f00_927);
and ( n10156 , n27977 , n27689 );
or ( n27978 , n10155 , n10156 );
xor ( n27979 , RI19aaa330_2494 , RI174972c0_999);
not ( n10157 , n27689 );
and ( n10158 , n10157 , RI174972c0_999);
and ( n10159 , n27979 , n27689 );
or ( n27980 , n10158 , n10159 );
xor ( n27981 , RI19aa12d0_2559 , RI175274a0_644);
not ( n10160 , n27689 );
and ( n10161 , n10160 , RI175274a0_644);
and ( n10162 , n27981 , n27689 );
or ( n27982 , n10161 , n10162 );
xor ( n27983 , n27980 , n27982 );
buf ( n27984 , RI173b1fa0_1888);
xor ( n27985 , n27983 , n27984 );
buf ( n27986 , RI173fac90_1533);
xor ( n27987 , n27985 , n27986 );
buf ( n27988 , RI1739b9f8_1997);
xor ( n27989 , n27987 , n27988 );
xor ( n27990 , n27978 , n27989 );
xor ( n27991 , RI19a8cb28_2706 , RI1746bb20_1211);
not ( n10163 , n27689 );
and ( n10164 , n10163 , RI1746bb20_1211);
and ( n10165 , n27991 , n27689 );
or ( n27992 , n10164 , n10165 );
xor ( n27993 , RI19abddb8_2351 , RI174b47f8_856);
not ( n10166 , n27689 );
and ( n10167 , n10166 , RI174b47f8_856);
and ( n10168 , n27993 , n27689 );
or ( n27994 , n10167 , n10168 );
xor ( n27995 , n27992 , n27994 );
buf ( n27996 , RI17345f58_2100);
xor ( n27997 , n27995 , n27996 );
buf ( n27998 , RI173cf820_1744);
xor ( n27999 , n27997 , n27998 );
buf ( n28000 , RI17447310_1389);
xor ( n28001 , n27999 , n28000 );
xor ( n28002 , n27990 , n28001 );
not ( n28003 , n28002 );
xor ( n28004 , RI19abcdc8_2360 , RI174b6580_847);
not ( n10169 , n27689 );
and ( n10170 , n10169 , RI174b6580_847);
and ( n10171 , n28004 , n27689 );
or ( n28005 , n10170 , n10171 );
xor ( n28006 , RI19ab3138_2431 , RI174a7fd0_917);
not ( n10172 , n27689 );
and ( n10173 , n10172 , RI174a7fd0_917);
and ( n10174 , n28006 , n27689 );
or ( n28007 , n10173 , n10174 );
buf ( n28008 , RI17339730_2161);
xor ( n28009 , n28007 , n28008 );
buf ( n28010 , RI173c2cb0_1806);
xor ( n28011 , n28009 , n28010 );
buf ( n28012 , RI1740b9a0_1451);
xor ( n28013 , n28011 , n28012 );
buf ( n28014 , RI173895f0_2086);
xor ( n28015 , n28013 , n28014 );
xor ( n28016 , n28005 , n28015 );
xor ( n28017 , RI19a93068_2661 , RI1747c830_1129);
not ( n10175 , n27689 );
and ( n10176 , n10175 , RI1747c830_1129);
and ( n10177 , n28017 , n27689 );
or ( n28018 , n10176 , n10177 );
xor ( n28019 , RI19ac3290_2305 , RI174cc9c0_774);
not ( n10178 , n27689 );
and ( n10179 , n10178 , RI174cc9c0_774);
and ( n10180 , n28019 , n27689 );
or ( n28020 , n10179 , n10180 );
xor ( n28021 , n28018 , n28020 );
buf ( n28022 , RI17397510_2018);
xor ( n28023 , n28021 , n28022 );
buf ( n28024 , RI173e0200_1663);
xor ( n28025 , n28023 , n28024 );
buf ( n28026 , RI17458020_1307);
xor ( n28027 , n28025 , n28026 );
xor ( n28028 , n28016 , n28027 );
and ( n28029 , n28003 , n28028 );
xor ( n28030 , n27976 , n28029 );
xor ( n28031 , n27952 , n28030 );
buf ( n28032 , RI1744fce0_1347);
xor ( n28033 , RI19a90188_2682 , RI17465f40_1239);
not ( n10181 , n27689 );
and ( n10182 , n10181 , RI17465f40_1239);
and ( n10183 , n28033 , n27689 );
or ( n28034 , n10182 , n10183 );
xor ( n28035 , RI19ac0860_2327 , RI174aec18_884);
not ( n10184 , n27689 );
and ( n10185 , n10184 , RI174aec18_884);
and ( n10186 , n28035 , n27689 );
or ( n28036 , n10185 , n10186 );
xor ( n28037 , n28034 , n28036 );
buf ( n28038 , RI17340378_2128);
xor ( n28039 , n28037 , n28038 );
buf ( n28040 , RI173c98f8_1773);
xor ( n28041 , n28039 , n28040 );
buf ( n28042 , RI17412930_1417);
xor ( n28043 , n28041 , n28042 );
xor ( n28044 , n28032 , n28043 );
xor ( n28045 , RI19aa3c88_2539 , RI17483478_1096);
not ( n10187 , n27689 );
and ( n10188 , n10187 , RI17483478_1096);
and ( n10189 , n28045 , n27689 );
or ( n28046 , n10188 , n10189 );
xor ( n28047 , RI19a85058_2759 , RI17508078_741);
not ( n10190 , n27689 );
and ( n10191 , n10190 , RI17508078_741);
and ( n10192 , n28047 , n27689 );
or ( n28048 , n10191 , n10192 );
xor ( n28049 , n28046 , n28048 );
buf ( n28050 , RI1739e158_1985);
xor ( n28051 , n28049 , n28050 );
buf ( n28052 , RI173e7190_1629);
xor ( n28053 , n28051 , n28052 );
buf ( n28054 , RI1745ec68_1274);
xor ( n28055 , n28053 , n28054 );
xor ( n28056 , n28044 , n28055 );
xor ( n28057 , RI19aa3238_2544 , RI174820c8_1102);
not ( n10193 , n27689 );
and ( n10194 , n10193 , RI174820c8_1102);
and ( n10195 , n28057 , n27689 );
or ( n28058 , n10194 , n10195 );
xor ( n28059 , RI19a998f0_2615 , RI174737d0_1173);
not ( n10196 , n27689 );
and ( n10197 , n10196 , RI174737d0_1173);
and ( n10198 , n28059 , n27689 );
or ( n28060 , n10197 , n10198 );
xor ( n28061 , RI19ac92a8_2261 , RI174bec08_817);
not ( n10199 , n27689 );
and ( n10200 , n10199 , RI174bec08_817);
and ( n10201 , n28061 , n27689 );
or ( n28062 , n10200 , n10201 );
xor ( n28063 , n28060 , n28062 );
buf ( n28064 , RI1738e7f8_2061);
xor ( n28065 , n28063 , n28064 );
buf ( n28066 , RI173d74e8_1706);
xor ( n28067 , n28065 , n28066 );
buf ( n28068 , RI1744efc0_1351);
xor ( n28069 , n28067 , n28068 );
xor ( n28070 , n28058 , n28069 );
xor ( n28071 , RI19aad648_2472 , RI17491050_1029);
not ( n10202 , n27689 );
and ( n10203 , n10202 , RI17491050_1029);
and ( n10204 , n28071 , n27689 );
or ( n28072 , n10203 , n10204 );
xor ( n28073 , RI19abf690_2337 , RI1751d9f0_674);
not ( n10205 , n27689 );
and ( n10206 , n10205 , RI1751d9f0_674);
and ( n10207 , n28073 , n27689 );
or ( n28074 , n10206 , n10207 );
xor ( n28075 , n28072 , n28074 );
buf ( n28076 , RI173abd30_1918);
xor ( n28077 , n28075 , n28076 );
buf ( n28078 , RI173f4a20_1563);
xor ( n28079 , n28077 , n28078 );
buf ( n28080 , RI17512aa0_708);
xor ( n28081 , n28079 , n28080 );
xor ( n28082 , n28070 , n28081 );
not ( n28083 , n28082 );
xor ( n28084 , RI19a23678_2793 , RI1751ab88_683);
not ( n10208 , n27689 );
and ( n10209 , n10208 , RI1751ab88_683);
and ( n10210 , n28084 , n27689 );
or ( n28085 , n10209 , n10210 );
xor ( n28086 , RI19aa48b8_2533 , RI17480688_1110);
not ( n10211 , n27689 );
and ( n10212 , n10211 , RI17480688_1110);
and ( n10213 , n28086 , n27689 );
or ( n28087 , n10212 , n10213 );
xor ( n28088 , RI19a85c10_2754 , RI175019d0_755);
not ( n10214 , n27689 );
and ( n10215 , n10214 , RI175019d0_755);
and ( n10216 , n28088 , n27689 );
or ( n28089 , n10215 , n10216 );
xor ( n28090 , n28087 , n28089 );
buf ( n28091 , RI1739b368_1999);
xor ( n28092 , n28090 , n28091 );
buf ( n28093 , RI173e4058_1644);
xor ( n28094 , n28092 , n28093 );
buf ( n28095 , RI1745be78_1288);
xor ( n28096 , n28094 , n28095 );
xor ( n28097 , n28085 , n28096 );
xor ( n28098 , RI19ab8b38_2390 , RI1749dbc0_967);
not ( n10217 , n27689 );
and ( n10218 , n10217 , RI1749dbc0_967);
and ( n10219 , n28098 , n27689 );
or ( n28099 , n10218 , n10219 );
buf ( n28100 , RI175319a0_612);
xor ( n28101 , n28099 , n28100 );
buf ( n28102 , RI173b8be8_1855);
xor ( n28103 , n28101 , n28102 );
buf ( n28104 , RI174018d8_1500);
xor ( n28105 , n28103 , n28104 );
buf ( n28106 , RI173ddaa0_1675);
xor ( n28107 , n28105 , n28106 );
xor ( n28108 , n28097 , n28107 );
and ( n28109 , n28083 , n28108 );
xor ( n28110 , n28056 , n28109 );
xor ( n28111 , n28031 , n28110 );
xor ( n28112 , n27767 , n28111 );
xor ( n28113 , RI19acb300_2246 , RI174b8650_837);
not ( n10220 , n27689 );
and ( n10221 , n10220 , RI174b8650_837);
and ( n10222 , n28113 , n27689 );
or ( n28114 , n10221 , n10222 );
xor ( n28115 , RI19a91e98_2669 , RI174613c8_1262);
not ( n10223 , n27689 );
and ( n10224 , n10223 , RI174613c8_1262);
and ( n10225 , n28115 , n27689 );
or ( n28116 , n10224 , n10225 );
xor ( n28117 , RI19ac21b0_2313 , RI174aa0a0_907);
not ( n10226 , n27689 );
and ( n10227 , n10226 , RI174aa0a0_907);
and ( n10228 , n28117 , n27689 );
or ( n28118 , n10227 , n10228 );
xor ( n28119 , n28116 , n28118 );
buf ( n28120 , RI1733b800_2151);
xor ( n28121 , n28119 , n28120 );
buf ( n28122 , RI173c4d80_1796);
xor ( n28123 , n28121 , n28122 );
buf ( n28124 , RI1740da70_1441);
xor ( n28125 , n28123 , n28124 );
xor ( n28126 , n28114 , n28125 );
xor ( n28127 , RI19aa5740_2526 , RI1747e5b8_1120);
not ( n10229 , n27689 );
and ( n10230 , n10229 , RI1747e5b8_1120);
and ( n10231 , n28127 , n27689 );
or ( n28128 , n10230 , n10231 );
xor ( n28129 , RI19a86c00_2747 , RI174cf828_765);
not ( n10232 , n27689 );
and ( n10233 , n10232 , RI174cf828_765);
and ( n10234 , n28129 , n27689 );
or ( n28130 , n10233 , n10234 );
xor ( n28131 , n28128 , n28130 );
buf ( n28132 , RI17399298_2009);
xor ( n28133 , n28131 , n28132 );
buf ( n28134 , RI173e1f88_1654);
xor ( n28135 , n28133 , n28134 );
buf ( n28136 , RI17459da8_1298);
xor ( n28137 , n28135 , n28136 );
xor ( n28138 , n28126 , n28137 );
buf ( n28139 , RI173a7848_1939);
xor ( n28140 , RI19a94238_2653 , RI1747df28_1122);
not ( n10235 , n27689 );
and ( n10236 , n10235 , RI1747df28_1122);
and ( n10237 , n28140 , n27689 );
or ( n28141 , n10236 , n10237 );
xor ( n28142 , n28141 , n27715 );
buf ( n28143 , RI17398c08_2011);
xor ( n28144 , n28142 , n28143 );
buf ( n28145 , RI173e18f8_1656);
xor ( n28146 , n28144 , n28145 );
buf ( n28147 , RI17459718_1300);
xor ( n28148 , n28146 , n28147 );
xor ( n28149 , n28139 , n28148 );
xor ( n28150 , RI19aafad8_2456 , RI1748cb68_1050);
not ( n10238 , n27689 );
and ( n10239 , n10238 , RI1748cb68_1050);
and ( n10240 , n28150 , n27689 );
or ( n28151 , n10239 , n10240 );
xor ( n28152 , RI19a85508_2757 , RI175172d0_694);
not ( n10241 , n27689 );
and ( n10242 , n10241 , RI175172d0_694);
and ( n10243 , n28152 , n27689 );
or ( n28153 , n10242 , n10243 );
xor ( n28154 , n28151 , n28153 );
buf ( n28155 , RI173a7b90_1938);
xor ( n28156 , n28154 , n28155 );
buf ( n28157 , RI173f0880_1583);
xor ( n28158 , n28156 , n28157 );
buf ( n28159 , RI174a9d58_908);
xor ( n28160 , n28158 , n28159 );
xor ( n28161 , n28149 , n28160 );
not ( n28162 , n28161 );
buf ( n28163 , RI173f9c28_1538);
xor ( n28164 , RI19a9fae8_2571 , RI17487618_1076);
not ( n10244 , n27689 );
and ( n10245 , n10244 , RI17487618_1076);
and ( n10246 , n28164 , n27689 );
or ( n28165 , n10245 , n10246 );
xor ( n28166 , RI19ace870_2221 , RI1750e798_721);
not ( n10247 , n27689 );
and ( n10248 , n10247 , RI1750e798_721);
and ( n10249 , n28166 , n27689 );
or ( n28167 , n10248 , n10249 );
xor ( n28168 , n28165 , n28167 );
buf ( n28169 , RI173a2640_1964);
xor ( n28170 , n28168 , n28169 );
buf ( n28171 , RI173eb330_1609);
xor ( n28172 , n28170 , n28171 );
buf ( n28173 , RI17475558_1164);
xor ( n28174 , n28172 , n28173 );
xor ( n28175 , n28163 , n28174 );
xor ( n28176 , RI19ab36d8_2428 , RI174a4b50_933);
not ( n10250 , n27689 );
and ( n10251 , n10250 , RI174a4b50_933);
and ( n10252 , n28176 , n27689 );
or ( n28177 , n10251 , n10252 );
buf ( n28178 , RI173365f8_2176);
xor ( n28179 , n28177 , n28178 );
buf ( n28180 , RI173bfb78_1821);
xor ( n28181 , n28179 , n28180 );
buf ( n28182 , RI17408868_1466);
xor ( n28183 , n28181 , n28182 );
buf ( n28184 , RI17453160_1331);
xor ( n28185 , n28183 , n28184 );
xor ( n28186 , n28175 , n28185 );
and ( n28187 , n28162 , n28186 );
xor ( n28188 , n28138 , n28187 );
buf ( n28189 , RI17335f68_2178);
xor ( n28190 , RI19aa9688_2500 , RI17495f10_1005);
not ( n10253 , n27689 );
and ( n10254 , n10253 , RI17495f10_1005);
and ( n10255 , n28190 , n27689 );
or ( n28191 , n10254 , n10255 );
xor ( n28192 , RI19a981f8_2625 , RI175255b0_650);
not ( n10256 , n27689 );
and ( n10257 , n10256 , RI175255b0_650);
and ( n10258 , n28192 , n27689 );
or ( n28193 , n10257 , n10258 );
xor ( n28194 , n28191 , n28193 );
buf ( n28195 , RI173b0bf0_1894);
xor ( n28196 , n28194 , n28195 );
buf ( n28197 , RI173f98e0_1539);
xor ( n28198 , n28196 , n28197 );
buf ( n28199 , RI1738e168_2063);
xor ( n28200 , n28198 , n28199 );
xor ( n28201 , n28189 , n28200 );
xor ( n28202 , RI19a8be08_2712 , RI1746a770_1217);
not ( n10259 , n27689 );
and ( n10260 , n10259 , RI1746a770_1217);
and ( n10261 , n28202 , n27689 );
or ( n28203 , n10260 , n10261 );
xor ( n28204 , RI19abd2f0_2357 , RI174b3448_862);
not ( n10262 , n27689 );
and ( n10263 , n10262 , RI174b3448_862);
and ( n10264 , n28204 , n27689 );
or ( n28205 , n10263 , n10264 );
xor ( n28206 , n28203 , n28205 );
buf ( n28207 , RI17344ba8_2106);
xor ( n28208 , n28206 , n28207 );
buf ( n28209 , RI173ce470_1750);
xor ( n28210 , n28208 , n28209 );
buf ( n28211 , RI17445f60_1395);
xor ( n28212 , n28210 , n28211 );
xor ( n28213 , n28201 , n28212 );
buf ( n28214 , RI17340a08_2126);
xor ( n28215 , RI19ab7f80_2395 , RI174a0668_954);
not ( n10265 , n27689 );
and ( n10266 , n10265 , RI174a0668_954);
and ( n10267 , n28215 , n27689 );
or ( n28216 , n10266 , n10267 );
buf ( n28217 , RI17535ca8_599);
xor ( n28218 , n28216 , n28217 );
buf ( n28219 , RI173bb690_1842);
xor ( n28220 , n28218 , n28219 );
buf ( n28221 , RI17404380_1487);
xor ( n28222 , n28220 , n28221 );
buf ( n28223 , RI173f8f08_1542);
xor ( n28224 , n28222 , n28223 );
xor ( n28225 , n28214 , n28224 );
xor ( n28226 , RI19a983d8_2624 , RI17474ec8_1166);
not ( n10268 , n27689 );
and ( n10269 , n10268 , RI17474ec8_1166);
and ( n10270 , n28226 , n27689 );
or ( n28227 , n10269 , n10270 );
xor ( n28228 , RI19ac7f70_2270 , RI174c1020_810);
not ( n10271 , n27689 );
and ( n10272 , n10271 , RI174c1020_810);
and ( n10273 , n28228 , n27689 );
or ( n28229 , n10272 , n10273 );
xor ( n28230 , n28227 , n28229 );
buf ( n28231 , RI1738fef0_2054);
xor ( n28232 , n28230 , n28231 );
buf ( n28233 , RI173d8be0_1699);
xor ( n28234 , n28232 , n28233 );
buf ( n28235 , RI174506b8_1344);
xor ( n28236 , n28234 , n28235 );
xor ( n28237 , n28225 , n28236 );
not ( n28238 , n28237 );
buf ( n28239 , RI173d39d8_1724);
xor ( n28240 , RI19a920f0_2668 , RI17461710_1261);
not ( n10274 , n27689 );
and ( n10275 , n10274 , RI17461710_1261);
and ( n10276 , n28240 , n27689 );
or ( n28241 , n10275 , n10276 );
xor ( n28242 , RI19ac2390_2312 , RI174aa3e8_906);
not ( n10277 , n27689 );
and ( n10278 , n10277 , RI174aa3e8_906);
and ( n10279 , n28242 , n27689 );
or ( n28243 , n10278 , n10279 );
xor ( n28244 , n28241 , n28243 );
buf ( n28245 , RI1733bb48_2150);
xor ( n28246 , n28244 , n28245 );
buf ( n28247 , RI173c50c8_1795);
xor ( n28248 , n28246 , n28247 );
buf ( n28249 , RI1740ddb8_1440);
xor ( n28250 , n28248 , n28249 );
xor ( n28251 , n28239 , n28250 );
xor ( n28252 , RI19aa5dd0_2524 , RI1747ec48_1118);
not ( n10280 , n27689 );
and ( n10281 , n10280 , RI1747ec48_1118);
and ( n10282 , n28252 , n27689 );
or ( n28253 , n10281 , n10282 );
xor ( n28254 , RI19a86fc0_2745 , RI174d0278_763);
not ( n10283 , n27689 );
and ( n10284 , n10283 , RI174d0278_763);
and ( n10285 , n28254 , n27689 );
or ( n28255 , n10284 , n10285 );
xor ( n28256 , n28253 , n28255 );
buf ( n28257 , RI17399928_2007);
xor ( n28258 , n28256 , n28257 );
buf ( n28259 , RI173e2618_1652);
xor ( n28260 , n28258 , n28259 );
buf ( n28261 , RI1745a438_1296);
xor ( n28262 , n28260 , n28261 );
xor ( n28263 , n28251 , n28262 );
and ( n28264 , n28238 , n28263 );
xor ( n28265 , n28213 , n28264 );
xor ( n28266 , n28188 , n28265 );
xor ( n28267 , RI19a831e0_2772 , RI17509518_737);
not ( n10286 , n27689 );
and ( n10287 , n10286 , RI17509518_737);
and ( n10288 , n28267 , n27689 );
or ( n28268 , n10287 , n10288 );
xor ( n28269 , RI19a98888_2622 , RI174758a0_1163);
not ( n10289 , n27689 );
and ( n10290 , n10289 , RI174758a0_1163);
and ( n10291 , n28269 , n27689 );
or ( n28270 , n10290 , n10291 );
xor ( n28271 , RI19ac8330_2268 , RI174c1f98_807);
not ( n10292 , n27689 );
and ( n10293 , n10292 , RI174c1f98_807);
and ( n10294 , n28271 , n27689 );
or ( n28272 , n10293 , n10294 );
xor ( n28273 , n28270 , n28272 );
buf ( n28274 , RI173908c8_2051);
xor ( n28275 , n28273 , n28274 );
buf ( n28276 , RI173d95b8_1696);
xor ( n28277 , n28275 , n28276 );
buf ( n28278 , RI17451090_1341);
xor ( n28279 , n28277 , n28278 );
xor ( n28280 , n28268 , n28279 );
xor ( n28281 , RI19aac838_2479 , RI17492dd8_1020);
not ( n10295 , n27689 );
and ( n10296 , n10295 , RI17492dd8_1020);
and ( n10297 , n28281 , n27689 );
or ( n28282 , n10296 , n10297 );
xor ( n28283 , RI19ab54d8_2414 , RI17520858_665);
not ( n10298 , n27689 );
and ( n10299 , n10298 , RI17520858_665);
and ( n10300 , n28283 , n27689 );
or ( n28284 , n10299 , n10300 );
xor ( n28285 , n28282 , n28284 );
buf ( n28286 , RI173adab8_1909);
xor ( n28287 , n28285 , n28286 );
buf ( n28288 , RI173f67a8_1554);
xor ( n28289 , n28287 , n28288 );
buf ( n28290 , RI17532918_609);
xor ( n28291 , n28289 , n28290 );
xor ( n28292 , n28280 , n28291 );
buf ( n28293 , RI173b1c58_1889);
xor ( n28294 , RI19aa05b0_2566 , RI17488680_1071);
not ( n10301 , n27689 );
and ( n10302 , n10301 , RI17488680_1071);
and ( n10303 , n28294 , n27689 );
or ( n28295 , n10302 , n10303 );
xor ( n28296 , RI19acf1d0_2217 , RI17510160_716);
not ( n10304 , n27689 );
and ( n10305 , n10304 , RI17510160_716);
and ( n10306 , n28296 , n27689 );
or ( n28297 , n10305 , n10306 );
xor ( n28298 , n28295 , n28297 );
buf ( n28299 , RI173a36a8_1959);
xor ( n28300 , n28298 , n28299 );
buf ( n28301 , RI173ec398_1604);
xor ( n28302 , n28300 , n28301 );
buf ( n28303 , RI1747e900_1119);
xor ( n28304 , n28302 , n28303 );
xor ( n28305 , n28293 , n28304 );
buf ( n28306 , RI17337660_2171);
xor ( n28307 , n27978 , n28306 );
buf ( n28308 , RI173c0be0_1816);
xor ( n28309 , n28307 , n28308 );
buf ( n28310 , RI174098d0_1461);
xor ( n28311 , n28309 , n28310 );
buf ( n28312 , RI1745c508_1286);
xor ( n28313 , n28311 , n28312 );
xor ( n28314 , n28305 , n28313 );
not ( n28315 , n28314 );
buf ( n28316 , RI17405730_1481);
xor ( n28317 , RI19aaca18_2478 , RI17493468_1018);
not ( n10307 , n27689 );
and ( n10308 , n10307 , RI17493468_1018);
and ( n10309 , n28317 , n27689 );
or ( n28318 , n10308 , n10309 );
xor ( n28319 , RI19ab6cc0_2403 , RI175212a8_663);
not ( n10310 , n27689 );
and ( n10311 , n10310 , RI175212a8_663);
and ( n10312 , n28319 , n27689 );
or ( n28320 , n10311 , n10312 );
xor ( n28321 , n28318 , n28320 );
buf ( n28322 , RI173ae148_1907);
xor ( n28323 , n28321 , n28322 );
buf ( n28324 , RI173f6e38_1552);
xor ( n28325 , n28323 , n28324 );
buf ( n28326 , RI17332458_2196);
xor ( n28327 , n28325 , n28326 );
xor ( n28328 , n28316 , n28327 );
xor ( n28329 , RI19a8efb8_2690 , RI17467980_1231);
not ( n10313 , n27689 );
and ( n10314 , n10313 , RI17467980_1231);
and ( n10315 , n28329 , n27689 );
or ( n28330 , n10314 , n10315 );
xor ( n28331 , RI19abfa50_2335 , RI174b0658_876);
not ( n10316 , n27689 );
and ( n10317 , n10316 , RI174b0658_876);
and ( n10318 , n28331 , n27689 );
or ( n28332 , n10317 , n10318 );
xor ( n28333 , n28330 , n28332 );
buf ( n28334 , RI17341db8_2120);
xor ( n28335 , n28333 , n28334 );
buf ( n28336 , RI173cb338_1765);
xor ( n28337 , n28335 , n28336 );
buf ( n28338 , RI17414370_1409);
xor ( n28339 , n28337 , n28338 );
xor ( n28340 , n28328 , n28339 );
and ( n28341 , n28315 , n28340 );
xor ( n28342 , n28292 , n28341 );
xor ( n28343 , n28266 , n28342 );
xor ( n28344 , RI19abaa28_2376 , RI174b68c8_846);
not ( n10319 , n27689 );
and ( n10320 , n10319 , RI174b68c8_846);
and ( n10321 , n28344 , n27689 );
or ( n28345 , n10320 , n10321 );
xor ( n28346 , RI19ab0e10_2447 , RI174a8318_916);
not ( n10322 , n27689 );
and ( n10323 , n10322 , RI174a8318_916);
and ( n10324 , n28346 , n27689 );
or ( n28347 , n10323 , n10324 );
buf ( n28348 , RI17339a78_2160);
xor ( n28349 , n28347 , n28348 );
buf ( n28350 , RI173c2ff8_1805);
xor ( n28351 , n28349 , n28350 );
buf ( n28352 , RI1740bce8_1450);
xor ( n28353 , n28351 , n28352 );
buf ( n28354 , RI173a0228_1975);
xor ( n28355 , n28353 , n28354 );
xor ( n28356 , n28345 , n28355 );
xor ( n28357 , RI19a932c0_2660 , RI1747cb78_1128);
not ( n10325 , n27689 );
and ( n10326 , n10325 , RI1747cb78_1128);
and ( n10327 , n28357 , n27689 );
or ( n28358 , n10326 , n10327 );
xor ( n28359 , RI19ac34e8_2304 , RI174ccee8_773);
not ( n10328 , n27689 );
and ( n10329 , n10328 , RI174ccee8_773);
and ( n10330 , n28359 , n27689 );
or ( n28360 , n10329 , n10330 );
xor ( n28361 , n28358 , n28360 );
buf ( n28362 , RI17397858_2017);
xor ( n28363 , n28361 , n28362 );
buf ( n28364 , RI173e0548_1662);
xor ( n28365 , n28363 , n28364 );
buf ( n28366 , RI17458368_1306);
xor ( n28367 , n28365 , n28366 );
xor ( n28368 , n28356 , n28367 );
buf ( n28369 , RI173915e8_2047);
xor ( n28370 , RI19a8f210_2689 , RI17468010_1229);
not ( n10331 , n27689 );
and ( n10332 , n10331 , RI17468010_1229);
and ( n10333 , n28370 , n27689 );
or ( n28371 , n10332 , n10333 );
xor ( n28372 , RI19abfc30_2334 , RI174b0ce8_874);
not ( n10334 , n27689 );
and ( n10335 , n10334 , RI174b0ce8_874);
and ( n10336 , n28372 , n27689 );
or ( n28373 , n10335 , n10336 );
xor ( n28374 , n28371 , n28373 );
buf ( n28375 , RI17342448_2118);
xor ( n28376 , n28374 , n28375 );
buf ( n28377 , RI173cb9c8_1763);
xor ( n28378 , n28376 , n28377 );
buf ( n28379 , RI17414a00_1407);
xor ( n28380 , n28378 , n28379 );
xor ( n28381 , n28369 , n28380 );
xor ( n28382 , RI19aa2e78_2546 , RI17485200_1087);
not ( n10337 , n27689 );
and ( n10338 , n10337 , RI17485200_1087);
and ( n10339 , n28382 , n27689 );
or ( n28383 , n10338 , n10339 );
xor ( n28384 , RI19a83f78_2766 , RI1750aee0_732);
not ( n10340 , n27689 );
and ( n10341 , n10340 , RI1750aee0_732);
and ( n10342 , n28384 , n27689 );
or ( n28385 , n10341 , n10342 );
xor ( n28386 , n28383 , n28385 );
buf ( n28387 , RI1739fee0_1976);
xor ( n28388 , n28386 , n28387 );
buf ( n28389 , RI173e8f18_1620);
xor ( n28390 , n28388 , n28389 );
buf ( n28391 , RI174609f0_1265);
xor ( n28392 , n28390 , n28391 );
xor ( n28393 , n28381 , n28392 );
not ( n28394 , n28393 );
buf ( n28395 , RI173e9f80_1615);
xor ( n28396 , RI19a976b8_2630 , RI17477628_1154);
not ( n10343 , n27689 );
and ( n10344 , n10343 , RI17477628_1154);
and ( n10345 , n28396 , n27689 );
or ( n28397 , n10344 , n10345 );
xor ( n28398 , RI19ac74a8_2275 , RI174c4e00_798);
not ( n10346 , n27689 );
and ( n10347 , n10346 , RI174c4e00_798);
and ( n10348 , n28398 , n27689 );
or ( n28399 , n10347 , n10348 );
xor ( n28400 , n28397 , n28399 );
buf ( n28401 , RI17392650_2042);
xor ( n28402 , n28400 , n28401 );
buf ( n28403 , RI173db340_1687);
xor ( n28404 , n28402 , n28403 );
buf ( n28405 , RI17452e18_1332);
xor ( n28406 , n28404 , n28405 );
xor ( n28407 , n28395 , n28406 );
xor ( n28408 , RI19aab410_2487 , RI17494ea8_1010);
not ( n10349 , n27689 );
and ( n10350 , n10349 , RI17494ea8_1010);
and ( n10351 , n28408 , n27689 );
or ( n28409 , n10350 , n10351 );
xor ( n28410 , RI19aaa858_2492 , RI17523be8_655);
not ( n10352 , n27689 );
and ( n10353 , n10352 , RI17523be8_655);
and ( n10354 , n28410 , n27689 );
or ( n28411 , n10353 , n10354 );
xor ( n28412 , n28409 , n28411 );
buf ( n28413 , RI173afb88_1899);
xor ( n28414 , n28412 , n28413 );
buf ( n28415 , RI173f8878_1544);
xor ( n28416 , n28414 , n28415 );
buf ( n28417 , RI17344518_2108);
xor ( n28418 , n28416 , n28417 );
xor ( n28419 , n28407 , n28418 );
and ( n28420 , n28394 , n28419 );
xor ( n28421 , n28368 , n28420 );
xor ( n28422 , n28343 , n28421 );
xor ( n28423 , RI19a23858_2792 , RI1751b0b0_682);
not ( n10355 , n27689 );
and ( n10356 , n10355 , RI1751b0b0_682);
and ( n10357 , n28423 , n27689 );
or ( n28424 , n10356 , n10357 );
xor ( n28425 , n28424 , n27964 );
xor ( n28426 , n28425 , n27975 );
buf ( n28427 , RI173c39d0_1802);
xor ( n28428 , RI19aa71f8_2515 , RI1749a3f8_984);
not ( n10358 , n27689 );
and ( n10359 , n10358 , RI1749a3f8_984);
and ( n10360 , n28428 , n27689 );
or ( n28429 , n10359 , n10360 );
xor ( n28430 , RI19a88460_2736 , RI1752c1f8_629);
not ( n10361 , n27689 );
and ( n10362 , n10361 , RI1752c1f8_629);
and ( n10363 , n28430 , n27689 );
or ( n28431 , n10362 , n10363 );
xor ( n28432 , n28429 , n28431 );
buf ( n28433 , RI173b50d8_1873);
xor ( n28434 , n28432 , n28433 );
buf ( n28435 , RI173fe110_1517);
xor ( n28436 , n28434 , n28435 );
buf ( n28437 , RI173b95c0_1852);
xor ( n28438 , n28436 , n28437 );
xor ( n28439 , n28427 , n28438 );
xor ( n28440 , RI19a89888_2727 , RI1746ec58_1196);
not ( n10364 , n27689 );
and ( n10365 , n10364 , RI1746ec58_1196);
and ( n10366 , n28440 , n27689 );
or ( n28441 , n10365 , n10366 );
xor ( n28442 , RI19abb5e0_2372 , RI174b7930_841);
not ( n10367 , n27689 );
and ( n10368 , n10367 , RI174b7930_841);
and ( n10369 , n28442 , n27689 );
or ( n28443 , n10368 , n10369 );
xor ( n28444 , n28441 , n28443 );
buf ( n28445 , RI17389c80_2084);
xor ( n28446 , n28444 , n28445 );
buf ( n28447 , RI173d2970_1729);
xor ( n28448 , n28446 , n28447 );
buf ( n28449 , RI1744a448_1374);
xor ( n28450 , n28448 , n28449 );
xor ( n28451 , n28439 , n28450 );
not ( n28452 , n28451 );
buf ( n28453 , RI173d2cb8_1728);
xor ( n28454 , RI19ab1860_2442 , RI174a9380_911);
not ( n10370 , n27689 );
and ( n10371 , n10370 , RI174a9380_911);
and ( n10372 , n28454 , n27689 );
or ( n28455 , n10371 , n10372 );
buf ( n28456 , RI1733aae0_2155);
xor ( n28457 , n28455 , n28456 );
buf ( n28458 , RI173c4060_1800);
xor ( n28459 , n28457 , n28458 );
buf ( n28460 , RI1740cd50_1445);
xor ( n28461 , n28459 , n28460 );
buf ( n28462 , RI17411f58_1420);
xor ( n28463 , n28461 , n28462 );
xor ( n28464 , n28453 , n28463 );
xor ( n28465 , n28464 , n27752 );
and ( n28466 , n28452 , n28465 );
xor ( n28467 , n28426 , n28466 );
xor ( n28468 , n28422 , n28467 );
xor ( n28469 , n28112 , n28468 );
xor ( n28470 , RI19aad828_2471 , RI17491398_1028);
not ( n10373 , n27689 );
and ( n10374 , n10373 , RI17491398_1028);
and ( n10375 , n28470 , n27689 );
or ( n28471 , n10374 , n10375 );
xor ( n28472 , RI19ac0a40_2326 , RI1751df18_673);
not ( n10376 , n27689 );
and ( n10377 , n10376 , RI1751df18_673);
and ( n10378 , n28472 , n27689 );
or ( n28473 , n10377 , n10378 );
xor ( n28474 , n28471 , n28473 );
buf ( n28475 , RI173ac078_1917);
xor ( n28476 , n28474 , n28475 );
buf ( n28477 , RI173f4d68_1562);
xor ( n28478 , n28476 , n28477 );
buf ( n28479 , RI17516358_697);
xor ( n28480 , n28478 , n28479 );
xor ( n28481 , n27693 , n28480 );
xor ( n28482 , n28481 , n27909 );
buf ( n28483 , RI1733be90_2149);
xor ( n28484 , RI19ab9a38_2383 , RI1749baf0_977);
not ( n10379 , n27689 );
and ( n10380 , n10379 , RI1749baf0_977);
and ( n10381 , n28484 , n27689 );
or ( n28485 , n10380 , n10381 );
buf ( n28486 , RI1752e610_622);
xor ( n28487 , n28485 , n28486 );
buf ( n28488 , RI173b67d0_1866);
xor ( n28489 , n28487 , n28488 );
buf ( n28490 , RI173ff808_1510);
xor ( n28491 , n28489 , n28490 );
buf ( n28492 , RI173c9268_1775);
xor ( n28493 , n28491 , n28492 );
xor ( n28494 , n28483 , n28493 );
xor ( n28495 , RI19a9c5f0_2595 , RI17470350_1189);
not ( n10382 , n27689 );
and ( n10383 , n10382 , RI17470350_1189);
and ( n10384 , n28495 , n27689 );
or ( n28496 , n10383 , n10384 );
xor ( n28497 , RI19acb828_2243 , RI174b9460_834);
not ( n10385 , n27689 );
and ( n10386 , n10385 , RI174b9460_834);
and ( n10387 , n28497 , n27689 );
or ( n28498 , n10386 , n10387 );
xor ( n28499 , n28496 , n28498 );
buf ( n28500 , RI1738b378_2077);
xor ( n28501 , n28499 , n28500 );
buf ( n28502 , RI173d4068_1722);
xor ( n28503 , n28501 , n28502 );
buf ( n28504 , RI1744bb40_1367);
xor ( n28505 , n28503 , n28504 );
xor ( n28506 , n28494 , n28505 );
not ( n28507 , n28506 );
buf ( n28508 , RI173dd410_1677);
xor ( n28509 , RI19a8c498_2709 , RI1746b148_1214);
not ( n10388 , n27689 );
and ( n10389 , n10388 , RI1746b148_1214);
and ( n10390 , n28509 , n27689 );
or ( n28510 , n10389 , n10390 );
xor ( n28511 , RI19abd890_2354 , RI174b3e20_859);
not ( n10391 , n27689 );
and ( n10392 , n10391 , RI174b3e20_859);
and ( n10393 , n28511 , n27689 );
or ( n28512 , n10392 , n10393 );
xor ( n28513 , n28510 , n28512 );
buf ( n28514 , RI17345580_2103);
xor ( n28515 , n28513 , n28514 );
buf ( n28516 , RI173cee48_1747);
xor ( n28517 , n28515 , n28516 );
buf ( n28518 , RI17446938_1392);
xor ( n28519 , n28517 , n28518 );
xor ( n28520 , n28508 , n28519 );
xor ( n28521 , n28520 , n28304 );
and ( n28522 , n28507 , n28521 );
xor ( n28523 , n28482 , n28522 );
xor ( n28524 , RI19ab1ef0_2440 , RI174a9a10_909);
not ( n10394 , n27689 );
and ( n10395 , n10394 , RI174a9a10_909);
and ( n10396 , n28524 , n27689 );
or ( n28525 , n10395 , n10396 );
buf ( n28526 , RI1733b170_2153);
xor ( n28527 , n28525 , n28526 );
buf ( n28528 , RI173c46f0_1798);
xor ( n28529 , n28527 , n28528 );
buf ( n28530 , RI1740d3e0_1443);
xor ( n28531 , n28529 , n28530 );
buf ( n28532 , RI175361d0_598);
xor ( n28533 , n28531 , n28532 );
xor ( n28534 , n27717 , n28533 );
xor ( n28535 , RI19a9bfd8_2598 , RI1746f978_1192);
not ( n10397 , n27689 );
and ( n10398 , n10397 , RI1746f978_1192);
and ( n10399 , n28535 , n27689 );
or ( n28536 , n10398 , n10399 );
xor ( n28537 , n28536 , n28114 );
buf ( n28538 , RI1738a9a0_2080);
xor ( n28539 , n28537 , n28538 );
buf ( n28540 , RI173d3690_1725);
xor ( n28541 , n28539 , n28540 );
buf ( n28542 , RI1744b168_1370);
xor ( n28543 , n28541 , n28542 );
xor ( n28544 , n28534 , n28543 );
xor ( n28545 , RI19ac6080_2284 , RI174c7c68_789);
not ( n10400 , n27689 );
and ( n10401 , n10400 , RI174c7c68_789);
and ( n10402 , n28545 , n27689 );
or ( n28546 , n10401 , n10402 );
xor ( n28547 , RI19a8c240_2710 , RI1746ae00_1215);
not ( n10403 , n27689 );
and ( n10404 , n10403 , RI1746ae00_1215);
and ( n10405 , n28547 , n27689 );
or ( n28548 , n10404 , n10405 );
xor ( n28549 , RI19abd6b0_2355 , RI174b3ad8_860);
not ( n10406 , n27689 );
and ( n10407 , n10406 , RI174b3ad8_860);
and ( n10408 , n28549 , n27689 );
or ( n28550 , n10407 , n10408 );
xor ( n28551 , n28548 , n28550 );
buf ( n28552 , RI17345238_2104);
xor ( n28553 , n28551 , n28552 );
buf ( n28554 , RI173ceb00_1748);
xor ( n28555 , n28553 , n28554 );
buf ( n28556 , RI174465f0_1393);
xor ( n28557 , n28555 , n28556 );
xor ( n28558 , n28546 , n28557 );
xor ( n28559 , RI19aa0358_2567 , RI17488338_1072);
not ( n10409 , n27689 );
and ( n10410 , n10409 , RI17488338_1072);
and ( n10411 , n28559 , n27689 );
or ( n28560 , n10410 , n10411 );
xor ( n28561 , RI19acef78_2218 , RI1750fc38_717);
not ( n10412 , n27689 );
and ( n10413 , n10412 , RI1750fc38_717);
and ( n10414 , n28561 , n27689 );
or ( n28562 , n10413 , n10414 );
xor ( n28563 , n28560 , n28562 );
buf ( n28564 , RI173a3360_1960);
xor ( n28565 , n28563 , n28564 );
buf ( n28566 , RI173ec050_1605);
xor ( n28567 , n28565 , n28566 );
buf ( n28568 , RI1747c4e8_1130);
xor ( n28569 , n28567 , n28568 );
xor ( n28570 , n28558 , n28569 );
not ( n28571 , n28570 );
buf ( n28572 , RI173a2cd0_1962);
xor ( n28573 , RI19a96038_2640 , RI174793b0_1145);
not ( n10415 , n27689 );
and ( n10416 , n10415 , RI174793b0_1145);
and ( n10417 , n28573 , n27689 );
or ( n28574 , n10416 , n10417 );
xor ( n28575 , RI19ac5e28_2285 , RI174c7740_790);
not ( n10418 , n27689 );
and ( n10419 , n10418 , RI174c7740_790);
and ( n10420 , n28575 , n27689 );
or ( n28576 , n10419 , n10420 );
xor ( n28577 , n28574 , n28576 );
buf ( n28578 , RI17394090_2034);
xor ( n28579 , n28577 , n28578 );
buf ( n28580 , RI173dcd80_1679);
xor ( n28581 , n28579 , n28580 );
buf ( n28582 , RI17454858_1324);
xor ( n28583 , n28581 , n28582 );
xor ( n28584 , n28572 , n28583 );
xor ( n28585 , RI19aa9d90_2497 , RI174968e8_1002);
not ( n10421 , n27689 );
and ( n10422 , n10421 , RI174968e8_1002);
and ( n10423 , n28585 , n27689 );
or ( n28586 , n10422 , n10423 );
xor ( n28587 , RI19a9cc08_2592 , RI17526528_647);
not ( n10424 , n27689 );
and ( n10425 , n10424 , RI17526528_647);
and ( n10426 , n28587 , n27689 );
or ( n28588 , n10425 , n10426 );
xor ( n28589 , n28586 , n28588 );
buf ( n28590 , RI173b15c8_1891);
xor ( n28591 , n28589 , n28590 );
buf ( n28592 , RI173fa2b8_1536);
xor ( n28593 , n28591 , n28592 );
buf ( n28594 , RI17394db0_2030);
xor ( n28595 , n28593 , n28594 );
xor ( n28596 , n28584 , n28595 );
and ( n28597 , n28571 , n28596 );
xor ( n28598 , n28544 , n28597 );
or ( n28599 , n27689 , RI17539830_589);
or ( n28600 , n28599 , RI17539218_590);
or ( n28601 , n28600 , RI175385e8_592);
or ( n28602 , n28601 , RI17537fd0_593);
or ( n28603 , n28602 , RI175379b8_594);
or ( n28604 , n28603 , RI17536770_597);
or ( n28605 , n28604 , RI17539e48_588);
xor ( n28606 , n28598 , n28605 );
xor ( n28607 , RI19aa2248_2551 , RI174844e0_1091);
not ( n10427 , n27689 );
and ( n10428 , n10427 , RI174844e0_1091);
and ( n10429 , n28607 , n27689 );
or ( n28608 , n10428 , n10429 );
xor ( n28609 , RI19a83438_2771 , RI17509a40_736);
not ( n10430 , n27689 );
and ( n10431 , n10430 , RI17509a40_736);
and ( n10432 , n28609 , n27689 );
or ( n28610 , n10431 , n10432 );
xor ( n28611 , n28608 , n28610 );
buf ( n28612 , RI1739f1c0_1980);
xor ( n28613 , n28611 , n28612 );
buf ( n28614 , RI173e81f8_1624);
xor ( n28615 , n28613 , n28614 );
buf ( n28616 , RI1745fcd0_1269);
xor ( n28617 , n28615 , n28616 );
xor ( n28618 , n28282 , n28617 );
xor ( n28619 , RI19ab63d8_2407 , RI174a1a18_948);
not ( n10433 , n27689 );
and ( n10434 , n10433 , RI174a1a18_948);
and ( n10435 , n28619 , n27689 );
or ( n28620 , n10434 , n10435 );
buf ( n28621 , RI173334c0_2191);
xor ( n28622 , n28620 , n28621 );
buf ( n28623 , RI173bca40_1836);
xor ( n28624 , n28622 , n28623 );
xor ( n28625 , n28624 , n28316 );
buf ( n28626 , RI174046c8_1486);
xor ( n28627 , n28625 , n28626 );
xor ( n28628 , n28618 , n28627 );
not ( n28629 , n28482 );
and ( n28630 , n28629 , n28506 );
xor ( n28631 , n28628 , n28630 );
xor ( n28632 , n28606 , n28631 );
xor ( n28633 , n28536 , n28125 );
xor ( n28634 , n28633 , n28137 );
xor ( n28635 , RI19a876c8_2742 , RI174d1208_760);
not ( n10436 , n27689 );
and ( n10437 , n10436 , RI174d1208_760);
and ( n10438 , n28635 , n27689 );
or ( n28636 , n10437 , n10438 );
xor ( n28637 , RI19a9ca28_2593 , RI174709e0_1187);
not ( n10439 , n27689 );
and ( n10440 , n10439 , RI174709e0_1187);
and ( n10441 , n28637 , n27689 );
or ( n28638 , n10440 , n10441 );
xor ( n28639 , RI19acbc60_2241 , RI174b9eb0_832);
not ( n10442 , n27689 );
and ( n10443 , n10442 , RI174b9eb0_832);
and ( n10444 , n28639 , n27689 );
or ( n28640 , n10443 , n10444 );
xor ( n28641 , n28638 , n28640 );
buf ( n28642 , RI1738ba08_2075);
xor ( n28643 , n28641 , n28642 );
buf ( n28644 , RI173d46f8_1720);
xor ( n28645 , n28643 , n28644 );
buf ( n28646 , RI1744c1d0_1365);
xor ( n28647 , n28645 , n28646 );
xor ( n28648 , n28636 , n28647 );
xor ( n28649 , RI19ab0870_2450 , RI1748df18_1044);
not ( n10445 , n27689 );
and ( n10446 , n10445 , RI1748df18_1044);
and ( n10447 , n28649 , n27689 );
or ( n28650 , n10446 , n10447 );
xor ( n28651 , RI19ac1d78_2315 , RI175191c0_688);
not ( n10448 , n27689 );
and ( n10449 , n10448 , RI175191c0_688);
and ( n10450 , n28651 , n27689 );
or ( n28652 , n10449 , n10450 );
xor ( n28653 , n28650 , n28652 );
buf ( n28654 , RI173a8f40_1932);
xor ( n28655 , n28653 , n28654 );
buf ( n28656 , RI173f1c30_1577);
xor ( n28657 , n28655 , n28656 );
buf ( n28658 , RI174b75e8_842);
xor ( n28659 , n28657 , n28658 );
xor ( n28660 , n28648 , n28659 );
not ( n28661 , n28660 );
buf ( n28662 , RI173ad0e0_1912);
xor ( n28663 , RI19aa1d20_2554 , RI17483b08_1094);
not ( n10451 , n27689 );
and ( n10452 , n10451 , RI17483b08_1094);
and ( n10453 , n28663 , n27689 );
or ( n28664 , n10452 , n10453 );
xor ( n28665 , RI19a82d30_2774 , RI17508ac8_739);
not ( n10454 , n27689 );
and ( n10455 , n10454 , RI17508ac8_739);
and ( n10456 , n28665 , n27689 );
or ( n28666 , n10455 , n10456 );
xor ( n28667 , n28664 , n28666 );
buf ( n28668 , RI1739e7e8_1983);
xor ( n28669 , n28667 , n28668 );
buf ( n28670 , RI173e7820_1627);
xor ( n28671 , n28669 , n28670 );
buf ( n28672 , RI1745f2f8_1272);
xor ( n28673 , n28671 , n28672 );
xor ( n28674 , n28662 , n28673 );
xor ( n28675 , RI19ab5d48_2410 , RI174a1040_951);
not ( n10457 , n27689 );
and ( n10458 , n10457 , RI174a1040_951);
and ( n10459 , n28675 , n27689 );
or ( n28676 , n10458 , n10459 );
buf ( n28677 , RI17332ae8_2194);
xor ( n28678 , n28676 , n28677 );
buf ( n28679 , RI173bc068_1839);
xor ( n28680 , n28678 , n28679 );
buf ( n28681 , RI17404d58_1484);
xor ( n28682 , n28680 , n28681 );
buf ( n28683 , RI173fda80_1519);
xor ( n28684 , n28682 , n28683 );
xor ( n28685 , n28674 , n28684 );
and ( n28686 , n28661 , n28685 );
xor ( n28687 , n28634 , n28686 );
xor ( n28688 , n28632 , n28687 );
xor ( n28689 , RI19ab5f28_2409 , RI174a1388_950);
not ( n10460 , n27689 );
and ( n10461 , n10460 , RI174a1388_950);
and ( n10462 , n28689 , n27689 );
or ( n28690 , n10461 , n10462 );
xor ( n28691 , n28690 , n27948 );
xor ( n28692 , RI19a8e8b0_2693 , RI174672f0_1233);
not ( n10463 , n27689 );
and ( n10464 , n10463 , RI174672f0_1233);
and ( n10465 , n28692 , n27689 );
or ( n28693 , n10464 , n10465 );
xor ( n28694 , RI19abf4b0_2338 , RI174affc8_878);
not ( n10466 , n27689 );
and ( n10467 , n10466 , RI174affc8_878);
and ( n10468 , n28694 , n27689 );
or ( n28695 , n10467 , n10468 );
xor ( n28696 , n28693 , n28695 );
buf ( n28697 , RI17341728_2122);
xor ( n28698 , n28696 , n28697 );
buf ( n28699 , RI173caca8_1767);
xor ( n28700 , n28698 , n28699 );
buf ( n28701 , RI17413ce0_1411);
xor ( n28702 , n28700 , n28701 );
xor ( n28703 , n28691 , n28702 );
xor ( n28704 , RI19abe6a0_2346 , RI174b1d50_869);
not ( n10469 , n27689 );
and ( n10470 , n10469 , RI174b1d50_869);
and ( n10471 , n28704 , n27689 );
or ( n28705 , n10470 , n10471 );
xor ( n28706 , RI19ab4dd0_2417 , RI174a3458_940);
not ( n10472 , n27689 );
and ( n10473 , n10472 , RI174a3458_940);
and ( n10474 , n28706 , n27689 );
or ( n28707 , n10473 , n10474 );
buf ( n28708 , RI17334f00_2183);
xor ( n28709 , n28707 , n28708 );
buf ( n28710 , RI173be480_1828);
xor ( n28711 , n28709 , n28710 );
buf ( n28712 , RI17407170_1473);
xor ( n28713 , n28711 , n28712 );
buf ( n28714 , RI174146b8_1408);
xor ( n28715 , n28713 , n28714 );
xor ( n28716 , n28705 , n28715 );
xor ( n28717 , RI19a97820_2629 , RI17478000_1151);
not ( n10475 , n27689 );
and ( n10476 , n10475 , RI17478000_1151);
and ( n10477 , n28717 , n27689 );
or ( n28718 , n10476 , n10477 );
xor ( n28719 , RI19ac7700_2274 , RI174c5850_796);
not ( n10478 , n27689 );
and ( n10479 , n10478 , RI174c5850_796);
and ( n10480 , n28719 , n27689 );
or ( n28720 , n10479 , n10480 );
xor ( n28721 , n28718 , n28720 );
buf ( n28722 , RI17392ce0_2040);
xor ( n28723 , n28721 , n28722 );
buf ( n28724 , RI173db9d0_1685);
xor ( n28725 , n28723 , n28724 );
buf ( n28726 , RI174534a8_1330);
xor ( n28727 , n28725 , n28726 );
xor ( n28728 , n28716 , n28727 );
not ( n28729 , n28728 );
buf ( n28730 , RI1738ca70_2070);
xor ( n28731 , RI19a90cc8_2677 , RI17463150_1253);
not ( n10481 , n27689 );
and ( n10482 , n10481 , RI17463150_1253);
and ( n10483 , n28731 , n27689 );
or ( n28732 , n10482 , n10483 );
xor ( n28733 , RI19ac1148_2322 , RI174abe28_898);
not ( n10484 , n27689 );
and ( n10485 , n10484 , RI174abe28_898);
and ( n10486 , n28733 , n27689 );
or ( n28734 , n10485 , n10486 );
xor ( n28735 , n28732 , n28734 );
buf ( n28736 , RI1733d588_2142);
xor ( n28737 , n28735 , n28736 );
buf ( n28738 , RI173c6b08_1787);
xor ( n28739 , n28737 , n28738 );
buf ( n28740 , RI1740f7f8_1432);
xor ( n28741 , n28739 , n28740 );
xor ( n28742 , n28730 , n28741 );
xor ( n28743 , n28742 , n28096 );
and ( n28744 , n28729 , n28743 );
xor ( n28745 , n28703 , n28744 );
xor ( n28746 , n28688 , n28745 );
xor ( n28747 , RI19a9e030_2584 , RI1748be48_1054);
not ( n10487 , n27689 );
and ( n10488 , n10487 , RI1748be48_1054);
and ( n10489 , n28747 , n27689 );
or ( n28748 , n10488 , n10489 );
xor ( n28749 , RI19a93d88_2655 , RI1747d898_1124);
not ( n10490 , n27689 );
and ( n10491 , n10490 , RI1747d898_1124);
and ( n10492 , n28749 , n27689 );
or ( n28750 , n10491 , n10492 );
xor ( n28751 , RI19ac40a0_2299 , RI174ce388_769);
not ( n10493 , n27689 );
and ( n10494 , n10493 , RI174ce388_769);
and ( n10495 , n28751 , n27689 );
or ( n28752 , n10494 , n10495 );
xor ( n28753 , n28750 , n28752 );
buf ( n28754 , RI17398578_2013);
xor ( n28755 , n28753 , n28754 );
buf ( n28756 , RI173e1268_1658);
xor ( n28757 , n28755 , n28756 );
buf ( n28758 , RI17459088_1302);
xor ( n28759 , n28757 , n28758 );
xor ( n28760 , n28748 , n28759 );
xor ( n28761 , RI19aa7c48_2511 , RI1749add0_981);
not ( n10496 , n27689 );
and ( n10497 , n10496 , RI1749add0_981);
and ( n10498 , n28761 , n27689 );
or ( n28762 , n10497 , n10498 );
xor ( n28763 , RI19a88e38_2732 , RI1752d170_626);
not ( n10499 , n27689 );
and ( n10500 , n10499 , RI1752d170_626);
and ( n10501 , n28763 , n27689 );
or ( n28764 , n10500 , n10501 );
xor ( n28765 , n28762 , n28764 );
buf ( n28766 , RI173b5ab0_1870);
xor ( n28767 , n28765 , n28766 );
buf ( n28768 , RI173feae8_1514);
xor ( n28769 , n28767 , n28768 );
buf ( n28770 , RI173c0208_1819);
xor ( n28771 , n28769 , n28770 );
xor ( n28772 , n28760 , n28771 );
xor ( n28773 , RI19a95048_2647 , RI1752a308_635);
not ( n10502 , n27689 );
and ( n10503 , n10502 , RI1752a308_635);
and ( n10504 , n28773 , n27689 );
or ( n28774 , n10503 , n10504 );
xor ( n28775 , RI19a9f548_2574 , RI1748a750_1061);
not ( n10505 , n27689 );
and ( n10506 , n10505 , RI1748a750_1061);
and ( n10507 , n28775 , n27689 );
or ( n28776 , n10506 , n10507 );
xor ( n28777 , RI19ace168_2224 , RI17513a18_705);
not ( n10508 , n27689 );
and ( n10509 , n10508 , RI17513a18_705);
and ( n10510 , n28777 , n27689 );
or ( n28778 , n10509 , n10510 );
xor ( n28779 , n28776 , n28778 );
buf ( n28780 , RI173a5778_1949);
xor ( n28781 , n28779 , n28780 );
buf ( n28782 , RI173ee468_1594);
xor ( n28783 , n28781 , n28782 );
buf ( n28784 , RI17493120_1019);
xor ( n28785 , n28783 , n28784 );
xor ( n28786 , n28774 , n28785 );
xor ( n28787 , n28786 , n28015 );
not ( n28788 , n28787 );
buf ( n28789 , RI173bee58_1825);
xor ( n28790 , RI19aab938_2485 , RI17495880_1007);
not ( n10511 , n27689 );
and ( n10512 , n10511 , RI17495880_1007);
and ( n10513 , n28790 , n27689 );
or ( n28791 , n10512 , n10513 );
xor ( n28792 , RI19aadb70_2470 , RI17524b60_652);
not ( n10514 , n27689 );
and ( n10515 , n10514 , RI17524b60_652);
and ( n10516 , n28792 , n27689 );
or ( n28793 , n10515 , n10516 );
xor ( n28794 , n28791 , n28793 );
buf ( n28795 , RI173b0560_1896);
xor ( n28796 , n28794 , n28795 );
buf ( n28797 , RI173f9250_1541);
xor ( n28798 , n28796 , n28797 );
buf ( n28799 , RI17389938_2085);
xor ( n28800 , n28798 , n28799 );
xor ( n28801 , n28789 , n28800 );
xor ( n28802 , RI19a8dfc8_2697 , RI17469d98_1220);
not ( n10517 , n27689 );
and ( n10518 , n10517 , RI17469d98_1220);
and ( n10519 , n28802 , n27689 );
or ( n28803 , n10518 , n10519 );
xor ( n28804 , RI19abeda8_2342 , RI174b2a70_865);
not ( n10520 , n27689 );
and ( n10521 , n10520 , RI174b2a70_865);
and ( n10522 , n28804 , n27689 );
or ( n28805 , n10521 , n10522 );
xor ( n28806 , n28803 , n28805 );
buf ( n28807 , RI173441d0_2109);
xor ( n28808 , n28806 , n28807 );
buf ( n28809 , RI173cd750_1754);
xor ( n28810 , n28808 , n28809 );
buf ( n28811 , RI17445588_1398);
xor ( n28812 , n28810 , n28811 );
xor ( n28813 , n28801 , n28812 );
and ( n28814 , n28788 , n28813 );
xor ( n28815 , n28772 , n28814 );
xor ( n28816 , n28746 , n28815 );
xor ( n28817 , n28523 , n28816 );
buf ( n28818 , RI173a3018_1961);
xor ( n28819 , RI19a96290_2639 , RI174796f8_1144);
not ( n10523 , n27689 );
and ( n10524 , n10523 , RI174796f8_1144);
and ( n10525 , n28819 , n27689 );
or ( n28820 , n10524 , n10525 );
xor ( n28821 , n28820 , n28546 );
buf ( n28822 , RI173943d8_2033);
xor ( n28823 , n28821 , n28822 );
buf ( n28824 , RI173dd0c8_1678);
xor ( n28825 , n28823 , n28824 );
buf ( n28826 , RI17454ba0_1323);
xor ( n28827 , n28825 , n28826 );
xor ( n28828 , n28818 , n28827 );
xor ( n28829 , RI19aa9f70_2496 , RI17496c30_1001);
not ( n10526 , n27689 );
and ( n10527 , n10526 , RI17496c30_1001);
and ( n10528 , n28829 , n27689 );
or ( n28830 , n10527 , n10528 );
xor ( n28831 , RI19a9e6c0_2581 , RI17526a50_646);
not ( n10529 , n27689 );
and ( n10530 , n10529 , RI17526a50_646);
and ( n10531 , n28831 , n27689 );
or ( n28832 , n10530 , n10531 );
xor ( n28833 , n28830 , n28832 );
buf ( n28834 , RI173b1910_1890);
xor ( n28835 , n28833 , n28834 );
buf ( n28836 , RI173fa600_1535);
xor ( n28837 , n28835 , n28836 );
buf ( n28838 , RI173971c8_2019);
xor ( n28839 , n28837 , n28838 );
xor ( n28840 , n28828 , n28839 );
buf ( n28841 , RI173f53f8_1560);
xor ( n28842 , n28841 , n27921 );
xor ( n28843 , RI19ab7da0_2396 , RI174a0320_955);
not ( n10532 , n27689 );
and ( n10533 , n10532 , RI174a0320_955);
and ( n10534 , n28843 , n27689 );
or ( n28844 , n10533 , n10534 );
buf ( n28845 , RI17535780_600);
xor ( n28846 , n28844 , n28845 );
buf ( n28847 , RI173bb348_1843);
xor ( n28848 , n28846 , n28847 );
buf ( n28849 , RI17404038_1488);
xor ( n28850 , n28848 , n28849 );
buf ( n28851 , RI173f6af0_1553);
xor ( n28852 , n28850 , n28851 );
xor ( n28853 , n28842 , n28852 );
not ( n28854 , n28853 );
buf ( n28855 , RI173e4a30_1641);
xor ( n28856 , RI19aaf628_2458 , RI1748ffe8_1034);
not ( n10535 , n27689 );
and ( n10536 , n10535 , RI1748ffe8_1034);
and ( n10537 , n28856 , n27689 );
or ( n28857 , n10536 , n10537 );
xor ( n28858 , RI19a23150_2796 , RI1751c028_679);
not ( n10538 , n27689 );
and ( n10539 , n10538 , RI1751c028_679);
and ( n10540 , n28858 , n27689 );
or ( n28859 , n10539 , n10540 );
xor ( n28860 , n28857 , n28859 );
buf ( n28861 , RI173aacc8_1923);
xor ( n28862 , n28860 , n28861 );
buf ( n28863 , RI173f39b8_1568);
xor ( n28864 , n28862 , n28863 );
buf ( n28865 , RI17502420_753);
xor ( n28866 , n28864 , n28865 );
xor ( n28867 , n28855 , n28866 );
xor ( n28868 , RI19a919e8_2671 , RI17464848_1246);
not ( n10541 , n27689 );
and ( n10542 , n10541 , RI17464848_1246);
and ( n10543 , n28868 , n27689 );
or ( n28869 , n10542 , n10543 );
xor ( n28870 , RI19ac1b98_2316 , RI174ad520_891);
not ( n10544 , n27689 );
and ( n10545 , n10544 , RI174ad520_891);
and ( n10546 , n28870 , n27689 );
or ( n28871 , n10545 , n10546 );
xor ( n28872 , n28869 , n28871 );
buf ( n28873 , RI1733ec80_2135);
xor ( n28874 , n28872 , n28873 );
buf ( n28875 , RI173c8200_1780);
xor ( n28876 , n28874 , n28875 );
buf ( n28877 , RI17410ef0_1425);
xor ( n28878 , n28876 , n28877 );
xor ( n28879 , n28867 , n28878 );
and ( n28880 , n28854 , n28879 );
xor ( n28881 , n28840 , n28880 );
buf ( n28882 , RI1733c1d8_2148);
xor ( n28883 , RI19ab9c18_2382 , RI1749be38_976);
not ( n10547 , n27689 );
and ( n10548 , n10547 , RI1749be38_976);
and ( n10549 , n28883 , n27689 );
or ( n28884 , n10548 , n10549 );
buf ( n28885 , RI1752eb38_621);
xor ( n28886 , n28884 , n28885 );
buf ( n28887 , RI173b6b18_1865);
xor ( n28888 , n28886 , n28887 );
buf ( n28889 , RI173ffb50_1509);
xor ( n28890 , n28888 , n28889 );
buf ( n28891 , RI173cb680_1764);
xor ( n28892 , n28890 , n28891 );
xor ( n28893 , n28882 , n28892 );
xor ( n28894 , RI19a9c848_2594 , RI17470698_1188);
not ( n10550 , n27689 );
and ( n10551 , n10550 , RI17470698_1188);
and ( n10552 , n28894 , n27689 );
or ( n28895 , n10551 , n10552 );
xor ( n28896 , RI19acba08_2242 , RI174b9988_833);
not ( n10553 , n27689 );
and ( n10554 , n10553 , RI174b9988_833);
and ( n10555 , n28896 , n27689 );
or ( n28897 , n10554 , n10555 );
xor ( n28898 , n28895 , n28897 );
buf ( n28899 , RI1738b6c0_2076);
xor ( n28900 , n28898 , n28899 );
buf ( n28901 , RI173d43b0_1721);
xor ( n28902 , n28900 , n28901 );
buf ( n28903 , RI1744be88_1366);
xor ( n28904 , n28902 , n28903 );
xor ( n28905 , n28893 , n28904 );
buf ( n28906 , RI173dd758_1676);
xor ( n28907 , RI19a8c6f0_2708 , RI1746b490_1213);
not ( n10556 , n27689 );
and ( n10557 , n10556 , RI1746b490_1213);
and ( n10558 , n28907 , n27689 );
or ( n28908 , n10557 , n10558 );
xor ( n28909 , RI19abd9f8_2353 , RI174b4168_858);
not ( n10559 , n27689 );
and ( n10560 , n10559 , RI174b4168_858);
and ( n10561 , n28909 , n27689 );
or ( n28910 , n10560 , n10561 );
xor ( n28911 , n28908 , n28910 );
buf ( n28912 , RI173458c8_2102);
xor ( n28913 , n28911 , n28912 );
buf ( n28914 , RI173cf190_1746);
xor ( n28915 , n28913 , n28914 );
buf ( n28916 , RI17446c80_1391);
xor ( n28917 , n28915 , n28916 );
xor ( n28918 , n28906 , n28917 );
xor ( n28919 , RI19aa0790_2565 , RI174889c8_1070);
not ( n10562 , n27689 );
and ( n10563 , n10562 , RI174889c8_1070);
and ( n10564 , n28919 , n27689 );
or ( n28920 , n10563 , n10564 );
xor ( n28921 , RI19acf428_2216 , RI17510688_715);
not ( n10565 , n27689 );
and ( n10566 , n10565 , RI17510688_715);
and ( n10567 , n28921 , n27689 );
or ( n28922 , n10566 , n10567 );
xor ( n28923 , n28920 , n28922 );
buf ( n28924 , RI173a39f0_1958);
xor ( n28925 , n28923 , n28924 );
buf ( n28926 , RI173ec6e0_1603);
xor ( n28927 , n28925 , n28926 );
buf ( n28928 , RI17480d18_1108);
xor ( n28929 , n28927 , n28928 );
xor ( n28930 , n28918 , n28929 );
not ( n28931 , n28930 );
buf ( n28932 , RI174a2dc8_942);
xor ( n28933 , n28932 , n28759 );
xor ( n28934 , n28933 , n28771 );
and ( n28935 , n28931 , n28934 );
xor ( n28936 , n28905 , n28935 );
xor ( n28937 , n28881 , n28936 );
buf ( n28938 , RI173ad428_1911);
xor ( n28939 , RI19aa1f00_2553 , RI17483e50_1093);
not ( n10568 , n27689 );
and ( n10569 , n10568 , RI17483e50_1093);
and ( n10570 , n28939 , n27689 );
or ( n28940 , n10569 , n10570 );
xor ( n28941 , n28940 , n27925 );
buf ( n28942 , RI1739eb30_1982);
xor ( n28943 , n28941 , n28942 );
buf ( n28944 , RI173e7b68_1626);
xor ( n28945 , n28943 , n28944 );
buf ( n28946 , RI1745f640_1271);
xor ( n28947 , n28945 , n28946 );
xor ( n28948 , n28938 , n28947 );
buf ( n28949 , RI17332e30_2193);
xor ( n28950 , n28690 , n28949 );
buf ( n28951 , RI173bc3b0_1838);
xor ( n28952 , n28950 , n28951 );
buf ( n28953 , RI174050a0_1483);
xor ( n28954 , n28952 , n28953 );
buf ( n28955 , RI173ffe98_1508);
xor ( n28956 , n28954 , n28955 );
xor ( n28957 , n28948 , n28956 );
buf ( n28958 , RI17400f00_1503);
xor ( n28959 , RI19aae7a0_2465 , RI1748ec38_1040);
not ( n10571 , n27689 );
and ( n10572 , n10571 , RI1748ec38_1040);
and ( n10573 , n28959 , n27689 );
or ( n28960 , n10572 , n10573 );
xor ( n28961 , RI19a23330_2795 , RI1751a138_685);
not ( n10574 , n27689 );
and ( n10575 , n10574 , RI1751a138_685);
and ( n10576 , n28961 , n27689 );
or ( n28962 , n10575 , n10576 );
xor ( n28963 , n28960 , n28962 );
buf ( n28964 , RI173a9918_1929);
xor ( n28965 , n28963 , n28964 );
buf ( n28966 , RI173f2608_1574);
xor ( n28967 , n28965 , n28966 );
buf ( n28968 , RI174be1b8_819);
xor ( n28969 , n28967 , n28968 );
xor ( n28970 , n28958 , n28969 );
xor ( n28971 , n28970 , n28741 );
not ( n28972 , n28971 );
buf ( n28973 , RI174118c8_1422);
xor ( n28974 , RI19ab73c8_2400 , RI1749f600_959);
not ( n10577 , n27689 );
and ( n10578 , n10577 , RI1749f600_959);
and ( n10579 , n28974 , n27689 );
or ( n28975 , n10578 , n10579 );
buf ( n28976 , RI175342e0_604);
xor ( n28977 , n28975 , n28976 );
buf ( n28978 , RI173ba628_1847);
xor ( n28979 , n28977 , n28978 );
buf ( n28980 , RI17403318_1492);
xor ( n28981 , n28979 , n28980 );
buf ( n28982 , RI173eda90_1597);
xor ( n28983 , n28981 , n28982 );
xor ( n28984 , n28973 , n28983 );
xor ( n28985 , RI19a99f80_2612 , RI17473e60_1171);
not ( n10580 , n27689 );
and ( n10581 , n10580 , RI17473e60_1171);
and ( n10582 , n28985 , n27689 );
or ( n28986 , n10581 , n10582 );
xor ( n28987 , RI19ac96e0_2259 , RI174bf658_815);
not ( n10583 , n27689 );
and ( n10584 , n10583 , RI174bf658_815);
and ( n10585 , n28987 , n27689 );
or ( n28988 , n10584 , n10585 );
xor ( n28989 , n28986 , n28988 );
buf ( n28990 , RI1738ee88_2059);
xor ( n28991 , n28989 , n28990 );
buf ( n28992 , RI173d7b78_1704);
xor ( n28993 , n28991 , n28992 );
buf ( n28994 , RI1744f650_1349);
xor ( n28995 , n28993 , n28994 );
xor ( n28996 , n28984 , n28995 );
and ( n28997 , n28972 , n28996 );
xor ( n28998 , n28957 , n28997 );
xor ( n28999 , n28937 , n28998 );
buf ( n29000 , RI1738cdb8_2069);
xor ( n29001 , RI19a90f20_2676 , RI174637e0_1251);
not ( n10586 , n27689 );
and ( n10587 , n10586 , RI174637e0_1251);
and ( n10588 , n29001 , n27689 );
or ( n29002 , n10587 , n10588 );
xor ( n29003 , RI19ac12b0_2321 , RI174ac4b8_896);
not ( n10589 , n27689 );
and ( n10590 , n10589 , RI174ac4b8_896);
and ( n10591 , n29003 , n27689 );
or ( n29004 , n10590 , n10591 );
xor ( n29005 , n29002 , n29004 );
buf ( n29006 , RI1733dc18_2140);
xor ( n29007 , n29005 , n29006 );
buf ( n29008 , RI173c7198_1785);
xor ( n29009 , n29007 , n29008 );
buf ( n29010 , RI1740fe88_1430);
xor ( n29011 , n29009 , n29010 );
xor ( n29012 , n29000 , n29011 );
xor ( n29013 , n29012 , n27964 );
buf ( n29014 , RI173e5750_1637);
xor ( n29015 , RI19a9bd80_2599 , RI17472df8_1176);
not ( n10592 , n27689 );
and ( n10593 , n10592 , RI17472df8_1176);
and ( n10594 , n29015 , n27689 );
or ( n29016 , n10593 , n10594 );
xor ( n29017 , RI19acb120_2247 , RI174bd768_821);
not ( n10595 , n27689 );
and ( n10596 , n10595 , RI174bd768_821);
and ( n10597 , n29017 , n27689 );
or ( n29018 , n10596 , n10597 );
xor ( n29019 , n29016 , n29018 );
buf ( n29020 , RI1738de20_2064);
xor ( n29021 , n29019 , n29020 );
buf ( n29022 , RI173d6b10_1709);
xor ( n29023 , n29021 , n29022 );
buf ( n29024 , RI1744e5e8_1354);
xor ( n29025 , n29023 , n29024 );
xor ( n29026 , n29014 , n29025 );
xor ( n29027 , RI19aad300_2474 , RI17490678_1032);
not ( n10598 , n27689 );
and ( n10599 , n10598 , RI17490678_1032);
and ( n10600 , n29027 , n27689 );
or ( n29028 , n10599 , n10600 );
xor ( n29029 , RI19abcfa8_2359 , RI1751ca78_677);
not ( n10601 , n27689 );
and ( n10602 , n10601 , RI1751ca78_677);
and ( n10603 , n29029 , n27689 );
or ( n29030 , n10602 , n10603 );
xor ( n29031 , n29028 , n29030 );
buf ( n29032 , RI173ab358_1921);
xor ( n29033 , n29031 , n29032 );
buf ( n29034 , RI173f4048_1566);
xor ( n29035 , n29033 , n29034 );
buf ( n29036 , RI1750b408_731);
xor ( n29037 , n29035 , n29036 );
xor ( n29038 , n29026 , n29037 );
not ( n29039 , n29038 );
buf ( n29040 , RI173b2630_1886);
xor ( n29041 , RI19a9d400_2589 , RI1748ade0_1059);
not ( n10604 , n27689 );
and ( n10605 , n10604 , RI1748ade0_1059);
and ( n10606 , n29041 , n27689 );
or ( n29042 , n10605 , n10606 );
xor ( n29043 , RI19acc200_2238 , RI17514468_703);
not ( n10607 , n27689 );
and ( n10608 , n10607 , RI17514468_703);
and ( n10609 , n29043 , n27689 );
or ( n29044 , n10608 , n10609 );
xor ( n29045 , n29042 , n29044 );
buf ( n29046 , RI173a5e08_1947);
xor ( n29047 , n29045 , n29046 );
buf ( n29048 , RI173eeaf8_1592);
xor ( n29049 , n29047 , n29048 );
buf ( n29050 , RI17497950_997);
xor ( n29051 , n29049 , n29050 );
xor ( n29052 , n29040 , n29051 );
xor ( n29053 , RI19ab0ff0_2446 , RI174a8660_915);
not ( n10610 , n27689 );
and ( n10611 , n10610 , RI174a8660_915);
and ( n10612 , n29053 , n27689 );
or ( n29054 , n10611 , n10612 );
buf ( n29055 , RI17339dc0_2159);
xor ( n29056 , n29054 , n29055 );
buf ( n29057 , RI173c3340_1804);
xor ( n29058 , n29056 , n29057 );
buf ( n29059 , RI1740c030_1449);
xor ( n29060 , n29058 , n29059 );
buf ( n29061 , RI173b6e60_1864);
xor ( n29062 , n29060 , n29061 );
xor ( n29063 , n29052 , n29062 );
and ( n29064 , n29039 , n29063 );
xor ( n29065 , n29013 , n29064 );
xor ( n29066 , n28999 , n29065 );
buf ( n29067 , RI173bf1a0_1824);
xor ( n29068 , n29067 , n27858 );
xor ( n29069 , n29068 , n27870 );
xor ( n29070 , RI19ab34f8_2429 , RI174a4808_934);
not ( n10613 , n27689 );
and ( n10614 , n10613 , RI174a4808_934);
and ( n10615 , n29070 , n27689 );
or ( n29071 , n10614 , n10615 );
buf ( n29072 , RI173362b0_2177);
xor ( n29073 , n29071 , n29072 );
buf ( n29074 , RI173bf830_1822);
xor ( n29075 , n29073 , n29074 );
buf ( n29076 , RI17408520_1467);
xor ( n29077 , n29075 , n29076 );
buf ( n29078 , RI17450d48_1342);
xor ( n29079 , n29077 , n29078 );
xor ( n29080 , n28209 , n29079 );
xor ( n29081 , n29080 , n28583 );
not ( n29082 , n29081 );
buf ( n29083 , RI1744b7f8_1368);
xor ( n29084 , RI19a922d0_2667 , RI17461a58_1260);
not ( n10616 , n27689 );
and ( n10617 , n10616 , RI17461a58_1260);
and ( n10618 , n29084 , n27689 );
or ( n29085 , n10617 , n10618 );
xor ( n29086 , RI19ac25e8_2311 , RI174aa730_905);
not ( n10619 , n27689 );
and ( n10620 , n10619 , RI174aa730_905);
and ( n10621 , n29086 , n27689 );
or ( n29087 , n10620 , n10621 );
xor ( n29088 , n29085 , n29087 );
xor ( n29089 , n29088 , n28483 );
buf ( n29090 , RI173c5410_1794);
xor ( n29091 , n29089 , n29090 );
buf ( n29092 , RI1740e100_1439);
xor ( n29093 , n29091 , n29092 );
xor ( n29094 , n29083 , n29093 );
xor ( n29095 , RI19aa5fb0_2523 , RI1747ef90_1117);
not ( n10622 , n27689 );
and ( n10623 , n10622 , RI1747ef90_1117);
and ( n10624 , n29095 , n27689 );
or ( n29096 , n10623 , n10624 );
xor ( n29097 , RI19a87218_2744 , RI174d07a0_762);
not ( n10625 , n27689 );
and ( n10626 , n10625 , RI174d07a0_762);
and ( n10627 , n29097 , n27689 );
or ( n29098 , n10626 , n10627 );
xor ( n29099 , n29096 , n29098 );
buf ( n29100 , RI17399c70_2006);
xor ( n29101 , n29099 , n29100 );
buf ( n29102 , RI173e2960_1651);
xor ( n29103 , n29101 , n29102 );
buf ( n29104 , RI1745a780_1295);
xor ( n29105 , n29103 , n29104 );
xor ( n29106 , n29094 , n29105 );
and ( n29107 , n29082 , n29106 );
xor ( n29108 , n29069 , n29107 );
xor ( n29109 , n29066 , n29108 );
xor ( n29110 , n28817 , n29109 );
not ( n29111 , n29110 );
buf ( n29112 , RI173acd98_1913);
xor ( n29113 , RI19aa3ee0_2538 , RI174837c0_1095);
not ( n10628 , n27689 );
and ( n10629 , n10628 , RI174837c0_1095);
and ( n10630 , n29113 , n27689 );
or ( n29114 , n10629 , n10630 );
xor ( n29115 , RI19a852b0_2758 , RI175085a0_740);
not ( n10631 , n27689 );
and ( n10632 , n10631 , RI175085a0_740);
and ( n10633 , n29115 , n27689 );
or ( n29116 , n10632 , n10633 );
xor ( n29117 , n29114 , n29116 );
buf ( n29118 , RI1739e4a0_1984);
xor ( n29119 , n29117 , n29118 );
buf ( n29120 , RI173e74d8_1628);
xor ( n29121 , n29119 , n29120 );
buf ( n29122 , RI1745efb0_1273);
xor ( n29123 , n29121 , n29122 );
xor ( n29124 , n29112 , n29123 );
xor ( n29125 , RI19ab5a00_2411 , RI174a0cf8_952);
not ( n10634 , n27689 );
and ( n10635 , n10634 , RI174a0cf8_952);
and ( n10636 , n29125 , n27689 );
or ( n29126 , n10635 , n10636 );
buf ( n29127 , RI173327a0_2195);
xor ( n29128 , n29126 , n29127 );
buf ( n29129 , RI173bbd20_1840);
xor ( n29130 , n29128 , n29129 );
buf ( n29131 , RI17404a10_1485);
xor ( n29132 , n29130 , n29131 );
buf ( n29133 , RI173fb668_1530);
xor ( n29134 , n29132 , n29133 );
xor ( n29135 , n29124 , n29134 );
buf ( n29136 , RI17400870_1505);
xor ( n29137 , n29136 , n28659 );
xor ( n29138 , RI19a92e10_2662 , RI17462ac0_1255);
not ( n10637 , n27689 );
and ( n10638 , n10637 , RI17462ac0_1255);
and ( n10639 , n29138 , n27689 );
or ( n29139 , n10638 , n10639 );
xor ( n29140 , RI19ac30b0_2306 , RI174ab798_900);
not ( n10640 , n27689 );
and ( n10641 , n10640 , RI174ab798_900);
and ( n10642 , n29140 , n27689 );
or ( n29141 , n10641 , n10642 );
xor ( n29142 , n29139 , n29141 );
buf ( n29143 , RI1733cef8_2144);
xor ( n29144 , n29142 , n29143 );
buf ( n29145 , RI173c6478_1789);
xor ( n29146 , n29144 , n29145 );
buf ( n29147 , RI1740f168_1434);
xor ( n29148 , n29146 , n29147 );
xor ( n29149 , n29137 , n29148 );
not ( n29150 , n29149 );
buf ( n29151 , RI17411238_1424);
xor ( n29152 , RI19ab7008_2402 , RI1749ef70_961);
not ( n10643 , n27689 );
and ( n10644 , n10643 , RI1749ef70_961);
and ( n10645 , n29152 , n27689 );
or ( n29153 , n10644 , n10645 );
buf ( n29154 , RI17533890_606);
xor ( n29155 , n29153 , n29154 );
buf ( n29156 , RI173b9f98_1849);
xor ( n29157 , n29155 , n29156 );
buf ( n29158 , RI17402c88_1494);
xor ( n29159 , n29157 , n29158 );
buf ( n29160 , RI173e9260_1619);
xor ( n29161 , n29159 , n29160 );
xor ( n29162 , n29151 , n29161 );
xor ( n29163 , n29162 , n28069 );
and ( n29164 , n29150 , n29163 );
xor ( n29165 , n29135 , n29164 );
xor ( n29166 , RI19a8bfe8_2711 , RI1746aab8_1216);
not ( n10646 , n27689 );
and ( n10647 , n10646 , RI1746aab8_1216);
and ( n10648 , n29166 , n27689 );
or ( n29167 , n10647 , n10648 );
xor ( n29168 , RI19abd4d0_2356 , RI174b3790_861);
not ( n10649 , n27689 );
and ( n10650 , n10649 , RI174b3790_861);
and ( n10651 , n29168 , n27689 );
or ( n29169 , n10650 , n10651 );
xor ( n29170 , n29167 , n29169 );
buf ( n29171 , RI17344ef0_2105);
xor ( n29172 , n29170 , n29171 );
buf ( n29173 , RI173ce7b8_1749);
xor ( n29174 , n29172 , n29173 );
buf ( n29175 , RI174462a8_1394);
xor ( n29176 , n29174 , n29175 );
xor ( n29177 , n28576 , n29176 );
xor ( n29178 , RI19aa0100_2568 , RI17487ff0_1073);
not ( n10652 , n27689 );
and ( n10653 , n10652 , RI17487ff0_1073);
and ( n10654 , n29178 , n27689 );
or ( n29179 , n10653 , n10654 );
xor ( n29180 , RI19aced20_2219 , RI1750f710_718);
not ( n10655 , n27689 );
and ( n10656 , n10655 , RI1750f710_718);
and ( n10657 , n29180 , n27689 );
or ( n29181 , n10656 , n10657 );
xor ( n29182 , n29179 , n29181 );
xor ( n29183 , n29182 , n28818 );
buf ( n29184 , RI173ebd08_1606);
xor ( n29185 , n29183 , n29184 );
buf ( n29186 , RI1747a0d0_1141);
xor ( n29187 , n29185 , n29186 );
xor ( n29188 , n29177 , n29187 );
xor ( n29189 , RI19a95de0_2641 , RI17479068_1146);
not ( n10658 , n27689 );
and ( n10659 , n10658 , RI17479068_1146);
and ( n10660 , n29189 , n27689 );
or ( n29190 , n10659 , n10660 );
xor ( n29191 , RI19ac5bd0_2286 , RI174c7218_791);
not ( n10661 , n27689 );
and ( n10662 , n10661 , RI174c7218_791);
and ( n10663 , n29191 , n27689 );
or ( n29192 , n10662 , n10663 );
xor ( n29193 , n29190 , n29192 );
buf ( n29194 , RI17393d48_2035);
xor ( n29195 , n29193 , n29194 );
buf ( n29196 , RI173dca38_1680);
xor ( n29197 , n29195 , n29196 );
buf ( n29198 , RI17454510_1325);
xor ( n29199 , n29197 , n29198 );
xor ( n29200 , n28169 , n29199 );
xor ( n29201 , RI19aa9bb0_2498 , RI174965a0_1003);
not ( n10664 , n27689 );
and ( n10665 , n10664 , RI174965a0_1003);
and ( n10666 , n29201 , n27689 );
or ( n29202 , n10665 , n10666 );
xor ( n29203 , RI19a9b420_2603 , RI17526000_648);
not ( n10667 , n27689 );
and ( n10668 , n10667 , RI17526000_648);
and ( n10669 , n29203 , n27689 );
or ( n29204 , n10668 , n10669 );
xor ( n29205 , n29202 , n29204 );
buf ( n29206 , RI173b1280_1892);
xor ( n29207 , n29205 , n29206 );
buf ( n29208 , RI173f9f70_1537);
xor ( n29209 , n29207 , n29208 );
buf ( n29210 , RI17392998_2041);
xor ( n29211 , n29209 , n29210 );
xor ( n29212 , n29200 , n29211 );
not ( n29213 , n29212 );
xor ( n29214 , RI19aa3580_2542 , RI17482758_1100);
not ( n10670 , n27689 );
and ( n10671 , n10670 , RI17482758_1100);
and ( n10672 , n29214 , n27689 );
or ( n29215 , n10671 , n10672 );
xor ( n29216 , RI19a84950_2762 , RI17506bd8_745);
not ( n10673 , n27689 );
and ( n10674 , n10673 , RI17506bd8_745);
and ( n10675 , n29216 , n27689 );
or ( n29217 , n10674 , n10675 );
xor ( n29218 , n29215 , n29217 );
buf ( n29219 , RI1739d438_1989);
xor ( n29220 , n29218 , n29219 );
buf ( n29221 , RI173e6470_1633);
xor ( n29222 , n29220 , n29221 );
buf ( n29223 , RI1745df48_1278);
xor ( n29224 , n29222 , n29223 );
xor ( n29225 , n28477 , n29224 );
xor ( n29226 , RI19ab7878_2398 , RI1749fc90_957);
not ( n10676 , n27689 );
and ( n10677 , n10676 , RI1749fc90_957);
and ( n10678 , n29226 , n27689 );
or ( n29227 , n10677 , n10678 );
buf ( n29228 , RI17534d30_602);
xor ( n29229 , n29227 , n29228 );
buf ( n29230 , RI173bacb8_1845);
xor ( n29231 , n29229 , n29230 );
buf ( n29232 , RI174039a8_1490);
xor ( n29233 , n29231 , n29232 );
buf ( n29234 , RI173f22c0_1575);
xor ( n29235 , n29233 , n29234 );
xor ( n29236 , n29225 , n29235 );
and ( n29237 , n29213 , n29236 );
xor ( n29238 , n29188 , n29237 );
xor ( n29239 , n28976 , n28081 );
xor ( n29240 , RI19ac04a0_2329 , RI174ae240_887);
not ( n10679 , n27689 );
and ( n10680 , n10679 , RI174ae240_887);
and ( n10681 , n29240 , n27689 );
or ( n29241 , n10680 , n10681 );
xor ( n29242 , n27690 , n29241 );
buf ( n29243 , RI1733f9a0_2131);
xor ( n29244 , n29242 , n29243 );
buf ( n29245 , RI173c8f20_1776);
xor ( n29246 , n29244 , n29245 );
buf ( n29247 , RI17411c10_1421);
xor ( n29248 , n29246 , n29247 );
xor ( n29249 , n29239 , n29248 );
xor ( n29250 , RI19ab98d0_2384 , RI1749b7a8_978);
not ( n10682 , n27689 );
and ( n10683 , n10682 , RI1749b7a8_978);
and ( n10684 , n29250 , n27689 );
or ( n29251 , n10683 , n10684 );
buf ( n29252 , RI1752e0e8_623);
xor ( n29253 , n29251 , n29252 );
buf ( n29254 , RI173b6488_1867);
xor ( n29255 , n29253 , n29254 );
buf ( n29256 , RI173ff4c0_1511);
xor ( n29257 , n29255 , n29256 );
buf ( n29258 , RI173c6e50_1786);
xor ( n29259 , n29257 , n29258 );
xor ( n29260 , n28245 , n29259 );
xor ( n29261 , RI19a9c398_2596 , RI17470008_1190);
not ( n10685 , n27689 );
and ( n10686 , n10685 , RI17470008_1190);
and ( n10687 , n29261 , n27689 );
or ( n29262 , n10686 , n10687 );
xor ( n29263 , RI19acb648_2244 , RI174b8f38_835);
not ( n10688 , n27689 );
and ( n10689 , n10688 , RI174b8f38_835);
and ( n10690 , n29263 , n27689 );
or ( n29264 , n10689 , n10690 );
xor ( n29265 , n29262 , n29264 );
buf ( n29266 , RI1738b030_2078);
xor ( n29267 , n29265 , n29266 );
buf ( n29268 , RI173d3d20_1723);
xor ( n29269 , n29267 , n29268 );
xor ( n29270 , n29269 , n29083 );
xor ( n29271 , n29260 , n29270 );
not ( n29272 , n29271 );
xor ( n29273 , n28824 , n28557 );
xor ( n29274 , n29273 , n28569 );
and ( n29275 , n29272 , n29274 );
xor ( n29276 , n29249 , n29275 );
xor ( n29277 , n29238 , n29276 );
xor ( n29278 , RI19a87470_2743 , RI174d0cc8_761);
not ( n10691 , n27689 );
and ( n10692 , n10691 , RI174d0cc8_761);
and ( n10693 , n29278 , n27689 );
or ( n29279 , n10692 , n10693 );
xor ( n29280 , n29279 , n28904 );
xor ( n29281 , RI19ab0528_2451 , RI1748dbd0_1045);
not ( n10694 , n27689 );
and ( n10695 , n10694 , RI1748dbd0_1045);
and ( n10696 , n29281 , n27689 );
or ( n29282 , n10695 , n10696 );
xor ( n29283 , RI19ab3a20_2426 , RI17518c98_689);
not ( n10697 , n27689 );
and ( n10698 , n10697 , RI17518c98_689);
and ( n10699 , n29283 , n27689 );
or ( n29284 , n10698 , n10699 );
xor ( n29285 , n29282 , n29284 );
buf ( n29286 , RI173a8bf8_1933);
xor ( n29287 , n29285 , n29286 );
buf ( n29288 , RI173f18e8_1578);
xor ( n29289 , n29287 , n29288 );
buf ( n29290 , RI174b51d0_853);
xor ( n29291 , n29289 , n29290 );
xor ( n29292 , n29280 , n29291 );
not ( n29293 , n29135 );
and ( n29294 , n29293 , n29149 );
xor ( n29295 , n29292 , n29294 );
xor ( n29296 , n29277 , n29295 );
xor ( n29297 , RI19ab4bf0_2418 , RI174a3110_941);
not ( n10700 , n27689 );
and ( n10701 , n10700 , RI174a3110_941);
and ( n10702 , n29297 , n27689 );
or ( n29298 , n10701 , n10702 );
buf ( n29299 , RI17334bb8_2184);
xor ( n29300 , n29298 , n29299 );
buf ( n29301 , RI173be138_1829);
xor ( n29302 , n29300 , n29301 );
buf ( n29303 , RI17406e28_1474);
xor ( n29304 , n29302 , n29303 );
buf ( n29305 , RI174122a0_1419);
xor ( n29306 , n29304 , n29305 );
xor ( n29307 , n27784 , n29306 );
xor ( n29308 , n29307 , n28406 );
buf ( n29309 , RI1738c728_2071);
xor ( n29310 , RI19a90a70_2678 , RI17462e08_1254);
not ( n10703 , n27689 );
and ( n10704 , n10703 , RI17462e08_1254);
and ( n10705 , n29310 , n27689 );
or ( n29311 , n10704 , n10705 );
xor ( n29312 , RI19ac0f68_2323 , RI174abae0_899);
not ( n10706 , n27689 );
and ( n10707 , n10706 , RI174abae0_899);
and ( n10708 , n29312 , n27689 );
or ( n29313 , n10707 , n10708 );
xor ( n29314 , n29311 , n29313 );
buf ( n29315 , RI1733d240_2143);
xor ( n29316 , n29314 , n29315 );
buf ( n29317 , RI173c67c0_1788);
xor ( n29318 , n29316 , n29317 );
buf ( n29319 , RI1740f4b0_1433);
xor ( n29320 , n29318 , n29319 );
xor ( n29321 , n29309 , n29320 );
xor ( n29322 , RI19aa46d8_2534 , RI17480340_1111);
not ( n10709 , n27689 );
and ( n10710 , n10709 , RI17480340_1111);
and ( n10711 , n29322 , n27689 );
or ( n29323 , n10710 , n10711 );
xor ( n29324 , RI19a859b8_2755 , RI175014a8_756);
not ( n10712 , n27689 );
and ( n10713 , n10712 , RI175014a8_756);
and ( n10714 , n29324 , n27689 );
or ( n29325 , n10713 , n10714 );
xor ( n29326 , n29323 , n29325 );
buf ( n29327 , RI1739b020_2000);
xor ( n29328 , n29326 , n29327 );
buf ( n29329 , RI173e3d10_1645);
xor ( n29330 , n29328 , n29329 );
buf ( n29331 , RI1745bb30_1289);
xor ( n29332 , n29330 , n29331 );
xor ( n29333 , n29321 , n29332 );
not ( n29334 , n29333 );
buf ( n29335 , RI173e50c0_1639);
xor ( n29336 , RI19a9b8d0_2601 , RI17472768_1178);
not ( n10715 , n27689 );
and ( n10716 , n10715 , RI17472768_1178);
and ( n10717 , n29336 , n27689 );
or ( n29337 , n10716 , n10717 );
xor ( n29338 , RI19acadd8_2249 , RI174bcd18_823);
not ( n10718 , n27689 );
and ( n10719 , n10718 , RI174bcd18_823);
and ( n10720 , n29338 , n27689 );
or ( n29339 , n10719 , n10720 );
xor ( n29340 , n29337 , n29339 );
buf ( n29341 , RI1738d790_2066);
xor ( n29342 , n29340 , n29341 );
buf ( n29343 , RI173d6480_1711);
xor ( n29344 , n29342 , n29343 );
buf ( n29345 , RI1744df58_1356);
xor ( n29346 , n29344 , n29345 );
xor ( n29347 , n29335 , n29346 );
xor ( n29348 , n29347 , n28866 );
and ( n29349 , n29334 , n29348 );
xor ( n29350 , n29308 , n29349 );
xor ( n29351 , n29296 , n29350 );
xor ( n29352 , RI19a93518_2659 , RI17529de0_636);
not ( n10721 , n27689 );
and ( n10722 , n10721 , RI17529de0_636);
and ( n10723 , n29352 , n27689 );
or ( n29353 , n10722 , n10723 );
xor ( n29354 , RI19a9f368_2575 , RI1748a408_1062);
not ( n10724 , n27689 );
and ( n10725 , n10724 , RI1748a408_1062);
and ( n10726 , n29354 , n27689 );
or ( n29355 , n10725 , n10726 );
xor ( n29356 , RI19acdf10_2225 , RI175134f0_706);
not ( n10727 , n27689 );
and ( n10728 , n10727 , RI175134f0_706);
and ( n10729 , n29356 , n27689 );
or ( n29357 , n10728 , n10729 );
xor ( n29358 , n29355 , n29357 );
buf ( n29359 , RI173a5430_1950);
xor ( n29360 , n29358 , n29359 );
buf ( n29361 , RI173ee120_1595);
xor ( n29362 , n29360 , n29361 );
buf ( n29363 , RI17490d08_1030);
xor ( n29364 , n29362 , n29363 );
xor ( n29365 , n29353 , n29364 );
xor ( n29366 , RI19ab2f58_2432 , RI174a7c88_918);
not ( n10730 , n27689 );
and ( n10731 , n10730 , RI174a7c88_918);
and ( n10732 , n29366 , n27689 );
or ( n29367 , n10731 , n10732 );
buf ( n29368 , RI173393e8_2162);
xor ( n29369 , n29367 , n29368 );
buf ( n29370 , RI173c2968_1807);
xor ( n29371 , n29369 , n29370 );
buf ( n29372 , RI1740b658_1452);
xor ( n29373 , n29371 , n29372 );
buf ( n29374 , RI17332110_2197);
xor ( n29375 , n29373 , n29374 );
xor ( n29376 , n29365 , n29375 );
xor ( n29377 , RI19aab5f0_2486 , RI174951f0_1009);
not ( n10733 , n27689 );
and ( n10734 , n10733 , RI174951f0_1009);
and ( n10735 , n29377 , n27689 );
or ( n29378 , n10734 , n10735 );
xor ( n29379 , RI19aac388_2481 , RI17524110_654);
not ( n10736 , n27689 );
and ( n10737 , n10736 , RI17524110_654);
and ( n10738 , n29379 , n27689 );
or ( n29380 , n10737 , n10738 );
xor ( n29381 , n29378 , n29380 );
buf ( n29382 , RI173afed0_1898);
xor ( n29383 , n29381 , n29382 );
buf ( n29384 , RI173f8bc0_1543);
xor ( n29385 , n29383 , n29384 );
buf ( n29386 , RI17346930_2097);
xor ( n29387 , n29385 , n29386 );
xor ( n29388 , n27880 , n29387 );
xor ( n29389 , RI19a8dd70_2698 , RI17469a50_1221);
not ( n10739 , n27689 );
and ( n10740 , n10739 , RI17469a50_1221);
and ( n10741 , n29389 , n27689 );
or ( n29390 , n10740 , n10741 );
xor ( n29391 , RI19abebc8_2343 , RI174b2728_866);
not ( n10742 , n27689 );
and ( n10743 , n10742 , RI174b2728_866);
and ( n10744 , n29391 , n27689 );
or ( n29392 , n10743 , n10744 );
xor ( n29393 , n29390 , n29392 );
buf ( n29394 , RI17343e88_2110);
xor ( n29395 , n29393 , n29394 );
buf ( n29396 , RI173cd408_1755);
xor ( n29397 , n29395 , n29396 );
buf ( n29398 , RI17445240_1399);
xor ( n29399 , n29397 , n29398 );
xor ( n29400 , n29388 , n29399 );
not ( n29401 , n29400 );
xor ( n29402 , RI19ab5820_2412 , RI174a4178_936);
not ( n10745 , n27689 );
and ( n10746 , n10745 , RI174a4178_936);
and ( n10747 , n29402 , n27689 );
or ( n29403 , n10746 , n10747 );
xor ( n29404 , n29403 , n27847 );
xor ( n29405 , n29404 , n29067 );
buf ( n29406 , RI17407e90_1469);
xor ( n29407 , n29405 , n29406 );
buf ( n29408 , RI1744c518_1364);
xor ( n29409 , n29407 , n29408 );
xor ( n29410 , n28809 , n29409 );
xor ( n29411 , RI19a95b88_2642 , RI17478d20_1147);
not ( n10748 , n27689 );
and ( n10749 , n10748 , RI17478d20_1147);
and ( n10750 , n29411 , n27689 );
or ( n29412 , n10749 , n10750 );
xor ( n29413 , RI19ac5978_2287 , RI174c6cf0_792);
not ( n10751 , n27689 );
and ( n10752 , n10751 , RI174c6cf0_792);
and ( n10753 , n29413 , n27689 );
or ( n29414 , n10752 , n10753 );
xor ( n29415 , n29412 , n29414 );
buf ( n29416 , RI17393a00_2036);
xor ( n29417 , n29415 , n29416 );
buf ( n29418 , RI173dc6f0_1681);
xor ( n29419 , n29417 , n29418 );
buf ( n29420 , RI174541c8_1326);
xor ( n29421 , n29419 , n29420 );
xor ( n29422 , n29410 , n29421 );
and ( n29423 , n29401 , n29422 );
xor ( n29424 , n29376 , n29423 );
xor ( n29425 , n29351 , n29424 );
xor ( n29426 , n29165 , n29425 );
buf ( n29427 , RI173f50b0_1561);
xor ( n29428 , RI19aa38c8_2541 , RI17482aa0_1099);
not ( n10754 , n27689 );
and ( n10755 , n10754 , RI17482aa0_1099);
and ( n10756 , n29428 , n27689 );
or ( n29429 , n10755 , n10756 );
xor ( n29430 , RI19a84ba8_2761 , RI17507100_744);
not ( n10757 , n27689 );
and ( n10758 , n10757 , RI17507100_744);
and ( n10759 , n29430 , n27689 );
or ( n29431 , n10758 , n10759 );
xor ( n29432 , n29429 , n29431 );
buf ( n29433 , RI1739d780_1988);
xor ( n29434 , n29432 , n29433 );
buf ( n29435 , RI173e67b8_1632);
xor ( n29436 , n29434 , n29435 );
buf ( n29437 , RI1745e290_1277);
xor ( n29438 , n29436 , n29437 );
xor ( n29439 , n29427 , n29438 );
xor ( n29440 , RI19ab7a58_2397 , RI1749ffd8_956);
not ( n10760 , n27689 );
and ( n10761 , n10760 , RI1749ffd8_956);
and ( n10762 , n29440 , n27689 );
or ( n29441 , n10761 , n10762 );
buf ( n29442 , RI17535258_601);
xor ( n29443 , n29441 , n29442 );
buf ( n29444 , RI173bb000_1844);
xor ( n29445 , n29443 , n29444 );
buf ( n29446 , RI17403cf0_1489);
xor ( n29447 , n29445 , n29446 );
buf ( n29448 , RI173f46d8_1564);
xor ( n29449 , n29447 , n29448 );
xor ( n29450 , n29439 , n29449 );
buf ( n29451 , RI173e22d0_1653);
xor ( n29452 , RI19aaf268_2460 , RI1748fca0_1035);
not ( n10763 , n27689 );
and ( n10764 , n10763 , RI1748fca0_1035);
and ( n10765 , n29452 , n27689 );
or ( n29453 , n10764 , n10765 );
xor ( n29454 , RI19a23c18_2790 , RI1751bb00_680);
not ( n10766 , n27689 );
and ( n10767 , n10766 , RI1751bb00_680);
and ( n10768 , n29454 , n27689 );
or ( n29455 , n10767 , n10768 );
xor ( n29456 , n29453 , n29455 );
buf ( n29457 , RI173aa980_1924);
xor ( n29458 , n29456 , n29457 );
buf ( n29459 , RI173f3670_1569);
xor ( n29460 , n29458 , n29459 );
buf ( n29461 , RI174cfd50_764);
xor ( n29462 , n29460 , n29461 );
xor ( n29463 , n29451 , n29462 );
xor ( n29464 , RI19a91808_2672 , RI17464500_1247);
not ( n10769 , n27689 );
and ( n10770 , n10769 , RI17464500_1247);
and ( n10771 , n29464 , n27689 );
or ( n29465 , n10770 , n10771 );
xor ( n29466 , RI19ac1a30_2317 , RI174ad1d8_892);
not ( n10772 , n27689 );
and ( n10773 , n10772 , RI174ad1d8_892);
and ( n10774 , n29466 , n27689 );
or ( n29467 , n10773 , n10774 );
xor ( n29468 , n29465 , n29467 );
buf ( n29469 , RI1733e938_2136);
xor ( n29470 , n29468 , n29469 );
buf ( n29471 , RI173c7eb8_1781);
xor ( n29472 , n29470 , n29471 );
buf ( n29473 , RI17410ba8_1426);
xor ( n29474 , n29472 , n29473 );
xor ( n29475 , n29463 , n29474 );
not ( n29476 , n29475 );
and ( n29477 , n29476 , n28544 );
xor ( n29478 , n29450 , n29477 );
buf ( n29479 , RI174a09b0_953);
xor ( n29480 , RI19a93ba8_2656 , RI1747d550_1125);
not ( n10775 , n27689 );
and ( n10776 , n10775 , RI1747d550_1125);
and ( n10777 , n29480 , n27689 );
or ( n29481 , n10776 , n10777 );
xor ( n29482 , RI19ac3d58_2300 , RI174cde60_770);
not ( n10778 , n27689 );
and ( n10779 , n10778 , RI174cde60_770);
and ( n10780 , n29482 , n27689 );
or ( n29483 , n10779 , n10780 );
xor ( n29484 , n29481 , n29483 );
buf ( n29485 , RI17398230_2014);
xor ( n29486 , n29484 , n29485 );
buf ( n29487 , RI173e0f20_1659);
xor ( n29488 , n29486 , n29487 );
buf ( n29489 , RI17458d40_1303);
xor ( n29490 , n29488 , n29489 );
xor ( n29491 , n29479 , n29490 );
xor ( n29492 , RI19aa7a68_2512 , RI1749aa88_982);
not ( n10781 , n27689 );
and ( n10782 , n10781 , RI1749aa88_982);
and ( n10783 , n29492 , n27689 );
or ( n29493 , n10782 , n10783 );
xor ( n29494 , RI19a88be0_2733 , RI1752cc48_627);
not ( n10784 , n27689 );
and ( n10785 , n10784 , RI1752cc48_627);
and ( n10786 , n29494 , n27689 );
or ( n29495 , n10785 , n10786 );
xor ( n29496 , n29493 , n29495 );
buf ( n29497 , RI173b5768_1871);
xor ( n29498 , n29496 , n29497 );
buf ( n29499 , RI173fe7a0_1515);
xor ( n29500 , n29498 , n29499 );
buf ( n29501 , RI173bddf0_1830);
xor ( n29502 , n29500 , n29501 );
xor ( n29503 , n29491 , n29502 );
not ( n29504 , n29503 );
and ( n29505 , n29504 , n28628 );
xor ( n29506 , n28521 , n29505 );
xor ( n29507 , n29478 , n29506 );
buf ( n29508 , RI17400bb8_1504);
xor ( n29509 , RI19ab0a50_2449 , RI1748e260_1043);
not ( n10787 , n27689 );
and ( n10788 , n10787 , RI1748e260_1043);
and ( n10789 , n29509 , n27689 );
or ( n29510 , n10788 , n10789 );
xor ( n29511 , RI19ad0238_2210 , RI175196e8_687);
not ( n10790 , n27689 );
and ( n10791 , n10790 , RI175196e8_687);
and ( n10792 , n29511 , n27689 );
or ( n29512 , n10791 , n10792 );
xor ( n29513 , n29510 , n29512 );
buf ( n29514 , RI173a9288_1931);
xor ( n29515 , n29513 , n29514 );
buf ( n29516 , RI173f1f78_1576);
xor ( n29517 , n29515 , n29516 );
buf ( n29518 , RI174ba3d8_831);
xor ( n29519 , n29517 , n29518 );
xor ( n29520 , n29508 , n29519 );
xor ( n29521 , n29520 , n29320 );
buf ( n29522 , RI17411580_1423);
xor ( n29523 , RI19ab71e8_2401 , RI1749f2b8_960);
not ( n10793 , n27689 );
and ( n10794 , n10793 , RI1749f2b8_960);
and ( n10795 , n29523 , n27689 );
or ( n29524 , n10794 , n10795 );
buf ( n29525 , RI17533db8_605);
xor ( n29526 , n29524 , n29525 );
buf ( n29527 , RI173ba2e0_1848);
xor ( n29528 , n29526 , n29527 );
buf ( n29529 , RI17402fd0_1493);
xor ( n29530 , n29528 , n29529 );
buf ( n29531 , RI173eb678_1608);
xor ( n29532 , n29530 , n29531 );
xor ( n29533 , n29522 , n29532 );
xor ( n29534 , RI19a99d28_2613 , RI17473b18_1172);
not ( n10796 , n27689 );
and ( n10797 , n10796 , RI17473b18_1172);
and ( n10798 , n29534 , n27689 );
or ( n29535 , n10797 , n10798 );
xor ( n29536 , RI19ac9500_2260 , RI174bf130_816);
not ( n10799 , n27689 );
and ( n10800 , n10799 , RI174bf130_816);
and ( n10801 , n29536 , n27689 );
or ( n29537 , n10800 , n10801 );
xor ( n29538 , n29535 , n29537 );
buf ( n29539 , RI1738eb40_2060);
xor ( n29540 , n29538 , n29539 );
buf ( n29541 , RI173d7830_1705);
xor ( n29542 , n29540 , n29541 );
buf ( n29543 , RI1744f308_1350);
xor ( n29544 , n29542 , n29543 );
xor ( n29545 , n29533 , n29544 );
not ( n29546 , n29545 );
and ( n29547 , n29546 , n28634 );
xor ( n29548 , n29521 , n29547 );
xor ( n29549 , n29507 , n29548 );
buf ( n29550 , RI173e5408_1638);
xor ( n29551 , RI19a9bb28_2600 , RI17472ab0_1177);
not ( n10802 , n27689 );
and ( n10803 , n10802 , RI17472ab0_1177);
and ( n10804 , n29551 , n27689 );
or ( n29552 , n10803 , n10804 );
xor ( n29553 , RI19acaf40_2248 , RI174bd240_822);
not ( n10805 , n27689 );
and ( n10806 , n10805 , RI174bd240_822);
and ( n10807 , n29553 , n27689 );
or ( n29554 , n10806 , n10807 );
xor ( n29555 , n29552 , n29554 );
buf ( n29556 , RI1738dad8_2065);
xor ( n29557 , n29555 , n29556 );
buf ( n29558 , RI173d67c8_1710);
xor ( n29559 , n29557 , n29558 );
buf ( n29560 , RI1744e2a0_1355);
xor ( n29561 , n29559 , n29560 );
xor ( n29562 , n29550 , n29561 );
xor ( n29563 , RI19aaf790_2457 , RI17490330_1033);
not ( n10808 , n27689 );
and ( n10809 , n10808 , RI17490330_1033);
and ( n10810 , n29563 , n27689 );
or ( n29564 , n10809 , n10810 );
xor ( n29565 , RI19a83b40_2768 , RI1751c550_678);
not ( n10811 , n27689 );
and ( n10812 , n10811 , RI1751c550_678);
and ( n10813 , n29565 , n27689 );
or ( n29566 , n10812 , n10813 );
xor ( n29567 , n29564 , n29566 );
buf ( n29568 , RI173ab010_1922);
xor ( n29569 , n29567 , n29568 );
buf ( n29570 , RI173f3d00_1567);
xor ( n29571 , n29569 , n29570 );
buf ( n29572 , RI17507b50_742);
xor ( n29573 , n29571 , n29572 );
xor ( n29574 , n29562 , n29573 );
buf ( n29575 , RI173b0218_1897);
xor ( n29576 , RI19a9f728_2573 , RI1748aa98_1060);
not ( n10814 , n27689 );
and ( n10815 , n10814 , RI1748aa98_1060);
and ( n10816 , n29576 , n27689 );
or ( n29577 , n10815 , n10816 );
xor ( n29578 , RI19ace3c0_2223 , RI17513f40_704);
not ( n10817 , n27689 );
and ( n10818 , n10817 , RI17513f40_704);
and ( n10819 , n29578 , n27689 );
or ( n29579 , n10818 , n10819 );
xor ( n29580 , n29577 , n29579 );
buf ( n29581 , RI173a5ac0_1948);
xor ( n29582 , n29580 , n29581 );
buf ( n29583 , RI173ee7b0_1593);
xor ( n29584 , n29582 , n29583 );
buf ( n29585 , RI17495538_1008);
xor ( n29586 , n29584 , n29585 );
xor ( n29587 , n29575 , n29586 );
xor ( n29588 , n29587 , n28355 );
not ( n29589 , n29588 );
and ( n29590 , n29589 , n28703 );
xor ( n29591 , n29574 , n29590 );
xor ( n29592 , n29549 , n29591 );
xor ( n29593 , RI19ab3318_2430 , RI174a44c0_935);
not ( n10820 , n27689 );
and ( n10821 , n10820 , RI174a44c0_935);
and ( n10822 , n29593 , n27689 );
or ( n29594 , n10821 , n10822 );
xor ( n29595 , n29594 , n28189 );
buf ( n29596 , RI173bf4e8_1823);
xor ( n29597 , n29595 , n29596 );
buf ( n29598 , RI174081d8_1468);
xor ( n29599 , n29597 , n29598 );
buf ( n29600 , RI1744e930_1353);
xor ( n29601 , n29599 , n29600 );
xor ( n29602 , n27867 , n29601 );
xor ( n29603 , n29602 , n29199 );
buf ( n29604 , RI1744b4b0_1369);
xor ( n29605 , n29604 , n28250 );
xor ( n29606 , n29605 , n28262 );
not ( n29607 , n29606 );
and ( n29608 , n29607 , n28772 );
xor ( n29609 , n29603 , n29608 );
xor ( n29610 , n29592 , n29609 );
xor ( n29611 , n29426 , n29610 );
and ( n29612 , n29111 , n29611 );
xor ( n29613 , n28469 , n29612 );
or ( n29614 , RI1753aa78_586 , n27689 );
not ( n10823 , n29614 );
and ( n10824 , n10823 , RI17465568_1242);
and ( n10825 , n29613 , n29614 );
or ( n29615 , n10824 , n10825 );
not ( n10826 , RI1754c610_2);
and ( n10827 , n10826 , n29615 );
and ( n10828 , C0 , RI1754c610_2);
or ( n29616 , n10827 , n10828 );
buf ( n29617 , n29616 );
xor ( n29618 , RI19a8a080_2724 , RI1746f2e8_1194);
not ( n10829 , n27689 );
and ( n10830 , n10829 , RI1746f2e8_1194);
and ( n10831 , n29618 , n27689 );
or ( n29619 , n10830 , n10831 );
xor ( n29620 , RI19abbc70_2369 , RI174b7fc0_839);
not ( n10832 , n27689 );
and ( n10833 , n10832 , RI174b7fc0_839);
and ( n10834 , n29620 , n27689 );
or ( n29621 , n10833 , n10834 );
xor ( n29622 , n29619 , n29621 );
buf ( n29623 , RI1738a310_2082);
xor ( n29624 , n29622 , n29623 );
buf ( n29625 , RI173d3000_1727);
xor ( n29626 , n29624 , n29625 );
buf ( n29627 , RI1744aad8_1372);
xor ( n29628 , n29626 , n29627 );
xor ( n29629 , n27745 , n29628 );
xor ( n29630 , RI19a9e468_2582 , RI1748c820_1051);
not ( n10835 , n27689 );
and ( n10836 , n10835 , RI1748c820_1051);
and ( n10837 , n29630 , n27689 );
or ( n29631 , n10836 , n10837 );
xor ( n29632 , RI19acd100_2231 , RI17516da8_695);
not ( n10838 , n27689 );
and ( n10839 , n10838 , RI17516da8_695);
and ( n10840 , n29632 , n27689 );
or ( n29633 , n10839 , n10840 );
xor ( n29634 , n29631 , n29633 );
xor ( n29635 , n29634 , n28139 );
buf ( n29636 , RI173f0538_1584);
xor ( n29637 , n29635 , n29636 );
buf ( n29638 , RI174a7940_919);
xor ( n29639 , n29637 , n29638 );
xor ( n29640 , n29629 , n29639 );
buf ( n29641 , RI173a6e70_1942);
xor ( n29642 , n29641 , n28759 );
xor ( n29643 , n29642 , n28771 );
not ( n29644 , n29643 );
xor ( n29645 , RI19aa19d8_2555 , RI17486f88_1078);
not ( n10841 , n27689 );
and ( n10842 , n10841 , RI17486f88_1078);
and ( n10843 , n29645 , n27689 );
or ( n29646 , n10842 , n10843 );
xor ( n29647 , RI19a82b50_2775 , RI1750dd48_723);
not ( n10844 , n27689 );
and ( n10845 , n10844 , RI1750dd48_723);
and ( n10846 , n29647 , n27689 );
or ( n29648 , n10845 , n10846 );
xor ( n29649 , n29646 , n29648 );
buf ( n29650 , RI173a1fb0_1966);
xor ( n29651 , n29649 , n29650 );
buf ( n29652 , RI173eaca0_1611);
xor ( n29653 , n29651 , n29652 );
buf ( n29654 , RI17470d28_1186);
xor ( n29655 , n29653 , n29654 );
xor ( n29656 , n27855 , n29655 );
xor ( n29657 , n29656 , n29601 );
and ( n29658 , n29644 , n29657 );
xor ( n29659 , n29640 , n29658 );
xor ( n29660 , RI19a8faf8_2685 , RI17465220_1243);
not ( n10847 , n27689 );
and ( n10848 , n10847 , RI17465220_1243);
and ( n10849 , n29660 , n27689 );
or ( n29661 , n10848 , n10849 );
xor ( n29662 , n29661 , n28983 );
xor ( n29663 , n29662 , n28995 );
not ( n29664 , n29640 );
and ( n29665 , n29664 , n29643 );
xor ( n29666 , n29663 , n29665 );
xor ( n29667 , n27980 , n28929 );
xor ( n29668 , RI19ab4560_2421 , RI174a6248_926);
not ( n10850 , n27689 );
and ( n10851 , n10850 , RI174a6248_926);
and ( n10852 , n29668 , n27689 );
or ( n29669 , n10851 , n10852 );
buf ( n29670 , RI173379a8_2170);
xor ( n29671 , n29669 , n29670 );
buf ( n29672 , RI173c0f28_1815);
xor ( n29673 , n29671 , n29672 );
buf ( n29674 , RI17409c18_1460);
xor ( n29675 , n29673 , n29674 );
buf ( n29676 , RI1745e920_1275);
xor ( n29677 , n29675 , n29676 );
xor ( n29678 , n29667 , n29677 );
buf ( n29679 , RI173358d8_2180);
xor ( n29680 , n29679 , n28800 );
xor ( n29681 , n29680 , n28812 );
not ( n29682 , n29681 );
xor ( n29683 , n28038 , n29449 );
xor ( n29684 , RI19a9a610_2609 , RI17474838_1168);
not ( n10853 , n27689 );
and ( n10854 , n10853 , RI17474838_1168);
and ( n10855 , n29684 , n27689 );
or ( n29685 , n10854 , n10855 );
xor ( n29686 , RI19ac9de8_2256 , RI174c05d0_812);
not ( n10856 , n27689 );
and ( n10857 , n10856 , RI174c05d0_812);
and ( n10858 , n29686 , n27689 );
or ( n29687 , n10857 , n10858 );
xor ( n29688 , n29685 , n29687 );
buf ( n29689 , RI1738f860_2056);
xor ( n29690 , n29688 , n29689 );
buf ( n29691 , RI173d8550_1701);
xor ( n29692 , n29690 , n29691 );
buf ( n29693 , RI17450028_1346);
xor ( n29694 , n29692 , n29693 );
xor ( n29695 , n29683 , n29694 );
and ( n29696 , n29682 , n29695 );
xor ( n29697 , n29678 , n29696 );
xor ( n29698 , n29666 , n29697 );
xor ( n29699 , n28986 , n29248 );
xor ( n29700 , n29699 , n29438 );
xor ( n29701 , n28666 , n28236 );
xor ( n29702 , RI19aac040_2482 , RI17492748_1022);
not ( n10859 , n27689 );
and ( n10860 , n10859 , RI17492748_1022);
and ( n10861 , n29702 , n27689 );
or ( n29703 , n10860 , n10861 );
xor ( n29704 , RI19ab2508_2437 , RI1751fe08_667);
not ( n10862 , n27689 );
and ( n10863 , n10862 , RI1751fe08_667);
and ( n10864 , n29704 , n27689 );
or ( n29705 , n10863 , n10864 );
xor ( n29706 , n29703 , n29705 );
xor ( n29707 , n29706 , n28938 );
buf ( n29708 , RI173f6118_1556);
xor ( n29709 , n29707 , n29708 );
buf ( n29710 , RI1752b7a8_631);
xor ( n29711 , n29709 , n29710 );
xor ( n29712 , n29701 , n29711 );
not ( n29713 , n29712 );
xor ( n29714 , n28590 , n29187 );
xor ( n29715 , RI19ab3de0_2424 , RI174a5870_929);
not ( n10865 , n27689 );
and ( n10866 , n10865 , RI174a5870_929);
and ( n10867 , n29715 , n27689 );
or ( n29716 , n10866 , n10867 );
buf ( n29717 , RI17336fd0_2173);
xor ( n29718 , n29716 , n29717 );
buf ( n29719 , RI173c0550_1818);
xor ( n29720 , n29718 , n29719 );
buf ( n29721 , RI17409240_1463);
xor ( n29722 , n29720 , n29721 );
buf ( n29723 , RI17457cd8_1308);
xor ( n29724 , n29722 , n29723 );
xor ( n29725 , n29714 , n29724 );
and ( n29726 , n29713 , n29725 );
xor ( n29727 , n29700 , n29726 );
xor ( n29728 , n29698 , n29727 );
xor ( n29729 , RI19ab4038_2423 , RI174a5bb8_928);
not ( n10868 , n27689 );
and ( n10869 , n10868 , RI174a5bb8_928);
and ( n10870 , n29729 , n27689 );
or ( n29730 , n10869 , n10870 );
xor ( n29731 , RI19aaa150_2495 , RI17496f78_1000);
not ( n10871 , n27689 );
and ( n10872 , n10871 , RI17496f78_1000);
and ( n10873 , n29731 , n27689 );
or ( n29732 , n10872 , n10873 );
xor ( n29733 , RI19a9fcc8_2570 , RI17526f78_645);
not ( n10874 , n27689 );
and ( n10875 , n10874 , RI17526f78_645);
and ( n10876 , n29733 , n27689 );
or ( n29734 , n10875 , n10876 );
xor ( n29735 , n29732 , n29734 );
xor ( n29736 , n29735 , n28293 );
buf ( n29737 , RI173fa948_1534);
xor ( n29738 , n29736 , n29737 );
buf ( n29739 , RI173995e0_2008);
xor ( n29740 , n29738 , n29739 );
xor ( n29741 , n29730 , n29740 );
xor ( n29742 , RI19a8c948_2707 , RI1746b7d8_1212);
not ( n10877 , n27689 );
and ( n10878 , n10877 , RI1746b7d8_1212);
and ( n10879 , n29742 , n27689 );
or ( n29743 , n10878 , n10879 );
xor ( n29744 , RI19abdbd8_2352 , RI174b44b0_857);
not ( n10880 , n27689 );
and ( n10881 , n10880 , RI174b44b0_857);
and ( n10882 , n29744 , n27689 );
or ( n29745 , n10881 , n10882 );
xor ( n29746 , n29743 , n29745 );
buf ( n29747 , RI17345c10_2101);
xor ( n29748 , n29746 , n29747 );
buf ( n29749 , RI173cf4d8_1745);
xor ( n29750 , n29748 , n29749 );
buf ( n29751 , RI17446fc8_1390);
xor ( n29752 , n29750 , n29751 );
xor ( n29753 , n29741 , n29752 );
xor ( n29754 , RI19abcbe8_2361 , RI174b6238_848);
not ( n10883 , n27689 );
and ( n10884 , n10883 , RI174b6238_848);
and ( n10885 , n29754 , n27689 );
or ( n29755 , n10884 , n10885 );
xor ( n29756 , n29755 , n29375 );
xor ( n29757 , RI19a95930_2643 , RI1747c1a0_1131);
not ( n10886 , n27689 );
and ( n10887 , n10886 , RI1747c1a0_1131);
and ( n10888 , n29757 , n27689 );
or ( n29758 , n10887 , n10888 );
xor ( n29759 , RI19ac5720_2288 , RI174cbf70_776);
not ( n10889 , n27689 );
and ( n10890 , n10889 , RI174cbf70_776);
and ( n10891 , n29759 , n27689 );
or ( n29760 , n10890 , n10891 );
xor ( n29761 , n29758 , n29760 );
buf ( n29762 , RI17396e80_2020);
xor ( n29763 , n29761 , n29762 );
buf ( n29764 , RI173dfb70_1665);
xor ( n29765 , n29763 , n29764 );
buf ( n29766 , RI17457648_1310);
xor ( n29767 , n29765 , n29766 );
xor ( n29768 , n29756 , n29767 );
not ( n29769 , n29768 );
buf ( n29770 , RI17390f58_2049);
xor ( n29771 , RI19a8ed60_2691 , RI17467638_1232);
not ( n10892 , n27689 );
and ( n10893 , n10892 , RI17467638_1232);
and ( n10894 , n29771 , n27689 );
or ( n29772 , n10893 , n10894 );
xor ( n29773 , RI19abf870_2336 , RI174b0310_877);
not ( n10895 , n27689 );
and ( n10896 , n10895 , RI174b0310_877);
and ( n10897 , n29773 , n27689 );
or ( n29774 , n10896 , n10897 );
xor ( n29775 , n29772 , n29774 );
buf ( n29776 , RI17341a70_2121);
xor ( n29777 , n29775 , n29776 );
buf ( n29778 , RI173caff0_1766);
xor ( n29779 , n29777 , n29778 );
buf ( n29780 , RI17414028_1410);
xor ( n29781 , n29779 , n29780 );
xor ( n29782 , n29770 , n29781 );
xor ( n29783 , RI19aa27e8_2549 , RI17484b70_1089);
not ( n10898 , n27689 );
and ( n10899 , n10898 , RI17484b70_1089);
and ( n10900 , n29783 , n27689 );
or ( n29784 , n10899 , n10900 );
xor ( n29785 , RI19a838e8_2769 , RI1750a490_734);
not ( n10901 , n27689 );
and ( n10902 , n10901 , RI1750a490_734);
and ( n10903 , n29785 , n27689 );
or ( n29786 , n10902 , n10903 );
xor ( n29787 , n29784 , n29786 );
buf ( n29788 , RI1739f850_1978);
xor ( n29789 , n29787 , n29788 );
buf ( n29790 , RI173e8888_1622);
xor ( n29791 , n29789 , n29790 );
buf ( n29792 , RI17460360_1267);
xor ( n29793 , n29791 , n29792 );
xor ( n29794 , n29782 , n29793 );
and ( n29795 , n29769 , n29794 );
xor ( n29796 , n29753 , n29795 );
xor ( n29797 , n29728 , n29796 );
xor ( n29798 , RI19aa3058_2545 , RI17481d80_1103);
not ( n10904 , n27689 );
and ( n10905 , n10904 , RI17481d80_1103);
and ( n10906 , n29798 , n27689 );
or ( n29799 , n10905 , n10906 );
xor ( n29800 , n29799 , n27807 );
xor ( n29801 , n29800 , n27819 );
xor ( n29802 , RI19a23510_2794 , RI1751a660_684);
not ( n10907 , n27689 );
and ( n10908 , n10907 , RI1751a660_684);
and ( n10909 , n29802 , n27689 );
or ( n29803 , n10908 , n10909 );
xor ( n29804 , n29803 , n29332 );
xor ( n29805 , RI19ab8958_2391 , RI1749d878_968);
not ( n10910 , n27689 );
and ( n10911 , n10910 , RI1749d878_968);
and ( n10912 , n29805 , n27689 );
or ( n29806 , n10911 , n10912 );
buf ( n29807 , RI17531478_613);
xor ( n29808 , n29806 , n29807 );
buf ( n29809 , RI173b88a0_1856);
xor ( n29810 , n29808 , n29809 );
buf ( n29811 , RI17401590_1501);
xor ( n29812 , n29810 , n29811 );
buf ( n29813 , RI173db688_1686);
xor ( n29814 , n29812 , n29813 );
xor ( n29815 , n29804 , n29814 );
not ( n29816 , n29815 );
xor ( n29817 , RI19aa6d48_2517 , RI17499a20_987);
not ( n10913 , n27689 );
and ( n10914 , n10913 , RI17499a20_987);
and ( n10915 , n29817 , n27689 );
or ( n29818 , n10914 , n10915 );
xor ( n29819 , RI19a88028_2738 , RI1752b280_632);
not ( n10916 , n27689 );
and ( n10917 , n10916 , RI1752b280_632);
and ( n10918 , n29819 , n27689 );
or ( n29820 , n10917 , n10918 );
xor ( n29821 , n29818 , n29820 );
buf ( n29822 , RI173b4700_1876);
xor ( n29823 , n29821 , n29822 );
buf ( n29824 , RI173fd738_1520);
xor ( n29825 , n29823 , n29824 );
buf ( n29826 , RI173b4a48_1875);
xor ( n29827 , n29825 , n29826 );
xor ( n29828 , n29057 , n29827 );
xor ( n29829 , RI19a894c8_2729 , RI1746e280_1199);
not ( n10919 , n27689 );
and ( n10920 , n10919 , RI1746e280_1199);
and ( n10921 , n29829 , n27689 );
or ( n29830 , n10920 , n10921 );
xor ( n29831 , RI19abaf50_2374 , RI174b6f58_844);
not ( n10922 , n27689 );
and ( n10923 , n10922 , RI174b6f58_844);
and ( n10924 , n29831 , n27689 );
or ( n29832 , n10923 , n10924 );
xor ( n29833 , n29830 , n29832 );
buf ( n29834 , RI173599e0_2088);
xor ( n29835 , n29833 , n29834 );
buf ( n29836 , RI173d1f98_1732);
xor ( n29837 , n29835 , n29836 );
buf ( n29838 , RI17449a70_1377);
xor ( n29839 , n29837 , n29838 );
xor ( n29840 , n29828 , n29839 );
and ( n29841 , n29816 , n29840 );
xor ( n29842 , n29801 , n29841 );
xor ( n29843 , n29797 , n29842 );
xor ( n29844 , n29659 , n29843 );
xor ( n29845 , RI19a9f908_2572 , RI174872d0_1077);
not ( n10925 , n27689 );
and ( n10926 , n10925 , RI174872d0_1077);
and ( n10927 , n29845 , n27689 );
or ( n29846 , n10926 , n10927 );
xor ( n29847 , RI19ace618_2222 , RI1750e270_722);
not ( n10928 , n27689 );
and ( n10929 , n10928 , RI1750e270_722);
and ( n10930 , n29847 , n27689 );
or ( n29848 , n10929 , n10930 );
xor ( n29849 , n29846 , n29848 );
buf ( n29850 , RI173a22f8_1965);
xor ( n29851 , n29849 , n29850 );
buf ( n29852 , RI173eafe8_1610);
xor ( n29853 , n29851 , n29852 );
buf ( n29854 , RI17473140_1175);
xor ( n29855 , n29853 , n29854 );
xor ( n29856 , n28197 , n29855 );
xor ( n29857 , n29856 , n29079 );
not ( n29858 , n29857 );
and ( n29859 , n29858 , n27792 );
xor ( n29860 , n27765 , n29859 );
buf ( n29861 , RI173406c0_2127);
xor ( n29862 , n29861 , n28852 );
xor ( n29863 , RI19a9a868_2608 , RI17474b80_1167);
not ( n10931 , n27689 );
and ( n10932 , n10931 , RI17474b80_1167);
and ( n10933 , n29863 , n27689 );
or ( n29864 , n10932 , n10933 );
xor ( n29865 , RI19aca040_2255 , RI174c0af8_811);
not ( n10934 , n27689 );
and ( n10935 , n10934 , RI174c0af8_811);
and ( n10936 , n29865 , n27689 );
or ( n29866 , n10935 , n10936 );
xor ( n29867 , n29864 , n29866 );
buf ( n29868 , RI1738fba8_2055);
xor ( n29869 , n29867 , n29868 );
buf ( n29870 , RI173d8898_1700);
xor ( n29871 , n29869 , n29870 );
buf ( n29872 , RI17450370_1345);
xor ( n29873 , n29871 , n29872 );
xor ( n29874 , n29862 , n29873 );
xor ( n29875 , n28540 , n28125 );
xor ( n29876 , n29875 , n28137 );
not ( n29877 , n29876 );
and ( n29878 , n29877 , n27820 );
xor ( n29879 , n29874 , n29878 );
xor ( n29880 , n29860 , n29879 );
xor ( n29881 , n28834 , n28569 );
buf ( n29882 , RI17337318_2172);
xor ( n29883 , n29730 , n29882 );
buf ( n29884 , RI173c0898_1817);
xor ( n29885 , n29883 , n29884 );
buf ( n29886 , RI17409588_1462);
xor ( n29887 , n29885 , n29886 );
buf ( n29888 , RI1745a0f0_1297);
xor ( n29889 , n29887 , n29888 );
xor ( n29890 , n29881 , n29889 );
buf ( n29891 , RI174053e8_1482);
xor ( n29892 , n29891 , n28291 );
xor ( n29893 , n29892 , n29781 );
not ( n29894 , n29893 );
and ( n29895 , n29894 , n27898 );
xor ( n29896 , n29890 , n29895 );
xor ( n29897 , n29880 , n29896 );
buf ( n29898 , RI173912a0_2048);
xor ( n29899 , n29898 , n28339 );
xor ( n29900 , RI19aa2c20_2547 , RI17484eb8_1088);
not ( n10937 , n27689 );
and ( n10938 , n10937 , RI17484eb8_1088);
and ( n10939 , n29900 , n27689 );
or ( n29901 , n10938 , n10939 );
xor ( n29902 , RI19a83d20_2767 , RI1750a9b8_733);
not ( n10940 , n27689 );
and ( n10941 , n10940 , RI1750a9b8_733);
and ( n10942 , n29902 , n27689 );
or ( n29903 , n10941 , n10942 );
xor ( n29904 , n29901 , n29903 );
buf ( n29905 , RI1739fb98_1977);
xor ( n29906 , n29904 , n29905 );
buf ( n29907 , RI173e8bd0_1621);
xor ( n29908 , n29906 , n29907 );
buf ( n29909 , RI174606a8_1266);
xor ( n29910 , n29908 , n29909 );
xor ( n29911 , n29899 , n29910 );
buf ( n29912 , RI173e9c38_1616);
xor ( n29913 , RI19a97460_2631 , RI174772e0_1155);
not ( n10943 , n27689 );
and ( n10944 , n10943 , RI174772e0_1155);
and ( n10945 , n29913 , n27689 );
or ( n29914 , n10944 , n10945 );
xor ( n29915 , RI19ac7250_2276 , RI174c48d8_799);
not ( n10946 , n27689 );
and ( n10947 , n10946 , RI174c48d8_799);
and ( n10948 , n29915 , n27689 );
or ( n29916 , n10947 , n10948 );
xor ( n29917 , n29914 , n29916 );
buf ( n29918 , RI17392308_2043);
xor ( n29919 , n29917 , n29918 );
buf ( n29920 , RI173daff8_1688);
xor ( n29921 , n29919 , n29920 );
buf ( n29922 , RI17452ad0_1333);
xor ( n29923 , n29921 , n29922 );
xor ( n29924 , n29912 , n29923 );
xor ( n29925 , RI19aab0c8_2488 , RI17494b60_1011);
not ( n10949 , n27689 );
and ( n10950 , n10949 , RI17494b60_1011);
and ( n10951 , n29925 , n27689 );
or ( n29926 , n10950 , n10951 );
xor ( n29927 , RI19aa8f80_2503 , RI175236c0_656);
not ( n10952 , n27689 );
and ( n10953 , n10952 , RI175236c0_656);
and ( n10954 , n29927 , n27689 );
or ( n29928 , n10953 , n10954 );
xor ( n29929 , n29926 , n29928 );
buf ( n29930 , RI173af840_1900);
xor ( n29931 , n29929 , n29930 );
buf ( n29932 , RI173f8530_1545);
xor ( n29933 , n29931 , n29932 );
buf ( n29934 , RI17342100_2119);
xor ( n29935 , n29933 , n29934 );
xor ( n29936 , n29924 , n29935 );
not ( n29937 , n29936 );
and ( n29938 , n29937 , n27976 );
xor ( n29939 , n29911 , n29938 );
xor ( n29940 , n29897 , n29939 );
buf ( n29941 , RI173c3688_1803);
xor ( n29942 , RI19aa7090_2516 , RI1749a0b0_985);
not ( n10955 , n27689 );
and ( n10956 , n10955 , RI1749a0b0_985);
and ( n10957 , n29942 , n27689 );
or ( n29943 , n10956 , n10957 );
xor ( n29944 , RI19a88208_2737 , RI1752bcd0_630);
not ( n10958 , n27689 );
and ( n10959 , n10958 , RI1752bcd0_630);
and ( n10960 , n29944 , n27689 );
or ( n29945 , n10959 , n10960 );
xor ( n29946 , n29943 , n29945 );
buf ( n29947 , RI173b4d90_1874);
xor ( n29948 , n29946 , n29947 );
buf ( n29949 , RI173fddc8_1518);
xor ( n29950 , n29948 , n29949 );
buf ( n29951 , RI173b71a8_1863);
xor ( n29952 , n29950 , n29951 );
xor ( n29953 , n29941 , n29952 );
xor ( n29954 , RI19a89720_2728 , RI1746e5c8_1198);
not ( n10961 , n27689 );
and ( n10962 , n10961 , RI1746e5c8_1198);
and ( n10963 , n29954 , n27689 );
or ( n29955 , n10962 , n10963 );
xor ( n29956 , RI19abb298_2373 , RI174b72a0_843);
not ( n10964 , n27689 );
and ( n10965 , n10964 , RI174b72a0_843);
and ( n10966 , n29956 , n27689 );
or ( n29957 , n10965 , n10966 );
xor ( n29958 , n29955 , n29957 );
buf ( n29959 , RI173892a8_2087);
xor ( n29960 , n29958 , n29959 );
buf ( n29961 , RI173d22e0_1731);
xor ( n29962 , n29960 , n29961 );
buf ( n29963 , RI17449db8_1376);
xor ( n29964 , n29962 , n29963 );
xor ( n29965 , n29953 , n29964 );
xor ( n29966 , RI19ab16f8_2443 , RI174a9038_912);
not ( n10967 , n27689 );
and ( n10968 , n10967 , RI174a9038_912);
and ( n10969 , n29966 , n27689 );
or ( n29967 , n10968 , n10969 );
buf ( n29968 , RI1733a798_2156);
xor ( n29969 , n29967 , n29968 );
buf ( n29970 , RI173c3d18_1801);
xor ( n29971 , n29969 , n29970 );
buf ( n29972 , RI1740ca08_1446);
xor ( n29973 , n29971 , n29972 );
buf ( n29974 , RI173fb320_1531);
xor ( n29975 , n29973 , n29974 );
xor ( n29976 , n28447 , n29975 );
xor ( n29977 , n29976 , n28759 );
not ( n29978 , n29977 );
and ( n29979 , n29978 , n28056 );
xor ( n29980 , n29965 , n29979 );
xor ( n29981 , n29940 , n29980 );
xor ( n29982 , n29844 , n29981 );
buf ( n29983 , RI173413e0_2123);
xor ( n29984 , n29983 , n28956 );
xor ( n29985 , RI19a98ae0_2621 , RI17475be8_1162);
not ( n10970 , n27689 );
and ( n10971 , n10970 , RI17475be8_1162);
and ( n10972 , n29985 , n27689 );
or ( n29986 , n10971 , n10972 );
xor ( n29987 , RI19ac8510_2267 , RI174c24c0_806);
not ( n10973 , n27689 );
and ( n10974 , n10973 , RI174c24c0_806);
and ( n10975 , n29987 , n27689 );
or ( n29988 , n10974 , n10975 );
xor ( n29989 , n29986 , n29988 );
buf ( n29990 , RI17390c10_2050);
xor ( n29991 , n29989 , n29990 );
buf ( n29992 , RI173d9900_1695);
xor ( n29993 , n29991 , n29992 );
buf ( n29994 , RI174513d8_1340);
xor ( n29995 , n29993 , n29994 );
xor ( n29996 , n29984 , n29995 );
xor ( n29997 , RI19a92708_2665 , RI174620e8_1258);
not ( n10976 , n27689 );
and ( n10977 , n10976 , RI174620e8_1258);
and ( n10978 , n29997 , n27689 );
or ( n29998 , n10977 , n10978 );
xor ( n29999 , RI19ac2a98_2309 , RI174aadc0_903);
not ( n10979 , n27689 );
and ( n10980 , n10979 , RI174aadc0_903);
and ( n10981 , n29999 , n27689 );
or ( n30000 , n10980 , n10981 );
xor ( n30001 , n29998 , n30000 );
buf ( n30002 , RI1733c520_2147);
xor ( n30003 , n30001 , n30002 );
buf ( n30004 , RI173c5aa0_1792);
xor ( n30005 , n30003 , n30004 );
buf ( n30006 , RI1740e790_1437);
xor ( n30007 , n30005 , n30006 );
xor ( n30008 , n28901 , n30007 );
xor ( n30009 , RI19aa62f8_2521 , RI1747f620_1115);
not ( n10982 , n27689 );
and ( n10983 , n10982 , RI1747f620_1115);
and ( n10984 , n30009 , n27689 );
or ( n30010 , n10983 , n10984 );
xor ( n30011 , n30010 , n28636 );
buf ( n30012 , RI1739a300_2004);
xor ( n30013 , n30011 , n30012 );
buf ( n30014 , RI173e2ff0_1649);
xor ( n30015 , n30013 , n30014 );
buf ( n30016 , RI1745ae10_1293);
xor ( n30017 , n30015 , n30016 );
xor ( n30018 , n30008 , n30017 );
not ( n30019 , n30018 );
xor ( n30020 , n29437 , n27712 );
xor ( n30021 , RI19aadfa8_2468 , RI17491a28_1026);
not ( n10985 , n27689 );
and ( n10986 , n10985 , RI17491a28_1026);
and ( n10987 , n30021 , n27689 );
or ( n30022 , n10986 , n10987 );
xor ( n30023 , RI19ac36c8_2303 , RI1751e968_671);
not ( n10988 , n27689 );
and ( n10989 , n10988 , RI1751e968_671);
and ( n10990 , n30023 , n27689 );
or ( n30024 , n10989 , n10990 );
xor ( n30025 , n30022 , n30024 );
buf ( n30026 , RI173ac708_1915);
xor ( n30027 , n30025 , n30026 );
xor ( n30028 , n30027 , n28841 );
buf ( n30029 , RI1751d4c8_675);
xor ( n30030 , n30028 , n30029 );
xor ( n30031 , n30020 , n30030 );
and ( n30032 , n30019 , n30031 );
xor ( n30033 , n29996 , n30032 );
xor ( n30034 , RI19a92528_2666 , RI17461da0_1259);
not ( n10991 , n27689 );
and ( n10992 , n10991 , RI17461da0_1259);
and ( n10993 , n30034 , n27689 );
or ( n30035 , n10992 , n10993 );
xor ( n30036 , RI19ac2840_2310 , RI174aaa78_904);
not ( n10994 , n27689 );
and ( n10995 , n10994 , RI174aaa78_904);
and ( n10996 , n30036 , n27689 );
or ( n30037 , n10995 , n10996 );
xor ( n30038 , n30035 , n30037 );
xor ( n30039 , n30038 , n28882 );
buf ( n30040 , RI173c5758_1793);
xor ( n30041 , n30039 , n30040 );
buf ( n30042 , RI1740e448_1438);
xor ( n30043 , n30041 , n30042 );
xor ( n30044 , n28498 , n30043 );
xor ( n30045 , RI19aa6190_2522 , RI1747f2d8_1116);
not ( n10997 , n27689 );
and ( n10998 , n10997 , RI1747f2d8_1116);
and ( n10999 , n30045 , n27689 );
or ( n30046 , n10998 , n10999 );
xor ( n30047 , n30046 , n29279 );
buf ( n30048 , RI17399fb8_2005);
xor ( n30049 , n30047 , n30048 );
buf ( n30050 , RI173e2ca8_1650);
xor ( n30051 , n30049 , n30050 );
buf ( n30052 , RI1745aac8_1294);
xor ( n30053 , n30051 , n30052 );
xor ( n30054 , n30044 , n30053 );
xor ( n30055 , n28257 , n29270 );
xor ( n30056 , RI19ab01e0_2453 , RI1748d540_1047);
not ( n11000 , n27689 );
and ( n11001 , n11000 , RI1748d540_1047);
and ( n11002 , n30056 , n27689 );
or ( n30057 , n11001 , n11002 );
xor ( n30058 , RI19a94df0_2648 , RI17518248_691);
not ( n11003 , n27689 );
and ( n11004 , n11003 , RI17518248_691);
and ( n11005 , n30058 , n27689 );
or ( n30059 , n11004 , n11005 );
xor ( n30060 , n30057 , n30059 );
buf ( n30061 , RI173a8568_1935);
xor ( n30062 , n30060 , n30061 );
buf ( n30063 , RI173f1258_1580);
xor ( n30064 , n30062 , n30063 );
buf ( n30065 , RI174b09a0_875);
xor ( n30066 , n30064 , n30065 );
xor ( n30067 , n30055 , n30066 );
not ( n30068 , n30067 );
xor ( n30069 , n28836 , n28569 );
xor ( n30070 , n30069 , n29889 );
and ( n30071 , n30068 , n30070 );
xor ( n30072 , n30054 , n30071 );
buf ( n30073 , RI17336940_2175);
xor ( n30074 , n30073 , n28595 );
xor ( n30075 , n30074 , n28519 );
not ( n30076 , n29996 );
and ( n30077 , n30076 , n30018 );
xor ( n30078 , n30075 , n30077 );
xor ( n30079 , n30072 , n30078 );
xor ( n30080 , RI19a98f90_2619 , RI17476278_1160);
not ( n11006 , n27689 );
and ( n11007 , n11006 , RI17476278_1160);
and ( n11008 , n30080 , n27689 );
or ( n30081 , n11007 , n11008 );
xor ( n30082 , RI19ac89c0_2265 , RI174c2f10_804);
not ( n11009 , n27689 );
and ( n11010 , n11009 , RI174c2f10_804);
and ( n11011 , n30082 , n27689 );
or ( n30083 , n11010 , n11011 );
xor ( n30084 , n30081 , n30083 );
xor ( n30085 , n30084 , n29898 );
buf ( n30086 , RI173d9f90_1693);
xor ( n30087 , n30085 , n30086 );
buf ( n30088 , RI17451a68_1338);
xor ( n30089 , n30087 , n30088 );
xor ( n30090 , n29786 , n30089 );
xor ( n30091 , RI19aacdd8_2476 , RI17493af8_1016);
not ( n11012 , n27689 );
and ( n11013 , n11012 , RI17493af8_1016);
and ( n11014 , n30091 , n27689 );
or ( n30092 , n11013 , n11014 );
xor ( n30093 , RI19ab9df8_2381 , RI17521cf8_661);
not ( n11015 , n27689 );
and ( n11016 , n11015 , RI17521cf8_661);
and ( n11017 , n30093 , n27689 );
or ( n30094 , n11016 , n11017 );
xor ( n30095 , n30092 , n30094 );
buf ( n30096 , RI173ae7d8_1905);
xor ( n30097 , n30095 , n30096 );
buf ( n30098 , RI173f74c8_1550);
xor ( n30099 , n30097 , n30098 );
buf ( n30100 , RI17336c88_2174);
xor ( n30101 , n30099 , n30100 );
xor ( n30102 , n30090 , n30101 );
buf ( n30103 , RI173b2978_1885);
xor ( n30104 , RI19a9e8a0_2580 , RI17489058_1068);
not ( n11018 , n27689 );
and ( n11019 , n11018 , RI17489058_1068);
and ( n11020 , n30104 , n27689 );
or ( n30105 , n11019 , n11020 );
xor ( n30106 , RI19acd358_2230 , RI175110d8_713);
not ( n11021 , n27689 );
and ( n11022 , n11021 , RI175110d8_713);
and ( n11023 , n30106 , n27689 );
or ( n30107 , n11022 , n11023 );
xor ( n30108 , n30105 , n30107 );
buf ( n30109 , RI173a4080_1956);
xor ( n30110 , n30108 , n30109 );
buf ( n30111 , RI173ecd70_1601);
xor ( n30112 , n30110 , n30111 );
buf ( n30113 , RI17485548_1086);
xor ( n30114 , n30112 , n30113 );
xor ( n30115 , n30103 , n30114 );
xor ( n30116 , RI19ab2328_2438 , RI174a68d8_924);
not ( n11024 , n27689 );
and ( n11025 , n11024 , RI174a68d8_924);
and ( n11026 , n30116 , n27689 );
or ( n30117 , n11025 , n11026 );
buf ( n30118 , RI17338038_2168);
xor ( n30119 , n30117 , n30118 );
buf ( n30120 , RI173c15b8_1813);
xor ( n30121 , n30119 , n30120 );
buf ( n30122 , RI1740a2a8_1458);
xor ( n30123 , n30121 , n30122 );
buf ( n30124 , RI17477970_1153);
xor ( n30125 , n30123 , n30124 );
xor ( n30126 , n30115 , n30125 );
not ( n30127 , n30126 );
buf ( n30128 , RI17406108_1478);
xor ( n30129 , RI19aad120_2475 , RI17493e40_1015);
not ( n11027 , n27689 );
and ( n11028 , n11027 , RI17493e40_1015);
and ( n11029 , n30129 , n27689 );
or ( n30130 , n11028 , n11029 );
xor ( n30131 , RI19abba90_2370 , RI17522220_660);
not ( n11030 , n27689 );
and ( n11031 , n11030 , RI17522220_660);
and ( n11032 , n30131 , n27689 );
or ( n30132 , n11031 , n11032 );
xor ( n30133 , n30130 , n30132 );
buf ( n30134 , RI173aeb20_1904);
xor ( n30135 , n30133 , n30134 );
buf ( n30136 , RI173f7810_1549);
xor ( n30137 , n30135 , n30136 );
buf ( n30138 , RI173390a0_2163);
xor ( n30139 , n30137 , n30138 );
xor ( n30140 , n30128 , n30139 );
xor ( n30141 , RI19a8cd80_2705 , RI174686a0_1227);
not ( n11033 , n27689 );
and ( n11034 , n11033 , RI174686a0_1227);
and ( n11035 , n30141 , n27689 );
or ( n30142 , n11034 , n11035 );
xor ( n30143 , RI19abdf98_2350 , RI174b1378_872);
not ( n11036 , n27689 );
and ( n11037 , n11036 , RI174b1378_872);
and ( n11038 , n30143 , n27689 );
or ( n30144 , n11037 , n11038 );
xor ( n30145 , n30142 , n30144 );
buf ( n30146 , RI17342ad8_2116);
xor ( n30147 , n30145 , n30146 );
buf ( n30148 , RI173cc058_1761);
xor ( n30149 , n30147 , n30148 );
buf ( n30150 , RI17415090_1405);
xor ( n30151 , n30149 , n30150 );
xor ( n30152 , n30140 , n30151 );
and ( n30153 , n30127 , n30152 );
xor ( n30154 , n30102 , n30153 );
xor ( n30155 , n30079 , n30154 );
xor ( n30156 , RI19ab1518_2444 , RI174a8cf0_913);
not ( n11039 , n27689 );
and ( n11040 , n11039 , RI174a8cf0_913);
and ( n11041 , n30156 , n27689 );
or ( n30157 , n11040 , n11041 );
buf ( n30158 , RI1733a450_2157);
xor ( n30159 , n30157 , n30158 );
xor ( n30160 , n30159 , n28427 );
buf ( n30161 , RI1740c6c0_1447);
xor ( n30162 , n30160 , n30161 );
buf ( n30163 , RI173e46e8_1642);
xor ( n30164 , n30162 , n30163 );
xor ( n30165 , n29957 , n30164 );
xor ( n30166 , n30165 , n29490 );
buf ( n30167 , RI17391fc0_2044);
xor ( n30168 , RI19a8cfd8_2704 , RI174689e8_1226);
not ( n11042 , n27689 );
and ( n11043 , n11042 , RI174689e8_1226);
and ( n11044 , n30168 , n27689 );
or ( n30169 , n11043 , n11044 );
xor ( n30170 , RI19abe100_2349 , RI174b16c0_871);
not ( n11045 , n27689 );
and ( n11046 , n11045 , RI174b16c0_871);
and ( n11047 , n30170 , n27689 );
or ( n30171 , n11046 , n11047 );
xor ( n30172 , n30169 , n30171 );
buf ( n30173 , RI17342e20_2115);
xor ( n30174 , n30172 , n30173 );
buf ( n30175 , RI173cc3a0_1760);
xor ( n30176 , n30174 , n30175 );
buf ( n30177 , RI174153d8_1404);
xor ( n30178 , n30176 , n30177 );
xor ( n30179 , n30167 , n30178 );
xor ( n30180 , RI19aa0f10_2561 , RI17485f20_1083);
not ( n11048 , n27689 );
and ( n11049 , n11048 , RI17485f20_1083);
and ( n11050 , n30180 , n27689 );
or ( n30181 , n11049 , n11050 );
xor ( n30182 , RI19acfd88_2212 , RI1750c380_728);
not ( n11051 , n27689 );
and ( n11052 , n11051 , RI1750c380_728);
and ( n11053 , n30182 , n27689 );
or ( n30183 , n11052 , n11053 );
xor ( n30184 , n30181 , n30183 );
buf ( n30185 , RI173a0f48_1971);
xor ( n30186 , n30184 , n30185 );
xor ( n30187 , n30186 , n29912 );
buf ( n30188 , RI174658b0_1241);
xor ( n30189 , n30187 , n30188 );
xor ( n30190 , n30179 , n30189 );
not ( n30191 , n30190 );
buf ( n30192 , RI173ea958_1612);
xor ( n30193 , n30192 , n27897 );
xor ( n30194 , n30193 , n27858 );
and ( n30195 , n30191 , n30194 );
xor ( n30196 , n30166 , n30195 );
xor ( n30197 , n30155 , n30196 );
xor ( n30198 , RI19aa5218_2529 , RI174816f0_1105);
not ( n11054 , n27689 );
and ( n11055 , n11054 , RI174816f0_1105);
and ( n11056 , n30198 , n27689 );
or ( n30199 , n11055 , n11056 );
xor ( n30200 , RI19a864f8_2750 , RI17503398_750);
not ( n11057 , n27689 );
and ( n11058 , n11057 , RI17503398_750);
and ( n11059 , n30200 , n27689 );
or ( n30201 , n11058 , n11059 );
xor ( n30202 , n30199 , n30201 );
buf ( n30203 , RI1739c3d0_1994);
xor ( n30204 , n30202 , n30203 );
xor ( n30205 , n30204 , n29550 );
buf ( n30206 , RI1745cee0_1283);
xor ( n30207 , n30205 , n30206 );
xor ( n30208 , n28859 , n30207 );
xor ( n30209 , RI19ab9498_2386 , RI1749ec28_962);
not ( n11060 , n27689 );
and ( n11061 , n11060 , RI1749ec28_962);
and ( n11062 , n30209 , n27689 );
or ( n30210 , n11061 , n11062 );
buf ( n30211 , RI17533368_607);
xor ( n30212 , n30210 , n30211 );
buf ( n30213 , RI173b9c50_1850);
xor ( n30214 , n30212 , n30213 );
buf ( n30215 , RI17402940_1495);
xor ( n30216 , n30214 , n30215 );
buf ( n30217 , RI173e6e48_1630);
xor ( n30218 , n30216 , n30217 );
xor ( n30219 , n30208 , n30218 );
buf ( n30220 , RI173c43a8_1799);
xor ( n30221 , n30220 , n28771 );
xor ( n30222 , n30221 , n27726 );
not ( n30223 , n30222 );
xor ( n30224 , RI19ab96f0_2385 , RI1749b460_979);
not ( n11063 , n27689 );
and ( n11064 , n11063 , RI1749b460_979);
and ( n11065 , n30224 , n27689 );
or ( n30225 , n11064 , n11065 );
buf ( n30226 , RI1752dbc0_624);
xor ( n30227 , n30225 , n30226 );
buf ( n30228 , RI173b6140_1868);
xor ( n30229 , n30227 , n30228 );
buf ( n30230 , RI173ff178_1512);
xor ( n30231 , n30229 , n30230 );
buf ( n30232 , RI173c4a38_1797);
xor ( n30233 , n30231 , n30232 );
xor ( n30234 , n28122 , n30233 );
xor ( n30235 , RI19a9c1b8_2597 , RI1746fcc0_1191);
not ( n11066 , n27689 );
and ( n11067 , n11066 , RI1746fcc0_1191);
and ( n11068 , n30235 , n27689 );
or ( n30236 , n11067 , n11068 );
xor ( n30237 , RI19acb4e0_2245 , RI174b8a10_836);
not ( n11069 , n27689 );
and ( n11070 , n11069 , RI174b8a10_836);
and ( n11071 , n30237 , n27689 );
or ( n30238 , n11070 , n11071 );
xor ( n30239 , n30236 , n30238 );
buf ( n30240 , RI1738ace8_2079);
xor ( n30241 , n30239 , n30240 );
xor ( n30242 , n30241 , n28239 );
xor ( n30243 , n30242 , n29604 );
xor ( n30244 , n30234 , n30243 );
and ( n30245 , n30223 , n30244 );
xor ( n30246 , n30219 , n30245 );
xor ( n30247 , n30197 , n30246 );
xor ( n30248 , n30033 , n30247 );
xor ( n30249 , n29737 , n28304 );
xor ( n30250 , n30249 , n28313 );
buf ( n30251 , RI1744a100_1375);
xor ( n30252 , n30251 , n28800 );
xor ( n30253 , n30252 , n28812 );
not ( n30254 , n30253 );
xor ( n30255 , RI19a8e220_2696 , RI17466918_1236);
not ( n11072 , n27689 );
and ( n11073 , n11072 , RI17466918_1236);
and ( n11074 , n30255 , n27689 );
or ( n30256 , n11073 , n11074 );
xor ( n30257 , n30256 , n29134 );
xor ( n30258 , n30257 , n27936 );
and ( n30259 , n30254 , n30258 );
xor ( n30260 , n30250 , n30259 );
xor ( n30261 , RI19a92960_2664 , RI17462430_1257);
not ( n11075 , n27689 );
and ( n11076 , n11075 , RI17462430_1257);
and ( n11077 , n30261 , n27689 );
or ( n30262 , n11076 , n11077 );
xor ( n30263 , RI19ac2cf0_2308 , RI174ab108_902);
not ( n11078 , n27689 );
and ( n11079 , n11078 , RI174ab108_902);
and ( n11080 , n30263 , n27689 );
or ( n30264 , n11079 , n11080 );
xor ( n30265 , n30262 , n30264 );
buf ( n30266 , RI1733c868_2146);
xor ( n30267 , n30265 , n30266 );
buf ( n30268 , RI173c5de8_1791);
xor ( n30269 , n30267 , n30268 );
buf ( n30270 , RI1740ead8_1436);
xor ( n30271 , n30269 , n30270 );
xor ( n30272 , n28644 , n30271 );
xor ( n30273 , RI19aa6640_2520 , RI1747f968_1114);
not ( n11081 , n27689 );
and ( n11082 , n11081 , RI1747f968_1114);
and ( n11083 , n30273 , n27689 );
or ( n30274 , n11082 , n11083 );
xor ( n30275 , RI19a87920_2741 , RI17500530_759);
not ( n11084 , n27689 );
and ( n11085 , n11084 , RI17500530_759);
and ( n11086 , n30275 , n27689 );
or ( n30276 , n11085 , n11086 );
xor ( n30277 , n30274 , n30276 );
buf ( n30278 , RI1739a648_2003);
xor ( n30279 , n30277 , n30278 );
buf ( n30280 , RI173e3338_1648);
xor ( n30281 , n30279 , n30280 );
buf ( n30282 , RI1745b158_1292);
xor ( n30283 , n30281 , n30282 );
xor ( n30284 , n30272 , n30283 );
xor ( n30285 , RI19a9a3b8_2610 , RI174744f0_1169);
not ( n11087 , n27689 );
and ( n11088 , n11087 , RI174744f0_1169);
and ( n11089 , n30285 , n27689 );
or ( n30286 , n11088 , n11089 );
xor ( n30287 , RI19ac9b90_2257 , RI174c00a8_813);
not ( n11090 , n27689 );
and ( n11091 , n11090 , RI174c00a8_813);
and ( n11092 , n30287 , n27689 );
or ( n30288 , n11091 , n11092 );
xor ( n30289 , n30286 , n30288 );
buf ( n30290 , RI1738f518_2057);
xor ( n30291 , n30289 , n30290 );
buf ( n30292 , RI173d8208_1702);
xor ( n30293 , n30291 , n30292 );
xor ( n30294 , n30293 , n28032 );
xor ( n30295 , n27920 , n30294 );
xor ( n30296 , RI19aae110_2467 , RI17491d70_1025);
not ( n11093 , n27689 );
and ( n11094 , n11093 , RI17491d70_1025);
and ( n11095 , n30296 , n27689 );
or ( n30297 , n11094 , n11095 );
xor ( n30298 , RI19ac4f28_2292 , RI1751ee90_670);
not ( n11096 , n27689 );
and ( n11097 , n11096 , RI1751ee90_670);
and ( n11098 , n30298 , n27689 );
or ( n30299 , n11097 , n11098 );
xor ( n30300 , n30297 , n30299 );
buf ( n30301 , RI173aca50_1914);
xor ( n30302 , n30300 , n30301 );
buf ( n30303 , RI173f5740_1559);
xor ( n30304 , n30302 , n30303 );
buf ( n30305 , RI17520d80_664);
xor ( n30306 , n30304 , n30305 );
xor ( n30307 , n30295 , n30306 );
not ( n30308 , n30307 );
xor ( n30309 , RI19aa8bc0_2505 , RI174989b8_992);
not ( n11099 , n27689 );
and ( n11100 , n11099 , RI174989b8_992);
and ( n11101 , n30309 , n27689 );
or ( n30310 , n11100 , n11101 );
xor ( n30311 , RI19a9f188_2576 , RI1748a0c0_1063);
not ( n11102 , n27689 );
and ( n11103 , n11102 , RI1748a0c0_1063);
and ( n11104 , n30311 , n27689 );
or ( n30312 , n11103 , n11104 );
xor ( n30313 , RI19acdcb8_2226 , RI17512fc8_707);
not ( n11105 , n27689 );
and ( n11106 , n11105 , RI17512fc8_707);
and ( n11107 , n30313 , n27689 );
or ( n30314 , n11106 , n11107 );
xor ( n30315 , n30312 , n30314 );
buf ( n30316 , RI173a50e8_1951);
xor ( n30317 , n30315 , n30316 );
buf ( n30318 , RI173eddd8_1596);
xor ( n30319 , n30317 , n30318 );
buf ( n30320 , RI1748e8f0_1041);
xor ( n30321 , n30319 , n30320 );
xor ( n30322 , n30310 , n30321 );
xor ( n30323 , RI19ab2d78_2433 , RI174a75f8_920);
not ( n11108 , n27689 );
and ( n11109 , n11108 , RI174a75f8_920);
and ( n11110 , n30323 , n27689 );
or ( n30324 , n11109 , n11110 );
buf ( n30325 , RI17338d58_2164);
xor ( n30326 , n30324 , n30325 );
buf ( n30327 , RI173c22d8_1809);
xor ( n30328 , n30326 , n30327 );
buf ( n30329 , RI1740afc8_1454);
xor ( n30330 , n30328 , n30329 );
buf ( n30331 , RI17512578_709);
xor ( n30332 , n30330 , n30331 );
xor ( n30333 , n30322 , n30332 );
and ( n30334 , n30308 , n30333 );
xor ( n30335 , n30284 , n30334 );
xor ( n30336 , n30260 , n30335 );
buf ( n30337 , RI17406450_1477);
xor ( n30338 , RI19aaaa38_2491 , RI17494188_1014);
not ( n11111 , n27689 );
and ( n11112 , n11111 , RI17494188_1014);
and ( n11113 , n30338 , n27689 );
or ( n30339 , n11112 , n11113 );
xor ( n30340 , RI19aa4318_2536 , RI17522748_659);
not ( n11114 , n27689 );
and ( n11115 , n11114 , RI17522748_659);
and ( n11116 , n30340 , n27689 );
or ( n30341 , n11115 , n11116 );
xor ( n30342 , n30339 , n30341 );
buf ( n30343 , RI173aee68_1903);
xor ( n30344 , n30342 , n30343 );
buf ( n30345 , RI173f7b58_1548);
xor ( n30346 , n30344 , n30345 );
buf ( n30347 , RI1733b4b8_2152);
xor ( n30348 , n30346 , n30347 );
xor ( n30349 , n30337 , n30348 );
xor ( n30350 , n30349 , n30178 );
xor ( n30351 , n29175 , n28185 );
xor ( n30352 , n30351 , n28827 );
not ( n30353 , n30352 );
xor ( n30354 , RI19a8e478_2695 , RI17466c60_1235);
not ( n11117 , n27689 );
and ( n11118 , n11117 , RI17466c60_1235);
and ( n11119 , n30354 , n27689 );
or ( n30355 , n11118 , n11119 );
xor ( n30356 , RI19abf0f0_2340 , RI174af938_880);
not ( n11120 , n27689 );
and ( n11121 , n11120 , RI174af938_880);
and ( n11122 , n30356 , n27689 );
or ( n30357 , n11121 , n11122 );
xor ( n30358 , n30355 , n30357 );
buf ( n30359 , RI17341098_2124);
xor ( n30360 , n30358 , n30359 );
buf ( n30361 , RI173ca618_1769);
xor ( n30362 , n30360 , n30361 );
buf ( n30363 , RI17413650_1413);
xor ( n30364 , n30362 , n30363 );
xor ( n30365 , n27927 , n30364 );
xor ( n30366 , RI19aa2068_2552 , RI17484198_1092);
not ( n11123 , n27689 );
and ( n11124 , n11123 , RI17484198_1092);
and ( n11125 , n30366 , n27689 );
or ( n30367 , n11124 , n11125 );
xor ( n30368 , n30367 , n28268 );
buf ( n30369 , RI1739ee78_1981);
xor ( n30370 , n30368 , n30369 );
buf ( n30371 , RI173e7eb0_1625);
xor ( n30372 , n30370 , n30371 );
buf ( n30373 , RI1745f988_1270);
xor ( n30374 , n30372 , n30373 );
xor ( n30375 , n30365 , n30374 );
and ( n30376 , n30353 , n30375 );
xor ( n30377 , n30350 , n30376 );
xor ( n30378 , n30336 , n30377 );
xor ( n30379 , RI19a98018_2626 , RI174789d8_1148);
not ( n11126 , n27689 );
and ( n11127 , n11126 , RI174789d8_1148);
and ( n11128 , n30379 , n27689 );
or ( n30380 , n11127 , n11128 );
xor ( n30381 , RI19ac7d90_2271 , RI174c67c8_793);
not ( n11129 , n27689 );
and ( n11130 , n11129 , RI174c67c8_793);
and ( n11131 , n30381 , n27689 );
or ( n30382 , n11130 , n11131 );
xor ( n30383 , n30380 , n30382 );
buf ( n30384 , RI173936b8_2037);
xor ( n30385 , n30383 , n30384 );
buf ( n30386 , RI173dc3a8_1682);
xor ( n30387 , n30385 , n30386 );
buf ( n30388 , RI17453e80_1327);
xor ( n30389 , n30387 , n30388 );
xor ( n30390 , n29652 , n30389 );
xor ( n30391 , n30390 , n28200 );
xor ( n30392 , RI19a841d0_2765 , RI17503de8_748);
not ( n11132 , n27689 );
and ( n11133 , n11132 , RI17503de8_748);
and ( n11134 , n30392 , n27689 );
or ( n30393 , n11133 , n11134 );
xor ( n30394 , n29799 , n30393 );
buf ( n30395 , RI1739ca60_1992);
xor ( n30396 , n30394 , n30395 );
buf ( n30397 , RI173e5a98_1636);
xor ( n30398 , n30396 , n30397 );
xor ( n30399 , n30398 , n27796 );
xor ( n30400 , n29036 , n30399 );
xor ( n30401 , n30400 , n29532 );
not ( n30402 , n30401 );
xor ( n30403 , RI19ab29b8_2435 , RI174a6f68_922);
not ( n11135 , n27689 );
and ( n11136 , n11135 , RI174a6f68_922);
and ( n11137 , n30403 , n27689 );
or ( n30404 , n11136 , n11137 );
xor ( n30405 , RI19aa8878_2506 , RI17498670_993);
not ( n11138 , n27689 );
and ( n11139 , n11138 , RI17498670_993);
and ( n11140 , n30405 , n27689 );
or ( n30406 , n11139 , n11140 );
xor ( n30407 , RI19a90368_2681 , RI17529390_638);
not ( n11141 , n27689 );
and ( n11142 , n11141 , RI17529390_638);
and ( n11143 , n30407 , n27689 );
or ( n30408 , n11142 , n11143 );
xor ( n30409 , n30406 , n30408 );
buf ( n30410 , RI173b3350_1882);
xor ( n30411 , n30409 , n30410 );
buf ( n30412 , RI173fc388_1526);
xor ( n30413 , n30411 , n30412 );
buf ( n30414 , RI173a71b8_1941);
xor ( n30415 , n30413 , n30414 );
xor ( n30416 , n30404 , n30415 );
xor ( n30417 , RI19a8af08_2718 , RI1746ced0_1205);
not ( n11144 , n27689 );
and ( n11145 , n11144 , RI1746ced0_1205);
and ( n11146 , n30417 , n27689 );
or ( n30418 , n11145 , n11146 );
xor ( n30419 , RI19abc8a0_2363 , RI174b5ba8_850);
not ( n11147 , n27689 );
and ( n11148 , n11147 , RI174b5ba8_850);
and ( n11149 , n30419 , n27689 );
or ( n30420 , n11148 , n11149 );
xor ( n30421 , n30418 , n30420 );
buf ( n30422 , RI17347308_2094);
xor ( n30423 , n30421 , n30422 );
buf ( n30424 , RI173d0bd0_1738);
xor ( n30425 , n30423 , n30424 );
buf ( n30426 , RI174486c0_1383);
xor ( n30427 , n30425 , n30426 );
xor ( n30428 , n30416 , n30427 );
and ( n30429 , n30402 , n30428 );
xor ( n30430 , n30391 , n30429 );
xor ( n30431 , n30378 , n30430 );
xor ( n30432 , n28247 , n29259 );
xor ( n30433 , n30432 , n29270 );
xor ( n30434 , RI19a8e6d0_2694 , RI17466fa8_1234);
not ( n11150 , n27689 );
and ( n11151 , n11150 , RI17466fa8_1234);
and ( n11152 , n30434 , n27689 );
or ( n30435 , n11151 , n11152 );
xor ( n30436 , RI19abf2d0_2339 , RI174afc80_879);
not ( n11153 , n27689 );
and ( n11154 , n11153 , RI174afc80_879);
and ( n11155 , n30436 , n27689 );
or ( n30437 , n11154 , n11155 );
xor ( n30438 , n30435 , n30437 );
xor ( n30439 , n30438 , n29983 );
buf ( n30440 , RI173ca960_1768);
xor ( n30441 , n30439 , n30440 );
buf ( n30442 , RI17413998_1412);
xor ( n30443 , n30441 , n30442 );
xor ( n30444 , n28278 , n30443 );
xor ( n30445 , n30444 , n28617 );
not ( n30446 , n30445 );
xor ( n30447 , n28046 , n29694 );
xor ( n30448 , RI19aae458_2466 , RI174920b8_1024);
not ( n11156 , n27689 );
and ( n11157 , n11156 , RI174920b8_1024);
and ( n11158 , n30448 , n27689 );
or ( n30449 , n11157 , n11158 );
xor ( n30450 , RI19ac6878_2281 , RI1751f3b8_669);
not ( n11159 , n27689 );
and ( n11160 , n11159 , RI1751f3b8_669);
and ( n11161 , n30450 , n27689 );
or ( n30451 , n11160 , n11161 );
xor ( n30452 , n30449 , n30451 );
xor ( n30453 , n30452 , n29112 );
buf ( n30454 , RI173f5a88_1558);
xor ( n30455 , n30453 , n30454 );
buf ( n30456 , RI17524638_653);
xor ( n30457 , n30455 , n30456 );
xor ( n30458 , n30447 , n30457 );
and ( n30459 , n30446 , n30458 );
xor ( n30460 , n30433 , n30459 );
xor ( n30461 , n30431 , n30460 );
xor ( n30462 , n30248 , n30461 );
not ( n30463 , n30462 );
buf ( n30464 , RI1740a5f0_1457);
xor ( n30465 , RI19aa8530_2507 , RI17498328_994);
not ( n11162 , n27689 );
and ( n11163 , n11162 , RI17498328_994);
and ( n11164 , n30465 , n27689 );
or ( n30466 , n11163 , n11164 );
xor ( n30467 , RI19a8eb08_2692 , RI17528e68_639);
not ( n11165 , n27689 );
and ( n11166 , n11165 , RI17528e68_639);
and ( n11167 , n30467 , n27689 );
or ( n30468 , n11166 , n11167 );
xor ( n30469 , n30466 , n30468 );
buf ( n30470 , RI173b3008_1883);
xor ( n30471 , n30469 , n30470 );
buf ( n30472 , RI173fc040_1527);
xor ( n30473 , n30471 , n30472 );
buf ( n30474 , RI173a4da0_1952);
xor ( n30475 , n30473 , n30474 );
xor ( n30476 , n30464 , n30475 );
xor ( n30477 , RI19a8acb0_2719 , RI1746cb88_1206);
not ( n11168 , n27689 );
and ( n11169 , n11168 , RI1746cb88_1206);
and ( n11170 , n30477 , n27689 );
or ( n30478 , n11169 , n11170 );
xor ( n30479 , RI19abc6c0_2364 , RI174b5860_851);
not ( n11171 , n27689 );
and ( n11172 , n11171 , RI174b5860_851);
and ( n11173 , n30479 , n27689 );
or ( n30480 , n11172 , n11173 );
xor ( n30481 , n30478 , n30480 );
buf ( n30482 , RI17346fc0_2095);
xor ( n30483 , n30481 , n30482 );
buf ( n30484 , RI173d0888_1739);
xor ( n30485 , n30483 , n30484 );
buf ( n30486 , RI17448378_1384);
xor ( n30487 , n30485 , n30486 );
xor ( n30488 , n30476 , n30487 );
xor ( n30489 , n28449 , n29975 );
xor ( n30490 , n30489 , n28759 );
not ( n30491 , n30490 );
xor ( n30492 , n28820 , n28557 );
xor ( n30493 , n30492 , n28569 );
and ( n30494 , n30491 , n30493 );
xor ( n30495 , n30488 , n30494 );
xor ( n30496 , n27916 , n30294 );
xor ( n30497 , n30496 , n30306 );
xor ( n30498 , n27761 , n29639 );
xor ( n30499 , n30498 , n30233 );
not ( n30500 , n30499 );
xor ( n30501 , RI19aa6b68_2518 , RI174996d8_988);
not ( n11174 , n27689 );
and ( n11175 , n11174 , RI174996d8_988);
and ( n11176 , n30501 , n27689 );
or ( n30502 , n11175 , n11176 );
xor ( n30503 , RI19a87dd0_2739 , RI1752ad58_633);
not ( n11177 , n27689 );
and ( n11178 , n11177 , RI1752ad58_633);
and ( n11179 , n30503 , n27689 );
or ( n30504 , n11178 , n11179 );
xor ( n30505 , n30502 , n30504 );
buf ( n30506 , RI173b43b8_1877);
xor ( n30507 , n30505 , n30506 );
buf ( n30508 , RI173fd3f0_1521);
xor ( n30509 , n30507 , n30508 );
xor ( n30510 , n30509 , n29040 );
xor ( n30511 , n28354 , n30510 );
xor ( n30512 , RI19a89270_2730 , RI1746df38_1200);
not ( n11180 , n27689 );
and ( n11181 , n11180 , RI1746df38_1200);
and ( n11182 , n30512 , n27689 );
or ( n30513 , n11181 , n11182 );
xor ( n30514 , RI19abad70_2375 , RI174b6c10_845);
not ( n11183 , n27689 );
and ( n11184 , n11183 , RI174b6c10_845);
and ( n11185 , n30514 , n27689 );
or ( n30515 , n11184 , n11185 );
xor ( n30516 , n30513 , n30515 );
buf ( n30517 , RI17359698_2089);
xor ( n30518 , n30516 , n30517 );
buf ( n30519 , RI173d1c50_1733);
xor ( n30520 , n30518 , n30519 );
buf ( n30521 , RI17449728_1378);
xor ( n30522 , n30520 , n30521 );
xor ( n30523 , n30511 , n30522 );
and ( n30524 , n30500 , n30523 );
xor ( n30525 , n30497 , n30524 );
xor ( n30526 , n28912 , n29889 );
xor ( n30527 , RI19a96bf0_2635 , RI1747a418_1140);
not ( n11186 , n27689 );
and ( n11187 , n11186 , RI1747a418_1140);
and ( n11188 , n30527 , n27689 );
or ( n30528 , n11187 , n11188 );
xor ( n30529 , RI19ac69e0_2280 , RI174c9108_785);
not ( n11189 , n27689 );
and ( n11190 , n11189 , RI174c9108_785);
and ( n11191 , n30529 , n27689 );
or ( n30530 , n11190 , n11191 );
xor ( n30531 , n30528 , n30530 );
buf ( n30532 , RI173950f8_2029);
xor ( n30533 , n30531 , n30532 );
buf ( n30534 , RI173ddde8_1674);
xor ( n30535 , n30533 , n30534 );
buf ( n30536 , RI174558c0_1319);
xor ( n30537 , n30535 , n30536 );
xor ( n30538 , n30526 , n30537 );
xor ( n30539 , RI19a90818_2679 , RI174665d0_1237);
not ( n11192 , n27689 );
and ( n11193 , n11192 , RI174665d0_1237);
and ( n11194 , n30539 , n27689 );
or ( n30540 , n11193 , n11194 );
xor ( n30541 , RI19ac0d88_2324 , RI174af2a8_882);
not ( n11195 , n27689 );
and ( n11196 , n11195 , RI174af2a8_882);
and ( n11197 , n30541 , n27689 );
or ( n30542 , n11196 , n11197 );
xor ( n30543 , n30540 , n30542 );
xor ( n30544 , n30543 , n28214 );
buf ( n30545 , RI173c9f88_1771);
xor ( n30546 , n30544 , n30545 );
buf ( n30547 , RI17412fc0_1415);
xor ( n30548 , n30546 , n30547 );
xor ( n30549 , n29870 , n30548 );
xor ( n30550 , n30549 , n28673 );
not ( n30551 , n30550 );
xor ( n30552 , n29654 , n30389 );
xor ( n30553 , n30552 , n28200 );
and ( n30554 , n30551 , n30553 );
xor ( n30555 , n30538 , n30554 );
xor ( n30556 , n30525 , n30555 );
xor ( n30557 , n30061 , n29105 );
xor ( n30558 , RI19aba050_2380 , RI1749c4c8_974);
not ( n11198 , n27689 );
and ( n11199 , n11198 , RI1749c4c8_974);
and ( n11200 , n30558 , n27689 );
or ( n30559 , n11199 , n11200 );
buf ( n30560 , RI1752f588_619);
xor ( n30561 , n30559 , n30560 );
buf ( n30562 , RI173b74f0_1862);
xor ( n30563 , n30561 , n30562 );
buf ( n30564 , RI174001e0_1507);
xor ( n30565 , n30563 , n30564 );
buf ( n30566 , RI173cdde0_1752);
xor ( n30567 , n30565 , n30566 );
xor ( n30568 , n30557 , n30567 );
not ( n30569 , n30488 );
and ( n30570 , n30569 , n30490 );
xor ( n30571 , n30568 , n30570 );
xor ( n30572 , n30556 , n30571 );
buf ( n30573 , RI173964a8_2023);
xor ( n30574 , n30573 , n30427 );
xor ( n30575 , n30574 , n29364 );
buf ( n30576 , RI173eee40_1591);
xor ( n30577 , n30576 , n28367 );
xor ( n30578 , n30577 , n29952 );
not ( n30579 , n30578 );
buf ( n30580 , RI1733fce8_2130);
xor ( n30581 , n30580 , n30189 );
xor ( n30582 , n30581 , n28715 );
and ( n30583 , n30579 , n30582 );
xor ( n30584 , n30575 , n30583 );
xor ( n30585 , n30572 , n30584 );
xor ( n30586 , n29527 , n27819 );
xor ( n30587 , RI19ac0338_2330 , RI174adef8_888);
not ( n11201 , n27689 );
and ( n11202 , n11201 , RI174adef8_888);
and ( n11203 , n30587 , n27689 );
or ( n30588 , n11202 , n11203 );
xor ( n30589 , n29661 , n30588 );
buf ( n30590 , RI1733f658_2132);
xor ( n30591 , n30589 , n30590 );
buf ( n30592 , RI173c8bd8_1777);
xor ( n30593 , n30591 , n30592 );
xor ( n30594 , n30593 , n28973 );
xor ( n30595 , n30586 , n30594 );
xor ( n30596 , n29245 , n27700 );
xor ( n30597 , n30596 , n27712 );
not ( n30598 , n30597 );
buf ( n30599 , RI17454ee8_1322);
xor ( n30600 , n30599 , n28519 );
xor ( n30601 , n30600 , n28304 );
and ( n30602 , n30598 , n30601 );
xor ( n30603 , n30595 , n30602 );
xor ( n30604 , n30585 , n30603 );
xor ( n30605 , n30495 , n30604 );
xor ( n30606 , n29061 , n29827 );
xor ( n30607 , n30606 , n29839 );
xor ( n30608 , RI19ab3840_2427 , RI174a4e98_932);
not ( n11204 , n27689 );
and ( n11205 , n11204 , RI174a4e98_932);
and ( n11206 , n30608 , n27689 );
or ( n30609 , n11205 , n11206 );
xor ( n30610 , n30609 , n30073 );
buf ( n30611 , RI173bfec0_1820);
xor ( n30612 , n30610 , n30611 );
buf ( n30613 , RI17408bb0_1465);
xor ( n30614 , n30612 , n30613 );
buf ( n30615 , RI17455578_1320);
xor ( n30616 , n30614 , n30615 );
xor ( n30617 , n28548 , n30616 );
xor ( n30618 , RI19a964e8_2638 , RI17479a40_1143);
not ( n11207 , n27689 );
and ( n11208 , n11207 , RI17479a40_1143);
and ( n11209 , n30618 , n27689 );
or ( n30619 , n11208 , n11209 );
xor ( n30620 , RI19ac63c8_2283 , RI174c8190_788);
not ( n11210 , n27689 );
and ( n11211 , n11210 , RI174c8190_788);
and ( n11212 , n30620 , n27689 );
or ( n30621 , n11211 , n11212 );
xor ( n30622 , n30619 , n30621 );
buf ( n30623 , RI17394720_2032);
xor ( n30624 , n30622 , n30623 );
xor ( n30625 , n30624 , n28508 );
xor ( n30626 , n30625 , n30599 );
xor ( n30627 , n30617 , n30626 );
not ( n30628 , n30627 );
xor ( n30629 , n29866 , n30548 );
xor ( n30630 , n30629 , n28673 );
and ( n30631 , n30628 , n30630 );
xor ( n30632 , n30607 , n30631 );
xor ( n30633 , n29854 , n29421 );
xor ( n30634 , RI19aa9868_2499 , RI17496258_1004);
not ( n11213 , n27689 );
and ( n11214 , n11213 , RI17496258_1004);
and ( n11215 , n30634 , n27689 );
or ( n30635 , n11214 , n11215 );
xor ( n30636 , RI19a99ad0_2614 , RI17525ad8_649);
not ( n11216 , n27689 );
and ( n11217 , n11216 , RI17525ad8_649);
and ( n11218 , n30636 , n27689 );
or ( n30637 , n11217 , n11218 );
xor ( n30638 , n30635 , n30637 );
buf ( n30639 , RI173b0f38_1893);
xor ( n30640 , n30638 , n30639 );
xor ( n30641 , n30640 , n28163 );
buf ( n30642 , RI17390580_2052);
xor ( n30643 , n30641 , n30642 );
xor ( n30644 , n30633 , n30643 );
xor ( n30645 , RI19aa6988_2519 , RI1747fcb0_1113);
not ( n11219 , n27689 );
and ( n11220 , n11219 , RI1747fcb0_1113);
and ( n11221 , n30645 , n27689 );
or ( n30646 , n11220 , n11221 );
xor ( n30647 , RI19a87b78_2740 , RI17500a58_758);
not ( n11222 , n27689 );
and ( n11223 , n11222 , RI17500a58_758);
and ( n11224 , n30647 , n27689 );
or ( n30648 , n11223 , n11224 );
xor ( n30649 , n30646 , n30648 );
buf ( n30650 , RI1739a990_2002);
xor ( n30651 , n30649 , n30650 );
buf ( n30652 , RI173e3680_1647);
xor ( n30653 , n30651 , n30652 );
buf ( n30654 , RI1745b4a0_1291);
xor ( n30655 , n30653 , n30654 );
xor ( n30656 , n29510 , n30655 );
xor ( n30657 , RI19ab82c8_2394 , RI1749d1e8_970);
not ( n11225 , n27689 );
and ( n11226 , n11225 , RI1749d1e8_970);
and ( n11227 , n30657 , n27689 );
or ( n30658 , n11226 , n11227 );
buf ( n30659 , RI17530a28_615);
xor ( n30660 , n30658 , n30659 );
buf ( n30661 , RI173b8210_1858);
xor ( n30662 , n30660 , n30661 );
xor ( n30663 , n30662 , n28958 );
buf ( n30664 , RI173d6e58_1708);
xor ( n30665 , n30663 , n30664 );
xor ( n30666 , n30656 , n30665 );
not ( n30667 , n30666 );
xor ( n30668 , n28526 , n27764 );
xor ( n30669 , n30668 , n28125 );
and ( n30670 , n30667 , n30669 );
xor ( n30671 , n30644 , n30670 );
xor ( n30672 , n30632 , n30671 );
buf ( n30673 , RI1744a790_1373);
xor ( n30674 , n30673 , n28463 );
xor ( n30675 , n30674 , n27752 );
xor ( n30676 , n30619 , n28519 );
xor ( n30677 , n30676 , n28304 );
not ( n30678 , n30677 );
xor ( n30679 , RI19acd5b0_2229 , RI17511600_712);
not ( n11228 , n27689 );
and ( n11229 , n11228 , RI17511600_712);
and ( n11230 , n30679 , n27689 );
or ( n30680 , n11229 , n11230 );
xor ( n30681 , RI19a946e8_2651 , RI1747adf0_1137);
not ( n11231 , n27689 );
and ( n11232 , n11231 , RI1747adf0_1137);
and ( n11233 , n30681 , n27689 );
or ( n30682 , n11232 , n11233 );
xor ( n30683 , RI19ac4910_2295 , RI174ca080_782);
not ( n11234 , n27689 );
and ( n11235 , n11234 , RI174ca080_782);
and ( n11236 , n30683 , n27689 );
or ( n30684 , n11235 , n11236 );
xor ( n30685 , n30682 , n30684 );
buf ( n30686 , RI17395ad0_2026);
xor ( n30687 , n30685 , n30686 );
buf ( n30688 , RI173de7c0_1671);
xor ( n30689 , n30687 , n30688 );
buf ( n30690 , RI17456298_1316);
xor ( n30691 , n30689 , n30690 );
xor ( n30692 , n30680 , n30691 );
xor ( n30693 , n30692 , n30475 );
and ( n30694 , n30678 , n30693 );
xor ( n30695 , n30675 , n30694 );
xor ( n30696 , n30672 , n30695 );
xor ( n30697 , RI19aa10f0_2560 , RI17486268_1082);
not ( n11237 , n27689 );
and ( n11238 , n11237 , RI17486268_1082);
and ( n11239 , n30697 , n27689 );
or ( n30698 , n11238 , n11239 );
xor ( n30699 , RI19acffe0_2211 , RI1750c8a8_727);
not ( n11240 , n27689 );
and ( n11241 , n11240 , RI1750c8a8_727);
and ( n11242 , n30699 , n27689 );
or ( n30700 , n11241 , n11242 );
xor ( n30701 , n30698 , n30700 );
buf ( n30702 , RI173a1290_1970);
xor ( n30703 , n30701 , n30702 );
xor ( n30704 , n30703 , n28395 );
buf ( n30705 , RI17467cc8_1230);
xor ( n30706 , n30704 , n30705 );
xor ( n30707 , n29934 , n30706 );
xor ( n30708 , RI19ab5118_2416 , RI174a37a0_939);
not ( n11243 , n27689 );
and ( n11244 , n11243 , RI174a37a0_939);
and ( n11245 , n30708 , n27689 );
or ( n30709 , n11244 , n11245 );
buf ( n30710 , RI17335248_2182);
xor ( n30711 , n30709 , n30710 );
buf ( n30712 , RI173be7c8_1827);
xor ( n30713 , n30711 , n30712 );
buf ( n30714 , RI174074b8_1472);
xor ( n30715 , n30713 , n30714 );
buf ( n30716 , RI174458d0_1397);
xor ( n30717 , n30715 , n30716 );
xor ( n30718 , n30707 , n30717 );
xor ( n30719 , RI19aba578_2378 , RI1749cb58_972);
not ( n11246 , n27689 );
and ( n11247 , n11246 , RI1749cb58_972);
and ( n11248 , n30719 , n27689 );
or ( n30720 , n11247 , n11248 );
xor ( n30721 , n30720 , n28659 );
xor ( n30722 , n30721 , n29148 );
not ( n30723 , n30722 );
xor ( n30724 , n28871 , n30218 );
xor ( n30725 , n30724 , n27807 );
and ( n30726 , n30723 , n30725 );
xor ( n30727 , n30718 , n30726 );
xor ( n30728 , n30696 , n30727 );
buf ( n30729 , RI17455230_1321);
xor ( n30730 , n30729 , n28917 );
xor ( n30731 , n30730 , n28929 );
xor ( n30732 , n28165 , n29199 );
xor ( n30733 , n30732 , n29211 );
not ( n30734 , n30733 );
xor ( n30735 , RI19aa7540_2514 , RI17523198_657);
not ( n11249 , n27689 );
and ( n11250 , n11249 , RI17523198_657);
and ( n11251 , n30735 , n27689 );
or ( n30736 , n11250 , n11251 );
xor ( n30737 , n30736 , n30189 );
xor ( n30738 , n30737 , n28715 );
and ( n30739 , n30734 , n30738 );
xor ( n30740 , n30731 , n30739 );
xor ( n30741 , n30728 , n30740 );
xor ( n30742 , n30605 , n30741 );
and ( n30743 , n30463 , n30742 );
xor ( n30744 , n29982 , n30743 );
not ( n11252 , n29614 );
and ( n11253 , n11252 , RI1733f310_2133);
and ( n11254 , n30744 , n29614 );
or ( n30745 , n11253 , n11254 );
not ( n11255 , RI1754c610_2);
and ( n11256 , n11255 , n30745 );
and ( n11257 , C0 , RI1754c610_2);
or ( n30746 , n11256 , n11257 );
buf ( n30747 , n30746 );
xor ( n30748 , n30213 , n29573 );
xor ( n30749 , RI19a8f648_2687 , RI17464b90_1245);
not ( n11258 , n27689 );
and ( n11259 , n11258 , RI17464b90_1245);
and ( n11260 , n30749 , n27689 );
or ( n30750 , n11259 , n11260 );
xor ( n30751 , RI19abff78_2332 , RI174ad868_890);
not ( n11261 , n27689 );
and ( n11262 , n11261 , RI174ad868_890);
and ( n11263 , n30751 , n27689 );
or ( n30752 , n11262 , n11263 );
xor ( n30753 , n30750 , n30752 );
buf ( n30754 , RI1733efc8_2134);
xor ( n30755 , n30753 , n30754 );
buf ( n30756 , RI173c8548_1779);
xor ( n30757 , n30755 , n30756 );
xor ( n30758 , n30757 , n29151 );
xor ( n30759 , n30748 , n30758 );
buf ( n30760 , RI173c8890_1778);
xor ( n30761 , n30760 , n29532 );
xor ( n30762 , n30761 , n29544 );
not ( n30763 , n30762 );
xor ( n30764 , n28582 , n29176 );
xor ( n30765 , n30764 , n29187 );
and ( n30766 , n30763 , n30765 );
xor ( n30767 , n30759 , n30766 );
xor ( n30768 , n27705 , n27909 );
xor ( n30769 , n30768 , n27921 );
xor ( n30770 , n29219 , n28995 );
xor ( n30771 , RI19aadd50_2469 , RI174916e0_1027);
not ( n11264 , n27689 );
and ( n11265 , n11264 , RI174916e0_1027);
and ( n11266 , n30771 , n27689 );
or ( n30772 , n11265 , n11266 );
xor ( n30773 , RI19ac1f58_2314 , RI1751e440_672);
not ( n11267 , n27689 );
and ( n11268 , n11267 , RI1751e440_672);
and ( n11269 , n30773 , n27689 );
or ( n30774 , n11268 , n11269 );
xor ( n30775 , n30772 , n30774 );
buf ( n30776 , RI173ac3c0_1916);
xor ( n30777 , n30775 , n30776 );
xor ( n30778 , n30777 , n29427 );
buf ( n30779 , RI17519c10_686);
xor ( n30780 , n30778 , n30779 );
xor ( n30781 , n30770 , n30780 );
not ( n30782 , n30781 );
xor ( n30783 , RI19accc50_2233 , RI17515e30_698);
not ( n11270 , n27689 );
and ( n11271 , n11270 , RI17515e30_698);
and ( n11272 , n30783 , n27689 );
or ( n30784 , n11271 , n11272 );
xor ( n30785 , n28748 , n30784 );
xor ( n30786 , n30785 , n29641 );
buf ( n30787 , RI173efb60_1587);
xor ( n30788 , n30786 , n30787 );
xor ( n30789 , n30788 , n28932 );
xor ( n30790 , n29499 , n30789 );
xor ( n30791 , RI19ab1ba8_2441 , RI174a96c8_910);
not ( n11273 , n27689 );
and ( n11274 , n11273 , RI174a96c8_910);
and ( n11275 , n30791 , n27689 );
or ( n30792 , n11274 , n11275 );
buf ( n30793 , RI1733ae28_2154);
xor ( n30794 , n30792 , n30793 );
xor ( n30795 , n30794 , n30220 );
buf ( n30796 , RI1740d098_1444);
xor ( n30797 , n30795 , n30796 );
buf ( n30798 , RI17457990_1309);
xor ( n30799 , n30797 , n30798 );
xor ( n30800 , n30790 , n30799 );
and ( n30801 , n30782 , n30800 );
xor ( n30802 , n30769 , n30801 );
xor ( n30803 , RI19aa7888_2513 , RI1749a740_983);
not ( n11276 , n27689 );
and ( n11277 , n11276 , RI1749a740_983);
and ( n11278 , n30803 , n27689 );
or ( n30804 , n11277 , n11278 );
xor ( n30805 , RI19a88a00_2734 , RI1752c720_628);
not ( n11279 , n27689 );
and ( n11280 , n11279 , RI1752c720_628);
and ( n11281 , n30805 , n27689 );
or ( n30806 , n11280 , n11281 );
xor ( n30807 , n30804 , n30806 );
buf ( n30808 , RI173b5420_1872);
xor ( n30809 , n30807 , n30808 );
buf ( n30810 , RI173fe458_1516);
xor ( n30811 , n30809 , n30810 );
buf ( n30812 , RI173bb9d8_1841);
xor ( n30813 , n30811 , n30812 );
xor ( n30814 , n29968 , n30813 );
xor ( n30815 , RI19a89bd0_2726 , RI1746efa0_1195);
not ( n11282 , n27689 );
and ( n11283 , n11282 , RI1746efa0_1195);
and ( n11284 , n30815 , n27689 );
or ( n30816 , n11283 , n11284 );
xor ( n30817 , RI19abb748_2371 , RI174b7c78_840);
not ( n11285 , n27689 );
and ( n11286 , n11285 , RI174b7c78_840);
and ( n11287 , n30817 , n27689 );
or ( n30818 , n11286 , n11287 );
xor ( n30819 , n30816 , n30818 );
buf ( n30820 , RI17389fc8_2083);
xor ( n30821 , n30819 , n30820 );
xor ( n30822 , n30821 , n28453 );
xor ( n30823 , n30822 , n30673 );
xor ( n30824 , n30814 , n30823 );
xor ( n30825 , n28552 , n30616 );
xor ( n30826 , n30825 , n30626 );
not ( n30827 , n30826 );
xor ( n30828 , n30292 , n28043 );
xor ( n30829 , n30828 , n28055 );
and ( n30830 , n30827 , n30829 );
xor ( n30831 , n30824 , n30830 );
xor ( n30832 , n30802 , n30831 );
xor ( n30833 , n28922 , n30537 );
xor ( n30834 , RI19aa29c8_2548 , RI175279c8_643);
not ( n11288 , n27689 );
and ( n11289 , n11288 , RI175279c8_643);
and ( n11290 , n30834 , n27689 );
or ( n30835 , n11289 , n11290 );
xor ( n30836 , n27822 , n30835 );
buf ( n30837 , RI173b22e8_1887);
xor ( n30838 , n30836 , n30837 );
buf ( n30839 , RI173fafd8_1532);
xor ( n30840 , n30838 , n30839 );
buf ( n30841 , RI1739de10_1986);
xor ( n30842 , n30840 , n30841 );
xor ( n30843 , n30833 , n30842 );
buf ( n30844 , RI173a7ed8_1937);
xor ( n30845 , n30844 , n28137 );
xor ( n30846 , n30845 , n28493 );
not ( n30847 , n30846 );
xor ( n30848 , RI19aa8080_2509 , RI17497c98_996);
not ( n11291 , n27689 );
and ( n11292 , n11291 , RI17497c98_996);
and ( n11293 , n30848 , n27689 );
or ( n30849 , n11292 , n11293 );
xor ( n30850 , RI19a8b958_2714 , RI17528418_641);
not ( n11294 , n27689 );
and ( n11295 , n11294 , RI17528418_641);
and ( n11296 , n30850 , n27689 );
or ( n30851 , n11295 , n11296 );
xor ( n30852 , n30849 , n30851 );
xor ( n30853 , n30852 , n30103 );
buf ( n30854 , RI173fb9b0_1529);
xor ( n30855 , n30853 , n30854 );
buf ( n30856 , RI173a0570_1974);
xor ( n30857 , n30855 , n30856 );
xor ( n30858 , n27841 , n30857 );
xor ( n30859 , RI19a8a878_2721 , RI1746c1b0_1209);
not ( n11297 , n27689 );
and ( n11298 , n11297 , RI1746c1b0_1209);
and ( n11299 , n30859 , n27689 );
or ( n30860 , n11298 , n11299 );
xor ( n30861 , RI19abc378_2366 , RI174b4e88_854);
not ( n11300 , n27689 );
and ( n11301 , n11300 , RI174b4e88_854);
and ( n11302 , n30861 , n27689 );
or ( n30862 , n11301 , n11302 );
xor ( n30863 , n30860 , n30862 );
buf ( n30864 , RI173465e8_2098);
xor ( n30865 , n30863 , n30864 );
buf ( n30866 , RI173cfeb0_1742);
xor ( n30867 , n30865 , n30866 );
buf ( n30868 , RI174479a0_1387);
xor ( n30869 , n30867 , n30868 );
xor ( n30870 , n30858 , n30869 );
and ( n30871 , n30847 , n30870 );
xor ( n30872 , n30843 , n30871 );
xor ( n30873 , n30832 , n30872 );
xor ( n30874 , RI19ac1670_2319 , RI174acb48_894);
not ( n11303 , n27689 );
and ( n11304 , n11303 , RI174acb48_894);
and ( n11305 , n30874 , n27689 );
or ( n30875 , n11304 , n11305 );
xor ( n30876 , n30875 , n27975 );
xor ( n30877 , n30876 , n29346 );
buf ( n30878 , RI17395e18_2025);
xor ( n30879 , RI19a8aad0_2720 , RI1746c840_1207);
not ( n11306 , n27689 );
and ( n11307 , n11306 , RI1746c840_1207);
and ( n11308 , n30879 , n27689 );
or ( n30880 , n11307 , n11308 );
xor ( n30881 , RI19abc4e0_2365 , RI174b5518_852);
not ( n11309 , n27689 );
and ( n11310 , n11309 , RI174b5518_852);
and ( n11311 , n30881 , n27689 );
or ( n30882 , n11310 , n11311 );
xor ( n30883 , n30880 , n30882 );
buf ( n30884 , RI17346c78_2096);
xor ( n30885 , n30883 , n30884 );
buf ( n30886 , RI173d0540_1740);
xor ( n30887 , n30885 , n30886 );
buf ( n30888 , RI17448030_1385);
xor ( n30889 , n30887 , n30888 );
xor ( n30890 , n30878 , n30889 );
xor ( n30891 , RI19a9efa8_2577 , RI17489a30_1065);
not ( n11312 , n27689 );
and ( n11313 , n11312 , RI17489a30_1065);
and ( n11314 , n30891 , n27689 );
or ( n30892 , n11313 , n11314 );
xor ( n30893 , RI19acda60_2227 , RI17512050_710);
not ( n11315 , n27689 );
and ( n11316 , n11315 , RI17512050_710);
and ( n11317 , n30893 , n27689 );
or ( n30894 , n11316 , n11317 );
xor ( n30895 , n30892 , n30894 );
buf ( n30896 , RI173a4a58_1953);
xor ( n30897 , n30895 , n30896 );
buf ( n30898 , RI173ed748_1598);
xor ( n30899 , n30897 , n30898 );
buf ( n30900 , RI1748c190_1053);
xor ( n30901 , n30899 , n30900 );
xor ( n30902 , n30890 , n30901 );
not ( n30903 , n30902 );
xor ( n30904 , n29583 , n29767 );
xor ( n30905 , n30904 , n30510 );
and ( n30906 , n30903 , n30905 );
xor ( n30907 , n30877 , n30906 );
xor ( n30908 , n30873 , n30907 );
xor ( n30909 , n30132 , n28392 );
xor ( n30910 , RI19ab4740_2420 , RI174a2738_944);
not ( n11318 , n27689 );
and ( n11319 , n11318 , RI174a2738_944);
and ( n11320 , n30910 , n27689 );
or ( n30911 , n11319 , n11320 );
buf ( n30912 , RI173341e0_2187);
xor ( n30913 , n30911 , n30912 );
buf ( n30914 , RI173bd760_1832);
xor ( n30915 , n30913 , n30914 );
xor ( n30916 , n30915 , n30337 );
buf ( n30917 , RI1740d728_1442);
xor ( n30918 , n30916 , n30917 );
xor ( n30919 , n30909 , n30918 );
not ( n30920 , n30759 );
and ( n30921 , n30920 , n30762 );
xor ( n30922 , n30919 , n30921 );
xor ( n30923 , n30908 , n30922 );
xor ( n30924 , n30767 , n30923 );
xor ( n30925 , RI19a9e288_2583 , RI1748c4d8_1052);
not ( n11321 , n27689 );
and ( n11322 , n11321 , RI1748c4d8_1052);
and ( n11323 , n30925 , n27689 );
or ( n30926 , n11322 , n11323 );
xor ( n30927 , RI19accea8_2232 , RI17516880_696);
not ( n11324 , n27689 );
and ( n11325 , n11324 , RI17516880_696);
and ( n11326 , n30927 , n27689 );
or ( n30928 , n11325 , n11326 );
xor ( n30929 , n30926 , n30928 );
xor ( n30930 , n30929 , n27741 );
buf ( n30931 , RI173f01f0_1585);
xor ( n30932 , n30930 , n30931 );
buf ( n30933 , RI174a5528_930);
xor ( n30934 , n30932 , n30933 );
xor ( n30935 , n28768 , n30934 );
xor ( n30936 , n30935 , n28533 );
xor ( n30937 , RI19aa9430_2501 , RI17499390_989);
not ( n11327 , n27689 );
and ( n11328 , n11327 , RI17499390_989);
and ( n11329 , n30937 , n27689 );
or ( n30938 , n11328 , n11329 );
xor ( n30939 , RI19a96998_2636 , RI1752a830_634);
not ( n11330 , n27689 );
and ( n11331 , n11330 , RI1752a830_634);
and ( n11332 , n30939 , n27689 );
or ( n30940 , n11331 , n11332 );
xor ( n30941 , n30938 , n30940 );
buf ( n30942 , RI173b4070_1878);
xor ( n30943 , n30941 , n30942 );
buf ( n30944 , RI173fd0a8_1522);
xor ( n30945 , n30943 , n30944 );
xor ( n30946 , n30945 , n29575 );
xor ( n30947 , n28014 , n30946 );
xor ( n30948 , RI19a89018_2731 , RI1746dbf0_1201);
not ( n11333 , n27689 );
and ( n11334 , n11333 , RI1746dbf0_1201);
and ( n11335 , n30948 , n27689 );
or ( n30949 , n11334 , n11335 );
xor ( n30950 , n30949 , n28345 );
buf ( n30951 , RI17359350_2090);
xor ( n30952 , n30950 , n30951 );
buf ( n30953 , RI173d1908_1734);
xor ( n30954 , n30952 , n30953 );
buf ( n30955 , RI174493e0_1379);
xor ( n30956 , n30954 , n30955 );
xor ( n30957 , n30947 , n30956 );
not ( n30958 , n30957 );
xor ( n30959 , n28203 , n29079 );
xor ( n30960 , n30959 , n28583 );
and ( n30961 , n30958 , n30960 );
xor ( n30962 , n30936 , n30961 );
xor ( n30963 , RI19a905c0_2680 , RI17466288_1238);
not ( n11336 , n27689 );
and ( n11337 , n11336 , RI17466288_1238);
and ( n11338 , n30963 , n27689 );
or ( n30964 , n11337 , n11338 );
xor ( n30965 , RI19ac0ba8_2325 , RI174aef60_883);
not ( n11339 , n27689 );
and ( n11340 , n11339 , RI174aef60_883);
and ( n11341 , n30965 , n27689 );
or ( n30966 , n11340 , n11341 );
xor ( n30967 , n30964 , n30966 );
xor ( n30968 , n30967 , n29861 );
buf ( n30969 , RI173c9c40_1772);
xor ( n30970 , n30968 , n30969 );
buf ( n30971 , RI17412c78_1416);
xor ( n30972 , n30970 , n30971 );
xor ( n30973 , n29691 , n30972 );
xor ( n30974 , n30973 , n29123 );
buf ( n30975 , RI1746e910_1197);
xor ( n30976 , n30975 , n27897 );
xor ( n30977 , n30976 , n27858 );
not ( n30978 , n30977 );
xor ( n30979 , n29282 , n30017 );
buf ( n30980 , RI1752ffd8_617);
xor ( n30981 , n30720 , n30980 );
buf ( n30982 , RI173b7b80_1860);
xor ( n30983 , n30981 , n30982 );
xor ( n30984 , n30983 , n29136 );
buf ( n30985 , RI173d2628_1730);
xor ( n30986 , n30984 , n30985 );
xor ( n30987 , n30979 , n30986 );
and ( n30988 , n30978 , n30987 );
xor ( n30989 , n30974 , n30988 );
xor ( n30990 , n30962 , n30989 );
xor ( n30991 , RI19aa81e8_2508 , RI17497fe0_995);
not ( n11342 , n27689 );
and ( n11343 , n11342 , RI17497fe0_995);
and ( n11344 , n30991 , n27689 );
or ( n30992 , n11343 , n11344 );
xor ( n30993 , RI19a8d230_2703 , RI17528940_640);
not ( n11345 , n27689 );
and ( n11346 , n11345 , RI17528940_640);
and ( n11347 , n30993 , n27689 );
or ( n30994 , n11346 , n11347 );
xor ( n30995 , n30992 , n30994 );
buf ( n30996 , RI173b2cc0_1884);
xor ( n30997 , n30995 , n30996 );
buf ( n30998 , RI173fbcf8_1528);
xor ( n30999 , n30997 , n30998 );
buf ( n31000 , RI173a2988_1963);
xor ( n31001 , n30999 , n31000 );
xor ( n31002 , n30122 , n31001 );
xor ( n31003 , n31002 , n30889 );
xor ( n31004 , n29963 , n30164 );
xor ( n31005 , n31004 , n29490 );
not ( n31006 , n31005 );
xor ( n31007 , n28574 , n29176 );
xor ( n31008 , n31007 , n29187 );
and ( n31009 , n31006 , n31008 );
xor ( n31010 , n31003 , n31009 );
xor ( n31011 , n30990 , n31010 );
xor ( n31012 , n29048 , n28027 );
xor ( n31013 , n31012 , n29827 );
xor ( n31014 , RI19aa0d30_2562 , RI17485bd8_1084);
not ( n11348 , n27689 );
and ( n11349 , n11348 , RI17485bd8_1084);
and ( n11350 , n31014 , n27689 );
or ( n31015 , n11349 , n11350 );
xor ( n31016 , RI19acfb30_2213 , RI1750be58_729);
not ( n11351 , n27689 );
and ( n11352 , n11351 , RI1750be58_729);
and ( n11353 , n31016 , n27689 );
or ( n31017 , n11352 , n11353 );
xor ( n31018 , n31015 , n31017 );
buf ( n31019 , RI173a0c00_1972);
xor ( n31020 , n31018 , n31019 );
buf ( n31021 , RI173e98f0_1617);
xor ( n31022 , n31020 , n31021 );
buf ( n31023 , RI17463498_1252);
xor ( n31024 , n31022 , n31023 );
xor ( n31025 , n27778 , n31024 );
xor ( n31026 , n31025 , n29306 );
not ( n31027 , n31026 );
xor ( n31028 , RI19ab03c0_2452 , RI1748d888_1046);
not ( n11354 , n27689 );
and ( n11355 , n11354 , RI1748d888_1046);
and ( n11356 , n31028 , n27689 );
or ( n31029 , n11355 , n11356 );
xor ( n31030 , RI19aa40c0_2537 , RI17518770_690);
not ( n11357 , n27689 );
and ( n11358 , n11357 , RI17518770_690);
and ( n11359 , n31030 , n27689 );
or ( n31031 , n11358 , n11359 );
xor ( n31032 , n31029 , n31031 );
buf ( n31033 , RI173a88b0_1934);
xor ( n31034 , n31032 , n31033 );
buf ( n31035 , RI173f15a0_1579);
xor ( n31036 , n31034 , n31035 );
buf ( n31037 , RI174b2db8_864);
xor ( n31038 , n31036 , n31037 );
xor ( n31039 , n30559 , n31038 );
xor ( n31040 , n31039 , n30271 );
and ( n31041 , n31027 , n31040 );
xor ( n31042 , n31013 , n31041 );
xor ( n31043 , n31011 , n31042 );
xor ( n31044 , n30592 , n28983 );
xor ( n31045 , n31044 , n28995 );
xor ( n31046 , n28826 , n28557 );
xor ( n31047 , n31046 , n28569 );
not ( n31048 , n31047 );
xor ( n31049 , n29646 , n30389 );
xor ( n31050 , n31049 , n28200 );
and ( n31051 , n31048 , n31050 );
xor ( n31052 , n31045 , n31051 );
xor ( n31053 , n31043 , n31052 );
xor ( n31054 , n30924 , n31053 );
xor ( n31055 , RI19aa24a0_2550 , RI17484828_1090);
not ( n11360 , n27689 );
and ( n11361 , n11360 , RI17484828_1090);
and ( n11362 , n31055 , n27689 );
or ( n31056 , n11361 , n11362 );
xor ( n31057 , RI19a83690_2770 , RI17509f68_735);
not ( n11363 , n27689 );
and ( n11364 , n11363 , RI17509f68_735);
and ( n11365 , n31057 , n27689 );
or ( n31058 , n11364 , n11365 );
xor ( n31059 , n31056 , n31058 );
buf ( n31060 , RI1739f508_1979);
xor ( n31061 , n31059 , n31060 );
buf ( n31062 , RI173e8540_1623);
xor ( n31063 , n31061 , n31062 );
buf ( n31064 , RI17460018_1268);
xor ( n31065 , n31063 , n31064 );
xor ( n31066 , n28324 , n31065 );
xor ( n31067 , RI19ab65b8_2406 , RI174a1d60_947);
not ( n11366 , n27689 );
and ( n11367 , n11366 , RI174a1d60_947);
and ( n11368 , n31067 , n27689 );
or ( n31068 , n11367 , n11368 );
buf ( n31069 , RI17333808_2190);
xor ( n31070 , n31068 , n31069 );
buf ( n31071 , RI173bcd88_1835);
xor ( n31072 , n31070 , n31071 );
buf ( n31073 , RI17405a78_1480);
xor ( n31074 , n31072 , n31073 );
buf ( n31075 , RI17406ae0_1475);
xor ( n31076 , n31074 , n31075 );
xor ( n31077 , n31066 , n31076 );
xor ( n31078 , n29448 , n30030 );
xor ( n31079 , n31078 , n30972 );
not ( n31080 , n31079 );
xor ( n31081 , RI19aba8c0_2377 , RI1749cea0_971);
not ( n11369 , n27689 );
and ( n11370 , n11369 , RI1749cea0_971);
and ( n11371 , n31081 , n27689 );
or ( n31082 , n11370 , n11371 );
buf ( n31083 , RI17530500_616);
xor ( n31084 , n31082 , n31083 );
buf ( n31085 , RI173b7ec8_1859);
xor ( n31086 , n31084 , n31085 );
xor ( n31087 , n31086 , n29508 );
buf ( n31088 , RI173d4a40_1719);
xor ( n31089 , n31087 , n31088 );
xor ( n31090 , n29139 , n31089 );
xor ( n31091 , RI19a9aac0_2607 , RI17471700_1183);
not ( n11372 , n27689 );
and ( n11373 , n11372 , RI17471700_1183);
and ( n11374 , n31091 , n27689 );
or ( n31092 , n11373 , n11374 );
xor ( n31093 , RI19aca298_2254 , RI174bb350_828);
not ( n11375 , n27689 );
and ( n11376 , n11375 , RI174bb350_828);
and ( n11377 , n31093 , n27689 );
or ( n31094 , n11376 , n11377 );
xor ( n31095 , n31092 , n31094 );
xor ( n31096 , n31095 , n29309 );
buf ( n31097 , RI173d5418_1716);
xor ( n31098 , n31096 , n31097 );
buf ( n31099 , RI1744cef0_1361);
xor ( n31100 , n31098 , n31099 );
xor ( n31101 , n31090 , n31100 );
and ( n31102 , n31080 , n31101 );
xor ( n31103 , n31077 , n31102 );
buf ( n31104 , RI173a4710_1954);
xor ( n31105 , RI19a94940_2650 , RI1747b138_1136);
not ( n11378 , n27689 );
and ( n11379 , n11378 , RI1747b138_1136);
and ( n11380 , n31105 , n27689 );
or ( n31106 , n11379 , n11380 );
xor ( n31107 , RI19ac4b68_2294 , RI174ca5a8_781);
not ( n11381 , n27689 );
and ( n11382 , n11381 , RI174ca5a8_781);
and ( n11383 , n31107 , n27689 );
or ( n31108 , n11382 , n11383 );
xor ( n31109 , n31106 , n31108 );
xor ( n31110 , n31109 , n30878 );
buf ( n31111 , RI173deb08_1670);
xor ( n31112 , n31110 , n31111 );
buf ( n31113 , RI174565e0_1315);
xor ( n31114 , n31112 , n31113 );
xor ( n31115 , n31104 , n31114 );
xor ( n31116 , n31115 , n30415 );
not ( n31117 , n31077 );
and ( n31118 , n31117 , n31079 );
xor ( n31119 , n31116 , n31118 );
xor ( n31120 , n29006 , n29814 );
xor ( n31121 , RI19a9b1c8_2604 , RI174720d8_1180);
not ( n11384 , n27689 );
and ( n11385 , n11384 , RI174720d8_1180);
and ( n11386 , n31121 , n27689 );
or ( n31122 , n11385 , n11386 );
xor ( n31123 , RI19aca9a0_2251 , RI174bc2c8_825);
not ( n11387 , n27689 );
and ( n11388 , n11387 , RI174bc2c8_825);
and ( n11389 , n31123 , n27689 );
or ( n31124 , n11388 , n11389 );
xor ( n31125 , n31122 , n31124 );
buf ( n31126 , RI1738d100_2068);
xor ( n31127 , n31125 , n31126 );
buf ( n31128 , RI173d5df0_1713);
xor ( n31129 , n31127 , n31128 );
buf ( n31130 , RI1744d8c8_1358);
xor ( n31131 , n31129 , n31130 );
xor ( n31132 , n31120 , n31131 );
buf ( n31133 , RI173df198_1668);
xor ( n31134 , n31133 , n30427 );
xor ( n31135 , n31134 , n29364 );
not ( n31136 , n31135 );
xor ( n31137 , n30052 , n28904 );
xor ( n31138 , n31137 , n29291 );
and ( n31139 , n31136 , n31138 );
xor ( n31140 , n31132 , n31139 );
xor ( n31141 , n31119 , n31140 );
xor ( n31142 , RI19aa0b50_2563 , RI17485890_1085);
not ( n11390 , n27689 );
and ( n11391 , n11390 , RI17485890_1085);
and ( n11392 , n31142 , n27689 );
or ( n31143 , n11391 , n11392 );
xor ( n31144 , RI19acf8d8_2214 , RI1750b930_730);
not ( n11393 , n27689 );
and ( n11394 , n11393 , RI1750b930_730);
and ( n11395 , n31144 , n27689 );
or ( n31145 , n11394 , n11395 );
xor ( n31146 , n31143 , n31145 );
buf ( n31147 , RI173a08b8_1973);
xor ( n31148 , n31146 , n31147 );
buf ( n31149 , RI173e95a8_1618);
xor ( n31150 , n31148 , n31149 );
buf ( n31151 , RI17461080_1263);
xor ( n31152 , n31150 , n31151 );
xor ( n31153 , n30343 , n31152 );
xor ( n31154 , RI19ab48a8_2419 , RI174a2a80_943);
not ( n11396 , n27689 );
and ( n11397 , n11396 , RI174a2a80_943);
and ( n11398 , n31154 , n27689 );
or ( n31155 , n11397 , n11398 );
buf ( n31156 , RI17334528_2186);
xor ( n31157 , n31155 , n31156 );
buf ( n31158 , RI173bdaa8_1831);
xor ( n31159 , n31157 , n31158 );
buf ( n31160 , RI17406798_1476);
xor ( n31161 , n31159 , n31160 );
xor ( n31162 , n31161 , n27768 );
xor ( n31163 , n31153 , n31162 );
xor ( n31164 , n30215 , n29573 );
xor ( n31165 , n31164 , n30758 );
not ( n31166 , n31165 );
xor ( n31167 , n30363 , n28684 );
xor ( n31168 , n31167 , n28279 );
and ( n31169 , n31166 , n31168 );
xor ( n31170 , n31163 , n31169 );
xor ( n31171 , n31141 , n31170 );
xor ( n31172 , RI19a8f8a0_2686 , RI17464ed8_1244);
not ( n11399 , n27689 );
and ( n11400 , n11399 , RI17464ed8_1244);
and ( n11401 , n31172 , n27689 );
or ( n31173 , n11400 , n11401 );
xor ( n31174 , RI19ac0158_2331 , RI174adbb0_889);
not ( n11402 , n27689 );
and ( n11403 , n11402 , RI174adbb0_889);
and ( n11404 , n31174 , n27689 );
or ( n31175 , n11403 , n11404 );
xor ( n31176 , n31173 , n31175 );
buf ( n31177 , RI1733f310_2133);
xor ( n31178 , n31176 , n31177 );
xor ( n31179 , n31178 , n30760 );
xor ( n31180 , n31179 , n29522 );
xor ( n31181 , n28064 , n31180 );
xor ( n31182 , RI19aa3418_2543 , RI17482410_1101);
not ( n11405 , n27689 );
and ( n11406 , n11405 , RI17482410_1101);
and ( n11407 , n31182 , n27689 );
or ( n31183 , n11406 , n11407 );
xor ( n31184 , RI19a846f8_2763 , RI175066b0_746);
not ( n11408 , n27689 );
and ( n11409 , n11408 , RI175066b0_746);
and ( n11410 , n31184 , n27689 );
or ( n31185 , n11409 , n11410 );
xor ( n31186 , n31183 , n31185 );
buf ( n31187 , RI1739d0f0_1990);
xor ( n31188 , n31186 , n31187 );
buf ( n31189 , RI173e6128_1634);
xor ( n31190 , n31188 , n31189 );
buf ( n31191 , RI1745dc00_1279);
xor ( n31192 , n31190 , n31191 );
xor ( n31193 , n31181 , n31192 );
xor ( n31194 , n28052 , n29694 );
xor ( n31195 , n31194 , n30457 );
not ( n31196 , n31195 );
xor ( n31197 , n27763 , n29639 );
xor ( n31198 , n31197 , n30233 );
and ( n31199 , n31196 , n31198 );
xor ( n31200 , n31193 , n31199 );
xor ( n31201 , n31171 , n31200 );
xor ( n31202 , n28308 , n27989 );
xor ( n31203 , n31202 , n28001 );
buf ( n31204 , RI173cfb68_1743);
xor ( n31205 , n31204 , n27844 );
xor ( n31206 , n31205 , n30691 );
not ( n31207 , n31206 );
buf ( n31208 , RI1744d238_1360);
xor ( n31209 , n31208 , n28741 );
xor ( n31210 , n31209 , n28096 );
and ( n31211 , n31207 , n31210 );
xor ( n31212 , n31203 , n31211 );
xor ( n31213 , n31201 , n31212 );
xor ( n31214 , n31103 , n31213 );
xor ( n31215 , n28851 , n30306 );
xor ( n31216 , n31215 , n30548 );
xor ( n31217 , n29311 , n30665 );
xor ( n31218 , RI19a9ad18_2606 , RI17471a48_1182);
not ( n11411 , n27689 );
and ( n11412 , n11411 , RI17471a48_1182);
and ( n11413 , n31218 , n27689 );
or ( n31219 , n11412 , n11413 );
xor ( n31220 , RI19aca4f0_2253 , RI174bb878_827);
not ( n11414 , n27689 );
and ( n11415 , n11414 , RI174bb878_827);
and ( n11416 , n31220 , n27689 );
or ( n31221 , n11415 , n11416 );
xor ( n31222 , n31219 , n31221 );
xor ( n31223 , n31222 , n28730 );
buf ( n31224 , RI173d5760_1715);
xor ( n31225 , n31223 , n31224 );
xor ( n31226 , n31225 , n31208 );
xor ( n31227 , n31217 , n31226 );
not ( n31228 , n31227 );
xor ( n31229 , RI19ac5108_2291 , RI174caff8_779);
not ( n11417 , n27689 );
and ( n11418 , n11417 , RI174caff8_779);
and ( n11419 , n31229 , n27689 );
or ( n31230 , n11418 , n11419 );
xor ( n31231 , n31230 , n30427 );
xor ( n31232 , n31231 , n29364 );
and ( n31233 , n31228 , n31232 );
xor ( n31234 , n31216 , n31233 );
xor ( n31235 , n30016 , n28647 );
xor ( n31236 , n31235 , n28659 );
xor ( n31237 , RI19aa1438_2558 , RI174865b0_1081);
not ( n11420 , n27689 );
and ( n11421 , n11420 , RI174865b0_1081);
and ( n11422 , n31237 , n27689 );
or ( n31238 , n11421 , n11422 );
xor ( n31239 , RI19a82538_2778 , RI1750cdd0_726);
not ( n11423 , n27689 );
and ( n11424 , n11423 , RI1750cdd0_726);
and ( n11425 , n31239 , n27689 );
or ( n31240 , n11424 , n11425 );
xor ( n31241 , n31238 , n31240 );
buf ( n31242 , RI173a15d8_1969);
xor ( n31243 , n31241 , n31242 );
buf ( n31244 , RI173ea2c8_1614);
xor ( n31245 , n31243 , n31244 );
buf ( n31246 , RI1746a0e0_1219);
xor ( n31247 , n31245 , n31246 );
xor ( n31248 , n28409 , n31247 );
xor ( n31249 , n31248 , n27885 );
not ( n31250 , n31249 );
xor ( n31251 , n28621 , n28327 );
xor ( n31252 , n31251 , n28339 );
and ( n31253 , n31250 , n31252 );
xor ( n31254 , n31236 , n31253 );
xor ( n31255 , n31234 , n31254 );
xor ( n31256 , n30442 , n28956 );
xor ( n31257 , n31256 , n29995 );
xor ( n31258 , n31219 , n28741 );
xor ( n31259 , n31258 , n28096 );
not ( n31260 , n31259 );
xor ( n31261 , n30201 , n29561 );
xor ( n31262 , n31261 , n29573 );
and ( n31263 , n31260 , n31262 );
xor ( n31264 , n31257 , n31263 );
xor ( n31265 , n31255 , n31264 );
xor ( n31266 , n28159 , n27738 );
xor ( n31267 , n31266 , n29259 );
xor ( n31268 , n28707 , n29935 );
xor ( n31269 , RI19a8d8c0_2700 , RI174693c0_1223);
not ( n11426 , n27689 );
and ( n11427 , n11426 , RI174693c0_1223);
and ( n11428 , n31269 , n27689 );
or ( n31270 , n11427 , n11428 );
xor ( n31271 , RI19abe808_2345 , RI174b2098_868);
not ( n11429 , n27689 );
and ( n11430 , n11429 , RI174b2098_868);
and ( n11431 , n31271 , n27689 );
or ( n31272 , n11430 , n11431 );
xor ( n31273 , n31270 , n31272 );
buf ( n31274 , RI173437f8_2112);
xor ( n31275 , n31273 , n31274 );
buf ( n31276 , RI173ccd78_1757);
xor ( n31277 , n31275 , n31276 );
buf ( n31278 , RI17444bb0_1401);
xor ( n31279 , n31277 , n31278 );
xor ( n31280 , n31268 , n31279 );
not ( n31281 , n31280 );
xor ( n31282 , n28512 , n29724 );
xor ( n31283 , RI19a96740_2637 , RI17479d88_1142);
not ( n11432 , n27689 );
and ( n11433 , n11432 , RI17479d88_1142);
and ( n11434 , n31283 , n27689 );
or ( n31284 , n11433 , n11434 );
xor ( n31285 , RI19ac6620_2282 , RI174c86b8_787);
not ( n11435 , n27689 );
and ( n11436 , n11435 , RI174c86b8_787);
and ( n11437 , n31285 , n27689 );
or ( n31286 , n11436 , n11437 );
xor ( n31287 , n31284 , n31286 );
buf ( n31288 , RI17394a68_2031);
xor ( n31289 , n31287 , n31288 );
xor ( n31290 , n31289 , n28906 );
xor ( n31291 , n31290 , n30729 );
xor ( n31292 , n31282 , n31291 );
and ( n31293 , n31281 , n31292 );
xor ( n31294 , n31267 , n31293 );
xor ( n31295 , n31265 , n31294 );
buf ( n31296 , RI1744d580_1359);
xor ( n31297 , n31296 , n29011 );
xor ( n31298 , n31297 , n27964 );
xor ( n31299 , RI19a9ce60_2591 , RI17471070_1185);
not ( n11438 , n27689 );
and ( n11439 , n11438 , RI17471070_1185);
and ( n11440 , n31299 , n27689 );
or ( n31300 , n11439 , n11440 );
xor ( n31301 , RI19acbe40_2240 , RI174ba900_830);
not ( n11441 , n27689 );
and ( n11442 , n11441 , RI174ba900_830);
and ( n11443 , n31301 , n27689 );
or ( n31302 , n11442 , n11443 );
xor ( n31303 , n31300 , n31302 );
buf ( n31304 , RI1738c098_2073);
xor ( n31305 , n31303 , n31304 );
buf ( n31306 , RI173d4d88_1718);
xor ( n31307 , n31305 , n31306 );
buf ( n31308 , RI1744c860_1363);
xor ( n31309 , n31307 , n31308 );
xor ( n31310 , n30274 , n31309 );
xor ( n31311 , n31310 , n29519 );
not ( n31312 , n31311 );
xor ( n31313 , n27757 , n29639 );
xor ( n31314 , n31313 , n30233 );
and ( n31315 , n31312 , n31314 );
xor ( n31316 , n31298 , n31315 );
xor ( n31317 , n31295 , n31316 );
xor ( n31318 , n31214 , n31317 );
not ( n31319 , n31318 );
not ( n31320 , n28628 );
and ( n31321 , n31320 , n28482 );
xor ( n31322 , n29503 , n31321 );
xor ( n31323 , n31322 , n29610 );
xor ( n31324 , n28116 , n30233 );
xor ( n31325 , n31324 , n30243 );
xor ( n31326 , n30621 , n28519 );
xor ( n31327 , n31326 , n28304 );
not ( n31328 , n31327 );
and ( n31329 , n31328 , n28840 );
xor ( n31330 , n31325 , n31329 );
or ( n31331 , RI1753a460_587 , RI17539218_590);
or ( n31332 , n31331 , RI175379b8_594);
or ( n31333 , n31332 , RI175373a0_595);
or ( n31334 , n31333 , RI17536770_597);
xor ( n31335 , n31330 , n31334 );
xor ( n31336 , n28318 , n31065 );
xor ( n31337 , n31336 , n31076 );
xor ( n31338 , n29228 , n30780 );
xor ( n31339 , n31338 , n28043 );
not ( n31340 , n31339 );
and ( n31341 , n31340 , n28905 );
xor ( n31342 , n31337 , n31341 );
xor ( n31343 , n31335 , n31342 );
xor ( n31344 , n30236 , n28250 );
xor ( n31345 , n31344 , n28262 );
xor ( n31346 , n30276 , n31309 );
xor ( n31347 , n31346 , n29519 );
not ( n31348 , n31347 );
and ( n31349 , n31348 , n28957 );
xor ( n31350 , n31345 , n31349 );
xor ( n31351 , n31343 , n31350 );
xor ( n31352 , RI19ab6090_2408 , RI174a16d0_949);
not ( n11444 , n27689 );
and ( n11445 , n11444 , RI174a16d0_949);
and ( n11446 , n31352 , n27689 );
or ( n31353 , n11445 , n11446 );
xor ( n31354 , n31353 , n28291 );
xor ( n31355 , n31354 , n29781 );
xor ( n31356 , n31272 , n30717 );
xor ( n31357 , RI19a97b68_2628 , RI17478348_1150);
not ( n11447 , n27689 );
and ( n11448 , n11447 , RI17478348_1150);
and ( n11449 , n31357 , n27689 );
or ( n31358 , n11448 , n11449 );
xor ( n31359 , RI19ac7958_2273 , RI174c5d78_795);
not ( n11450 , n27689 );
and ( n11451 , n11450 , RI174c5d78_795);
and ( n11452 , n31359 , n27689 );
or ( n31360 , n11451 , n11452 );
xor ( n31361 , n31358 , n31360 );
buf ( n31362 , RI17393028_2039);
xor ( n31363 , n31361 , n31362 );
buf ( n31364 , RI173dbd18_1684);
xor ( n31365 , n31363 , n31364 );
buf ( n31366 , RI174537f0_1329);
xor ( n31367 , n31365 , n31366 );
xor ( n31368 , n31356 , n31367 );
not ( n31369 , n31368 );
and ( n31370 , n31369 , n29013 );
xor ( n31371 , n31355 , n31370 );
xor ( n31372 , n31351 , n31371 );
xor ( n31373 , n30926 , n27752 );
xor ( n31374 , n31373 , n27764 );
xor ( n31375 , n30940 , n29586 );
xor ( n31376 , n31375 , n28355 );
not ( n31377 , n31376 );
and ( n31378 , n31377 , n29069 );
xor ( n31379 , n31374 , n31378 );
xor ( n31380 , n31372 , n31379 );
xor ( n31381 , n31323 , n31380 );
and ( n31382 , n31319 , n31381 );
xor ( n31383 , n31054 , n31382 );
not ( n11453 , n29614 );
and ( n11454 , n11453 , RI17336940_2175);
and ( n11455 , n31383 , n29614 );
or ( n31384 , n11454 , n11455 );
not ( n11456 , RI1754c610_2);
and ( n11457 , n11456 , n31384 );
and ( n11458 , C0 , RI1754c610_2);
or ( n31385 , n11457 , n11458 );
buf ( n31386 , n31385 );
buf ( n31387 , RI17514990_702);
xor ( n31388 , n28889 , n30066 );
xor ( n31389 , n31388 , n30007 );
buf ( n31390 , RI17410860_1427);
xor ( n31391 , RI19ab8f70_2388 , RI1749e250_965);
not ( n11459 , n27689 );
and ( n11460 , n11459 , RI1749e250_965);
and ( n11461 , n31391 , n27689 );
or ( n31392 , n11460 , n11461 );
buf ( n31393 , RI175323f0_610);
xor ( n31394 , n31392 , n31393 );
buf ( n31395 , RI173b9278_1853);
xor ( n31396 , n31394 , n31395 );
buf ( n31397 , RI17401f68_1498);
xor ( n31398 , n31396 , n31397 );
xor ( n31399 , n31398 , n29451 );
xor ( n31400 , n31390 , n31399 );
xor ( n31401 , n31400 , n29561 );
not ( n31402 , n31401 );
xor ( n31403 , n29481 , n28450 );
xor ( n31404 , n31403 , n30789 );
and ( n31405 , n31402 , n31404 );
xor ( n31406 , n31389 , n31405 );
buf ( n31407 , RI173a1c68_1967);
xor ( n31408 , n31407 , n27897 );
xor ( n31409 , n31408 , n27858 );
xor ( n31410 , n29034 , n30399 );
xor ( n31411 , n31410 , n29532 );
not ( n31412 , n31411 );
buf ( n31413 , RI173d9270_1697);
xor ( n31414 , RI19aae980_2464 , RI1748ef80_1039);
not ( n11462 , n27689 );
and ( n11463 , n11462 , RI1748ef80_1039);
and ( n11464 , n31414 , n27689 );
or ( n31415 , n11463 , n11464 );
xor ( n31416 , n31415 , n29803 );
buf ( n31417 , RI173a9c60_1928);
xor ( n31418 , n31416 , n31417 );
buf ( n31419 , RI173f2950_1573);
xor ( n31420 , n31418 , n31419 );
buf ( n31421 , RI174c1a70_808);
xor ( n31422 , n31420 , n31421 );
xor ( n31423 , n31413 , n31422 );
xor ( n31424 , n31423 , n29011 );
and ( n31425 , n31412 , n31424 );
xor ( n31426 , n31409 , n31425 );
xor ( n31427 , n29623 , n30799 );
xor ( n31428 , n31427 , n28148 );
xor ( n31429 , n29418 , n27870 );
xor ( n31430 , n31429 , n28174 );
not ( n31431 , n31430 );
xor ( n31432 , n29050 , n28027 );
xor ( n31433 , n31432 , n29827 );
and ( n31434 , n31431 , n31433 );
xor ( n31435 , n31428 , n31434 );
xor ( n31436 , n31426 , n31435 );
xor ( n31437 , n30776 , n29438 );
xor ( n31438 , n31437 , n29449 );
not ( n31439 , n31389 );
and ( n31440 , n31439 , n31401 );
xor ( n31441 , n31438 , n31440 );
xor ( n31442 , n31436 , n31441 );
xor ( n31443 , n28642 , n30271 );
xor ( n31444 , n31443 , n30283 );
xor ( n31445 , RI19a9af70_2605 , RI17471d90_1181);
not ( n11465 , n27689 );
and ( n11466 , n11465 , RI17471d90_1181);
and ( n11467 , n31445 , n27689 );
or ( n31446 , n11466 , n11467 );
xor ( n31447 , RI19aca748_2252 , RI174bbda0_826);
not ( n11468 , n27689 );
and ( n11469 , n11468 , RI174bbda0_826);
and ( n11470 , n31447 , n27689 );
or ( n31448 , n11469 , n11470 );
xor ( n31449 , n31446 , n31448 );
xor ( n31450 , n31449 , n29000 );
buf ( n31451 , RI173d5aa8_1714);
xor ( n31452 , n31450 , n31451 );
xor ( n31453 , n31452 , n31296 );
xor ( n31454 , n28093 , n31453 );
xor ( n31455 , RI19aaeea8_2462 , RI1748f610_1037);
not ( n11471 , n27689 );
and ( n11472 , n11471 , RI1748f610_1037);
and ( n11473 , n31455 , n27689 );
or ( n31456 , n11472 , n11473 );
xor ( n31457 , n31456 , n28424 );
buf ( n31458 , RI173aa2f0_1926);
xor ( n31459 , n31457 , n31458 );
buf ( n31460 , RI173f2fe0_1571);
xor ( n31461 , n31459 , n31460 );
xor ( n31462 , n31461 , n27953 );
xor ( n31463 , n31454 , n31462 );
not ( n31464 , n31463 );
xor ( n31465 , n30414 , n30901 );
xor ( n31466 , RI19ab2b98_2434 , RI174a72b0_921);
not ( n11474 , n27689 );
and ( n11475 , n11474 , RI174a72b0_921);
and ( n11476 , n31466 , n27689 );
or ( n31467 , n11475 , n11476 );
buf ( n31468 , RI17338a10_2165);
xor ( n31469 , n31467 , n31468 );
buf ( n31470 , RI173c1f90_1810);
xor ( n31471 , n31469 , n31470 );
buf ( n31472 , RI1740ac80_1455);
xor ( n31473 , n31471 , n31472 );
buf ( n31474 , RI174bdc90_820);
xor ( n31475 , n31473 , n31474 );
xor ( n31476 , n31465 , n31475 );
and ( n31477 , n31464 , n31476 );
xor ( n31478 , n31444 , n31477 );
xor ( n31479 , n31442 , n31478 );
xor ( n31480 , RI19aaad80_2489 , RI17494818_1012);
not ( n11477 , n27689 );
and ( n11478 , n11477 , RI17494818_1012);
and ( n11479 , n31480 , n27689 );
or ( n31481 , n11478 , n11479 );
xor ( n31482 , n31481 , n30736 );
buf ( n31483 , RI173af4f8_1901);
xor ( n31484 , n31482 , n31483 );
buf ( n31485 , RI173f81e8_1546);
xor ( n31486 , n31484 , n31485 );
xor ( n31487 , n31486 , n30580 );
xor ( n31488 , n29301 , n31487 );
xor ( n31489 , RI19a8d668_2701 , RI17469078_1224);
not ( n11480 , n27689 );
and ( n11481 , n11480 , RI17469078_1224);
and ( n11482 , n31489 , n27689 );
or ( n31490 , n11481 , n11482 );
xor ( n31491 , n31490 , n28705 );
buf ( n31492 , RI173434b0_2113);
xor ( n31493 , n31491 , n31492 );
buf ( n31494 , RI173cca30_1758);
xor ( n31495 , n31493 , n31494 );
buf ( n31496 , RI17415a68_1402);
xor ( n31497 , n31495 , n31496 );
xor ( n31498 , n31488 , n31497 );
xor ( n31499 , n31276 , n30717 );
xor ( n31500 , n31499 , n31367 );
not ( n31501 , n31500 );
xor ( n31502 , n28758 , n30823 );
xor ( n31503 , n31502 , n30934 );
and ( n31504 , n31501 , n31503 );
xor ( n31505 , n31498 , n31504 );
xor ( n31506 , n31479 , n31505 );
xor ( n31507 , n31406 , n31506 );
xor ( n31508 , RI19aaeb60_2463 , RI1748f2c8_1038);
not ( n11483 , n27689 );
and ( n11484 , n11483 , RI1748f2c8_1038);
and ( n11485 , n31508 , n27689 );
or ( n31509 , n11484 , n11485 );
xor ( n31510 , n31509 , n28085 );
buf ( n31511 , RI173a9fa8_1927);
xor ( n31512 , n31510 , n31511 );
buf ( n31513 , RI173f2c98_1572);
xor ( n31514 , n31512 , n31513 );
buf ( n31515 , RI174c5328_797);
xor ( n31516 , n31514 , n31515 );
xor ( n31517 , n29813 , n31516 );
xor ( n31518 , RI19a91100_2675 , RI17463b28_1250);
not ( n11486 , n27689 );
and ( n11487 , n11486 , RI17463b28_1250);
and ( n11488 , n31518 , n27689 );
or ( n31519 , n11487 , n11488 );
xor ( n31520 , RI19ac1490_2320 , RI174ac800_895);
not ( n11489 , n27689 );
and ( n11490 , n11489 , RI174ac800_895);
and ( n11491 , n31520 , n27689 );
or ( n31521 , n11490 , n11491 );
xor ( n31522 , n31519 , n31521 );
buf ( n31523 , RI1733df60_2139);
xor ( n31524 , n31522 , n31523 );
buf ( n31525 , RI173c74e0_1784);
xor ( n31526 , n31524 , n31525 );
buf ( n31527 , RI174101d0_1429);
xor ( n31528 , n31526 , n31527 );
xor ( n31529 , n31517 , n31528 );
xor ( n31530 , n28441 , n29975 );
xor ( n31531 , n31530 , n28759 );
not ( n31532 , n31531 );
xor ( n31533 , n29414 , n27870 );
xor ( n31534 , n31533 , n28174 );
and ( n31535 , n31532 , n31534 );
xor ( n31536 , n31529 , n31535 );
buf ( n31537 , RI17499d68_986);
xor ( n31538 , n31537 , n28367 );
xor ( n31539 , n31538 , n29952 );
xor ( n31540 , RI19aabcf8_2483 , RI17492400_1023);
not ( n11492 , n27689 );
and ( n11493 , n11492 , RI17492400_1023);
and ( n11494 , n31540 , n27689 );
or ( n31541 , n11493 , n11494 );
xor ( n31542 , n31541 , n28673 );
xor ( n31543 , n31542 , n28684 );
not ( n31544 , n31543 );
xor ( n31545 , n29154 , n29037 );
xor ( n31546 , n31545 , n31180 );
and ( n31547 , n31544 , n31546 );
xor ( n31548 , n31539 , n31547 );
xor ( n31549 , n31536 , n31548 );
xor ( n31550 , RI19ab92b8_2387 , RI1749e8e0_963);
not ( n11495 , n27689 );
and ( n11496 , n11495 , RI1749e8e0_963);
and ( n11497 , n31550 , n27689 );
or ( n31551 , n11496 , n11497 );
buf ( n31552 , RI17532e40_608);
xor ( n31553 , n31551 , n31552 );
buf ( n31554 , RI173b9908_1851);
xor ( n31555 , n31553 , n31554 );
buf ( n31556 , RI174025f8_1496);
xor ( n31557 , n31555 , n31556 );
xor ( n31558 , n31557 , n28855 );
xor ( n31559 , n29473 , n31558 );
xor ( n31560 , n31559 , n29025 );
xor ( n31561 , n28750 , n30823 );
xor ( n31562 , n31561 , n30934 );
not ( n31563 , n31562 );
xor ( n31564 , n28255 , n29270 );
xor ( n31565 , n31564 , n30066 );
and ( n31566 , n31563 , n31565 );
xor ( n31567 , n31560 , n31566 );
xor ( n31568 , n31549 , n31567 );
buf ( n31569 , RI173a95d0_1930);
xor ( n31570 , n31569 , n30321 );
xor ( n31571 , n31570 , n30332 );
xor ( n31572 , n28216 , n30457 );
xor ( n31573 , RI19abef88_2341 , RI174af5f0_881);
not ( n11498 , n27689 );
and ( n11499 , n11498 , RI174af5f0_881);
and ( n11500 , n31573 , n27689 );
or ( n31574 , n11499 , n11500 );
xor ( n31575 , n30256 , n31574 );
buf ( n31576 , RI17340d50_2125);
xor ( n31577 , n31575 , n31576 );
buf ( n31578 , RI173ca2d0_1770);
xor ( n31579 , n31577 , n31578 );
buf ( n31580 , RI17413308_1414);
xor ( n31581 , n31579 , n31580 );
xor ( n31582 , n31572 , n31581 );
not ( n31583 , n31582 );
xor ( n31584 , n30144 , n30918 );
xor ( n31585 , RI19a97208_2632 , RI17476f98_1156);
not ( n11501 , n27689 );
and ( n11502 , n11501 , RI17476f98_1156);
and ( n11503 , n31585 , n27689 );
or ( n31586 , n11502 , n11503 );
xor ( n31587 , RI19ac6ff8_2277 , RI174c43b0_800);
not ( n11504 , n27689 );
and ( n11505 , n11504 , RI174c43b0_800);
and ( n11506 , n31587 , n27689 );
or ( n31588 , n11505 , n11506 );
xor ( n31589 , n31586 , n31588 );
xor ( n31590 , n31589 , n30167 );
buf ( n31591 , RI173dacb0_1689);
xor ( n31592 , n31590 , n31591 );
buf ( n31593 , RI17452788_1334);
xor ( n31594 , n31592 , n31593 );
xor ( n31595 , n31584 , n31594 );
and ( n31596 , n31583 , n31595 );
xor ( n31597 , n31571 , n31596 );
xor ( n31598 , n31568 , n31597 );
xor ( n31599 , n27751 , n29628 );
xor ( n31600 , n31599 , n29639 );
xor ( n31601 , RI19a9d9a0_2587 , RI1748b470_1057);
not ( n11507 , n27689 );
and ( n11508 , n11507 , RI1748b470_1057);
and ( n11509 , n31601 , n27689 );
or ( n31602 , n11508 , n11509 );
xor ( n31603 , RI19a936f8_2658 , RI1747cec0_1127);
not ( n11510 , n27689 );
and ( n11511 , n11510 , RI1747cec0_1127);
and ( n11512 , n31603 , n27689 );
or ( n31604 , n11511 , n11512 );
xor ( n31605 , RI19ac3920_2302 , RI174cd410_772);
not ( n11513 , n27689 );
and ( n11514 , n11513 , RI174cd410_772);
and ( n11515 , n31605 , n27689 );
or ( n31606 , n11514 , n11515 );
xor ( n31607 , n31604 , n31606 );
buf ( n31608 , RI17397ba0_2016);
xor ( n31609 , n31607 , n31608 );
buf ( n31610 , RI173e0890_1661);
xor ( n31611 , n31609 , n31610 );
buf ( n31612 , RI174586b0_1305);
xor ( n31613 , n31611 , n31612 );
xor ( n31614 , n31602 , n31613 );
xor ( n31615 , n31614 , n28438 );
not ( n31616 , n31615 );
xor ( n31617 , n30408 , n30901 );
xor ( n31618 , n31617 , n31475 );
and ( n31619 , n31616 , n31618 );
xor ( n31620 , n31600 , n31619 );
xor ( n31621 , n31598 , n31620 );
xor ( n31622 , n31507 , n31621 );
xor ( n31623 , RI19aba398_2379 , RI1749c810_973);
not ( n11516 , n27689 );
and ( n11517 , n11516 , RI1749c810_973);
and ( n11518 , n31623 , n27689 );
or ( n31624 , n11517 , n11518 );
xor ( n31625 , n31624 , n29291 );
xor ( n31626 , RI19a92bb8_2663 , RI17462778_1256);
not ( n11519 , n27689 );
and ( n11520 , n11519 , RI17462778_1256);
and ( n11521 , n31626 , n27689 );
or ( n31627 , n11520 , n11521 );
xor ( n31628 , RI19ac2f48_2307 , RI174ab450_901);
not ( n11522 , n27689 );
and ( n11523 , n11522 , RI174ab450_901);
and ( n11524 , n31628 , n27689 );
or ( n31629 , n11523 , n11524 );
xor ( n31630 , n31627 , n31629 );
buf ( n31631 , RI1733cbb0_2145);
xor ( n31632 , n31630 , n31631 );
buf ( n31633 , RI173c6130_1790);
xor ( n31634 , n31632 , n31633 );
buf ( n31635 , RI1740ee20_1435);
xor ( n31636 , n31634 , n31635 );
xor ( n31637 , n31625 , n31636 );
not ( n31638 , n31637 );
xor ( n31639 , n29467 , n31558 );
xor ( n31640 , n31639 , n29025 );
and ( n31641 , n31638 , n31640 );
xor ( n31642 , n30582 , n31641 );
not ( n31643 , n30523 );
xor ( n31644 , n29167 , n28185 );
xor ( n31645 , n31644 , n28827 );
and ( n31646 , n31643 , n31645 );
xor ( n31647 , n30499 , n31646 );
not ( n31648 , n30553 );
xor ( n31649 , n28650 , n30283 );
xor ( n31650 , n31649 , n31089 );
and ( n31651 , n31648 , n31650 );
xor ( n31652 , n30550 , n31651 );
xor ( n31653 , n31647 , n31652 );
xor ( n31654 , n31653 , n30495 );
not ( n31655 , n30582 );
and ( n31656 , n31655 , n31637 );
xor ( n31657 , n30578 , n31656 );
xor ( n31658 , n31654 , n31657 );
not ( n31659 , n30601 );
xor ( n31660 , n29846 , n29421 );
xor ( n31661 , n31660 , n30643 );
and ( n31662 , n31659 , n31661 );
xor ( n31663 , n30597 , n31662 );
xor ( n31664 , n31658 , n31663 );
xor ( n31665 , n31642 , n31664 );
not ( n31666 , n30630 );
xor ( n31667 , n28050 , n29694 );
xor ( n31668 , n31667 , n30457 );
and ( n31669 , n31666 , n31668 );
xor ( n31670 , n30627 , n31669 );
not ( n31671 , n30669 );
xor ( n31672 , n29747 , n28313 );
xor ( n31673 , RI19a96e48_2634 , RI1747a760_1139);
not ( n11525 , n27689 );
and ( n11526 , n11525 , RI1747a760_1139);
and ( n11527 , n31673 , n27689 );
or ( n31674 , n11526 , n11527 );
xor ( n31675 , RI19ac6bc0_2279 , RI174c9630_784);
not ( n11528 , n27689 );
and ( n11529 , n11528 , RI174c9630_784);
and ( n11530 , n31675 , n27689 );
or ( n31676 , n11529 , n11530 );
xor ( n31677 , n31674 , n31676 );
buf ( n31678 , RI17395440_2028);
xor ( n31679 , n31677 , n31678 );
buf ( n31680 , RI173de130_1673);
xor ( n31681 , n31679 , n31680 );
buf ( n31682 , RI17455c08_1318);
xor ( n31683 , n31681 , n31682 );
xor ( n31684 , n31672 , n31683 );
and ( n31685 , n31671 , n31684 );
xor ( n31686 , n30666 , n31685 );
xor ( n31687 , n31670 , n31686 );
not ( n31688 , n30693 );
xor ( n31689 , n31033 , n30053 );
buf ( n31690 , RI1752fab0_618);
xor ( n31691 , n31624 , n31690 );
buf ( n31692 , RI173b7838_1861);
xor ( n31693 , n31691 , n31692 );
buf ( n31694 , RI17400528_1506);
xor ( n31695 , n31693 , n31694 );
buf ( n31696 , RI173d01f8_1741);
xor ( n31697 , n31695 , n31696 );
xor ( n31698 , n31689 , n31697 );
and ( n31699 , n31688 , n31698 );
xor ( n31700 , n30677 , n31699 );
xor ( n31701 , n31687 , n31700 );
not ( n31702 , n30725 );
buf ( n31703 , RI173967f0_2022);
xor ( n31704 , RI19a8b250_2717 , RI1746d218_1204);
not ( n11531 , n27689 );
and ( n11532 , n11531 , RI1746d218_1204);
and ( n11533 , n31704 , n27689 );
or ( n31705 , n11532 , n11533 );
xor ( n31706 , RI19abca80_2362 , RI174b5ef0_849);
not ( n11534 , n27689 );
and ( n11535 , n11534 , RI174b5ef0_849);
and ( n11536 , n31706 , n27689 );
or ( n31707 , n11535 , n11536 );
xor ( n31708 , n31705 , n31707 );
buf ( n31709 , RI17347650_2093);
xor ( n31710 , n31708 , n31709 );
buf ( n31711 , RI173d0f18_1737);
xor ( n31712 , n31710 , n31711 );
buf ( n31713 , RI17448a08_1382);
xor ( n31714 , n31712 , n31713 );
xor ( n31715 , n31703 , n31714 );
xor ( n31716 , n31715 , n28785 );
and ( n31717 , n31702 , n31716 );
xor ( n31718 , n30722 , n31717 );
xor ( n31719 , n31701 , n31718 );
not ( n31720 , n30738 );
xor ( n31721 , n28978 , n28081 );
xor ( n31722 , n31721 , n29248 );
and ( n31723 , n31720 , n31722 );
xor ( n31724 , n30733 , n31723 );
xor ( n31725 , n31719 , n31724 );
xor ( n31726 , n31665 , n31725 );
not ( n31727 , n31726 );
xor ( n31728 , RI19a9ed50_2578 , RI174896e8_1066);
not ( n11537 , n27689 );
and ( n11538 , n11537 , RI174896e8_1066);
and ( n11539 , n31728 , n27689 );
or ( n31729 , n11538 , n11539 );
xor ( n31730 , n31729 , n31114 );
xor ( n31731 , n31730 , n30415 );
xor ( n31732 , n28588 , n29187 );
xor ( n31733 , n31732 , n29724 );
not ( n31734 , n31733 );
buf ( n31735 , RI173bc6f8_1837);
xor ( n31736 , n31735 , n28291 );
xor ( n31737 , n31736 , n29781 );
and ( n31738 , n31734 , n31737 );
xor ( n31739 , n31731 , n31738 );
xor ( n31740 , RI19ab0000_2454 , RI1748d1f8_1048);
not ( n11540 , n27689 );
and ( n11541 , n11540 , RI1748d1f8_1048);
and ( n11542 , n31740 , n27689 );
or ( n31741 , n11541 , n11542 );
xor ( n31742 , RI19a887a8_2735 , RI17517d20_692);
not ( n11543 , n27689 );
and ( n11544 , n11543 , RI17517d20_692);
and ( n11545 , n31742 , n27689 );
or ( n31743 , n11544 , n11545 );
xor ( n31744 , n31741 , n31743 );
buf ( n31745 , RI173a8220_1936);
xor ( n31746 , n31744 , n31745 );
buf ( n31747 , RI173f0f10_1581);
xor ( n31748 , n31746 , n31747 );
buf ( n31749 , RI174ae588_886);
xor ( n31750 , n31748 , n31749 );
xor ( n31751 , n28492 , n31750 );
xor ( n31752 , n31751 , n30043 );
xor ( n31753 , n30418 , n31475 );
xor ( n31754 , RI19a954f8_2645 , RI1747bb10_1133);
not ( n11546 , n27689 );
and ( n11547 , n11546 , RI1747bb10_1133);
and ( n11548 , n31754 , n27689 );
or ( n31755 , n11547 , n11548 );
xor ( n31756 , RI19ac52e8_2290 , RI174cb520_778);
not ( n11549 , n27689 );
and ( n11550 , n11549 , RI174cb520_778);
and ( n11551 , n31756 , n27689 );
or ( n31757 , n11550 , n11551 );
xor ( n31758 , n31755 , n31757 );
xor ( n31759 , n31758 , n31703 );
buf ( n31760 , RI173df4e0_1667);
xor ( n31761 , n31759 , n31760 );
buf ( n31762 , RI17456fb8_1312);
xor ( n31763 , n31761 , n31762 );
xor ( n31764 , n31753 , n31763 );
not ( n31765 , n31764 );
xor ( n31766 , RI19ac6e18_2278 , RI174c3e88_801);
not ( n11552 , n27689 );
and ( n11553 , n11552 , RI174c3e88_801);
and ( n11554 , n31766 , n27689 );
or ( n31767 , n11553 , n11554 );
xor ( n31768 , n31767 , n30151 );
xor ( n31769 , n31768 , n31024 );
and ( n31770 , n31765 , n31769 );
xor ( n31771 , n31752 , n31770 );
buf ( n31772 , RI17487960_1075);
xor ( n31773 , n31772 , n30691 );
xor ( n31774 , n31773 , n30475 );
xor ( n31775 , n29028 , n30399 );
xor ( n31776 , n31775 , n29532 );
not ( n31777 , n31776 );
xor ( n31778 , n30659 , n28969 );
xor ( n31779 , n31778 , n28741 );
and ( n31780 , n31777 , n31779 );
xor ( n31781 , n31774 , n31780 );
xor ( n31782 , n31771 , n31781 );
xor ( n31783 , n31635 , n30986 );
xor ( n31784 , RI19a9d1a8_2590 , RI174713b8_1184);
not ( n11555 , n27689 );
and ( n11556 , n11555 , RI174713b8_1184);
and ( n11557 , n31784 , n27689 );
or ( n31785 , n11556 , n11557 );
xor ( n31786 , RI19acc020_2239 , RI174bae28_829);
not ( n11558 , n27689 );
and ( n11559 , n11558 , RI174bae28_829);
and ( n11560 , n31786 , n27689 );
or ( n31787 , n11559 , n11560 );
xor ( n31788 , n31785 , n31787 );
buf ( n31789 , RI1738c3e0_2072);
xor ( n31790 , n31788 , n31789 );
buf ( n31791 , RI173d50d0_1717);
xor ( n31792 , n31790 , n31791 );
buf ( n31793 , RI1744cba8_1362);
xor ( n31794 , n31792 , n31793 );
xor ( n31795 , n31783 , n31794 );
xor ( n31796 , n31755 , n31714 );
xor ( n31797 , n31796 , n28785 );
not ( n31798 , n31797 );
xor ( n31799 , RI19acc5c0_2236 , RI17514eb8_701);
not ( n11561 , n27689 );
and ( n11562 , n11561 , RI17514eb8_701);
and ( n11563 , n31799 , n27689 );
or ( n31800 , n11562 , n11563 );
xor ( n31801 , n31800 , n31613 );
xor ( n31802 , n31801 , n28438 );
and ( n31803 , n31798 , n31802 );
xor ( n31804 , n31795 , n31803 );
xor ( n31805 , n31782 , n31804 );
xor ( n31806 , n28838 , n28569 );
xor ( n31807 , n31806 , n29889 );
xor ( n31808 , n30210 , n29573 );
xor ( n31809 , n31808 , n30758 );
not ( n31810 , n31809 );
xor ( n31811 , n31574 , n29134 );
xor ( n31812 , n31811 , n27936 );
and ( n31813 , n31810 , n31812 );
xor ( n31814 , n31807 , n31813 );
xor ( n31815 , n31805 , n31814 );
buf ( n31816 , RI17457300_1311);
xor ( n31817 , RI19a8b4a8_2716 , RI1746d560_1203);
not ( n11564 , n27689 );
and ( n11565 , n11564 , RI1746d560_1203);
and ( n11566 , n31817 , n27689 );
or ( n31818 , n11565 , n11566 );
xor ( n31819 , n31818 , n29755 );
buf ( n31820 , RI17358cc0_2092);
xor ( n31821 , n31819 , n31820 );
buf ( n31822 , RI173d1278_1736);
xor ( n31823 , n31821 , n31822 );
buf ( n31824 , RI17448d50_1381);
xor ( n31825 , n31823 , n31824 );
xor ( n31826 , n31816 , n31825 );
xor ( n31827 , n31826 , n29586 );
not ( n31828 , n31731 );
and ( n31829 , n31828 , n31733 );
xor ( n31830 , n31827 , n31829 );
xor ( n31831 , n31815 , n31830 );
xor ( n31832 , n31739 , n31831 );
xor ( n31833 , n31588 , n30178 );
xor ( n31834 , n31833 , n30189 );
xor ( n31835 , RI19a97028_2633 , RI17476c50_1157);
not ( n11567 , n27689 );
and ( n11568 , n11567 , RI17476c50_1157);
and ( n11569 , n31835 , n27689 );
or ( n31836 , n11568 , n11569 );
xor ( n31837 , n31836 , n31767 );
buf ( n31838 , RI17391c78_2045);
xor ( n31839 , n31837 , n31838 );
buf ( n31840 , RI173da968_1690);
xor ( n31841 , n31839 , n31840 );
buf ( n31842 , RI17452440_1335);
xor ( n31843 , n31841 , n31842 );
xor ( n31844 , n31147 , n31843 );
xor ( n31845 , n31844 , n27779 );
not ( n31846 , n31845 );
xor ( n31847 , n31513 , n28096 );
xor ( n31848 , n31847 , n28107 );
and ( n31849 , n31846 , n31848 );
xor ( n31850 , n31834 , n31849 );
buf ( n31851 , RI17530f50_614);
xor ( n31852 , n31851 , n31422 );
xor ( n31853 , n31852 , n29011 );
xor ( n31854 , n30951 , n28355 );
xor ( n31855 , n31854 , n28367 );
not ( n31856 , n31855 );
xor ( n31857 , n29920 , n27791 );
xor ( n31858 , n31857 , n30706 );
and ( n31859 , n31856 , n31858 );
xor ( n31860 , n31853 , n31859 );
xor ( n31861 , n31850 , n31860 );
xor ( n31862 , RI19acc818_2235 , RI175153e0_700);
not ( n11570 , n27689 );
and ( n11571 , n11570 , RI175153e0_700);
and ( n11572 , n31862 , n27689 );
or ( n31863 , n11571 , n11572 );
xor ( n31864 , RI19a93950_2657 , RI1747d208_1126);
not ( n11573 , n27689 );
and ( n11574 , n11573 , RI1747d208_1126);
and ( n11575 , n31864 , n27689 );
or ( n31865 , n11574 , n11575 );
xor ( n31866 , RI19ac3b00_2301 , RI174cd938_771);
not ( n11576 , n27689 );
and ( n11577 , n11576 , RI174cd938_771);
and ( n11578 , n31866 , n27689 );
or ( n31867 , n11577 , n11578 );
xor ( n31868 , n31865 , n31867 );
buf ( n31869 , RI17397ee8_2015);
xor ( n31870 , n31868 , n31869 );
buf ( n31871 , RI173e0bd8_1660);
xor ( n31872 , n31870 , n31871 );
buf ( n31873 , RI174589f8_1304);
xor ( n31874 , n31872 , n31873 );
xor ( n31875 , n31863 , n31874 );
xor ( n31876 , n31875 , n30813 );
xor ( n31877 , n28861 , n30207 );
xor ( n31878 , n31877 , n30218 );
not ( n31879 , n31878 );
xor ( n31880 , n28460 , n29502 );
xor ( n31881 , n31880 , n29628 );
and ( n31882 , n31879 , n31881 );
xor ( n31883 , n31876 , n31882 );
xor ( n31884 , n31861 , n31883 );
xor ( n31885 , n30357 , n28684 );
xor ( n31886 , n31885 , n28279 );
xor ( n31887 , n28143 , n27726 );
xor ( n31888 , n31887 , n27738 );
not ( n31889 , n31888 );
xor ( n31890 , n30050 , n28904 );
xor ( n31891 , n31890 , n29291 );
and ( n31892 , n31889 , n31891 );
xor ( n31893 , n31886 , n31892 );
xor ( n31894 , n31884 , n31893 );
xor ( n31895 , n28832 , n28569 );
xor ( n31896 , n31895 , n29889 );
xor ( n31897 , n28623 , n28327 );
xor ( n31898 , n31897 , n28339 );
not ( n31899 , n31898 );
xor ( n31900 , RI19ab6900_2405 , RI174a20a8_946);
not ( n11579 , n27689 );
and ( n11580 , n11579 , RI174a20a8_946);
and ( n11581 , n31900 , n27689 );
or ( n31901 , n11580 , n11581 );
buf ( n31902 , RI17333b50_2189);
xor ( n31903 , n31901 , n31902 );
buf ( n31904 , RI173bd0d0_1834);
xor ( n31905 , n31903 , n31904 );
buf ( n31906 , RI17405dc0_1479);
xor ( n31907 , n31905 , n31906 );
buf ( n31908 , RI17408ef8_1464);
xor ( n31909 , n31907 , n31908 );
xor ( n31910 , n28377 , n31909 );
xor ( n31911 , RI19a99440_2617 , RI17476908_1158);
not ( n11582 , n27689 );
and ( n11583 , n11582 , RI17476908_1158);
and ( n11584 , n31911 , n27689 );
or ( n31912 , n11583 , n11584 );
xor ( n31913 , RI19ac8e70_2263 , RI174c3960_802);
not ( n11585 , n27689 );
and ( n11586 , n11585 , RI174c3960_802);
and ( n11587 , n31913 , n27689 );
or ( n31914 , n11586 , n11587 );
xor ( n31915 , n31912 , n31914 );
buf ( n31916 , RI17391930_2046);
xor ( n31917 , n31915 , n31916 );
buf ( n31918 , RI173da620_1691);
xor ( n31919 , n31917 , n31918 );
buf ( n31920 , RI174520f8_1336);
xor ( n31921 , n31919 , n31920 );
xor ( n31922 , n31910 , n31921 );
and ( n31923 , n31899 , n31922 );
xor ( n31924 , n31896 , n31923 );
xor ( n31925 , n31894 , n31924 );
xor ( n31926 , n31832 , n31925 );
and ( n31927 , n31727 , n31926 );
xor ( n31928 , n31622 , n31927 );
not ( n11588 , n29614 );
and ( n11589 , n11588 , RI173a0f48_1971);
and ( n11590 , n31928 , n29614 );
or ( n31929 , n11589 , n11590 );
not ( n11591 , RI1754c610_2);
and ( n11592 , n11591 , n31929 );
and ( n11593 , C0 , RI1754c610_2);
or ( n31930 , n11592 , n11593 );
buf ( n31931 , n31930 );
xor ( n31932 , n30856 , n30114 );
xor ( n31933 , n31932 , n30125 );
xor ( n31934 , n27692 , n28480 );
xor ( n31935 , n31934 , n27909 );
not ( n31936 , n31935 );
xor ( n31937 , n29774 , n28627 );
xor ( n31938 , n31937 , n30089 );
and ( n31939 , n31936 , n31938 );
xor ( n31940 , n31933 , n31939 );
xor ( n31941 , RI19aa4ed0_2530 , RI174813a8_1106);
not ( n11594 , n27689 );
and ( n11595 , n11594 , RI174813a8_1106);
and ( n11596 , n31941 , n27689 );
or ( n31942 , n11595 , n11596 );
xor ( n31943 , RI19a86318_2751 , RI17502e70_751);
not ( n11597 , n27689 );
and ( n11598 , n11597 , RI17502e70_751);
and ( n11599 , n31943 , n27689 );
or ( n31944 , n11598 , n11599 );
xor ( n31945 , n31942 , n31944 );
buf ( n31946 , RI1739c088_1995);
xor ( n31947 , n31945 , n31946 );
xor ( n31948 , n31947 , n29335 );
buf ( n31949 , RI1745cb98_1284);
xor ( n31950 , n31948 , n31949 );
xor ( n31951 , n29459 , n31950 );
xor ( n31952 , n31951 , n31558 );
xor ( n31953 , n30985 , n28659 );
xor ( n31954 , n31953 , n29148 );
not ( n31955 , n31954 );
xor ( n31956 , n30949 , n28355 );
xor ( n31957 , n31956 , n28367 );
and ( n31958 , n31955 , n31957 );
xor ( n31959 , n31952 , n31958 );
xor ( n31960 , RI19a8db18_2699 , RI17469708_1222);
not ( n11600 , n27689 );
and ( n11601 , n11600 , RI17469708_1222);
and ( n11602 , n31960 , n27689 );
or ( n31961 , n11601 , n11602 );
xor ( n31962 , RI19abe9e8_2344 , RI174b23e0_867);
not ( n11603 , n27689 );
and ( n11604 , n11603 , RI174b23e0_867);
and ( n11605 , n31962 , n27689 );
or ( n31963 , n11604 , n11605 );
xor ( n31964 , n31961 , n31963 );
buf ( n31965 , RI17343b40_2111);
xor ( n31966 , n31964 , n31965 );
buf ( n31967 , RI173cd0c0_1756);
xor ( n31968 , n31966 , n31967 );
xor ( n31969 , n31968 , n27875 );
xor ( n31970 , n31364 , n31969 );
xor ( n31971 , RI19aa17f8_2556 , RI17486c40_1079);
not ( n11606 , n27689 );
and ( n11607 , n11606 , RI17486c40_1079);
and ( n11608 , n31971 , n27689 );
or ( n31972 , n11607 , n11608 );
xor ( n31973 , RI19a82970_2776 , RI1750d820_724);
not ( n11609 , n27689 );
and ( n11610 , n11609 , RI1750d820_724);
and ( n11611 , n31973 , n27689 );
or ( n31974 , n11610 , n11611 );
xor ( n31975 , n31972 , n31974 );
xor ( n31976 , n31975 , n31407 );
xor ( n31977 , n31976 , n30192 );
xor ( n31978 , n31977 , n30975 );
xor ( n31979 , n31970 , n31978 );
xor ( n31980 , n29363 , n31763 );
xor ( n31981 , RI19aa90e8_2502 , RI17499048_990);
not ( n11612 , n27689 );
and ( n11613 , n11612 , RI17499048_990);
and ( n11614 , n31981 , n27689 );
or ( n31982 , n11613 , n11614 );
xor ( n31983 , n31982 , n28774 );
buf ( n31984 , RI173b3d28_1879);
xor ( n31985 , n31983 , n31984 );
buf ( n31986 , RI173fcd60_1523);
xor ( n31987 , n31985 , n31986 );
buf ( n31988 , RI173ade00_1908);
xor ( n31989 , n31987 , n31988 );
xor ( n31990 , n31980 , n31989 );
not ( n31991 , n31990 );
xor ( n31992 , n30772 , n29438 );
xor ( n31993 , n31992 , n29449 );
and ( n31994 , n31991 , n31993 );
xor ( n31995 , n31979 , n31994 );
xor ( n31996 , n31959 , n31995 );
xor ( n31997 , n30230 , n28160 );
xor ( n31998 , n31997 , n28250 );
xor ( n31999 , n29010 , n29814 );
xor ( n32000 , n31999 , n31131 );
not ( n32001 , n32000 );
xor ( n32002 , n28358 , n30522 );
xor ( n32003 , n31602 , n31800 );
buf ( n32004 , RI173a6498_1945);
xor ( n32005 , n32003 , n32004 );
buf ( n32006 , RI173ef188_1590);
xor ( n32007 , n32005 , n32006 );
buf ( n32008 , RI1749c180_975);
xor ( n32009 , n32007 , n32008 );
xor ( n32010 , n32002 , n32009 );
and ( n32011 , n32001 , n32010 );
xor ( n32012 , n31998 , n32011 );
xor ( n32013 , n31996 , n32012 );
xor ( n32014 , n30652 , n31794 );
xor ( n32015 , n32014 , n28969 );
not ( n32016 , n31933 );
and ( n32017 , n32016 , n31935 );
xor ( n32018 , n32015 , n32017 );
xor ( n32019 , n32013 , n32018 );
xor ( n32020 , n30175 , n31162 );
xor ( n32021 , n32020 , n29923 );
xor ( n32022 , n31612 , n29839 );
xor ( n32023 , RI19a9dbf8_2586 , RI1748b7b8_1056);
not ( n11615 , n27689 );
and ( n11616 , n11615 , RI1748b7b8_1056);
and ( n11617 , n32023 , n27689 );
or ( n32024 , n11616 , n11617 );
xor ( n32025 , n32024 , n31863 );
buf ( n32026 , RI173a67e0_1944);
xor ( n32027 , n32025 , n32026 );
buf ( n32028 , RI173ef4d0_1589);
xor ( n32029 , n32027 , n32028 );
buf ( n32030 , RI1749e598_964);
xor ( n32031 , n32029 , n32030 );
xor ( n32032 , n32022 , n32031 );
not ( n32033 , n32032 );
xor ( n32034 , RI19a95750_2644 , RI1747be58_1132);
not ( n11618 , n27689 );
and ( n11619 , n11618 , RI1747be58_1132);
and ( n11620 , n32034 , n27689 );
or ( n32035 , n11619 , n11620 );
xor ( n32036 , RI19ac5540_2289 , RI174cba48_777);
not ( n11621 , n27689 );
and ( n11622 , n11621 , RI174cba48_777);
and ( n11623 , n32036 , n27689 );
or ( n32037 , n11622 , n11623 );
xor ( n32038 , n32035 , n32037 );
buf ( n32039 , RI17396b38_2021);
xor ( n32040 , n32038 , n32039 );
buf ( n32041 , RI173df828_1666);
xor ( n32042 , n32040 , n32041 );
xor ( n32043 , n32042 , n31816 );
xor ( n32044 , n28776 , n32043 );
xor ( n32045 , n32044 , n30946 );
and ( n32046 , n32033 , n32045 );
xor ( n32047 , n32021 , n32046 );
xor ( n32048 , n32019 , n32047 );
xor ( n32049 , n31940 , n32048 );
xor ( n32050 , n30513 , n29062 );
xor ( n32051 , n32050 , n31613 );
xor ( n32052 , n31360 , n31969 );
xor ( n32053 , n32052 , n31978 );
not ( n32054 , n32053 );
xor ( n32055 , n31242 , n28727 );
xor ( n32056 , n32055 , n29387 );
and ( n32057 , n32054 , n32056 );
xor ( n32058 , n32051 , n32057 );
xor ( n32059 , n30022 , n27921 );
xor ( n32060 , n32059 , n28852 );
xor ( n32061 , n31393 , n29462 );
xor ( n32062 , n32061 , n29474 );
not ( n32063 , n32062 );
xor ( n32064 , n28445 , n29975 );
xor ( n32065 , n32064 , n28759 );
and ( n32066 , n32063 , n32065 );
xor ( n32067 , n32060 , n32066 );
xor ( n32068 , n32058 , n32067 );
xor ( n32069 , n31604 , n29839 );
xor ( n32070 , n32069 , n32031 );
xor ( n32071 , n29633 , n28148 );
xor ( n32072 , n32071 , n28160 );
not ( n32073 , n32072 );
xor ( n32074 , n28076 , n31192 );
xor ( n32075 , n32074 , n27700 );
and ( n32076 , n32073 , n32075 );
xor ( n32077 , n32070 , n32076 );
xor ( n32078 , n32068 , n32077 );
xor ( n32079 , n29227 , n30780 );
xor ( n32080 , n32079 , n28043 );
xor ( n32081 , n28332 , n31076 );
xor ( n32082 , RI19a991e8_2618 , RI174765c0_1159);
not ( n11624 , n27689 );
and ( n11625 , n11624 , RI174765c0_1159);
and ( n11626 , n32082 , n27689 );
or ( n32083 , n11625 , n11626 );
xor ( n32084 , RI19ac8c18_2264 , RI174c3438_803);
not ( n11627 , n27689 );
and ( n11628 , n11627 , RI174c3438_803);
and ( n11629 , n32084 , n27689 );
or ( n32085 , n11628 , n11629 );
xor ( n32086 , n32083 , n32085 );
xor ( n32087 , n32086 , n28369 );
buf ( n32088 , RI173da2d8_1692);
xor ( n32089 , n32087 , n32088 );
buf ( n32090 , RI17451db0_1337);
xor ( n32091 , n32089 , n32090 );
xor ( n32092 , n32081 , n32091 );
not ( n32093 , n32092 );
xor ( n32094 , n28500 , n30043 );
xor ( n32095 , n32094 , n30053 );
and ( n32096 , n32093 , n32095 );
xor ( n32097 , n32080 , n32096 );
xor ( n32098 , n32078 , n32097 );
xor ( n32099 , n29577 , n29767 );
xor ( n32100 , n32099 , n30510 );
xor ( n32101 , n30851 , n30114 );
xor ( n32102 , n32101 , n30125 );
not ( n32103 , n32102 );
xor ( n32104 , n30914 , n30348 );
xor ( n32105 , n32104 , n30178 );
and ( n32106 , n32103 , n32105 );
xor ( n32107 , n32100 , n32106 );
xor ( n32108 , n32098 , n32107 );
xor ( n32109 , n32049 , n32108 );
xor ( n32110 , n27729 , n28543 );
xor ( n32111 , RI19aafcb8_2455 , RI1748ceb0_1049);
not ( n11630 , n27689 );
and ( n11631 , n11630 , RI1748ceb0_1049);
and ( n11632 , n32111 , n27689 );
or ( n32112 , n11631 , n11632 );
xor ( n32113 , RI19a86de0_2746 , RI175177f8_693);
not ( n11633 , n27689 );
and ( n11634 , n11633 , RI175177f8_693);
and ( n11635 , n32113 , n27689 );
or ( n32114 , n11634 , n11635 );
xor ( n32115 , n32112 , n32114 );
xor ( n32116 , n32115 , n30844 );
buf ( n32117 , RI173f0bc8_1582);
xor ( n32118 , n32116 , n32117 );
buf ( n32119 , RI174ac170_897);
xor ( n32120 , n32118 , n32119 );
xor ( n32121 , n32110 , n32120 );
xor ( n32122 , RI19a9d658_2588 , RI1748b128_1058);
not ( n11636 , n27689 );
and ( n11637 , n11636 , RI1748b128_1058);
and ( n11638 , n32122 , n27689 );
or ( n32123 , n11637 , n11638 );
xor ( n32124 , RI19acc3e0_2237 , RI17514990_702);
not ( n11639 , n27689 );
and ( n11640 , n11639 , RI17514990_702);
and ( n11641 , n32124 , n27689 );
or ( n32125 , n11640 , n11641 );
xor ( n32126 , n32123 , n32125 );
buf ( n32127 , RI173a6150_1946);
xor ( n32128 , n32126 , n32127 );
xor ( n32129 , n32128 , n30576 );
xor ( n32130 , n32129 , n31537 );
xor ( n32131 , n29820 , n32130 );
xor ( n32132 , RI19ab11d0_2445 , RI174a89a8_914);
not ( n11642 , n27689 );
and ( n11643 , n11642 , RI174a89a8_914);
and ( n11644 , n32132 , n27689 );
or ( n32133 , n11643 , n11644 );
buf ( n32134 , RI1733a108_2158);
xor ( n32135 , n32133 , n32134 );
xor ( n32136 , n32135 , n29941 );
buf ( n32137 , RI1740c378_1448);
xor ( n32138 , n32136 , n32137 );
buf ( n32139 , RI173cda98_1753);
xor ( n32140 , n32138 , n32139 );
xor ( n32141 , n32131 , n32140 );
not ( n32142 , n32141 );
xor ( n32143 , n29074 , n30643 );
xor ( n32144 , n32143 , n29176 );
and ( n32145 , n32142 , n32144 );
xor ( n32146 , n32121 , n32145 );
xor ( n32147 , n29160 , n29037 );
xor ( n32148 , n32147 , n31180 );
xor ( n32149 , n29085 , n28493 );
xor ( n32150 , n32149 , n28505 );
not ( n32151 , n32150 );
xor ( n32152 , n30530 , n29752 );
xor ( n32153 , n32152 , n27833 );
and ( n32154 , n32151 , n32153 );
xor ( n32155 , n32148 , n32154 );
xor ( n32156 , n29638 , n28148 );
xor ( n32157 , n32156 , n28160 );
xor ( n32158 , n30092 , n29910 );
xor ( n32159 , RI19ab6ae0_2404 , RI174a23f0_945);
not ( n11645 , n27689 );
and ( n11646 , n11645 , RI174a23f0_945);
and ( n11647 , n32159 , n27689 );
or ( n32160 , n11646 , n11647 );
buf ( n32161 , RI17333e98_2188);
xor ( n32162 , n32160 , n32161 );
buf ( n32163 , RI173bd418_1833);
xor ( n32164 , n32162 , n32163 );
xor ( n32165 , n32164 , n30128 );
buf ( n32166 , RI1740b310_1453);
xor ( n32167 , n32165 , n32166 );
xor ( n32168 , n32158 , n32167 );
not ( n32169 , n32168 );
xor ( n32170 , n28845 , n30306 );
xor ( n32171 , n32170 , n30548 );
and ( n32172 , n32169 , n32171 );
xor ( n32173 , n32157 , n32172 );
xor ( n32174 , n32155 , n32173 );
xor ( n32175 , n27908 , n29235 );
xor ( n32176 , n32175 , n30294 );
xor ( n32177 , n28496 , n30043 );
xor ( n32178 , n32177 , n30053 );
not ( n32179 , n32178 );
xor ( n32180 , RI19a85760_2756 , RI17500f80_757);
not ( n11648 , n27689 );
and ( n11649 , n11648 , RI17500f80_757);
and ( n11650 , n32180 , n27689 );
or ( n32181 , n11649 , n11650 );
xor ( n32182 , n32181 , n31100 );
xor ( n32183 , n32182 , n31422 );
and ( n32184 , n32179 , n32183 );
xor ( n32185 , n32176 , n32184 );
xor ( n32186 , n32174 , n32185 );
xor ( n32187 , n29951 , n32009 );
xor ( n32188 , n32187 , n30164 );
xor ( n32189 , RI19aacbf8_2477 , RI174937b0_1017);
not ( n11651 , n27689 );
and ( n11652 , n11651 , RI174937b0_1017);
and ( n11653 , n32189 , n27689 );
or ( n32190 , n11652 , n11653 );
xor ( n32191 , RI19ab8778_2392 , RI175217d0_662);
not ( n11654 , n27689 );
and ( n11655 , n11654 , RI175217d0_662);
and ( n11656 , n32191 , n27689 );
or ( n32192 , n11655 , n11656 );
xor ( n32193 , n32190 , n32192 );
buf ( n32194 , RI173ae490_1906);
xor ( n32195 , n32193 , n32194 );
buf ( n32196 , RI173f7180_1551);
xor ( n32197 , n32195 , n32196 );
buf ( n32198 , RI17334870_2185);
xor ( n32199 , n32197 , n32198 );
xor ( n32200 , n31068 , n32199 );
xor ( n32201 , n32200 , n28380 );
not ( n32202 , n32201 );
xor ( n32203 , RI19ab5640_2413 , RI174a3e30_937);
not ( n11657 , n27689 );
and ( n11658 , n11657 , RI174a3e30_937);
and ( n11659 , n32203 , n27689 );
or ( n32204 , n11658 , n11659 );
xor ( n32205 , n32204 , n29679 );
xor ( n32206 , n32205 , n28789 );
buf ( n32207 , RI17407b48_1470);
xor ( n32208 , n32206 , n32207 );
xor ( n32209 , n32208 , n30251 );
xor ( n32210 , n29392 , n32209 );
xor ( n32211 , n32210 , n30389 );
and ( n32212 , n32202 , n32211 );
xor ( n32213 , n32188 , n32212 );
xor ( n32214 , n32186 , n32213 );
xor ( n32215 , n28903 , n30007 );
xor ( n32216 , n32215 , n30017 );
not ( n32217 , n32121 );
and ( n32218 , n32217 , n32141 );
xor ( n32219 , n32216 , n32218 );
xor ( n32220 , n32214 , n32219 );
xor ( n32221 , n32146 , n32220 );
xor ( n32222 , n31676 , n28001 );
xor ( n32223 , n32222 , n30114 );
xor ( n32224 , n28924 , n30537 );
xor ( n32225 , n32224 , n30842 );
not ( n32226 , n32225 );
buf ( n32227 , RI173f5dd0_1557);
xor ( n32228 , n32227 , n28673 );
xor ( n32229 , n32228 , n28684 );
and ( n32230 , n32226 , n32229 );
xor ( n32231 , n32223 , n32230 );
xor ( n32232 , n28217 , n30457 );
xor ( n32233 , n32232 , n31581 );
xor ( n32234 , n31631 , n30986 );
xor ( n32235 , n32234 , n31794 );
not ( n32236 , n32235 );
buf ( n32237 , RI173de478_1672);
xor ( n32238 , RI19a8a530_2722 , RI1746be68_1210);
not ( n11660 , n27689 );
and ( n11661 , n11660 , RI1746be68_1210);
and ( n11662 , n32238 , n27689 );
or ( n32239 , n11661 , n11662 );
xor ( n32240 , RI19abc198_2367 , RI174b4b40_855);
not ( n11663 , n27689 );
and ( n11664 , n11663 , RI174b4b40_855);
and ( n11665 , n32240 , n27689 );
or ( n32241 , n11664 , n11665 );
xor ( n32242 , n32239 , n32241 );
buf ( n32243 , RI173462a0_2099);
xor ( n32244 , n32242 , n32243 );
xor ( n32245 , n32244 , n31204 );
buf ( n32246 , RI17447658_1388);
xor ( n32247 , n32245 , n32246 );
xor ( n32248 , n32237 , n32247 );
xor ( n32249 , RI19a9eaf8_2579 , RI174893a0_1067);
not ( n11666 , n27689 );
and ( n11667 , n11666 , RI174893a0_1067);
and ( n11668 , n32249 , n27689 );
or ( n32250 , n11667 , n11668 );
xor ( n32251 , n32250 , n30680 );
buf ( n32252 , RI173a43c8_1955);
xor ( n32253 , n32251 , n32252 );
buf ( n32254 , RI173ed0b8_1600);
xor ( n32255 , n32253 , n32254 );
xor ( n32256 , n32255 , n31772 );
xor ( n32257 , n32248 , n32256 );
and ( n32258 , n32236 , n32257 );
xor ( n32259 , n32233 , n32258 );
xor ( n32260 , n32231 , n32259 );
xor ( n32261 , n29325 , n31226 );
xor ( n32262 , n32261 , n31516 );
xor ( n32263 , n28322 , n31065 );
xor ( n32264 , n32263 , n31076 );
not ( n32265 , n32264 );
xor ( n32266 , n28104 , n31462 );
xor ( n32267 , RI19a91358_2674 , RI17463e70_1249);
not ( n11669 , n27689 );
and ( n11670 , n11669 , RI17463e70_1249);
and ( n11671 , n32267 , n27689 );
or ( n32268 , n11670 , n11671 );
xor ( n32269 , n32268 , n30875 );
buf ( n32270 , RI1733e2a8_2138);
xor ( n32271 , n32269 , n32270 );
buf ( n32272 , RI173c7828_1783);
xor ( n32273 , n32271 , n32272 );
buf ( n32274 , RI17410518_1428);
xor ( n32275 , n32273 , n32274 );
xor ( n32276 , n32266 , n32275 );
and ( n32277 , n32265 , n32276 );
xor ( n32278 , n32262 , n32277 );
xor ( n32279 , n32260 , n32278 );
xor ( n32280 , n28805 , n29409 );
xor ( n32281 , n32280 , n29421 );
xor ( n32282 , RI19a915b0_2673 , RI174641b8_1248);
not ( n11672 , n27689 );
and ( n11673 , n11672 , RI174641b8_1248);
and ( n11674 , n32282 , n27689 );
or ( n32283 , n11673 , n11674 );
xor ( n32284 , RI19ac1850_2318 , RI174ace90_893);
not ( n11675 , n27689 );
and ( n11676 , n11675 , RI174ace90_893);
and ( n11677 , n32284 , n27689 );
or ( n32285 , n11676 , n11677 );
xor ( n32286 , n32283 , n32285 );
buf ( n32287 , RI1733e5f0_2137);
xor ( n32288 , n32286 , n32287 );
buf ( n32289 , RI173c7b70_1782);
xor ( n32290 , n32288 , n32289 );
xor ( n32291 , n32290 , n31390 );
xor ( n32292 , n29341 , n32291 );
xor ( n32293 , n32292 , n30207 );
not ( n32294 , n32293 );
xor ( n32295 , n31189 , n29544 );
xor ( n32296 , n32295 , n28480 );
and ( n32297 , n32294 , n32296 );
xor ( n32298 , n32281 , n32297 );
xor ( n32299 , n32279 , n32298 );
xor ( n32300 , n29945 , n32009 );
xor ( n32301 , n32300 , n30164 );
xor ( n32302 , n28180 , n29211 );
xor ( n32303 , n32302 , n28557 );
not ( n32304 , n32303 );
xor ( n32305 , n28516 , n29724 );
xor ( n32306 , n32305 , n31291 );
and ( n32307 , n32304 , n32306 );
xor ( n32308 , n32301 , n32307 );
xor ( n32309 , n32299 , n32308 );
xor ( n32310 , n32221 , n32309 );
not ( n32311 , n32310 );
xor ( n32312 , n30083 , n28339 );
xor ( n32313 , n32312 , n29910 );
xor ( n32314 , RI19a98d38_2620 , RI17475f30_1161);
not ( n11678 , n27689 );
and ( n11679 , n11678 , RI17475f30_1161);
and ( n11680 , n32314 , n27689 );
or ( n32315 , n11679 , n11680 );
xor ( n32316 , RI19ac8768_2266 , RI174c29e8_805);
not ( n11681 , n27689 );
and ( n11682 , n11681 , RI174c29e8_805);
and ( n11683 , n32316 , n27689 );
or ( n32317 , n11682 , n11683 );
xor ( n32318 , n32315 , n32317 );
xor ( n32319 , n32318 , n29770 );
buf ( n32320 , RI173d9c48_1694);
xor ( n32321 , n32319 , n32320 );
buf ( n32322 , RI17451720_1339);
xor ( n32323 , n32321 , n32322 );
xor ( n32324 , n31060 , n32323 );
xor ( n32325 , n32324 , n32199 );
not ( n32326 , n32325 );
xor ( n32327 , n28656 , n30283 );
xor ( n32328 , n32327 , n31089 );
and ( n32329 , n32326 , n32328 );
xor ( n32330 , n32313 , n32329 );
xor ( n32331 , n30860 , n30125 );
xor ( n32332 , n32331 , n31114 );
not ( n32333 , n32313 );
and ( n32334 , n32333 , n32325 );
xor ( n32335 , n32332 , n32334 );
xor ( n32336 , n29453 , n31950 );
xor ( n32337 , n32336 , n31558 );
xor ( n32338 , n31690 , n29291 );
xor ( n32339 , n32338 , n31636 );
not ( n32340 , n32339 );
xor ( n32341 , n30422 , n31475 );
xor ( n32342 , n32341 , n31763 );
and ( n32343 , n32340 , n32342 );
xor ( n32344 , n32337 , n32343 );
xor ( n32345 , n32335 , n32344 );
xor ( n32346 , n31106 , n30889 );
xor ( n32347 , n32346 , n30901 );
xor ( n32348 , n29579 , n29767 );
xor ( n32349 , n32348 , n30510 );
not ( n32350 , n32349 );
xor ( n32351 , n31511 , n28096 );
xor ( n32352 , n32351 , n28107 );
and ( n32353 , n32350 , n32352 );
xor ( n32354 , n32347 , n32353 );
xor ( n32355 , n32345 , n32354 );
xor ( n32356 , RI19aaf088_2461 , RI1748f958_1036);
not ( n11684 , n27689 );
and ( n11685 , n11684 , RI1748f958_1036);
and ( n11686 , n32356 , n27689 );
or ( n32357 , n11685 , n11686 );
xor ( n32358 , RI19a23a38_2791 , RI1751b5d8_681);
not ( n11687 , n27689 );
and ( n11688 , n11687 , RI1751b5d8_681);
and ( n11689 , n32358 , n27689 );
or ( n32359 , n11688 , n11689 );
xor ( n32360 , n32357 , n32359 );
buf ( n32361 , RI173aa638_1925);
xor ( n32362 , n32360 , n32361 );
buf ( n32363 , RI173f3328_1570);
xor ( n32364 , n32362 , n32363 );
buf ( n32365 , RI174cc498_775);
xor ( n32366 , n32364 , n32365 );
xor ( n32367 , n27967 , n32366 );
xor ( n32368 , n32367 , n32291 );
xor ( n32369 , n28036 , n29449 );
xor ( n32370 , n32369 , n29694 );
not ( n32371 , n32370 );
xor ( n32372 , n31869 , n29964 );
xor ( n32373 , RI19a9de50_2585 , RI1748bb00_1055);
not ( n11690 , n27689 );
and ( n11691 , n11690 , RI1748bb00_1055);
and ( n11692 , n32373 , n27689 );
or ( n32374 , n11691 , n11692 );
xor ( n32375 , RI19acc9f8_2234 , RI17515908_699);
not ( n11693 , n27689 );
and ( n11694 , n11693 , RI17515908_699);
and ( n11695 , n32375 , n27689 );
or ( n32376 , n11694 , n11695 );
xor ( n32377 , n32374 , n32376 );
buf ( n32378 , RI173a6b28_1943);
xor ( n32379 , n32377 , n32378 );
buf ( n32380 , RI173ef818_1588);
xor ( n32381 , n32379 , n32380 );
xor ( n32382 , n32381 , n29479 );
xor ( n32383 , n32372 , n32382 );
and ( n32384 , n32371 , n32383 );
xor ( n32385 , n32368 , n32384 );
xor ( n32386 , n32355 , n32385 );
xor ( n32387 , n27824 , n31683 );
xor ( n32388 , n32387 , n30857 );
xor ( n32389 , n28193 , n29855 );
xor ( n32390 , n32389 , n29079 );
not ( n32391 , n32390 );
xor ( n32392 , RI19ab0c30_2448 , RI1751f8e0_668);
not ( n11696 , n27689 );
and ( n11697 , n11696 , RI1751f8e0_668);
and ( n11698 , n32392 , n27689 );
or ( n32393 , n11697 , n11698 );
xor ( n32394 , n31541 , n32393 );
xor ( n32395 , n32394 , n28662 );
xor ( n32396 , n32395 , n32227 );
buf ( n32397 , RI17527ef0_642);
xor ( n32398 , n32396 , n32397 );
xor ( n32399 , n29129 , n32398 );
xor ( n32400 , n32399 , n30364 );
and ( n32401 , n32391 , n32400 );
xor ( n32402 , n32388 , n32401 );
xor ( n32403 , n32386 , n32402 );
xor ( n32404 , n32330 , n32403 );
xor ( n32405 , n29788 , n30089 );
xor ( n32406 , n32405 , n30101 );
xor ( n32407 , n29516 , n30655 );
xor ( n32408 , n32407 , n30665 );
not ( n32409 , n32408 );
xor ( n32410 , n30232 , n28160 );
xor ( n32411 , n32410 , n28250 );
and ( n32412 , n32409 , n32411 );
xor ( n32413 , n32406 , n32412 );
xor ( n32414 , n31709 , n30332 );
xor ( n32415 , n32414 , n32043 );
xor ( n32416 , RI19a8f3f0_2688 , RI17468358_1228);
not ( n11699 , n27689 );
and ( n11700 , n11699 , RI17468358_1228);
and ( n11701 , n32416 , n27689 );
or ( n32417 , n11700 , n11701 );
xor ( n32418 , RI19abfd98_2333 , RI174b1030_873);
not ( n11702 , n27689 );
and ( n11703 , n11702 , RI174b1030_873);
and ( n11704 , n32418 , n27689 );
or ( n32419 , n11703 , n11704 );
xor ( n32420 , n32417 , n32419 );
buf ( n32421 , RI17342790_2117);
xor ( n32422 , n32420 , n32421 );
buf ( n32423 , RI173cbd10_1762);
xor ( n32424 , n32422 , n32423 );
buf ( n32425 , RI17414d48_1406);
xor ( n32426 , n32424 , n32425 );
xor ( n32427 , n31918 , n32426 );
xor ( n32428 , n32427 , n31152 );
not ( n32429 , n32428 );
xor ( n32430 , n27832 , n31683 );
xor ( n32431 , n32430 , n30857 );
and ( n32432 , n32429 , n32431 );
xor ( n32433 , n32415 , n32432 );
xor ( n32434 , n32413 , n32433 );
xor ( n32435 , n31458 , n27964 );
xor ( n32436 , n32435 , n27975 );
xor ( n32437 , n32137 , n29952 );
xor ( n32438 , n32437 , n29964 );
not ( n32439 , n32438 );
xor ( n32440 , n30006 , n30567 );
xor ( n32441 , n32440 , n28647 );
and ( n32442 , n32439 , n32441 );
xor ( n32443 , n32436 , n32442 );
xor ( n32444 , n32434 , n32443 );
xor ( n32445 , n29485 , n28450 );
xor ( n32446 , n32445 , n30789 );
xor ( n32447 , n28134 , n30243 );
xor ( n32448 , n32447 , n31750 );
not ( n32449 , n32448 );
xor ( n32450 , RI19a9ff20_2569 , RI17487ca8_1074);
not ( n11705 , n27689 );
and ( n11706 , n11705 , RI17487ca8_1074);
and ( n11707 , n32450 , n27689 );
or ( n32451 , n11706 , n11707 );
xor ( n32452 , RI19aceac8_2220 , RI1750f1e8_719);
not ( n11708 , n27689 );
and ( n11709 , n11708 , RI1750f1e8_719);
and ( n11710 , n32452 , n27689 );
or ( n32453 , n11709 , n11710 );
xor ( n32454 , n32451 , n32453 );
xor ( n32455 , n32454 , n28572 );
buf ( n32456 , RI173eb9c0_1607);
xor ( n32457 , n32455 , n32456 );
buf ( n32458 , RI17477cb8_1152);
xor ( n32459 , n32457 , n32458 );
xor ( n32460 , n29210 , n32459 );
xor ( n32461 , n32460 , n30616 );
and ( n32462 , n32449 , n32461 );
xor ( n32463 , n32446 , n32462 );
xor ( n32464 , n32444 , n32463 );
xor ( n32465 , n28679 , n29711 );
xor ( n32466 , n32465 , n30443 );
buf ( n32467 , RI17333178_2192);
xor ( n32468 , n31353 , n32467 );
xor ( n32469 , n32468 , n31735 );
xor ( n32470 , n32469 , n29891 );
buf ( n32471 , RI174022b0_1497);
xor ( n32472 , n32470 , n32471 );
xor ( n32473 , n28699 , n32472 );
xor ( n32474 , n32473 , n32323 );
not ( n32475 , n32474 );
buf ( n32476 , RI17456c70_1313);
xor ( n32477 , n32476 , n30427 );
xor ( n32478 , n32477 , n29364 );
and ( n32479 , n32475 , n32478 );
xor ( n32480 , n32466 , n32479 );
xor ( n32481 , n32464 , n32480 );
xor ( n32482 , n32404 , n32481 );
and ( n32483 , n32311 , n32482 );
xor ( n32484 , n32109 , n32483 );
not ( n11711 , n29614 );
and ( n11712 , n11711 , RI173b2978_1885);
and ( n11713 , n32484 , n29614 );
or ( n32485 , n11712 , n11713 );
not ( n11714 , RI1754c610_2);
and ( n11715 , n11714 , n32485 );
and ( n11716 , C0 , RI1754c610_2);
or ( n32486 , n11715 , n11716 );
buf ( n32487 , n32486 );
not ( n11717 , n27683 );
and ( n11718 , n11717 , RI19a8d8c0_2700);
and ( n11719 , RI19a97820_2629 , n27683 );
or ( n32488 , n11718 , n11719 );
not ( n11720 , RI1754c610_2);
and ( n11721 , n11720 , n32488 );
and ( n11722 , C0 , RI1754c610_2);
or ( n32489 , n11721 , n11722 );
buf ( n32490 , n32489 );
not ( n11723 , n27683 );
and ( n11724 , n11723 , RI19aa3aa8_2540);
and ( n11725 , RI19aadfa8_2468 , n27683 );
or ( n32491 , n11724 , n11725 );
not ( n11726 , RI1754c610_2);
and ( n11727 , n11726 , n32491 );
and ( n11728 , C0 , RI1754c610_2);
or ( n32492 , n11727 , n11728 );
buf ( n32493 , n32492 );
xor ( n32494 , n30345 , n31152 );
xor ( n32495 , n32494 , n31162 );
xor ( n32496 , n28683 , n29711 );
xor ( n32497 , n32496 , n30443 );
not ( n32498 , n32497 );
xor ( n32499 , n31519 , n28107 );
xor ( n32500 , RI19a9b678_2602 , RI17472420_1179);
not ( n11729 , n27689 );
and ( n11730 , n11729 , RI17472420_1179);
and ( n11731 , n32500 , n27689 );
or ( n32501 , n11730 , n11731 );
xor ( n32502 , RI19acabf8_2250 , RI174bc7f0_824);
not ( n11732 , n27689 );
and ( n11733 , n11732 , RI174bc7f0_824);
and ( n11734 , n32502 , n27689 );
or ( n32503 , n11733 , n11734 );
xor ( n32504 , n32501 , n32503 );
buf ( n32505 , RI1738d448_2067);
xor ( n32506 , n32504 , n32505 );
buf ( n32507 , RI173d6138_1712);
xor ( n32508 , n32506 , n32507 );
buf ( n32509 , RI1744dc10_1357);
xor ( n32510 , n32508 , n32509 );
xor ( n32511 , n32499 , n32510 );
and ( n32512 , n32498 , n32511 );
xor ( n32513 , n32495 , n32512 );
xor ( n32514 , n28780 , n32043 );
xor ( n32515 , n32514 , n30946 );
not ( n32516 , n32495 );
and ( n32517 , n32516 , n32497 );
xor ( n32518 , n32515 , n32517 );
xor ( n32519 , n29469 , n31558 );
xor ( n32520 , n32519 , n29025 );
xor ( n32521 , n28024 , n30956 );
xor ( n32522 , n32521 , n32130 );
not ( n32523 , n32522 );
buf ( n32524 , RI1745b7e8_1290);
xor ( n32525 , n32524 , n31100 );
xor ( n32526 , n32525 , n31422 );
and ( n32527 , n32523 , n32526 );
xor ( n32528 , n32520 , n32527 );
xor ( n32529 , n32518 , n32528 );
xor ( n32530 , n28413 , n31247 );
xor ( n32531 , n32530 , n27885 );
xor ( n32532 , n27697 , n28480 );
xor ( n32533 , n32532 , n27909 );
not ( n32534 , n32533 );
xor ( n32535 , n28338 , n31076 );
xor ( n32536 , n32535 , n32091 );
and ( n32537 , n32534 , n32536 );
xor ( n32538 , n32531 , n32537 );
xor ( n32539 , n32529 , n32538 );
xor ( n32540 , n30290 , n28043 );
xor ( n32541 , n32540 , n28055 );
xor ( n32542 , n30371 , n28279 );
xor ( n32543 , n32542 , n28291 );
not ( n32544 , n32543 );
xor ( n32545 , n30065 , n29105 );
xor ( n32546 , n32545 , n30567 );
and ( n32547 , n32544 , n32546 );
xor ( n32548 , n32541 , n32547 );
xor ( n32549 , n32539 , n32548 );
buf ( n32550 , RI173c1900_1812);
xor ( n32551 , n32550 , n30475 );
xor ( n32552 , n32551 , n30487 );
xor ( n32553 , n30424 , n31475 );
xor ( n32554 , n32553 , n31763 );
not ( n32555 , n32554 );
xor ( n32556 , n29345 , n32291 );
xor ( n32557 , n32556 , n30207 );
and ( n32558 , n32555 , n32557 );
xor ( n32559 , n32552 , n32558 );
xor ( n32560 , n32549 , n32559 );
xor ( n32561 , n32513 , n32560 );
xor ( n32562 , n28955 , n27948 );
xor ( n32563 , n32562 , n28702 );
xor ( n32564 , n32268 , n27975 );
xor ( n32565 , n32564 , n29346 );
not ( n32566 , n32565 );
xor ( n32567 , n28020 , n30956 );
xor ( n32568 , n32567 , n32130 );
and ( n32569 , n32566 , n32568 );
xor ( n32570 , n32563 , n32569 );
xor ( n32571 , n29331 , n31226 );
xor ( n32572 , n32571 , n31516 );
xor ( n32573 , n28191 , n29855 );
xor ( n32574 , n32573 , n29079 );
not ( n32575 , n32574 );
xor ( n32576 , n30912 , n30348 );
xor ( n32577 , n32576 , n30178 );
and ( n32578 , n32575 , n32577 );
xor ( n32579 , n32572 , n32578 );
xor ( n32580 , n32570 , n32579 );
xor ( n32581 , n28379 , n31909 );
xor ( n32582 , n32581 , n31921 );
xor ( n32583 , n29337 , n32291 );
xor ( n32584 , n32583 , n30207 );
not ( n32585 , n32584 );
xor ( n32586 , n31185 , n29544 );
xor ( n32587 , n32586 , n28480 );
and ( n32588 , n32585 , n32587 );
xor ( n32589 , n32582 , n32588 );
xor ( n32590 , n32580 , n32589 );
xor ( n32591 , n31037 , n30053 );
xor ( n32592 , n32591 , n31697 );
xor ( n32593 , n29403 , n27858 );
xor ( n32594 , n32593 , n27870 );
not ( n32595 , n32594 );
xor ( n32596 , n32241 , n27844 );
xor ( n32597 , n32596 , n30691 );
and ( n32598 , n32595 , n32597 );
xor ( n32599 , n32592 , n32598 );
xor ( n32600 , n32590 , n32599 );
xor ( n32601 , n29560 , n29474 );
xor ( n32602 , RI19aa53f8_2528 , RI17481a38_1104);
not ( n11735 , n27689 );
and ( n11736 , n11735 , RI17481a38_1104);
and ( n11737 , n32602 , n27689 );
or ( n32603 , n11736 , n11737 );
xor ( n32604 , RI19a86750_2749 , RI175038c0_749);
not ( n11738 , n27689 );
and ( n11739 , n11738 , RI175038c0_749);
and ( n11740 , n32604 , n27689 );
or ( n32605 , n11739 , n11740 );
xor ( n32606 , n32603 , n32605 );
buf ( n32607 , RI1739c718_1993);
xor ( n32608 , n32606 , n32607 );
xor ( n32609 , n32608 , n29014 );
buf ( n32610 , RI1745d228_1282);
xor ( n32611 , n32609 , n32610 );
xor ( n32612 , n32601 , n32611 );
xor ( n32613 , n28087 , n31453 );
xor ( n32614 , n32613 , n31462 );
not ( n32615 , n32614 );
xor ( n32616 , n30059 , n29105 );
xor ( n32617 , n32616 , n30567 );
and ( n32618 , n32615 , n32617 );
xor ( n32619 , n32612 , n32618 );
xor ( n32620 , n32600 , n32619 );
xor ( n32621 , n32561 , n32620 );
xor ( n32622 , n27737 , n28543 );
xor ( n32623 , n32622 , n32120 );
xor ( n32624 , n30130 , n28392 );
xor ( n32625 , n32624 , n30918 );
not ( n32626 , n32625 );
and ( n32627 , n32626 , n32233 );
xor ( n32628 , n32623 , n32627 );
xor ( n32629 , n29531 , n27819 );
xor ( n32630 , n32629 , n30594 );
not ( n32631 , n32630 );
xor ( n32632 , n30035 , n28892 );
xor ( n32633 , n32632 , n28904 );
and ( n32634 , n32631 , n32633 );
xor ( n32635 , n32229 , n32634 );
not ( n32636 , n32623 );
and ( n32637 , n32636 , n32625 );
xor ( n32638 , n32257 , n32637 );
xor ( n32639 , n32635 , n32638 );
xor ( n32640 , n28042 , n29449 );
xor ( n32641 , n32640 , n29694 );
not ( n32642 , n32641 );
xor ( n32643 , n28895 , n30007 );
xor ( n32644 , n32643 , n30017 );
and ( n32645 , n32642 , n32644 );
xor ( n32646 , n32276 , n32645 );
xor ( n32647 , n32639 , n32646 );
xor ( n32648 , n28437 , n32031 );
xor ( n32649 , n32648 , n29975 );
not ( n32650 , n32649 );
xor ( n32651 , n31901 , n30101 );
xor ( n32652 , n32651 , n32426 );
and ( n32653 , n32650 , n32652 );
xor ( n32654 , n32296 , n32653 );
xor ( n32655 , n32647 , n32654 );
xor ( n32656 , n28646 , n30271 );
xor ( n32657 , n32656 , n30283 );
not ( n32658 , n32657 );
xor ( n32659 , n28128 , n30243 );
xor ( n32660 , n32659 , n31750 );
and ( n32661 , n32658 , n32660 );
xor ( n32662 , n32306 , n32661 );
xor ( n32663 , n32655 , n32662 );
xor ( n32664 , n32628 , n32663 );
xor ( n32665 , n29998 , n30567 );
xor ( n32666 , n32665 , n28647 );
xor ( n32667 , RI19ac46b8_2296 , RI174c9b58_783);
not ( n11741 , n27689 );
and ( n11742 , n11741 , RI174c9b58_783);
and ( n11743 , n32667 , n27689 );
or ( n32668 , n11742 , n11743 );
xor ( n32669 , n32668 , n32247 );
xor ( n32670 , n32669 , n32256 );
not ( n32671 , n32670 );
xor ( n32672 , n27828 , n31683 );
xor ( n32673 , n32672 , n30857 );
and ( n32674 , n32671 , n32673 );
xor ( n32675 , n32666 , n32674 );
xor ( n32676 , n30339 , n31152 );
xor ( n32677 , n32676 , n31162 );
xor ( n32678 , n29127 , n32398 );
xor ( n32679 , n32678 , n30364 );
not ( n32680 , n32679 );
xor ( n32681 , n29143 , n31089 );
xor ( n32682 , n32681 , n31100 );
and ( n32683 , n32680 , n32682 );
xor ( n32684 , n32677 , n32683 );
xor ( n32685 , n32675 , n32684 );
xor ( n32686 , n28638 , n30271 );
xor ( n32687 , n32686 , n30283 );
xor ( n32688 , n28089 , n31453 );
xor ( n32689 , n32688 , n31462 );
not ( n32690 , n32689 );
xor ( n32691 , n32194 , n29793 );
xor ( n32692 , n32691 , n31909 );
and ( n32693 , n32690 , n32692 );
xor ( n32694 , n32687 , n32693 );
xor ( n32695 , n32685 , n32694 );
xor ( n32696 , n32160 , n30139 );
xor ( n32697 , n32696 , n30151 );
xor ( n32698 , n27863 , n29601 );
xor ( n32699 , n32698 , n29199 );
not ( n32700 , n32699 );
xor ( n32701 , n29556 , n29474 );
xor ( n32702 , n32701 , n32611 );
and ( n32703 , n32700 , n32702 );
xor ( n32704 , n32697 , n32703 );
xor ( n32705 , n32695 , n32704 );
xor ( n32706 , n28253 , n29270 );
xor ( n32707 , n32706 , n30066 );
xor ( n32708 , n28431 , n32031 );
xor ( n32709 , n32708 , n29975 );
not ( n32710 , n32709 );
xor ( n32711 , n30611 , n28595 );
xor ( n32712 , n32711 , n28519 );
and ( n32713 , n32710 , n32712 );
xor ( n32714 , n32707 , n32713 );
xor ( n32715 , n32705 , n32714 );
xor ( n32716 , n32664 , n32715 );
not ( n32717 , n32716 );
xor ( n32718 , RI19a94b98_2649 , RI1747b480_1135);
not ( n11744 , n27689 );
and ( n11745 , n11744 , RI1747b480_1135);
and ( n11746 , n32718 , n27689 );
or ( n32719 , n11745 , n11746 );
xor ( n32720 , n32719 , n30487 );
xor ( n32721 , n32720 , n30321 );
xor ( n32722 , n29044 , n28027 );
xor ( n32723 , n32722 , n29827 );
not ( n32724 , n32723 );
and ( n32725 , n32724 , n32436 );
xor ( n32726 , n32721 , n32725 );
xor ( n32727 , RI19ab2670_2436 , RI174a6c20_923);
not ( n11747 , n27689 );
and ( n11748 , n11747 , RI174a6c20_923);
and ( n11749 , n32727 , n27689 );
or ( n32728 , n11748 , n11749 );
buf ( n32729 , RI17338380_2167);
xor ( n32730 , n32728 , n32729 );
xor ( n32731 , n32730 , n32550 );
xor ( n32732 , n32731 , n30464 );
buf ( n32733 , RI1748e5a8_1042);
xor ( n32734 , n32732 , n32733 );
xor ( n32735 , n30880 , n32734 );
xor ( n32736 , RI19ac4dc0_2293 , RI174caad0_780);
not ( n11750 , n27689 );
and ( n11751 , n11750 , RI174caad0_780);
and ( n11752 , n32736 , n27689 );
or ( n32737 , n11751 , n11752 );
xor ( n32738 , n32719 , n32737 );
buf ( n32739 , RI17396160_2024);
xor ( n32740 , n32738 , n32739 );
buf ( n32741 , RI173dee50_1669);
xor ( n32742 , n32740 , n32741 );
buf ( n32743 , RI17456928_1314);
xor ( n32744 , n32742 , n32743 );
xor ( n32745 , n32735 , n32744 );
not ( n32746 , n32745 );
xor ( n32747 , n32085 , n28380 );
xor ( n32748 , n32747 , n28392 );
and ( n32749 , n32746 , n32748 );
xor ( n32750 , n32411 , n32749 );
xor ( n32751 , n28857 , n30207 );
xor ( n32752 , n32751 , n30218 );
not ( n32753 , n32752 );
xor ( n32754 , n30980 , n28659 );
xor ( n32755 , n32754 , n29148 );
and ( n32756 , n32753 , n32755 );
xor ( n32757 , n32431 , n32756 );
xor ( n32758 , n32750 , n32757 );
not ( n32759 , n32721 );
and ( n32760 , n32759 , n32723 );
xor ( n32761 , n32441 , n32760 );
xor ( n32762 , n32758 , n32761 );
xor ( n32763 , n31392 , n29462 );
xor ( n32764 , n32763 , n29474 );
not ( n32765 , n32764 );
xor ( n32766 , n30966 , n28852 );
xor ( n32767 , n32766 , n29873 );
and ( n32768 , n32765 , n32767 );
xor ( n32769 , n32461 , n32768 );
xor ( n32770 , n32762 , n32769 );
xor ( n32771 , RI19a94490_2652 , RI1747aaa8_1138);
not ( n11753 , n27689 );
and ( n11754 , n11753 , RI1747aaa8_1138);
and ( n11755 , n32771 , n27689 );
or ( n32772 , n11754 , n11755 );
xor ( n32773 , n32772 , n32668 );
buf ( n32774 , RI17395788_2027);
xor ( n32775 , n32773 , n32774 );
xor ( n32776 , n32775 , n32237 );
buf ( n32777 , RI17455f50_1317);
xor ( n32778 , n32776 , n32777 );
xor ( n32779 , n30105 , n32778 );
xor ( n32780 , n32779 , n31001 );
not ( n32781 , n32780 );
xor ( n32782 , n30637 , n28174 );
xor ( n32783 , n32782 , n28185 );
and ( n32784 , n32781 , n32783 );
xor ( n32785 , n32478 , n32784 );
xor ( n32786 , n32770 , n32785 );
xor ( n32787 , n32726 , n32786 );
xor ( n32788 , n31914 , n32426 );
xor ( n32789 , n32788 , n31152 );
xor ( n32790 , n29905 , n32091 );
xor ( n32791 , n32790 , n30139 );
not ( n32792 , n32791 );
xor ( n32793 , RI19aa44f8_2535 , RI1747fff8_1112);
not ( n11756 , n27689 );
and ( n11757 , n11756 , RI1747fff8_1112);
and ( n11758 , n32793 , n27689 );
or ( n32794 , n11757 , n11758 );
xor ( n32795 , n32794 , n32181 );
buf ( n32796 , RI1739acd8_2001);
xor ( n32797 , n32795 , n32796 );
buf ( n32798 , RI173e39c8_1646);
xor ( n32799 , n32797 , n32798 );
xor ( n32800 , n32799 , n32524 );
xor ( n32801 , n28966 , n32800 );
xor ( n32802 , RI19ab8430_2393 , RI1749d530_969);
not ( n11759 , n27689 );
and ( n11760 , n11759 , RI1749d530_969);
and ( n11761 , n32802 , n27689 );
or ( n32803 , n11760 , n11761 );
xor ( n32804 , n32803 , n31851 );
buf ( n32805 , RI173b8558_1857);
xor ( n32806 , n32804 , n32805 );
buf ( n32807 , RI17401248_1502);
xor ( n32808 , n32806 , n32807 );
xor ( n32809 , n32808 , n31413 );
xor ( n32810 , n32801 , n32809 );
and ( n32811 , n32792 , n32810 );
xor ( n32812 , n32789 , n32811 );
xor ( n32813 , n31083 , n29519 );
xor ( n32814 , n32813 , n29320 );
xor ( n32815 , n31820 , n29375 );
xor ( n32816 , n32815 , n29767 );
not ( n32817 , n32816 );
xor ( n32818 , n31840 , n30151 );
xor ( n32819 , n32818 , n31024 );
and ( n32820 , n32817 , n32819 );
xor ( n32821 , n32814 , n32820 );
xor ( n32822 , n32812 , n32821 );
xor ( n32823 , n32125 , n28367 );
xor ( n32824 , n32823 , n29952 );
xor ( n32825 , RI19aa4cf0_2531 , RI17481060_1107);
not ( n11762 , n27689 );
and ( n11763 , n11762 , RI17481060_1107);
and ( n11764 , n32825 , n27689 );
or ( n32826 , n11763 , n11764 );
xor ( n32827 , RI19a860c0_2752 , RI17502948_752);
not ( n11765 , n27689 );
and ( n11766 , n11765 , RI17502948_752);
and ( n11767 , n32827 , n27689 );
or ( n32828 , n11766 , n11767 );
xor ( n32829 , n32826 , n32828 );
buf ( n32830 , RI1739bd40_1996);
xor ( n32831 , n32829 , n32830 );
buf ( n32832 , RI173e4d78_1640);
xor ( n32833 , n32831 , n32832 );
buf ( n32834 , RI1745c850_1285);
xor ( n32835 , n32833 , n32834 );
xor ( n32836 , n32361 , n32835 );
xor ( n32837 , n32836 , n31399 );
not ( n32838 , n32837 );
xor ( n32839 , n30161 , n28438 );
xor ( n32840 , n32839 , n28450 );
and ( n32841 , n32838 , n32840 );
xor ( n32842 , n32824 , n32841 );
xor ( n32843 , n32822 , n32842 );
xor ( n32844 , n30542 , n28224 );
xor ( n32845 , n32844 , n28236 );
xor ( n32846 , n28754 , n30823 );
xor ( n32847 , n32846 , n30934 );
not ( n32848 , n32847 );
xor ( n32849 , n28259 , n29270 );
xor ( n32850 , n32849 , n30066 );
and ( n32851 , n32848 , n32850 );
xor ( n32852 , n32845 , n32851 );
xor ( n32853 , n32843 , n32852 );
xor ( n32854 , n29204 , n32459 );
xor ( n32855 , n32854 , n30616 );
xor ( n32856 , n28951 , n27948 );
xor ( n32857 , n32856 , n28702 );
not ( n32858 , n32857 );
xor ( n32859 , n29778 , n28627 );
xor ( n32860 , n32859 , n30089 );
and ( n32861 , n32858 , n32860 );
xor ( n32862 , n32855 , n32861 );
xor ( n32863 , n32853 , n32862 );
xor ( n32864 , n32787 , n32863 );
and ( n32865 , n32717 , n32864 );
xor ( n32866 , n32621 , n32865 );
not ( n11768 , n29614 );
and ( n11769 , n11768 , RI174b47f8_856);
and ( n11770 , n32866 , n29614 );
or ( n32867 , n11769 , n11770 );
not ( n11771 , RI1754c610_2);
and ( n11772 , n11771 , n32867 );
and ( n11773 , C0 , RI1754c610_2);
or ( n32868 , n11772 , n11773 );
buf ( n32869 , n32868 );
not ( n11774 , n27683 );
and ( n11775 , n11774 , RI19abe100_2349);
and ( n11776 , RI19ac6ff8_2277 , n27683 );
or ( n32870 , n11775 , n11776 );
not ( n11777 , RI1754c610_2);
and ( n11778 , n11777 , n32870 );
and ( n11779 , C0 , RI1754c610_2);
or ( n32871 , n11778 , n11779 );
buf ( n32872 , n32871 );
buf ( n32873 , RI1747f2d8_1116);
xor ( n32874 , n28136 , n30243 );
xor ( n32875 , n32874 , n31750 );
not ( n32876 , n32677 );
and ( n32877 , n32876 , n32679 );
xor ( n32878 , n32875 , n32877 );
xor ( n32879 , n29708 , n28947 );
xor ( n32880 , n32879 , n28956 );
xor ( n32881 , n28982 , n28081 );
xor ( n32882 , n32881 , n29248 );
not ( n32883 , n32882 );
and ( n32884 , n32883 , n32666 );
xor ( n32885 , n32880 , n32884 );
xor ( n32886 , n30688 , n30869 );
xor ( n32887 , RI19acd808_2228 , RI17511b28_711);
not ( n11780 , n27689 );
and ( n11781 , n11780 , RI17511b28_711);
and ( n11782 , n32887 , n27689 );
or ( n32888 , n11781 , n11782 );
xor ( n32889 , n31729 , n32888 );
xor ( n32890 , n32889 , n31104 );
buf ( n32891 , RI173ed400_1599);
xor ( n32892 , n32890 , n32891 );
buf ( n32893 , RI17489d78_1064);
xor ( n32894 , n32892 , n32893 );
xor ( n32895 , n32886 , n32894 );
not ( n32896 , n32875 );
and ( n32897 , n32896 , n32677 );
xor ( n32898 , n32895 , n32897 );
xor ( n32899 , n32885 , n32898 );
xor ( n32900 , n27972 , n32366 );
xor ( n32901 , n32900 , n32291 );
xor ( n32902 , n30971 , n28852 );
xor ( n32903 , n32902 , n29873 );
not ( n32904 , n32903 );
and ( n32905 , n32904 , n32687 );
xor ( n32906 , n32901 , n32905 );
xor ( n32907 , n32899 , n32906 );
xor ( n32908 , n29221 , n28995 );
xor ( n32909 , n32908 , n30780 );
xor ( n32910 , n30812 , n32382 );
xor ( n32911 , n32910 , n28463 );
not ( n32912 , n32911 );
and ( n32913 , n32912 , n32697 );
xor ( n32914 , n32909 , n32913 );
xor ( n32915 , n32907 , n32914 );
xor ( n32916 , n28914 , n29889 );
xor ( n32917 , n32916 , n30537 );
xor ( n32918 , n31308 , n31636 );
xor ( n32919 , n32918 , n30655 );
not ( n32920 , n32919 );
and ( n32921 , n32920 , n32707 );
xor ( n32922 , n32917 , n32921 );
xor ( n32923 , n32915 , n32922 );
xor ( n32924 , n32878 , n32923 );
xor ( n32925 , n30262 , n31697 );
xor ( n32926 , n32925 , n31309 );
xor ( n32927 , n30684 , n30869 );
xor ( n32928 , n32927 , n32894 );
not ( n32929 , n32928 );
xor ( n32930 , n30109 , n32778 );
xor ( n32931 , n32930 , n31001 );
and ( n32932 , n32929 , n32931 );
xor ( n32933 , n32926 , n32932 );
xor ( n32934 , n27770 , n31024 );
xor ( n32935 , n32934 , n29306 );
xor ( n32936 , n28677 , n29711 );
xor ( n32937 , n32936 , n30443 );
not ( n32938 , n32937 );
xor ( n32939 , n29315 , n30665 );
xor ( n32940 , n32939 , n31226 );
and ( n32941 , n32938 , n32940 );
xor ( n32942 , n32935 , n32941 );
xor ( n32943 , n32933 , n32942 );
xor ( n32944 , n31300 , n31636 );
xor ( n32945 , n32944 , n30655 );
xor ( n32946 , n27957 , n31131 );
xor ( n32947 , n32946 , n32366 );
not ( n32948 , n32947 );
xor ( n32949 , n30096 , n29910 );
xor ( n32950 , n32949 , n32167 );
and ( n32951 , n32948 , n32950 );
xor ( n32952 , n32945 , n32951 );
xor ( n32953 , n32943 , n32952 );
xor ( n32954 , n30911 , n30348 );
xor ( n32955 , n32954 , n30178 );
xor ( n32956 , n28205 , n29079 );
xor ( n32957 , n32956 , n28583 );
not ( n32958 , n32957 );
xor ( n32959 , n29020 , n28878 );
xor ( n32960 , n32959 , n30399 );
and ( n32961 , n32958 , n32960 );
xor ( n32962 , n32955 , n32961 );
xor ( n32963 , n32953 , n32962 );
xor ( n32964 , n29096 , n28505 );
xor ( n32965 , n32964 , n31038 );
xor ( n32966 , n30806 , n32382 );
xor ( n32967 , n32966 , n28463 );
not ( n32968 , n32967 );
xor ( n32969 , n29719 , n28839 );
xor ( n32970 , n32969 , n28917 );
and ( n32971 , n32968 , n32970 );
xor ( n32972 , n32965 , n32971 );
xor ( n32973 , n32963 , n32972 );
xor ( n32974 , n32924 , n32973 );
xor ( n32975 , RI19a952a0_2646 , RI1747b7c8_1134);
not ( n11783 , n27689 );
and ( n11784 , n11783 , RI1747b7c8_1134);
and ( n11785 , n32975 , n27689 );
or ( n32976 , n11784 , n11785 );
xor ( n32977 , n32976 , n30427 );
xor ( n32978 , n32977 , n29364 );
not ( n32979 , n32824 );
and ( n32980 , n32979 , n32837 );
xor ( n32981 , n32978 , n32980 );
xor ( n32982 , n29258 , n32120 );
xor ( n32983 , n32982 , n29093 );
buf ( n32984 , RI173386c8_2166);
xor ( n32985 , n30404 , n32984 );
buf ( n32986 , RI173c1c48_1811);
xor ( n32987 , n32985 , n32986 );
buf ( n32988 , RI1740a938_1456);
xor ( n32989 , n32987 , n32988 );
buf ( n32990 , RI174a51e0_931);
xor ( n32991 , n32989 , n32990 );
xor ( n32992 , n30478 , n32991 );
xor ( n32993 , n32976 , n31230 );
xor ( n32994 , n32993 , n30573 );
xor ( n32995 , n32994 , n31133 );
xor ( n32996 , n32995 , n32476 );
xor ( n32997 , n32992 , n32996 );
not ( n32998 , n32997 );
and ( n32999 , n32998 , n32789 );
xor ( n33000 , n32983 , n32999 );
xor ( n33001 , n30113 , n32778 );
xor ( n33002 , n33001 , n31001 );
xor ( n33003 , n29564 , n32611 );
xor ( n33004 , n33003 , n29161 );
not ( n33005 , n33004 );
and ( n33006 , n33005 , n32814 );
xor ( n33007 , n33002 , n33006 );
xor ( n33008 , n33000 , n33007 );
xor ( n33009 , n30270 , n31697 );
xor ( n33010 , n33009 , n31309 );
not ( n33011 , n32978 );
and ( n33012 , n33011 , n32824 );
xor ( n33013 , n33010 , n33012 );
xor ( n33014 , n33008 , n33013 );
xor ( n33015 , n28594 , n29187 );
xor ( n33016 , n33015 , n29724 );
xor ( n33017 , n31551 , n28866 );
xor ( n33018 , n33017 , n28878 );
not ( n33019 , n33018 );
and ( n33020 , n33019 , n32845 );
xor ( n33021 , n33016 , n33020 );
xor ( n33022 , n33014 , n33021 );
xor ( n33023 , n31762 , n31714 );
xor ( n33024 , n33023 , n28785 );
xor ( n33025 , n32250 , n30691 );
xor ( n33026 , n33025 , n30475 );
not ( n33027 , n33026 );
and ( n33028 , n33027 , n32855 );
xor ( n33029 , n33024 , n33028 );
xor ( n33030 , n33022 , n33029 );
xor ( n33031 , n32981 , n33030 );
xor ( n33032 , n28387 , n31921 );
xor ( n33033 , n33032 , n30348 );
not ( n33034 , n33033 );
xor ( n33035 , n31419 , n29332 );
xor ( n33036 , n33035 , n29814 );
and ( n33037 , n33034 , n33036 );
xor ( n33038 , n31769 , n33037 );
buf ( n33039 , RI17359008_2091);
xor ( n33040 , n33039 , n28015 );
xor ( n33041 , n33040 , n28027 );
not ( n33042 , n33041 );
xor ( n33043 , n31591 , n30178 );
xor ( n33044 , n33043 , n30189 );
and ( n33045 , n33042 , n33044 );
xor ( n33046 , n31779 , n33045 );
xor ( n33047 , n33038 , n33046 );
xor ( n33048 , n29457 , n31950 );
xor ( n33049 , n33048 , n31558 );
not ( n33050 , n33049 );
xor ( n33051 , n29972 , n30813 );
xor ( n33052 , n33051 , n30823 );
and ( n33053 , n33050 , n33052 );
xor ( n33054 , n31802 , n33053 );
xor ( n33055 , n33047 , n33054 );
xor ( n33056 , n27747 , n29628 );
xor ( n33057 , n33056 , n29639 );
not ( n33058 , n33057 );
xor ( n33059 , n29102 , n28505 );
xor ( n33060 , n33059 , n31038 );
and ( n33061 , n33058 , n33060 );
xor ( n33062 , n31812 , n33061 );
xor ( n33063 , n33055 , n33062 );
not ( n33064 , n31737 );
xor ( n33065 , n28336 , n31076 );
xor ( n33066 , n33065 , n32091 );
and ( n33067 , n33064 , n33066 );
xor ( n33068 , n31733 , n33067 );
xor ( n33069 , n33063 , n33068 );
xor ( n33070 , n33031 , n33069 );
not ( n33071 , n33070 );
xor ( n33072 , n28243 , n29259 );
xor ( n33073 , n33072 , n29270 );
xor ( n33074 , n30384 , n28812 );
xor ( n33075 , n33074 , n29855 );
not ( n33076 , n33075 );
xor ( n33077 , n28566 , n30626 );
xor ( n33078 , n33077 , n29740 );
and ( n33079 , n33076 , n33078 );
xor ( n33080 , n33073 , n33079 );
xor ( n33081 , n28330 , n31076 );
xor ( n33082 , n33081 , n32091 );
xor ( n33083 , n31221 , n28741 );
xor ( n33084 , n33083 , n28096 );
not ( n33085 , n33084 );
xor ( n33086 , n32796 , n31100 );
xor ( n33087 , n33086 , n31422 );
and ( n33088 , n33085 , n33087 );
xor ( n33089 , n33082 , n33088 );
xor ( n33090 , n29818 , n32130 );
xor ( n33091 , n33090 , n32140 );
xor ( n33092 , n30118 , n31001 );
xor ( n33093 , n33092 , n30889 );
not ( n33094 , n33093 );
xor ( n33095 , n30146 , n30918 );
xor ( n33096 , n33095 , n31594 );
and ( n33097 , n33094 , n33096 );
xor ( n33098 , n33091 , n33097 );
xor ( n33099 , n33089 , n33098 );
xor ( n33100 , n32083 , n28380 );
xor ( n33101 , n33100 , n28392 );
xor ( n33102 , n30700 , n28406 );
xor ( n33103 , n33102 , n28418 );
not ( n33104 , n33103 );
xor ( n33105 , n31984 , n28785 );
xor ( n33106 , n33105 , n28015 );
and ( n33107 , n33104 , n33106 );
xor ( n33108 , n33101 , n33107 );
xor ( n33109 , n33099 , n33108 );
xor ( n33110 , n28347 , n30510 );
xor ( n33111 , n33110 , n30522 );
not ( n33112 , n33073 );
and ( n33113 , n33112 , n33075 );
xor ( n33114 , n33111 , n33113 );
xor ( n33115 , n33109 , n33114 );
xor ( n33116 , n28608 , n29995 );
xor ( n33117 , n33116 , n28327 );
xor ( n33118 , n30774 , n29438 );
xor ( n33119 , n33118 , n29449 );
not ( n33120 , n33119 );
xor ( n33121 , n30562 , n31038 );
xor ( n33122 , n33121 , n30271 );
and ( n33123 , n33120 , n33122 );
xor ( n33124 , n33117 , n33123 );
xor ( n33125 , n33115 , n33124 );
xor ( n33126 , n33080 , n33125 );
xor ( n33127 , n29327 , n31226 );
xor ( n33128 , n33127 , n31516 );
xor ( n33129 , n30412 , n30901 );
xor ( n33130 , n33129 , n31475 );
not ( n33131 , n33130 );
xor ( n33132 , n29723 , n28839 );
xor ( n33133 , n33132 , n28917 );
and ( n33134 , n33131 , n33133 );
xor ( n33135 , n33128 , n33134 );
xor ( n33136 , n30173 , n31162 );
xor ( n33137 , n33136 , n29923 );
xor ( n33138 , n31128 , n31528 );
xor ( n33139 , n33138 , n32835 );
not ( n33140 , n33139 );
xor ( n33141 , n28616 , n29995 );
xor ( n33142 , n33141 , n28327 );
and ( n33143 , n33140 , n33142 );
xor ( n33144 , n33137 , n33143 );
xor ( n33145 , n33135 , n33144 );
xor ( n33146 , n30942 , n29586 );
xor ( n33147 , n33146 , n28355 );
xor ( n33148 , n32207 , n28800 );
xor ( n33149 , n33148 , n28812 );
not ( n33150 , n33149 );
xor ( n33151 , n32246 , n27844 );
xor ( n33152 , n33151 , n30691 );
and ( n33153 , n33150 , n33152 );
xor ( n33154 , n33147 , n33153 );
xor ( n33155 , n33145 , n33154 );
xor ( n33156 , n29416 , n27870 );
xor ( n33157 , n33156 , n28174 );
xor ( n33158 , n28301 , n31291 );
xor ( n33159 , n33158 , n27989 );
not ( n33160 , n33159 );
xor ( n33161 , n30305 , n28055 );
xor ( n33162 , n33161 , n28224 );
and ( n33163 , n33160 , n33162 );
xor ( n33164 , n33157 , n33163 );
xor ( n33165 , n33155 , n33164 );
xor ( n33166 , n31692 , n29291 );
xor ( n33167 , n33166 , n31636 );
xor ( n33168 , n29145 , n31089 );
xor ( n33169 , n33168 , n31100 );
not ( n33170 , n33169 );
xor ( n33171 , n31842 , n30151 );
xor ( n33172 , n33171 , n31024 );
and ( n33173 , n33170 , n33172 );
xor ( n33174 , n33167 , n33173 );
xor ( n33175 , n33165 , n33174 );
xor ( n33176 , n33126 , n33175 );
and ( n33177 , n33071 , n33176 );
xor ( n33178 , n32974 , n33177 );
not ( n11786 , n29614 );
and ( n11787 , n11786 , RI174c9b58_783);
and ( n11788 , n33178 , n29614 );
or ( n33179 , n11787 , n11788 );
not ( n11789 , RI1754c610_2);
and ( n11790 , n11789 , n33179 );
and ( n11791 , C0 , RI1754c610_2);
or ( n33180 , n11790 , n11791 );
buf ( n33181 , n33180 );
xor ( n33182 , n27774 , n31024 );
xor ( n33183 , n33182 , n29306 );
not ( n33184 , n33183 );
xor ( n33185 , n29158 , n29037 );
xor ( n33186 , n33185 , n31180 );
and ( n33187 , n33184 , n33186 );
xor ( n33188 , n31262 , n33187 );
not ( n33189 , n31232 );
xor ( n33190 , n30896 , n32744 );
xor ( n33191 , RI19a91c40_2670 , RI175298b8_637);
not ( n11792 , n27689 );
and ( n11793 , n11792 , RI175298b8_637);
and ( n11794 , n33191 , n27689 );
or ( n33192 , n11793 , n11794 );
xor ( n33193 , n30310 , n33192 );
buf ( n33194 , RI173b3698_1881);
xor ( n33195 , n33193 , n33194 );
buf ( n33196 , RI173fc6d0_1525);
xor ( n33197 , n33195 , n33196 );
xor ( n33198 , n33197 , n31569 );
xor ( n33199 , n33190 , n33198 );
and ( n33200 , n33189 , n33199 );
xor ( n33201 , n31227 , n33200 );
not ( n33202 , n31252 );
xor ( n33203 , n31523 , n28107 );
xor ( n33204 , n33203 , n32510 );
and ( n33205 , n33202 , n33204 );
xor ( n33206 , n31249 , n33205 );
xor ( n33207 , n33201 , n33206 );
not ( n33208 , n31262 );
and ( n33209 , n33208 , n33183 );
xor ( n33210 , n31259 , n33209 );
xor ( n33211 , n33207 , n33210 );
not ( n33212 , n31292 );
xor ( n33213 , n29539 , n30594 );
xor ( n33214 , n33213 , n29224 );
and ( n33215 , n33212 , n33214 );
xor ( n33216 , n31280 , n33215 );
xor ( n33217 , n33211 , n33216 );
not ( n33218 , n31314 );
xor ( n33219 , n29672 , n30842 );
xor ( n33220 , n33219 , n32247 );
and ( n33221 , n33218 , n33220 );
xor ( n33222 , n31311 , n33221 );
xor ( n33223 , n33217 , n33222 );
xor ( n33224 , n33188 , n33223 );
xor ( n33225 , n30316 , n32996 );
xor ( n33226 , RI19aa8da0_2504 , RI17498d00_991);
not ( n11795 , n27689 );
and ( n11796 , n11795 , RI17498d00_991);
and ( n11797 , n33226 , n27689 );
or ( n33227 , n11796 , n11797 );
xor ( n33228 , n33227 , n29353 );
buf ( n33229 , RI173b39e0_1880);
xor ( n33230 , n33228 , n33229 );
buf ( n33231 , RI173fca18_1524);
xor ( n33232 , n33230 , n33231 );
buf ( n33233 , RI173ab9e8_1919);
xor ( n33234 , n33232 , n33233 );
xor ( n33235 , n33225 , n33234 );
xor ( n33236 , n30098 , n29910 );
xor ( n33237 , n33236 , n32167 );
not ( n33238 , n33237 );
xor ( n33239 , n28223 , n30457 );
xor ( n33240 , n33239 , n31581 );
and ( n33241 , n33238 , n33240 );
xor ( n33242 , n33235 , n33241 );
xor ( n33243 , n32270 , n27975 );
xor ( n33244 , n33243 , n29346 );
xor ( n33245 , n32041 , n31825 );
xor ( n33246 , n33245 , n29586 );
not ( n33247 , n33246 );
xor ( n33248 , n30282 , n31309 );
xor ( n33249 , n33248 , n29519 );
and ( n33250 , n33247 , n33249 );
xor ( n33251 , n33244 , n33250 );
xor ( n33252 , n33242 , n33251 );
xor ( n33253 , n31483 , n30189 );
xor ( n33254 , n33253 , n28715 );
xor ( n33255 , n29529 , n27819 );
xor ( n33256 , n33255 , n30594 );
not ( n33257 , n33256 );
xor ( n33258 , n28701 , n32472 );
xor ( n33259 , n33258 , n32323 );
and ( n33260 , n33257 , n33259 );
xor ( n33261 , n33254 , n33260 );
xor ( n33262 , n33252 , n33261 );
xor ( n33263 , n28990 , n29248 );
xor ( n33264 , n33263 , n29438 );
xor ( n33265 , n28670 , n28236 );
xor ( n33266 , n33265 , n29711 );
not ( n33267 , n33266 );
xor ( n33268 , n32119 , n28137 );
xor ( n33269 , n33268 , n28493 );
and ( n33270 , n33267 , n33269 );
xor ( n33271 , n33264 , n33270 );
xor ( n33272 , n33262 , n33271 );
xor ( n33273 , n27839 , n30857 );
xor ( n33274 , n33273 , n30869 );
xor ( n33275 , n30886 , n32734 );
xor ( n33276 , n33275 , n32744 );
not ( n33277 , n33276 );
xor ( n33278 , n31130 , n31528 );
xor ( n33279 , n33278 , n32835 );
and ( n33280 , n33277 , n33279 );
xor ( n33281 , n33274 , n33280 );
xor ( n33282 , n33272 , n33281 );
xor ( n33283 , n33224 , n33282 );
xor ( n33284 , n29868 , n30548 );
xor ( n33285 , n33284 , n28673 );
xor ( n33286 , n31062 , n32323 );
xor ( n33287 , n33286 , n32199 );
not ( n33288 , n33287 );
xor ( n33289 , n29290 , n30017 );
xor ( n33290 , n33289 , n30986 );
and ( n33291 , n33288 , n33290 );
xor ( n33292 , n33285 , n33291 );
xor ( n33293 , n28360 , n30522 );
xor ( n33294 , n33293 , n32009 );
xor ( n33295 , n29046 , n28027 );
xor ( n33296 , n33295 , n29827 );
not ( n33297 , n33296 );
xor ( n33298 , n31485 , n30189 );
xor ( n33299 , n33298 , n28715 );
and ( n33300 , n33297 , n33299 );
xor ( n33301 , n33294 , n33300 );
xor ( n33302 , n31156 , n27779 );
xor ( n33303 , n33302 , n27791 );
xor ( n33304 , n30754 , n29161 );
xor ( n33305 , n33304 , n28069 );
not ( n33306 , n33305 );
xor ( n33307 , n31610 , n29839 );
xor ( n33308 , n33307 , n32031 );
and ( n33309 , n33306 , n33308 );
xor ( n33310 , n33303 , n33309 );
xor ( n33311 , n33301 , n33310 );
xor ( n33312 , n29217 , n28995 );
xor ( n33313 , n33312 , n30780 );
xor ( n33314 , n28795 , n31978 );
xor ( n33315 , n33314 , n29409 );
not ( n33316 , n33315 );
xor ( n33317 , n29446 , n30030 );
xor ( n33318 , n33317 , n30972 );
and ( n33319 , n33316 , n33318 );
xor ( n33320 , n33313 , n33319 );
xor ( n33321 , n33311 , n33320 );
xor ( n33322 , n30862 , n30125 );
xor ( n33323 , n33322 , n31114 );
not ( n33324 , n33285 );
and ( n33325 , n33324 , n33287 );
xor ( n33326 , n33323 , n33325 );
xor ( n33327 , n33321 , n33326 );
xor ( n33328 , n31031 , n30053 );
xor ( n33329 , n33328 , n31697 );
xor ( n33330 , n31470 , n33198 );
xor ( n33331 , n33330 , n31714 );
not ( n33332 , n33331 );
xor ( n33333 , n31822 , n29375 );
xor ( n33334 , n33333 , n29767 );
and ( n33335 , n33332 , n33334 );
xor ( n33336 , n33329 , n33335 );
xor ( n33337 , n33327 , n33336 );
xor ( n33338 , n33292 , n33337 );
xor ( n33339 , n29932 , n30706 );
xor ( n33340 , n33339 , n30717 );
xor ( n33341 , n28626 , n28327 );
xor ( n33342 , n33341 , n28339 );
not ( n33343 , n33342 );
xor ( n33344 , n29465 , n31558 );
xor ( n33345 , n33344 , n29025 );
and ( n33346 , n33343 , n33345 );
xor ( n33347 , n33340 , n33346 );
xor ( n33348 , n31871 , n29964 );
xor ( n33349 , n33348 , n32382 );
xor ( n33350 , n27963 , n31131 );
xor ( n33351 , n33350 , n32366 );
not ( n33352 , n33351 );
xor ( n33353 , n29202 , n32459 );
xor ( n33354 , n33353 , n30616 );
and ( n33355 , n33352 , n33354 );
xor ( n33356 , n33349 , n33355 );
xor ( n33357 , n33347 , n33356 );
xor ( n33358 , n28849 , n30306 );
xor ( n33359 , n33358 , n30548 );
xor ( n33360 , n30150 , n30918 );
xor ( n33361 , n33360 , n31594 );
not ( n33362 , n33361 );
xor ( n33363 , n29016 , n28878 );
xor ( n33364 , n33363 , n30399 );
and ( n33365 , n33362 , n33364 );
xor ( n33366 , n33359 , n33365 );
xor ( n33367 , n33357 , n33366 );
xor ( n33368 , n29790 , n30089 );
xor ( n33369 , n33368 , n30101 );
xor ( n33370 , n28658 , n30283 );
xor ( n33371 , n33370 , n31089 );
not ( n33372 , n33371 );
xor ( n33373 , n29071 , n30643 );
xor ( n33374 , n33373 , n29176 );
and ( n33375 , n33372 , n33374 );
xor ( n33376 , n33369 , n33375 );
xor ( n33377 , n33367 , n33376 );
buf ( n33378 , RI173d15c0_1735);
xor ( n33379 , n33378 , n28015 );
xor ( n33380 , n33379 , n28027 );
xor ( n33381 , n27806 , n30758 );
xor ( n33382 , RI19a843b0_2764 , RI17506188_747);
not ( n11798 , n27689 );
and ( n11799 , n11798 , RI17506188_747);
and ( n11800 , n33382 , n27689 );
or ( n33383 , n11799 , n11800 );
xor ( n33384 , n28058 , n33383 );
buf ( n33385 , RI1739cda8_1991);
xor ( n33386 , n33384 , n33385 );
buf ( n33387 , RI173e5de0_1635);
xor ( n33388 , n33386 , n33387 );
buf ( n33389 , RI1745d8b8_1280);
xor ( n33390 , n33388 , n33389 );
xor ( n33391 , n33381 , n33390 );
not ( n33392 , n33391 );
xor ( n33393 , n32826 , n32510 );
xor ( n33394 , n33393 , n29462 );
and ( n33395 , n33392 , n33394 );
xor ( n33396 , n33380 , n33395 );
xor ( n33397 , n33377 , n33396 );
xor ( n33398 , n33338 , n33397 );
not ( n33399 , n33398 );
xor ( n33400 , n32423 , n32167 );
xor ( n33401 , n33400 , n31843 );
xor ( n33402 , n28026 , n30956 );
xor ( n33403 , n33402 , n32130 );
not ( n33404 , n33403 );
xor ( n33405 , n30312 , n32996 );
xor ( n33406 , n33405 , n33234 );
and ( n33407 , n33404 , n33406 );
xor ( n33408 , n33401 , n33407 );
xor ( n33409 , n31019 , n31594 );
xor ( n33410 , n33409 , n31487 );
xor ( n33411 , n31460 , n27964 );
xor ( n33412 , n33411 , n27975 );
not ( n33413 , n33412 );
xor ( n33414 , n30566 , n31038 );
xor ( n33415 , n33414 , n30271 );
and ( n33416 , n33413 , n33415 );
xor ( n33417 , n33410 , n33416 );
xor ( n33418 , n30517 , n29062 );
xor ( n33419 , n33418 , n31613 );
xor ( n33420 , n28403 , n31497 );
xor ( n33421 , n33420 , n31247 );
not ( n33422 , n33421 );
xor ( n33423 , n30900 , n32744 );
xor ( n33424 , n33423 , n33198 );
and ( n33425 , n33422 , n33424 );
xor ( n33426 , n33419 , n33425 );
xor ( n33427 , n33417 , n33426 );
xor ( n33428 , n29568 , n32611 );
xor ( n33429 , n33428 , n29161 );
xor ( n33430 , n30796 , n28771 );
xor ( n33431 , n33430 , n27726 );
not ( n33432 , n33431 );
xor ( n33433 , n29319 , n30665 );
xor ( n33434 , n33433 , n31226 );
and ( n33435 , n33432 , n33434 );
xor ( n33436 , n33429 , n33435 );
xor ( n33437 , n33427 , n33436 );
xor ( n33438 , n28538 , n28125 );
xor ( n33439 , n33438 , n28137 );
xor ( n33440 , n30014 , n28647 );
xor ( n33441 , n33440 , n28659 );
not ( n33442 , n33441 );
xor ( n33443 , n27988 , n28929 );
xor ( n33444 , n33443 , n29677 );
and ( n33445 , n33442 , n33444 );
xor ( n33446 , n33439 , n33445 );
xor ( n33447 , n33437 , n33446 );
xor ( n33448 , n31071 , n32199 );
xor ( n33449 , n33448 , n28380 );
not ( n33450 , n33401 );
and ( n33451 , n33450 , n33403 );
xor ( n33452 , n33449 , n33451 );
xor ( n33453 , n33447 , n33452 );
xor ( n33454 , n33408 , n33453 );
xor ( n33455 , n31696 , n29291 );
xor ( n33456 , n33455 , n31636 );
xor ( n33457 , RI19a8b700_2715 , RI1746d8a8_1202);
not ( n11801 , n27689 );
and ( n11802 , n11801 , RI1746d8a8_1202);
and ( n11803 , n33457 , n27689 );
or ( n33458 , n11802 , n11803 );
xor ( n33459 , n33458 , n28015 );
xor ( n33460 , n33459 , n28027 );
not ( n33461 , n33460 );
xor ( n33462 , n28399 , n31497 );
xor ( n33463 , n33462 , n31247 );
and ( n33464 , n33461 , n33463 );
xor ( n33465 , n33456 , n33464 );
xor ( n33466 , n30320 , n32996 );
xor ( n33467 , n33466 , n33234 );
xor ( n33468 , n28471 , n29224 );
xor ( n33469 , n33468 , n29235 );
not ( n33470 , n33469 );
xor ( n33471 , n28100 , n31462 );
xor ( n33472 , n33471 , n32275 );
and ( n33473 , n33470 , n33472 );
xor ( n33474 , n33467 , n33473 );
xor ( n33475 , n33465 , n33474 );
xor ( n33476 , n28740 , n32809 );
xor ( n33477 , n33476 , n31453 );
xor ( n33478 , n28018 , n30956 );
xor ( n33479 , n33478 , n32130 );
not ( n33480 , n33479 );
xor ( n33481 , n30784 , n28759 );
xor ( n33482 , n33481 , n28771 );
and ( n33483 , n33480 , n33482 );
xor ( n33484 , n33477 , n33483 );
xor ( n33485 , n33475 , n33484 );
xor ( n33486 , n30841 , n27833 );
xor ( n33487 , n33486 , n27844 );
xor ( n33488 , n28975 , n28081 );
xor ( n33489 , n33488 , n29248 );
not ( n33490 , n33489 );
xor ( n33491 , n28695 , n32472 );
xor ( n33492 , n33491 , n32323 );
and ( n33493 , n33490 , n33492 );
xor ( n33494 , n33487 , n33493 );
xor ( n33495 , n33485 , n33494 );
xor ( n33496 , n28366 , n30522 );
xor ( n33497 , n33496 , n32009 );
xor ( n33498 , n29355 , n31763 );
xor ( n33499 , n33498 , n31989 );
not ( n33500 , n33499 );
xor ( n33501 , n27982 , n28929 );
xor ( n33502 , n33501 , n29677 );
and ( n33503 , n33500 , n33502 );
xor ( n33504 , n33497 , n33503 );
xor ( n33505 , n33495 , n33504 );
xor ( n33506 , n33454 , n33505 );
and ( n33507 , n33399 , n33506 );
xor ( n33508 , n33283 , n33507 );
not ( n11804 , n29614 );
and ( n11805 , n11804 , RI173f01f0_1585);
and ( n11806 , n33508 , n29614 );
or ( n33509 , n11805 , n11806 );
not ( n11807 , RI1754c610_2);
and ( n11808 , n11807 , n33509 );
and ( n11809 , C0 , RI1754c610_2);
or ( n33510 , n11808 , n11809 );
buf ( n33511 , n33510 );
xor ( n33512 , n29194 , n28212 );
xor ( n33513 , n33512 , n32459 );
xor ( n33514 , n28926 , n30537 );
xor ( n33515 , n33514 , n30842 );
not ( n33516 , n33515 );
xor ( n33517 , n30456 , n29123 );
xor ( n33518 , n33517 , n29134 );
and ( n33519 , n33516 , n33518 );
xor ( n33520 , n33513 , n33519 );
xor ( n33521 , n31124 , n31528 );
xor ( n33522 , n33521 , n32835 );
xor ( n33523 , n28091 , n31453 );
xor ( n33524 , n33523 , n31462 );
not ( n33525 , n33524 );
xor ( n33526 , n33196 , n30321 );
xor ( n33527 , n33526 , n30332 );
and ( n33528 , n33525 , n33527 );
xor ( n33529 , n33522 , n33528 );
xor ( n33530 , n32984 , n30415 );
xor ( n33531 , n33530 , n30427 );
xor ( n33532 , n27786 , n29306 );
xor ( n33533 , n33532 , n28406 );
not ( n33534 , n33533 );
xor ( n33535 , n32507 , n32275 );
xor ( n33536 , n33535 , n31950 );
and ( n33537 , n33534 , n33536 );
xor ( n33538 , n33531 , n33537 );
xor ( n33539 , n33529 , n33538 );
xor ( n33540 , RI19a82790_2777 , RI1750d2f8_725);
not ( n11810 , n27689 );
and ( n11811 , n11810 , RI1750d2f8_725);
and ( n11812 , n33540 , n27689 );
or ( n33541 , n11811 , n11812 );
xor ( n33542 , n33541 , n31367 );
xor ( n33543 , n33542 , n28800 );
xor ( n33544 , n30506 , n29051 );
xor ( n33545 , n33544 , n29062 );
not ( n33546 , n33545 );
xor ( n33547 , n29406 , n27858 );
xor ( n33548 , n33547 , n27870 );
and ( n33549 , n33546 , n33548 );
xor ( n33550 , n33543 , n33549 );
xor ( n33551 , n33539 , n33550 );
xor ( n33552 , n30037 , n28892 );
xor ( n33553 , n33552 , n28904 );
not ( n33554 , n33513 );
and ( n33555 , n33554 , n33515 );
xor ( n33556 , n33553 , n33555 );
xor ( n33557 , n33551 , n33556 );
xor ( n33558 , n30299 , n28055 );
xor ( n33559 , n33558 , n28224 );
xor ( n33560 , n30982 , n28659 );
xor ( n33561 , n33560 , n29148 );
not ( n33562 , n33561 );
xor ( n33563 , n29317 , n30665 );
xor ( n33564 , n33563 , n31226 );
and ( n33565 , n33562 , n33564 );
xor ( n33566 , n33559 , n33565 );
xor ( n33567 , n33557 , n33566 );
xor ( n33568 , n33520 , n33567 );
xor ( n33569 , n33231 , n29364 );
xor ( n33570 , n33569 , n29375 );
xor ( n33571 , n28312 , n27989 );
xor ( n33572 , n33571 , n28001 );
not ( n33573 , n33572 );
xor ( n33574 , n30142 , n30918 );
xor ( n33575 , n33574 , n31594 );
and ( n33576 , n33573 , n33575 );
xor ( n33577 , n33570 , n33576 );
xor ( n33578 , n29343 , n32291 );
xor ( n33579 , n33578 , n30207 );
xor ( n33580 , n29792 , n30089 );
xor ( n33581 , n33580 , n30101 );
not ( n33582 , n33581 );
xor ( n33583 , n30804 , n32382 );
xor ( n33584 , n33583 , n28463 );
and ( n33585 , n33582 , n33584 );
xor ( n33586 , n33579 , n33585 );
xor ( n33587 , n33577 , n33586 );
xor ( n33588 , n29598 , n28200 );
xor ( n33589 , n33588 , n28212 );
xor ( n33590 , n30888 , n32734 );
xor ( n33591 , n33590 , n32744 );
not ( n33592 , n33591 );
xor ( n33593 , n31586 , n30178 );
xor ( n33594 , n33593 , n30189 );
and ( n33595 , n33592 , n33594 );
xor ( n33596 , n33589 , n33595 );
xor ( n33597 , n33587 , n33596 );
xor ( n33598 , n27830 , n31683 );
xor ( n33599 , n33598 , n30857 );
xor ( n33600 , n32397 , n28673 );
xor ( n33601 , n33600 , n28684 );
not ( n33602 , n33601 );
xor ( n33603 , n30157 , n28438 );
xor ( n33604 , n33603 , n28450 );
and ( n33605 , n33602 , n33604 );
xor ( n33606 , n33599 , n33605 );
xor ( n33607 , n33597 , n33606 );
xor ( n33608 , n28738 , n32809 );
xor ( n33609 , n33608 , n31453 );
xor ( n33610 , n29922 , n27791 );
xor ( n33611 , n33610 , n30706 );
not ( n33612 , n33611 );
xor ( n33613 , n29901 , n32091 );
xor ( n33614 , n33613 , n30139 );
and ( n33615 , n33612 , n33614 );
xor ( n33616 , n33609 , n33615 );
xor ( n33617 , n33607 , n33616 );
xor ( n33618 , n33568 , n33617 );
xor ( n33619 , n30866 , n30125 );
xor ( n33620 , n33619 , n31114 );
not ( n33621 , n31298 );
and ( n33622 , n33621 , n31311 );
xor ( n33623 , n33620 , n33622 );
xor ( n33624 , n32196 , n29793 );
xor ( n33625 , n33624 , n31909 );
not ( n33626 , n33625 );
and ( n33627 , n33626 , n31216 );
xor ( n33628 , n33199 , n33627 );
xor ( n33629 , n31760 , n31714 );
xor ( n33630 , n33629 , n28785 );
not ( n33631 , n33630 );
and ( n33632 , n33631 , n31236 );
xor ( n33633 , n33204 , n33632 );
xor ( n33634 , n33628 , n33633 );
not ( n33635 , n33186 );
and ( n33636 , n33635 , n31257 );
xor ( n33637 , n33183 , n33636 );
xor ( n33638 , n33634 , n33637 );
xor ( n33639 , n29120 , n29873 );
xor ( n33640 , n33639 , n32398 );
not ( n33641 , n33640 );
and ( n33642 , n33641 , n31267 );
xor ( n33643 , n33214 , n33642 );
xor ( n33644 , n33638 , n33643 );
not ( n33645 , n33620 );
and ( n33646 , n33645 , n31298 );
xor ( n33647 , n33220 , n33646 );
xor ( n33648 , n33644 , n33647 );
xor ( n33649 , n33623 , n33648 );
xor ( n33650 , n28732 , n32809 );
xor ( n33651 , n33650 , n31453 );
not ( n33652 , n33651 );
xor ( n33653 , n31757 , n31714 );
xor ( n33654 , n33653 , n28785 );
and ( n33655 , n33652 , n33654 );
xor ( n33656 , n33240 , n33655 );
xor ( n33657 , RI19aa1618_2557 , RI174868f8_1080);
not ( n11813 , n27689 );
and ( n11814 , n11813 , RI174868f8_1080);
and ( n11815 , n33657 , n27689 );
or ( n33658 , n11814 , n11815 );
xor ( n33659 , n33658 , n33541 );
buf ( n33660 , RI173a1920_1968);
xor ( n33661 , n33659 , n33660 );
buf ( n33662 , RI173ea610_1613);
xor ( n33663 , n33661 , n33662 );
buf ( n33664 , RI1746c4f8_1208);
xor ( n33665 , n33663 , n33664 );
xor ( n33666 , n29378 , n33665 );
xor ( n33667 , n33666 , n32209 );
not ( n33668 , n33667 );
xor ( n33669 , n31069 , n32199 );
xor ( n33670 , n33669 , n28380 );
and ( n33671 , n33668 , n33670 );
xor ( n33672 , n33249 , n33671 );
xor ( n33673 , n33656 , n33672 );
xor ( n33674 , n31446 , n29011 );
xor ( n33675 , n33674 , n27964 );
not ( n33676 , n33675 );
xor ( n33677 , n32605 , n29025 );
xor ( n33678 , n33677 , n29037 );
and ( n33679 , n33676 , n33678 );
xor ( n33680 , n33259 , n33679 );
xor ( n33681 , n33673 , n33680 );
xor ( n33682 , n30709 , n28418 );
xor ( n33683 , n33682 , n31969 );
not ( n33684 , n33683 );
xor ( n33685 , n28910 , n29889 );
xor ( n33686 , n33685 , n30537 );
and ( n33687 , n33684 , n33686 );
xor ( n33688 , n33269 , n33687 );
xor ( n33689 , n33681 , n33688 );
xor ( n33690 , n30646 , n31794 );
xor ( n33691 , n33690 , n28969 );
not ( n33692 , n33691 );
xor ( n33693 , n28153 , n27738 );
xor ( n33694 , n33693 , n29259 );
and ( n33695 , n33692 , n33694 );
xor ( n33696 , n33279 , n33695 );
xor ( n33697 , n33689 , n33696 );
xor ( n33698 , n33649 , n33697 );
not ( n33699 , n33698 );
xor ( n33700 , n28157 , n27738 );
xor ( n33701 , n33700 , n29259 );
not ( n33702 , n30607 );
and ( n33703 , n33702 , n30627 );
xor ( n33704 , n33701 , n33703 );
xor ( n33705 , n28233 , n31581 );
xor ( n33706 , n33705 , n28947 );
not ( n33707 , n30644 );
and ( n33708 , n33707 , n30666 );
xor ( n33709 , n33706 , n33708 );
xor ( n33710 , n33704 , n33709 );
xor ( n33711 , n32988 , n30415 );
xor ( n33712 , n33711 , n30427 );
not ( n33713 , n30675 );
and ( n33714 , n33713 , n30677 );
xor ( n33715 , n33712 , n33714 );
xor ( n33716 , n33710 , n33715 );
xor ( n33717 , n32006 , n31613 );
xor ( n33718 , n33717 , n28438 );
not ( n33719 , n30718 );
and ( n33720 , n33719 , n30722 );
xor ( n33721 , n33718 , n33720 );
xor ( n33722 , n33716 , n33721 );
xor ( n33723 , n27906 , n29235 );
xor ( n33724 , n33723 , n30294 );
not ( n33725 , n30731 );
and ( n33726 , n33725 , n30733 );
xor ( n33727 , n33724 , n33726 );
xor ( n33728 , n33722 , n33727 );
xor ( n33729 , n30632 , n33728 );
xor ( n33730 , n28510 , n29724 );
xor ( n33731 , n33730 , n31291 );
xor ( n33732 , n28229 , n31581 );
xor ( n33733 , n33732 , n28947 );
not ( n33734 , n33733 );
xor ( n33735 , n29118 , n29873 );
xor ( n33736 , n33735 , n32398 );
and ( n33737 , n33734 , n33736 );
xor ( n33738 , n33731 , n33737 );
xor ( n33739 , n28960 , n32800 );
xor ( n33740 , n33739 , n32809 );
xor ( n33741 , n30226 , n28160 );
xor ( n33742 , n33741 , n28250 );
not ( n33743 , n33742 );
xor ( n33744 , n27996 , n29677 );
xor ( n33745 , n33744 , n32778 );
and ( n33746 , n33743 , n33745 );
xor ( n33747 , n33740 , n33746 );
xor ( n33748 , n33738 , n33747 );
xor ( n33749 , n31284 , n28917 );
xor ( n33750 , n33749 , n28929 );
xor ( n33751 , n32888 , n31114 );
xor ( n33752 , n33751 , n30415 );
not ( n33753 , n33752 );
xor ( n33754 , n29286 , n30017 );
xor ( n33755 , n33754 , n30986 );
and ( n33756 , n33753 , n33755 );
xor ( n33757 , n33750 , n33756 );
xor ( n33758 , n33748 , n33757 );
xor ( n33759 , n31082 , n29519 );
xor ( n33760 , n33759 , n29320 );
xor ( n33761 , n30752 , n29161 );
xor ( n33762 , n33761 , n28069 );
not ( n33763 , n33762 );
xor ( n33764 , n32039 , n31825 );
xor ( n33765 , n33764 , n29586 );
and ( n33766 , n33763 , n33765 );
xor ( n33767 , n33760 , n33766 );
xor ( n33768 , n33758 , n33767 );
xor ( n33769 , n32451 , n28583 );
xor ( n33770 , n33769 , n28595 );
xor ( n33771 , n29928 , n30706 );
xor ( n33772 , n33771 , n30717 );
not ( n33773 , n33772 );
xor ( n33774 , n27695 , n28480 );
xor ( n33775 , n33774 , n27909 );
and ( n33776 , n33773 , n33775 );
xor ( n33777 , n33770 , n33776 );
xor ( n33778 , n33768 , n33777 );
xor ( n33779 , n33729 , n33778 );
and ( n33780 , n33699 , n33779 );
xor ( n33781 , n33618 , n33780 );
not ( n11816 , n29614 );
and ( n11817 , n11816 , RI173f4048_1566);
and ( n11818 , n33781 , n29614 );
or ( n33782 , n11817 , n11818 );
not ( n11819 , RI1754c610_2);
and ( n11820 , n11819 , n33782 );
and ( n11821 , C0 , RI1754c610_2);
or ( n33783 , n11820 , n11821 );
buf ( n33784 , n33783 );
xor ( n33785 , n32088 , n28380 );
xor ( n33786 , n33785 , n28392 );
xor ( n33787 , n28928 , n30537 );
xor ( n33788 , n33787 , n30842 );
not ( n33789 , n33788 );
and ( n33790 , n33789 , n32337 );
xor ( n33791 , n33786 , n33790 );
not ( n33792 , n32328 );
xor ( n33793 , n28532 , n27764 );
xor ( n33794 , n33793 , n28125 );
and ( n33795 , n33792 , n33794 );
xor ( n33796 , n32325 , n33795 );
not ( n33797 , n33786 );
and ( n33798 , n33797 , n33788 );
xor ( n33799 , n32342 , n33798 );
xor ( n33800 , n33796 , n33799 );
xor ( n33801 , n29059 , n29827 );
xor ( n33802 , n33801 , n29839 );
not ( n33803 , n33802 );
xor ( n33804 , n30042 , n28892 );
xor ( n33805 , n33804 , n28904 );
and ( n33806 , n33803 , n33805 );
xor ( n33807 , n32352 , n33806 );
xor ( n33808 , n33800 , n33807 );
xor ( n33809 , n27735 , n28543 );
xor ( n33810 , n33809 , n32120 );
not ( n33811 , n33810 );
xor ( n33812 , n30642 , n28174 );
xor ( n33813 , n33812 , n28185 );
and ( n33814 , n33811 , n33813 );
xor ( n33815 , n32383 , n33814 );
xor ( n33816 , n33808 , n33815 );
xor ( n33817 , n30440 , n28956 );
xor ( n33818 , n33817 , n29995 );
not ( n33819 , n33818 );
xor ( n33820 , n32743 , n30487 );
xor ( n33821 , n33820 , n30321 );
and ( n33822 , n33819 , n33821 );
xor ( n33823 , n32400 , n33822 );
xor ( n33824 , n33816 , n33823 );
xor ( n33825 , n33791 , n33824 );
xor ( n33826 , n33825 , n32786 );
xor ( n33827 , n30486 , n32991 );
xor ( n33828 , n33827 , n32996 );
xor ( n33829 , n29914 , n27791 );
xor ( n33830 , n33829 , n30706 );
not ( n33831 , n33830 );
xor ( n33832 , n29648 , n30389 );
xor ( n33833 , n33832 , n28200 );
and ( n33834 , n33831 , n33833 );
xor ( n33835 , n33828 , n33834 );
xor ( n33836 , n31986 , n28785 );
xor ( n33837 , n33836 , n28015 );
xor ( n33838 , n29676 , n30842 );
xor ( n33839 , n33838 , n32247 );
not ( n33840 , n33839 );
xor ( n33841 , n30169 , n31162 );
xor ( n33842 , n33841 , n29923 );
and ( n33843 , n33840 , n33842 );
xor ( n33844 , n33837 , n33843 );
xor ( n33845 , n29558 , n29474 );
xor ( n33846 , n33845 , n32611 );
xor ( n33847 , n29909 , n32091 );
xor ( n33848 , n33847 , n30139 );
not ( n33849 , n33848 );
xor ( n33850 , n29493 , n30789 );
xor ( n33851 , n33850 , n30799 );
and ( n33852 , n33849 , n33851 );
xor ( n33853 , n33846 , n33852 );
xor ( n33854 , n33844 , n33853 );
xor ( n33855 , n29076 , n30643 );
xor ( n33856 , n33855 , n29176 );
not ( n33857 , n33828 );
and ( n33858 , n33857 , n33830 );
xor ( n33859 , n33856 , n33858 );
xor ( n33860 , n33854 , n33859 );
xor ( n33861 , n30111 , n32778 );
xor ( n33862 , n33861 , n31001 );
xor ( n33863 , n29710 , n28947 );
xor ( n33864 , n33863 , n28956 );
not ( n33865 , n33864 );
xor ( n33866 , n29967 , n30813 );
xor ( n33867 , n33866 , n30823 );
and ( n33868 , n33865 , n33867 );
xor ( n33869 , n33862 , n33868 );
xor ( n33870 , n33860 , n33869 );
xor ( n33871 , n29008 , n29814 );
xor ( n33872 , n33871 , n31131 );
xor ( n33873 , n28405 , n31497 );
xor ( n33874 , n33873 , n31247 );
not ( n33875 , n33874 );
xor ( n33876 , n28383 , n31921 );
xor ( n33877 , n33876 , n30348 );
and ( n33878 , n33875 , n33877 );
xor ( n33879 , n33872 , n33878 );
xor ( n33880 , n33870 , n33879 );
xor ( n33881 , n33835 , n33880 );
xor ( n33882 , n27782 , n29306 );
xor ( n33883 , n33882 , n28406 );
xor ( n33884 , n29554 , n29474 );
xor ( n33885 , n33884 , n32611 );
not ( n33886 , n33885 );
xor ( n33887 , n31946 , n29346 );
xor ( n33888 , n33887 , n28866 );
and ( n33889 , n33886 , n33888 );
xor ( n33890 , n33883 , n33889 );
xor ( n33891 , n28762 , n30934 );
xor ( n33892 , n33891 , n28533 );
xor ( n33893 , n29368 , n31989 );
xor ( n33894 , n33458 , n28005 );
xor ( n33895 , n33894 , n33039 );
xor ( n33896 , n33895 , n33378 );
buf ( n33897 , RI17449098_1380);
xor ( n33898 , n33896 , n33897 );
xor ( n33899 , n33893 , n33898 );
not ( n33900 , n33899 );
xor ( n33901 , n31965 , n27885 );
xor ( n33902 , n33901 , n27897 );
and ( n33903 , n33900 , n33902 );
xor ( n33904 , n33892 , n33903 );
xor ( n33905 , n33890 , n33904 );
xor ( n33906 , n28397 , n31497 );
xor ( n33907 , n33906 , n31247 );
xor ( n33908 , n29848 , n29421 );
xor ( n33909 , n33908 , n30643 );
not ( n33910 , n33909 );
xor ( n33911 , n28433 , n32031 );
xor ( n33912 , n33911 , n29975 );
and ( n33913 , n33910 , n33912 );
xor ( n33914 , n33907 , n33913 );
xor ( n33915 , n33905 , n33914 );
xor ( n33916 , n28455 , n29502 );
xor ( n33917 , n33916 , n29628 );
xor ( n33918 , n31629 , n30986 );
xor ( n33919 , n33918 , n31794 );
not ( n33920 , n33919 );
xor ( n33921 , n30623 , n28519 );
xor ( n33922 , n33921 , n28304 );
and ( n33923 , n33920 , n33922 );
xor ( n33924 , n33917 , n33923 );
xor ( n33925 , n33915 , n33924 );
xor ( n33926 , n31143 , n31843 );
xor ( n33927 , n33926 , n27779 );
xor ( n33928 , n29705 , n28947 );
xor ( n33929 , n33928 , n28956 );
not ( n33930 , n33929 );
xor ( n33931 , n32805 , n31422 );
xor ( n33932 , n33931 , n29011 );
and ( n33933 , n33930 , n33932 );
xor ( n33934 , n33927 , n33933 );
xor ( n33935 , n33925 , n33934 );
xor ( n33936 , n33881 , n33935 );
not ( n33937 , n33936 );
xor ( n33938 , n30792 , n28771 );
xor ( n33939 , n33938 , n27726 );
xor ( n33940 , n29141 , n31089 );
xor ( n33941 , n33940 , n31100 );
not ( n33942 , n33941 );
xor ( n33943 , n31288 , n28917 );
xor ( n33944 , n33943 , n28929 );
and ( n33945 , n33942 , n33944 );
xor ( n33946 , n33939 , n33945 );
xor ( n33947 , n30124 , n31001 );
xor ( n33948 , n33947 , n30889 );
xor ( n33949 , n31490 , n28715 );
xor ( n33950 , n33949 , n28727 );
not ( n33951 , n33950 );
xor ( n33952 , n29018 , n28878 );
xor ( n33953 , n33952 , n30399 );
and ( n33954 , n33951 , n33953 );
xor ( n33955 , n33948 , n33954 );
xor ( n33956 , n31151 , n31843 );
xor ( n33957 , n33956 , n27779 );
xor ( n33958 , n27755 , n29639 );
xor ( n33959 , n33958 , n30233 );
not ( n33960 , n33959 );
xor ( n33961 , n28008 , n30946 );
xor ( n33962 , n33961 , n30956 );
and ( n33963 , n33960 , n33962 );
xor ( n33964 , n33957 , n33963 );
xor ( n33965 , n33955 , n33964 );
xor ( n33966 , n31713 , n30332 );
xor ( n33967 , n33966 , n32043 );
xor ( n33968 , n28718 , n31279 );
xor ( n33969 , n33968 , n33665 );
not ( n33970 , n33969 );
xor ( n33971 , n28167 , n29199 );
xor ( n33972 , n33971 , n29211 );
and ( n33973 , n33970 , n33972 );
xor ( n33974 , n33967 , n33973 );
xor ( n33975 , n33965 , n33974 );
xor ( n33976 , n28290 , n28617 );
xor ( n33977 , n33976 , n28627 );
not ( n33978 , n33939 );
and ( n33979 , n33978 , n33941 );
xor ( n33980 , n33977 , n33979 );
xor ( n33981 , n33975 , n33980 );
xor ( n33982 , n31366 , n31969 );
xor ( n33983 , n33982 , n31978 );
xor ( n33984 , n31015 , n31594 );
xor ( n33985 , n33984 , n31487 );
not ( n33986 , n33985 );
xor ( n33987 , n27941 , n30374 );
xor ( n33988 , n33987 , n32472 );
and ( n33989 , n33986 , n33988 );
xor ( n33990 , n33983 , n33989 );
xor ( n33991 , n33981 , n33990 );
xor ( n33992 , n33946 , n33991 );
xor ( n33993 , n27800 , n30758 );
xor ( n33994 , n33993 , n33390 );
xor ( n33995 , n32607 , n29025 );
xor ( n33996 , n33995 , n29037 );
not ( n33997 , n33996 );
xor ( n33998 , n29824 , n32130 );
xor ( n33999 , n33998 , n32140 );
and ( n34000 , n33997 , n33999 );
xor ( n34001 , n33994 , n34000 );
xor ( n34002 , n28348 , n30510 );
xor ( n34003 , n34002 , n30522 );
xor ( n34004 , n28807 , n29409 );
xor ( n34005 , n34004 , n29421 );
not ( n34006 , n34005 );
xor ( n34007 , n28066 , n31180 );
xor ( n34008 , n34007 , n31192 );
and ( n34009 , n34006 , n34008 );
xor ( n34010 , n34003 , n34009 );
xor ( n34011 , n34001 , n34010 );
xor ( n34012 , n32453 , n28583 );
xor ( n34013 , n34012 , n28595 );
xor ( n34014 , n29497 , n30789 );
xor ( n34015 , n34014 , n30799 );
not ( n34016 , n34015 );
xor ( n34017 , n29721 , n28839 );
xor ( n34018 , n34017 , n28917 );
and ( n34019 , n34016 , n34018 );
xor ( n34020 , n34013 , n34019 );
xor ( n34021 , n34011 , n34020 );
xor ( n34022 , n29313 , n30665 );
xor ( n34023 , n34022 , n31226 );
xor ( n34024 , n30532 , n29752 );
xor ( n34025 , n34024 , n27833 );
not ( n34026 , n34025 );
xor ( n34027 , n30898 , n32744 );
xor ( n34028 , n34027 , n33198 );
and ( n34029 , n34026 , n34028 );
xor ( n34030 , n34023 , n34029 );
xor ( n34031 , n34021 , n34030 );
xor ( n34032 , n28284 , n28617 );
xor ( n34033 , n34032 , n28627 );
xor ( n34034 , n28102 , n31462 );
xor ( n34035 , n34034 , n32275 );
not ( n34036 , n34035 );
xor ( n34037 , n32289 , n31399 );
xor ( n34038 , n34037 , n29561 );
and ( n34039 , n34036 , n34038 );
xor ( n34040 , n34033 , n34039 );
xor ( n34041 , n34031 , n34040 );
xor ( n34042 , n33992 , n34041 );
and ( n34043 , n33937 , n34042 );
xor ( n34044 , n33826 , n34043 );
not ( n11822 , n29614 );
and ( n11823 , n11822 , RI174586b0_1305);
and ( n11824 , n34044 , n29614 );
or ( n34045 , n11823 , n11824 );
not ( n11825 , RI1754c610_2);
and ( n11826 , n11825 , n34045 );
and ( n11827 , C0 , RI1754c610_2);
or ( n34046 , n11826 , n11827 );
buf ( n34047 , n34046 );
xor ( n34048 , n31274 , n30717 );
xor ( n34049 , n34048 , n31367 );
not ( n34050 , n33846 );
and ( n34051 , n34050 , n33848 );
xor ( n34052 , n34049 , n34051 );
xor ( n34053 , n29339 , n32291 );
xor ( n34054 , n34053 , n30207 );
xor ( n34055 , n32830 , n32510 );
xor ( n34056 , n34055 , n29462 );
not ( n34057 , n34056 );
and ( n34058 , n34057 , n33837 );
xor ( n34059 , n34054 , n34058 );
xor ( n34060 , n30325 , n33234 );
xor ( n34061 , n34060 , n31825 );
not ( n34062 , n34049 );
and ( n34063 , n34062 , n33846 );
xor ( n34064 , n34061 , n34063 );
xor ( n34065 , n34059 , n34064 );
xor ( n34066 , n29947 , n32009 );
xor ( n34067 , n34066 , n30164 );
not ( n34068 , n34067 );
and ( n34069 , n34068 , n33856 );
xor ( n34070 , n33833 , n34069 );
xor ( n34071 , n34065 , n34070 );
xor ( n34072 , n30264 , n31697 );
xor ( n34073 , n34072 , n31309 );
xor ( n34074 , n28822 , n28557 );
xor ( n34075 , n34074 , n28569 );
not ( n34076 , n34075 );
and ( n34077 , n34076 , n33862 );
xor ( n34078 , n34073 , n34077 );
xor ( n34079 , n34071 , n34078 );
xor ( n34080 , n32393 , n28673 );
xor ( n34081 , n34080 , n28684 );
xor ( n34082 , n30661 , n28969 );
xor ( n34083 , n34082 , n28741 );
not ( n34084 , n34083 );
and ( n34085 , n34084 , n33872 );
xor ( n34086 , n34081 , n34085 );
xor ( n34087 , n34079 , n34086 );
xor ( n34088 , n34052 , n34087 );
xor ( n34089 , n30944 , n29586 );
xor ( n34090 , n34089 , n28355 );
xor ( n34091 , n27843 , n30857 );
xor ( n34092 , n34091 , n30869 );
not ( n34093 , n34092 );
and ( n34094 , n34093 , n33883 );
xor ( n34095 , n34090 , n34094 );
xor ( n34096 , n29022 , n28878 );
xor ( n34097 , n34096 , n30399 );
xor ( n34098 , n28391 , n31921 );
xor ( n34099 , n34098 , n30348 );
not ( n34100 , n34099 );
and ( n34101 , n34100 , n33892 );
xor ( n34102 , n34097 , n34101 );
xor ( n34103 , n34095 , n34102 );
xor ( n34104 , n28182 , n29211 );
xor ( n34105 , n34104 , n28557 );
xor ( n34106 , n30426 , n31475 );
xor ( n34107 , n34106 , n31763 );
not ( n34108 , n34107 );
and ( n34109 , n34108 , n33907 );
xor ( n34110 , n34105 , n34109 );
xor ( n34111 , n34103 , n34110 );
xor ( n34112 , n32254 , n30691 );
xor ( n34113 , n34112 , n30475 );
xor ( n34114 , n27947 , n30374 );
xor ( n34115 , n34114 , n32472 );
not ( n34116 , n34115 );
and ( n34117 , n34116 , n33917 );
xor ( n34118 , n34113 , n34117 );
xor ( n34119 , n34111 , n34118 );
xor ( n34120 , n31525 , n28107 );
xor ( n34121 , n34120 , n32510 );
xor ( n34122 , n28726 , n31279 );
xor ( n34123 , n34122 , n33665 );
not ( n34124 , n34123 );
and ( n34125 , n34124 , n33927 );
xor ( n34126 , n34121 , n34125 );
xor ( n34127 , n34119 , n34126 );
xor ( n34128 , n34088 , n34127 );
not ( n34129 , n31795 );
and ( n34130 , n34129 , n31797 );
xor ( n34131 , n33052 , n34130 );
not ( n34132 , n33036 );
and ( n34133 , n34132 , n31752 );
xor ( n34134 , n33033 , n34133 );
not ( n34135 , n33044 );
and ( n34136 , n34135 , n31774 );
xor ( n34137 , n33041 , n34136 );
xor ( n34138 , n34134 , n34137 );
not ( n34139 , n33052 );
and ( n34140 , n34139 , n31795 );
xor ( n34141 , n33049 , n34140 );
xor ( n34142 , n34138 , n34141 );
not ( n34143 , n33060 );
and ( n34144 , n34143 , n31807 );
xor ( n34145 , n33057 , n34144 );
xor ( n34146 , n34142 , n34145 );
not ( n34147 , n33066 );
and ( n34148 , n34147 , n31827 );
xor ( n34149 , n31737 , n34148 );
xor ( n34150 , n34146 , n34149 );
xor ( n34151 , n34131 , n34150 );
xor ( n34152 , n28891 , n30066 );
xor ( n34153 , n34152 , n30007 );
xor ( n34154 , n31705 , n30332 );
xor ( n34155 , n34154 , n32043 );
not ( n34156 , n34155 );
and ( n34157 , n34156 , n31834 );
xor ( n34158 , n34153 , n34157 );
xor ( n34159 , n32893 , n31114 );
xor ( n34160 , n34159 , n30415 );
xor ( n34161 , n27810 , n33390 );
xor ( n34162 , n34161 , n28983 );
not ( n34163 , n34162 );
and ( n34164 , n34163 , n31853 );
xor ( n34165 , n34160 , n34164 );
xor ( n34166 , n34158 , n34165 );
xor ( n34167 , n29147 , n31089 );
xor ( n34168 , n34167 , n31100 );
xor ( n34169 , n32035 , n31825 );
xor ( n34170 , n34169 , n29586 );
not ( n34171 , n34170 );
and ( n34172 , n34171 , n31876 );
xor ( n34173 , n34168 , n34172 );
xor ( n34174 , n34166 , n34173 );
xor ( n34175 , n29739 , n28304 );
xor ( n34176 , n34175 , n28313 );
xor ( n34177 , n29153 , n29037 );
xor ( n34178 , n34177 , n31180 );
not ( n34179 , n34178 );
and ( n34180 , n34179 , n31886 );
xor ( n34181 , n34176 , n34180 );
xor ( n34182 , n34174 , n34181 );
xor ( n34183 , n29766 , n33898 );
xor ( n34184 , n34183 , n29051 );
xor ( n34185 , n30892 , n32744 );
xor ( n34186 , n34185 , n33198 );
not ( n34187 , n34186 );
and ( n34188 , n34187 , n31896 );
xor ( n34189 , n34184 , n34188 );
xor ( n34190 , n34182 , n34189 );
xor ( n34191 , n34151 , n34190 );
not ( n34192 , n34191 );
xor ( n34193 , n30508 , n29051 );
xor ( n34194 , n34193 , n29062 );
not ( n34195 , n33948 );
and ( n34196 , n34195 , n33950 );
xor ( n34197 , n34194 , n34196 );
xor ( n34198 , n27804 , n30758 );
xor ( n34199 , n34198 , n33390 );
not ( n34200 , n33957 );
and ( n34201 , n34200 , n33959 );
xor ( n34202 , n34199 , n34201 );
xor ( n34203 , n34197 , n34202 );
xor ( n34204 , n30613 , n28595 );
xor ( n34205 , n34204 , n28519 );
not ( n34206 , n33967 );
and ( n34207 , n34206 , n33969 );
xor ( n34208 , n34205 , n34207 );
xor ( n34209 , n34203 , n34208 );
xor ( n34210 , n32891 , n31114 );
xor ( n34211 , n34210 , n30415 );
not ( n34212 , n33977 );
and ( n34213 , n34212 , n33939 );
xor ( n34214 , n34211 , n34213 );
xor ( n34215 , n34209 , n34214 );
xor ( n34216 , n32272 , n27975 );
xor ( n34217 , n34216 , n29346 );
not ( n34218 , n33983 );
and ( n34219 , n34218 , n33985 );
xor ( n34220 , n34217 , n34219 );
xor ( n34221 , n34215 , n34220 );
xor ( n34222 , n33980 , n34221 );
xor ( n34223 , n31270 , n30717 );
xor ( n34224 , n34223 , n31367 );
not ( n34225 , n33994 );
and ( n34226 , n34225 , n33996 );
xor ( n34227 , n34224 , n34226 );
xor ( n34228 , n28151 , n27738 );
xor ( n34229 , n34228 , n29259 );
not ( n34230 , n34003 );
and ( n34231 , n34230 , n34005 );
xor ( n34232 , n34229 , n34231 );
xor ( n34233 , n34227 , n34232 );
xor ( n34234 , n31358 , n31969 );
xor ( n34235 , n34234 , n31978 );
not ( n34236 , n34013 );
and ( n34237 , n34236 , n34015 );
xor ( n34238 , n34235 , n34237 );
xor ( n34239 , n34233 , n34238 );
xor ( n34240 , n28525 , n27764 );
xor ( n34241 , n34240 , n28125 );
not ( n34242 , n34023 );
and ( n34243 , n34242 , n34025 );
xor ( n34244 , n34241 , n34243 );
xor ( n34245 , n34239 , n34244 );
xor ( n34246 , n30181 , n29923 );
xor ( n34247 , n34246 , n29935 );
not ( n34248 , n34033 );
and ( n34249 , n34248 , n34035 );
xor ( n34250 , n34247 , n34249 );
xor ( n34251 , n34245 , n34250 );
xor ( n34252 , n34222 , n34251 );
and ( n34253 , n34192 , n34252 );
xor ( n34254 , n34128 , n34253 );
not ( n11828 , n29614 );
and ( n11829 , n11828 , RI17390c10_2050);
and ( n11830 , n34254 , n29614 );
or ( n34255 , n11829 , n11830 );
not ( n11831 , RI1754c610_2);
and ( n11832 , n11831 , n34255 );
and ( n11833 , C0 , RI1754c610_2);
or ( n34256 , n11832 , n11833 );
buf ( n34257 , n34256 );
not ( n11834 , n27683 );
and ( n11835 , n11834 , RI19acf680_2215);
and ( n11836 , RI19aa29c8_2548 , n27683 );
or ( n34258 , n11835 , n11836 );
not ( n11837 , RI1754c610_2);
and ( n11838 , n11837 , n34258 );
and ( n11839 , C0 , RI1754c610_2);
or ( n34259 , n11838 , n11839 );
buf ( n34260 , n34259 );
xor ( n34261 , n28130 , n30243 );
xor ( n34262 , n34261 , n31750 );
not ( n34263 , n34262 );
and ( n34264 , n34263 , n31438 );
xor ( n34265 , n31404 , n34264 );
xor ( n34266 , n29955 , n30164 );
xor ( n34267 , n34266 , n29490 );
not ( n34268 , n34267 );
xor ( n34269 , n30382 , n28812 );
xor ( n34270 , n34269 , n29855 );
and ( n34271 , n34268 , n34270 );
xor ( n34272 , n31424 , n34271 );
xor ( n34273 , n30449 , n29123 );
xor ( n34274 , n34273 , n29134 );
not ( n34275 , n34274 );
xor ( n34276 , n30211 , n29573 );
xor ( n34277 , n34276 , n30758 );
and ( n34278 , n34275 , n34277 );
xor ( n34279 , n31433 , n34278 );
xor ( n34280 , n34272 , n34279 );
not ( n34281 , n31404 );
and ( n34282 , n34281 , n34262 );
xor ( n34283 , n31401 , n34282 );
xor ( n34284 , n34280 , n34283 );
xor ( n34285 , n28844 , n30306 );
xor ( n34286 , n34285 , n30548 );
not ( n34287 , n34286 );
xor ( n34288 , n32419 , n32167 );
xor ( n34289 , n34288 , n31843 );
and ( n34290 , n34287 , n34289 );
xor ( n34291 , n31476 , n34290 );
xor ( n34292 , n34284 , n34291 );
xor ( n34293 , n32123 , n28367 );
xor ( n34294 , n34293 , n29952 );
not ( n34295 , n34294 );
xor ( n34296 , n30468 , n32894 );
xor ( n34297 , n34296 , n32991 );
and ( n34298 , n34295 , n34297 );
xor ( n34299 , n31503 , n34298 );
xor ( n34300 , n34292 , n34299 );
xor ( n34301 , n34265 , n34300 );
xor ( n34302 , n29650 , n30389 );
xor ( n34303 , n34302 , n28200 );
not ( n34304 , n34303 );
xor ( n34305 , n27816 , n33390 );
xor ( n34306 , n34305 , n28983 );
and ( n34307 , n34304 , n34306 );
xor ( n34308 , n31534 , n34307 );
xor ( n34309 , n27721 , n28533 );
xor ( n34310 , n34309 , n28543 );
not ( n34311 , n34310 );
xor ( n34312 , n29196 , n28212 );
xor ( n34313 , n34312 , n32459 );
and ( n34314 , n34311 , n34313 );
xor ( n34315 , n31546 , n34314 );
xor ( n34316 , n34308 , n34315 );
xor ( n34317 , n30026 , n27921 );
xor ( n34318 , n34317 , n28852 );
not ( n34319 , n34318 );
xor ( n34320 , n30564 , n31038 );
xor ( n34321 , n34320 , n30271 );
and ( n34322 , n34319 , n34321 );
xor ( n34323 , n31565 , n34322 );
xor ( n34324 , n34316 , n34323 );
xor ( n34325 , n31304 , n31636 );
xor ( n34326 , n34325 , n30655 );
not ( n34327 , n34326 );
xor ( n34328 , n27961 , n31131 );
xor ( n34329 , n34328 , n32366 );
and ( n34330 , n34327 , n34329 );
xor ( n34331 , n31595 , n34330 );
xor ( n34332 , n34324 , n34331 );
xor ( n34333 , n28710 , n29935 );
xor ( n34334 , n34333 , n31279 );
not ( n34335 , n34334 );
xor ( n34336 , n31967 , n27885 );
xor ( n34337 , n34336 , n27897 );
and ( n34338 , n34335 , n34337 );
xor ( n34339 , n31618 , n34338 );
xor ( n34340 , n34332 , n34339 );
xor ( n34341 , n34301 , n34340 );
xor ( n34342 , n28734 , n32809 );
xor ( n34343 , n34342 , n31453 );
xor ( n34344 , n31678 , n28001 );
xor ( n34345 , n34344 , n30114 );
not ( n34346 , n34345 );
xor ( n34347 , n30318 , n32996 );
xor ( n34348 , n34347 , n33234 );
and ( n34349 , n34346 , n34348 );
xor ( n34350 , n34343 , n34349 );
xor ( n34351 , n31961 , n27885 );
xor ( n34352 , n34351 , n27897 );
xor ( n34353 , n28062 , n31180 );
xor ( n34354 , n34353 , n31192 );
not ( n34355 , n34354 );
xor ( n34356 , n30395 , n27807 );
xor ( n34357 , n34356 , n27819 );
and ( n34358 , n34355 , n34357 );
xor ( n34359 , n34352 , n34358 );
xor ( n34360 , n32112 , n28137 );
xor ( n34361 , n34360 , n28493 );
xor ( n34362 , n29055 , n29827 );
xor ( n34363 , n34362 , n29839 );
not ( n34364 , n34363 );
xor ( n34365 , n27865 , n29601 );
xor ( n34366 , n34365 , n29199 );
and ( n34367 , n34364 , n34366 );
xor ( n34368 , n34361 , n34367 );
xor ( n34369 , n34359 , n34368 );
xor ( n34370 , n27888 , n29399 );
xor ( n34371 , n34370 , n29655 );
xor ( n34372 , n29181 , n28827 );
xor ( n34373 , n34372 , n28839 );
not ( n34374 , n34373 );
xor ( n34375 , n28766 , n30934 );
xor ( n34376 , n34375 , n28533 );
and ( n34377 , n34374 , n34376 );
xor ( n34378 , n34371 , n34377 );
xor ( n34379 , n34369 , n34378 );
xor ( n34380 , n30225 , n28160 );
xor ( n34381 , n34380 , n28250 );
not ( n34382 , n34343 );
and ( n34383 , n34382 , n34345 );
xor ( n34384 , n34381 , n34383 );
xor ( n34385 , n34379 , n34384 );
xor ( n34386 , n30698 , n28406 );
xor ( n34387 , n34386 , n28418 );
xor ( n34388 , n28320 , n31065 );
xor ( n34389 , n34388 , n31076 );
not ( n34390 , n34389 );
xor ( n34391 , n27970 , n32366 );
xor ( n34392 , n34391 , n32291 );
and ( n34393 , n34390 , n34392 );
xor ( n34394 , n34387 , n34393 );
xor ( n34395 , n34385 , n34394 );
xor ( n34396 , n34350 , n34395 );
xor ( n34397 , n33385 , n28069 );
xor ( n34398 , n34397 , n28081 );
xor ( n34399 , n28435 , n32031 );
xor ( n34400 , n34399 , n29975 );
not ( n34401 , n34400 );
xor ( n34402 , n31474 , n33198 );
xor ( n34403 , n34402 , n31714 );
and ( n34404 , n34401 , n34403 );
xor ( n34405 , n34398 , n34404 );
xor ( n34406 , n28207 , n29079 );
xor ( n34407 , n34406 , n28583 );
xor ( n34408 , n28992 , n29248 );
xor ( n34409 , n34408 , n29438 );
not ( n34410 , n34409 );
xor ( n34411 , n30705 , n28406 );
xor ( n34412 , n34411 , n28418 );
and ( n34413 , n34410 , n34412 );
xor ( n34414 , n34407 , n34413 );
xor ( n34415 , n34405 , n34414 );
xor ( n34416 , n27759 , n29639 );
xor ( n34417 , n34416 , n30233 );
xor ( n34418 , n28310 , n27989 );
xor ( n34419 , n34418 , n28001 );
not ( n34420 , n34419 );
xor ( n34421 , n30955 , n28355 );
xor ( n34422 , n34421 , n28367 );
and ( n34423 , n34420 , n34422 );
xor ( n34424 , n34417 , n34423 );
xor ( n34425 , n34415 , n34424 );
xor ( n34426 , n32774 , n32247 );
xor ( n34427 , n34426 , n32256 );
xor ( n34428 , n29361 , n31763 );
xor ( n34429 , n34428 , n31989 );
not ( n34430 , n34429 );
xor ( n34431 , n30100 , n29910 );
xor ( n34432 , n34431 , n32167 );
and ( n34433 , n34430 , n34432 );
xor ( n34434 , n34427 , n34433 );
xor ( n34435 , n34425 , n34434 );
xor ( n34436 , n31395 , n29462 );
xor ( n34437 , n34436 , n29474 );
xor ( n34438 , n28875 , n30218 );
xor ( n34439 , n34438 , n27807 );
not ( n34440 , n34439 );
xor ( n34441 , n29420 , n27870 );
xor ( n34442 , n34441 , n28174 );
and ( n34443 , n34440 , n34442 );
xor ( n34444 , n34437 , n34443 );
xor ( n34445 , n34435 , n34444 );
xor ( n34446 , n34396 , n34445 );
not ( n34447 , n34446 );
not ( n34448 , n31922 );
and ( n34449 , n34448 , n34184 );
xor ( n34450 , n31898 , n34449 );
xor ( n34451 , n34450 , n31925 );
not ( n34452 , n33415 );
xor ( n34453 , n31818 , n29375 );
xor ( n34454 , n34453 , n29767 );
and ( n34455 , n34452 , n34454 );
xor ( n34456 , n33412 , n34455 );
not ( n34457 , n33424 );
xor ( n34458 , n28072 , n31192 );
xor ( n34459 , n34458 , n27700 );
and ( n34460 , n34457 , n34459 );
xor ( n34461 , n33421 , n34460 );
xor ( n34462 , n34456 , n34461 );
not ( n34463 , n33434 );
xor ( n34464 , n29758 , n33898 );
xor ( n34465 , n34464 , n29051 );
and ( n34466 , n34463 , n34465 );
xor ( n34467 , n33431 , n34466 );
xor ( n34468 , n34462 , n34467 );
not ( n34469 , n33444 );
xor ( n34470 , n29524 , n27819 );
xor ( n34471 , n34470 , n30594 );
and ( n34472 , n34469 , n34471 );
xor ( n34473 , n33441 , n34472 );
xor ( n34474 , n34468 , n34473 );
xor ( n34475 , n34474 , n33408 );
xor ( n34476 , n34451 , n34475 );
and ( n34477 , n34447 , n34476 );
xor ( n34478 , n34341 , n34477 );
not ( n11840 , n29614 );
and ( n11841 , n11840 , RI17514468_703);
and ( n11842 , n34478 , n29614 );
or ( n34479 , n11841 , n11842 );
not ( n11843 , RI1754c610_2);
and ( n11844 , n11843 , n34479 );
and ( n11845 , C0 , RI1754c610_2);
or ( n34480 , n11844 , n11845 );
buf ( n34481 , n34480 );
not ( n34482 , n28544 );
and ( n34483 , n34482 , n28570 );
xor ( n34484 , n29475 , n34483 );
xor ( n34485 , n34484 , n31322 );
not ( n34486 , n28634 );
and ( n34487 , n34486 , n28660 );
xor ( n34488 , n29545 , n34487 );
xor ( n34489 , n34485 , n34488 );
not ( n34490 , n28703 );
and ( n34491 , n34490 , n28728 );
xor ( n34492 , n29588 , n34491 );
xor ( n34493 , n34489 , n34492 );
not ( n34494 , n28772 );
and ( n34495 , n34494 , n28787 );
xor ( n34496 , n29606 , n34495 );
xor ( n34497 , n34493 , n34496 );
xor ( n34498 , n28815 , n34497 );
not ( n34499 , n28840 );
and ( n34500 , n34499 , n28853 );
xor ( n34501 , n31327 , n34500 );
not ( n34502 , n28905 );
and ( n34503 , n34502 , n28930 );
xor ( n34504 , n31339 , n34503 );
xor ( n34505 , n34501 , n34504 );
not ( n34506 , n28957 );
and ( n34507 , n34506 , n28971 );
xor ( n34508 , n31347 , n34507 );
xor ( n34509 , n34505 , n34508 );
not ( n34510 , n29013 );
and ( n34511 , n34510 , n29038 );
xor ( n34512 , n31368 , n34511 );
xor ( n34513 , n34509 , n34512 );
not ( n34514 , n29069 );
and ( n34515 , n34514 , n29081 );
xor ( n34516 , n31376 , n34515 );
xor ( n34517 , n34513 , n34516 );
xor ( n34518 , n34498 , n34517 );
xor ( n34519 , n28272 , n30443 );
xor ( n34520 , n34519 , n28617 );
xor ( n34521 , n28942 , n27936 );
xor ( n34522 , n34521 , n27948 );
not ( n34523 , n34522 );
xor ( n34524 , n30063 , n29105 );
xor ( n34525 , n34524 , n30567 );
and ( n34526 , n34523 , n34525 );
xor ( n34527 , n34520 , n34526 );
xor ( n34528 , n29743 , n28313 );
xor ( n34529 , n34528 , n31683 );
not ( n34530 , n34520 );
and ( n34531 , n34530 , n34522 );
xor ( n34532 , n34529 , n34531 );
xor ( n34533 , n31509 , n28096 );
xor ( n34534 , n34533 , n28107 );
xor ( n34535 , n28486 , n31750 );
xor ( n34536 , n34535 , n30043 );
not ( n34537 , n34536 );
xor ( n34538 , n30864 , n30125 );
xor ( n34539 , n34538 , n31114 );
and ( n34540 , n34537 , n34539 );
xor ( n34541 , n34534 , n34540 );
xor ( n34542 , n34532 , n34541 );
xor ( n34543 , n31674 , n28001 );
xor ( n34544 , n34543 , n30114 );
xor ( n34545 , n30314 , n32996 );
xor ( n34546 , n34545 , n33234 );
not ( n34547 , n34546 );
xor ( n34548 , n29514 , n30655 );
xor ( n34549 , n34548 , n30665 );
and ( n34550 , n34547 , n34549 );
xor ( n34551 , n34544 , n34550 );
xor ( n34552 , n34542 , n34551 );
xor ( n34553 , n32803 , n31422 );
xor ( n34554 , n34553 , n29011 );
xor ( n34555 , n30588 , n28983 );
xor ( n34556 , n34555 , n28995 );
not ( n34557 , n34556 );
xor ( n34558 , n28022 , n30956 );
xor ( n34559 , n34558 , n32130 );
and ( n34560 , n34557 , n34559 );
xor ( n34561 , n34554 , n34560 );
xor ( n34562 , n34552 , n34561 );
xor ( n34563 , n28560 , n30626 );
xor ( n34564 , n34563 , n29740 );
xor ( n34565 , n29380 , n33665 );
xor ( n34566 , n34565 , n32209 );
not ( n34567 , n34566 );
xor ( n34568 , n29444 , n30030 );
xor ( n34569 , n34568 , n30972 );
and ( n34570 , n34567 , n34569 );
xor ( n34571 , n34564 , n34570 );
xor ( n34572 , n34562 , n34571 );
xor ( n34573 , n34527 , n34572 );
xor ( n34574 , n30369 , n28279 );
xor ( n34575 , n34574 , n28291 );
xor ( n34576 , n31035 , n30053 );
xor ( n34577 , n34576 , n31697 );
not ( n34578 , n34577 );
xor ( n34579 , n28462 , n29502 );
xor ( n34580 , n34579 , n29628 );
and ( n34581 , n34578 , n34580 );
xor ( n34582 , n34575 , n34581 );
xor ( n34583 , n30884 , n32734 );
xor ( n34584 , n34583 , n32744 );
xor ( n34585 , n32320 , n29781 );
xor ( n34586 , n34585 , n29793 );
not ( n34587 , n34586 );
xor ( n34588 , n28568 , n30626 );
xor ( n34589 , n34588 , n29740 );
and ( n34590 , n34587 , n34589 );
xor ( n34591 , n34584 , n34590 );
xor ( n34592 , n34582 , n34591 );
xor ( n34593 , n28964 , n32800 );
xor ( n34594 , n34593 , n32809 );
xor ( n34595 , n28012 , n30946 );
xor ( n34596 , n34595 , n30956 );
not ( n34597 , n34596 );
xor ( n34598 , n28249 , n29259 );
xor ( n34599 , n34598 , n29270 );
and ( n34600 , n34597 , n34599 );
xor ( n34601 , n34594 , n34600 );
xor ( n34602 , n34592 , n34601 );
xor ( n34603 , n28362 , n30522 );
xor ( n34604 , n34603 , n32009 );
xor ( n34605 , n30931 , n27752 );
xor ( n34606 , n34605 , n27764 );
not ( n34607 , n34606 );
xor ( n34608 , n27857 , n29655 );
xor ( n34609 , n34608 , n29601 );
and ( n34610 , n34607 , n34609 );
xor ( n34611 , n34604 , n34610 );
xor ( n34612 , n34602 , n34611 );
xor ( n34613 , n28847 , n30306 );
xor ( n34614 , n34613 , n30548 );
xor ( n34615 , n31578 , n29134 );
xor ( n34616 , n34615 , n27936 );
not ( n34617 , n34616 );
xor ( n34618 , n30690 , n30869 );
xor ( n34619 , n34618 , n32894 );
and ( n34620 , n34617 , n34619 );
xor ( n34621 , n34614 , n34620 );
xor ( n34622 , n34612 , n34621 );
xor ( n34623 , n34573 , n34622 );
not ( n34624 , n34623 );
not ( n34625 , n32819 );
and ( n34626 , n34625 , n33002 );
xor ( n34627 , n32816 , n34626 );
xor ( n34628 , n34627 , n32863 );
not ( n34629 , n31752 );
and ( n34630 , n34629 , n31764 );
xor ( n34631 , n33036 , n34630 );
not ( n34632 , n31774 );
and ( n34633 , n34632 , n31776 );
xor ( n34634 , n33044 , n34633 );
xor ( n34635 , n34631 , n34634 );
xor ( n34636 , n34635 , n34131 );
not ( n34637 , n31807 );
and ( n34638 , n34637 , n31809 );
xor ( n34639 , n33060 , n34638 );
xor ( n34640 , n34636 , n34639 );
not ( n34641 , n31827 );
and ( n34642 , n34641 , n31731 );
xor ( n34643 , n33066 , n34642 );
xor ( n34644 , n34640 , n34643 );
xor ( n34645 , n34628 , n34644 );
and ( n34646 , n34624 , n34645 );
xor ( n34647 , n34518 , n34646 );
not ( n11846 , n29614 );
and ( n11847 , n11846 , RI173c0898_1817);
and ( n11848 , n34647 , n29614 );
or ( n34648 , n11847 , n11848 );
not ( n11849 , RI1754c610_2);
and ( n11850 , n11849 , n34648 );
and ( n11851 , C0 , RI1754c610_2);
or ( n34649 , n11850 , n11851 );
buf ( n34650 , n34649 );
not ( n34651 , n33024 );
and ( n34652 , n34651 , n33026 );
xor ( n34653 , n32860 , n34652 );
not ( n34654 , n32810 );
and ( n34655 , n34654 , n32983 );
xor ( n34656 , n32791 , n34655 );
xor ( n34657 , n34656 , n34627 );
not ( n34658 , n32840 );
and ( n34659 , n34658 , n33010 );
xor ( n34660 , n32837 , n34659 );
xor ( n34661 , n34657 , n34660 );
not ( n34662 , n32850 );
and ( n34663 , n34662 , n33016 );
xor ( n34664 , n32847 , n34663 );
xor ( n34665 , n34661 , n34664 );
not ( n34666 , n32860 );
and ( n34667 , n34666 , n33024 );
xor ( n34668 , n32857 , n34667 );
xor ( n34669 , n34665 , n34668 );
xor ( n34670 , n34653 , n34669 );
xor ( n34671 , n34670 , n31831 );
xor ( n34672 , n30716 , n28418 );
xor ( n34673 , n34672 , n31969 );
xor ( n34674 , n30964 , n28852 );
xor ( n34675 , n34674 , n29873 );
not ( n34676 , n34675 );
xor ( n34677 , n29264 , n29093 );
xor ( n34678 , n34677 , n29105 );
and ( n34679 , n34676 , n34678 );
xor ( n34680 , n34673 , n34679 );
xor ( n34681 , n28592 , n29187 );
xor ( n34682 , n34681 , n29724 );
not ( n34683 , n34673 );
and ( n34684 , n34683 , n34675 );
xor ( n34685 , n34682 , n34684 );
xor ( n34686 , n28502 , n30043 );
xor ( n34687 , n34686 , n30053 );
xor ( n34688 , n29223 , n28995 );
xor ( n34689 , n34688 , n30780 );
not ( n34690 , n34689 );
xor ( n34691 , n30466 , n32894 );
xor ( n34692 , n34691 , n32991 );
and ( n34693 , n34690 , n34692 );
xor ( n34694 , n34687 , n34693 );
xor ( n34695 , n34685 , n34694 );
xor ( n34696 , n31906 , n30101 );
xor ( n34697 , n34696 , n32426 );
xor ( n34698 , n27869 , n29601 );
xor ( n34699 , n34698 , n29199 );
not ( n34700 , n34699 );
xor ( n34701 , n29864 , n30548 );
xor ( n34702 , n34701 , n28673 );
and ( n34703 , n34700 , n34702 );
xor ( n34704 , n34697 , n34703 );
xor ( n34705 , n34695 , n34704 );
xor ( n34706 , n33662 , n31367 );
xor ( n34707 , n34706 , n28800 );
xor ( n34708 , n28865 , n30207 );
xor ( n34709 , n34708 , n30218 );
not ( n34710 , n34709 );
xor ( n34711 , n30117 , n31001 );
xor ( n34712 , n34711 , n30889 );
and ( n34713 , n34710 , n34712 );
xor ( n34714 , n34707 , n34713 );
xor ( n34715 , n34705 , n34714 );
xor ( n34716 , n27723 , n28533 );
xor ( n34717 , n34716 , n28543 );
xor ( n34718 , n28235 , n31581 );
xor ( n34719 , n34718 , n28947 );
not ( n34720 , n34719 );
xor ( n34721 , n29429 , n27712 );
xor ( n34722 , n34721 , n30030 );
and ( n34723 , n34720 , n34722 );
xor ( n34724 , n34717 , n34723 );
xor ( n34725 , n34715 , n34724 );
xor ( n34726 , n34680 , n34725 );
xor ( n34727 , n30540 , n28224 );
xor ( n34728 , n34727 , n28236 );
not ( n34729 , n30054 );
and ( n34730 , n34729 , n30067 );
xor ( n34731 , n34728 , n34730 );
xor ( n34732 , n30406 , n30901 );
xor ( n34733 , n34732 , n31475 );
not ( n34734 , n30075 );
and ( n34735 , n34734 , n29996 );
xor ( n34736 , n34733 , n34735 );
xor ( n34737 , n34731 , n34736 );
xor ( n34738 , n28227 , n31581 );
xor ( n34739 , n34738 , n28947 );
not ( n34740 , n30102 );
and ( n34741 , n34740 , n30126 );
xor ( n34742 , n34739 , n34741 );
xor ( n34743 , n34737 , n34742 );
xor ( n34744 , n32728 , n30475 );
xor ( n34745 , n34744 , n30487 );
not ( n34746 , n30166 );
and ( n34747 , n34746 , n30190 );
xor ( n34748 , n34745 , n34747 );
xor ( n34749 , n34743 , n34748 );
xor ( n34750 , n27912 , n30294 );
xor ( n34751 , n34750 , n30306 );
not ( n34752 , n30219 );
and ( n34753 , n34752 , n30222 );
xor ( n34754 , n34751 , n34753 );
xor ( n34755 , n34749 , n34754 );
xor ( n34756 , n34726 , n34755 );
not ( n34757 , n34756 );
xor ( n34758 , n28429 , n32031 );
xor ( n34759 , n34758 , n29975 );
not ( n34760 , n33531 );
and ( n34761 , n34760 , n33533 );
xor ( n34762 , n34759 , n34761 );
xor ( n34763 , n29888 , n29740 );
xor ( n34764 , n34763 , n29752 );
xor ( n34765 , n32417 , n32167 );
xor ( n34766 , n34765 , n31843 );
not ( n34767 , n34766 );
and ( n34768 , n34767 , n33522 );
xor ( n34769 , n34764 , n34768 );
xor ( n34770 , n31064 , n32323 );
xor ( n34771 , n34770 , n32199 );
not ( n34772 , n34759 );
and ( n34773 , n34772 , n33531 );
xor ( n34774 , n34771 , n34773 );
xor ( n34775 , n34769 , n34774 );
xor ( n34776 , n30868 , n30125 );
xor ( n34777 , n34776 , n31114 );
xor ( n34778 , n31836 , n30151 );
xor ( n34779 , n34778 , n31024 );
not ( n34780 , n34779 );
and ( n34781 , n34780 , n33543 );
xor ( n34782 , n34777 , n34781 );
xor ( n34783 , n34775 , n34782 );
xor ( n34784 , n32133 , n29952 );
xor ( n34785 , n34784 , n29964 );
not ( n34786 , n34785 );
and ( n34787 , n34786 , n33553 );
xor ( n34788 , n33518 , n34787 );
xor ( n34789 , n34783 , n34788 );
xor ( n34790 , n31593 , n30178 );
xor ( n34791 , n34790 , n30189 );
xor ( n34792 , n29784 , n30089 );
xor ( n34793 , n34792 , n30101 );
not ( n34794 , n34793 );
and ( n34795 , n34794 , n33559 );
xor ( n34796 , n34791 , n34795 );
xor ( n34797 , n34789 , n34796 );
xor ( n34798 , n34762 , n34797 );
xor ( n34799 , n32503 , n32275 );
xor ( n34800 , n34799 , n31950 );
xor ( n34801 , n27959 , n31131 );
xor ( n34802 , n34801 , n32366 );
not ( n34803 , n34802 );
and ( n34804 , n34803 , n33570 );
xor ( n34805 , n34800 , n34804 );
xor ( n34806 , n31468 , n33198 );
xor ( n34807 , n34806 , n31714 );
xor ( n34808 , n31492 , n28715 );
xor ( n34809 , n34808 , n28727 );
not ( n34810 , n34809 );
and ( n34811 , n34810 , n33579 );
xor ( n34812 , n34807 , n34811 );
xor ( n34813 , n34805 , n34812 );
xor ( n34814 , n31974 , n27897 );
xor ( n34815 , n34814 , n27858 );
xor ( n34816 , n29822 , n32130 );
xor ( n34817 , n34816 , n32140 );
not ( n34818 , n34817 );
and ( n34819 , n34818 , n33589 );
xor ( n34820 , n34815 , n34819 );
xor ( n34821 , n34813 , n34820 );
xor ( n34822 , n30000 , n30567 );
xor ( n34823 , n34822 , n28647 );
xor ( n34824 , n28578 , n29176 );
xor ( n34825 , n34824 , n29187 );
not ( n34826 , n34825 );
and ( n34827 , n34826 , n33599 );
xor ( n34828 , n34823 , n34827 );
xor ( n34829 , n34821 , n34828 );
xor ( n34830 , n30451 , n29123 );
xor ( n34831 , n34830 , n29134 );
xor ( n34832 , n31085 , n29519 );
xor ( n34833 , n34832 , n29320 );
not ( n34834 , n34833 );
and ( n34835 , n34834 , n33609 );
xor ( n34836 , n34831 , n34835 );
xor ( n34837 , n34829 , n34836 );
xor ( n34838 , n34798 , n34837 );
and ( n34839 , n34757 , n34838 );
xor ( n34840 , n34671 , n34839 );
not ( n11852 , n29614 );
and ( n11853 , n11852 , RI1740c6c0_1447);
and ( n11854 , n34840 , n29614 );
or ( n34841 , n11853 , n11854 );
not ( n11855 , RI1754c610_2);
and ( n11856 , n11855 , n34841 );
and ( n11857 , C0 , RI1754c610_2);
or ( n34842 , n11856 , n11857 );
buf ( n34843 , n34842 );
and ( n34844 , RI1754a5b8_71 , RI1754a630_70 , RI1754a6a8_69);
and ( n34845 , RI1754bad0_26 , n34844 );
not ( n34846 , RI1754a5b8_71);
and ( n34847 , n34846 , RI1754a630_70 , RI1754a6a8_69);
and ( n34848 , RI1754bad0_26 , n34847 );
not ( n34849 , RI1754a630_70);
and ( n34850 , RI1754a5b8_71 , n34849 , RI1754a6a8_69);
and ( n34851 , RI1754bad0_26 , n34850 );
and ( n34852 , n34846 , n34849 , RI1754a6a8_69);
and ( n34853 , RI1754bad0_26 , n34852 );
nor ( n34854 , n34846 , n34849 , RI1754a6a8_69);
and ( n34855 , RI1754bad0_26 , n34854 );
nor ( n34856 , RI1754a5b8_71 , n34849 , RI1754a6a8_69);
buf ( n34857 , n34856 );
or ( n34858 , n34845 , n34848 , n34851 , n34853 , n34855 , n34857 , C0 , C0 );
not ( n34859 , RI1754a720_68);
not ( n11858 , n34859 );
and ( n11859 , n11858 , n34858 );
and ( n11860 , RI1754bad0_26 , n34859 );
or ( n34860 , n11859 , n11860 );
not ( n11861 , RI19a22f70_2797);
and ( n11862 , n11861 , n34860 );
and ( n11863 , C0 , RI19a22f70_2797);
or ( n34861 , n11862 , n11863 );
not ( n11864 , n27683 );
and ( n11865 , n11864 , RI19aa29c8_2548);
and ( n11866 , n34861 , n27683 );
or ( n34862 , n11865 , n11866 );
not ( n11867 , RI1754c610_2);
and ( n11868 , n11867 , n34862 );
and ( n11869 , C0 , RI1754c610_2);
or ( n34863 , n11868 , n11869 );
buf ( n34864 , n34863 );
xor ( n34865 , n30004 , n30567 );
xor ( n34866 , n34865 , n28647 );
xor ( n34867 , n30088 , n28339 );
xor ( n34868 , n34867 , n29910 );
not ( n34869 , n34868 );
xor ( n34870 , n28940 , n27936 );
xor ( n34871 , n34870 , n27948 );
and ( n34872 , n34869 , n34871 );
xor ( n34873 , n34866 , n34872 );
xor ( n34874 , n30278 , n31309 );
xor ( n34875 , n34874 , n29519 );
xor ( n34876 , n30854 , n30114 );
xor ( n34877 , n34876 , n30125 );
not ( n34878 , n34877 );
xor ( n34879 , n29078 , n30643 );
xor ( n34880 , n34879 , n29176 );
and ( n34881 , n34878 , n34880 );
xor ( n34882 , n34875 , n34881 );
xor ( n34883 , n28375 , n31909 );
xor ( n34884 , n34883 , n31921 );
xor ( n34885 , n31097 , n29320 );
xor ( n34886 , n34885 , n29332 );
not ( n34887 , n34886 );
xor ( n34888 , n28672 , n28236 );
xor ( n34889 , n34888 , n29711 );
and ( n34890 , n34887 , n34889 );
xor ( n34891 , n34884 , n34890 );
xor ( n34892 , n34882 , n34891 );
xor ( n34893 , n33194 , n30321 );
xor ( n34894 , n34893 , n30332 );
xor ( n34895 , n28712 , n29935 );
xor ( n34896 , n34895 , n31279 );
not ( n34897 , n34896 );
xor ( n34898 , n28916 , n29889 );
xor ( n34899 , n34898 , n30537 );
and ( n34900 , n34897 , n34899 );
xor ( n34901 , n34894 , n34900 );
xor ( n34902 , n34892 , n34901 );
xor ( n34903 , n31362 , n31969 );
xor ( n34904 , n34903 , n31978 );
xor ( n34905 , n32456 , n28583 );
xor ( n34906 , n34905 , n28595 );
not ( n34907 , n34906 );
xor ( n34908 , n28479 , n29224 );
xor ( n34909 , n34908 , n29235 );
and ( n34910 , n34907 , n34909 );
xor ( n34911 , n34904 , n34910 );
xor ( n34912 , n34902 , n34911 );
xor ( n34913 , n28488 , n31750 );
xor ( n34914 , n34913 , n30043 );
not ( n34915 , n34866 );
and ( n34916 , n34915 , n34868 );
xor ( n34917 , n34914 , n34916 );
xor ( n34918 , n34912 , n34917 );
xor ( n34919 , n34873 , n34918 );
xor ( n34920 , n28184 , n29211 );
xor ( n34921 , n34920 , n28557 );
xor ( n34922 , n29772 , n28627 );
xor ( n34923 , n34922 , n30089 );
not ( n34924 , n34923 );
xor ( n34925 , n31094 , n29320 );
xor ( n34926 , n34925 , n29332 );
and ( n34927 , n34924 , n34926 );
xor ( n34928 , n34921 , n34927 );
xor ( n34929 , n28946 , n27936 );
xor ( n34930 , n34929 , n27948 );
xor ( n34931 , n30502 , n29051 );
xor ( n34932 , n34931 , n29062 );
not ( n34933 , n34932 );
xor ( n34934 , n27837 , n30857 );
xor ( n34935 , n34934 , n30869 );
and ( n34936 , n34933 , n34935 );
xor ( n34937 , n34930 , n34936 );
xor ( n34938 , n34928 , n34937 );
xor ( n34939 , n29751 , n28313 );
xor ( n34940 , n34939 , n31683 );
xor ( n34941 , n30081 , n28339 );
xor ( n34942 , n34941 , n29910 );
not ( n34943 , n34942 );
xor ( n34944 , n30183 , n29923 );
xor ( n34945 , n34944 , n29935 );
and ( n34946 , n34943 , n34945 );
xor ( n34947 , n34940 , n34946 );
xor ( n34948 , n34938 , n34947 );
xor ( n34949 , n30779 , n29438 );
xor ( n34950 , n34949 , n29449 );
xor ( n34951 , n28007 , n30946 );
xor ( n34952 , n34951 , n30956 );
not ( n34953 , n34952 );
xor ( n34954 , n28118 , n30233 );
xor ( n34955 , n34954 , n30243 );
and ( n34956 , n34953 , n34955 );
xor ( n34957 , n34950 , n34956 );
xor ( n34958 , n34948 , n34957 );
xor ( n34959 , n32090 , n28380 );
xor ( n34960 , n34959 , n28392 );
xor ( n34961 , n30367 , n28279 );
xor ( n34962 , n34961 , n28291 );
not ( n34963 , n34962 );
xor ( n34964 , n28473 , n29224 );
xor ( n34965 , n34964 , n29235 );
and ( n34966 , n34963 , n34965 );
xor ( n34967 , n34960 , n34966 );
xor ( n34968 , n34958 , n34967 );
xor ( n34969 , n34919 , n34968 );
xor ( n34970 , n27974 , n32366 );
xor ( n34971 , n34970 , n32291 );
xor ( n34972 , n29619 , n30799 );
xor ( n34973 , n34972 , n28148 );
not ( n34974 , n34973 );
and ( n34975 , n34974 , n29188 );
xor ( n34976 , n34971 , n34975 );
not ( n34977 , n34971 );
and ( n34978 , n34977 , n34973 );
xor ( n34979 , n29236 , n34978 );
xor ( n34980 , n32030 , n31874 );
xor ( n34981 , n34980 , n30813 );
not ( n34982 , n34981 );
xor ( n34983 , n27939 , n30374 );
xor ( n34984 , n34983 , n32472 );
and ( n34985 , n34982 , n34984 );
xor ( n34986 , n29274 , n34985 );
xor ( n34987 , n34979 , n34986 );
not ( n34988 , n29163 );
xor ( n34989 , n28141 , n27726 );
xor ( n34990 , n34989 , n27738 );
and ( n34991 , n34988 , n34990 );
xor ( n34992 , n29149 , n34991 );
xor ( n34993 , n34987 , n34992 );
xor ( n34994 , n31988 , n28785 );
xor ( n34995 , n34994 , n28015 );
not ( n34996 , n34995 );
xor ( n34997 , n28676 , n29711 );
xor ( n34998 , n34997 , n30443 );
and ( n34999 , n34996 , n34998 );
xor ( n35000 , n29348 , n34999 );
xor ( n35001 , n34993 , n35000 );
xor ( n35002 , n28542 , n28125 );
xor ( n35003 , n35002 , n28137 );
not ( n35004 , n35003 );
xor ( n35005 , n32374 , n29490 );
xor ( n35006 , n35005 , n29502 );
and ( n35007 , n35004 , n35006 );
xor ( n35008 , n29422 , n35007 );
xor ( n35009 , n35001 , n35008 );
xor ( n35010 , n34976 , n35009 );
xor ( n35011 , n35010 , n28816 );
not ( n35012 , n35011 );
xor ( n35013 , n29926 , n30706 );
xor ( n35014 , n35013 , n30717 );
xor ( n35015 , n32467 , n28291 );
xor ( n35016 , n35015 , n29781 );
not ( n35017 , n35016 );
and ( n35018 , n35017 , n31132 );
xor ( n35019 , n35014 , n35018 );
not ( n35020 , n31101 );
xor ( n35021 , n32737 , n30487 );
xor ( n35022 , n35021 , n30321 );
and ( n35023 , n35020 , n35022 );
xor ( n35024 , n31079 , n35023 );
not ( n35025 , n35014 );
and ( n35026 , n35025 , n35016 );
xor ( n35027 , n31138 , n35026 );
xor ( n35028 , n35024 , n35027 );
xor ( n35029 , n31092 , n29320 );
xor ( n35030 , n35029 , n29332 );
not ( n35031 , n35030 );
xor ( n35032 , n31944 , n29346 );
xor ( n35033 , n35032 , n28866 );
and ( n35034 , n35031 , n35033 );
xor ( n35035 , n31168 , n35034 );
xor ( n35036 , n35028 , n35035 );
xor ( n35037 , n29298 , n31487 );
xor ( n35038 , n35037 , n31497 );
not ( n35039 , n35038 );
xor ( n35040 , n28550 , n30616 );
xor ( n35041 , n35040 , n30626 );
and ( n35042 , n35039 , n35041 );
xor ( n35043 , n31198 , n35042 );
xor ( n35044 , n35036 , n35043 );
xor ( n35045 , n30010 , n28647 );
xor ( n35046 , n35045 , n28659 );
not ( n35047 , n35046 );
xor ( n35048 , n28764 , n30934 );
xor ( n35049 , n35048 , n28533 );
and ( n35050 , n35047 , n35049 );
xor ( n35051 , n31210 , n35050 );
xor ( n35052 , n35044 , n35051 );
xor ( n35053 , n35019 , n35052 );
not ( n35054 , n33199 );
and ( n35055 , n35054 , n33625 );
xor ( n35056 , n31232 , n35055 );
not ( n35057 , n33204 );
and ( n35058 , n35057 , n33630 );
xor ( n35059 , n31252 , n35058 );
xor ( n35060 , n35056 , n35059 );
xor ( n35061 , n35060 , n33188 );
not ( n35062 , n33214 );
and ( n35063 , n35062 , n33640 );
xor ( n35064 , n31292 , n35063 );
xor ( n35065 , n35061 , n35064 );
not ( n35066 , n33220 );
and ( n35067 , n35066 , n33620 );
xor ( n35068 , n31314 , n35067 );
xor ( n35069 , n35065 , n35068 );
xor ( n35070 , n35053 , n35069 );
and ( n35071 , n35012 , n35070 );
xor ( n35072 , n34969 , n35071 );
not ( n11870 , n29614 );
and ( n11871 , n11870 , RI17407170_1473);
and ( n11872 , n35072 , n29614 );
or ( n35073 , n11871 , n11872 );
not ( n11873 , RI1754c610_2);
and ( n11874 , n11873 , n35073 );
and ( n11875 , C0 , RI1754c610_2);
or ( n35074 , n11874 , n11875 );
buf ( n35075 , n35074 );
not ( n35076 , n33694 );
and ( n35077 , n35076 , n33274 );
xor ( n35078 , n33691 , n35077 );
xor ( n35079 , n35078 , n33697 );
xor ( n35080 , n32037 , n31825 );
xor ( n35081 , n35080 , n29586 );
xor ( n35082 , n29359 , n31763 );
xor ( n35083 , n35082 , n31989 );
not ( n35084 , n35083 );
xor ( n35085 , n30136 , n28392 );
xor ( n35086 , n35085 , n30918 );
and ( n35087 , n35084 , n35086 );
xor ( n35088 , n35081 , n35087 );
xor ( n35089 , n31902 , n30101 );
xor ( n35090 , n35089 , n32426 );
xor ( n35091 , n32287 , n31399 );
xor ( n35092 , n35091 , n29561 );
not ( n35093 , n35092 );
xor ( n35094 , n29764 , n33898 );
xor ( n35095 , n35094 , n29051 );
and ( n35096 , n35093 , n35095 );
xor ( n35097 , n35090 , n35096 );
xor ( n35098 , n35088 , n35097 );
xor ( n35099 , n30393 , n27807 );
xor ( n35100 , n35099 , n27819 );
xor ( n35101 , n29930 , n30706 );
xor ( n35102 , n35101 , n30717 );
not ( n35103 , n35102 );
xor ( n35104 , n28980 , n28081 );
xor ( n35105 , n35104 , n29248 );
and ( n35106 , n35103 , n35105 );
xor ( n35107 , n35100 , n35106 );
xor ( n35108 , n35098 , n35107 );
xor ( n35109 , n29745 , n28313 );
xor ( n35110 , n35109 , n31683 );
xor ( n35111 , n27707 , n27909 );
xor ( n35112 , n35111 , n27921 );
not ( n35113 , n35112 );
xor ( n35114 , n28944 , n27936 );
xor ( n35115 , n35114 , n27948 );
and ( n35116 , n35113 , n35115 );
xor ( n35117 , n35110 , n35116 );
xor ( n35118 , n35108 , n35117 );
xor ( n35119 , n32114 , n28137 );
xor ( n35120 , n35119 , n28493 );
xor ( n35121 , n30120 , n31001 );
xor ( n35122 , n35121 , n30889 );
not ( n35123 , n35122 );
xor ( n35124 , n30484 , n32991 );
xor ( n35125 , n35124 , n32996 );
and ( n35126 , n35123 , n35125 );
xor ( n35127 , n35120 , n35126 );
xor ( n35128 , n35118 , n35127 );
xor ( n35129 , n35079 , n35128 );
xor ( n35130 , n28720 , n31279 );
xor ( n35131 , n35130 , n33665 );
xor ( n35132 , n30702 , n28406 );
xor ( n35133 , n35132 , n28418 );
not ( n35134 , n35133 );
and ( n35135 , n35134 , n31952 );
xor ( n35136 , n35131 , n35135 );
not ( n35137 , n35131 );
and ( n35138 , n35137 , n35133 );
xor ( n35139 , n31957 , n35138 );
or ( n35140 , RI1753a460_587 , RI17539830_589);
or ( n35141 , n35140 , RI17539218_590);
or ( n35142 , n35141 , RI17538c00_591);
or ( n35143 , n35142 , RI17537fd0_593);
or ( n35144 , n35143 , RI175379b8_594);
or ( n35145 , n35144 , RI17536770_597);
xor ( n35146 , n35139 , n35145 );
xor ( n35147 , n27968 , n32366 );
xor ( n35148 , n35147 , n32291 );
not ( n35149 , n35148 );
xor ( n35150 , n29959 , n30164 );
xor ( n35151 , n35150 , n29490 );
and ( n35152 , n35149 , n35151 );
xor ( n35153 , n31993 , n35152 );
xor ( n35154 , n35146 , n35153 );
xor ( n35155 , n30928 , n27752 );
xor ( n35156 , n35155 , n27764 );
not ( n35157 , n35156 );
xor ( n35158 , n27814 , n33390 );
xor ( n35159 , n35158 , n28983 );
and ( n35160 , n35157 , n35159 );
xor ( n35161 , n32010 , n35160 );
xor ( n35162 , n35154 , n35161 );
not ( n35163 , n31938 );
xor ( n35164 , n29266 , n29093 );
xor ( n35165 , n35164 , n29105 );
and ( n35166 , n35163 , n35165 );
xor ( n35167 , n31935 , n35166 );
xor ( n35168 , n35162 , n35167 );
xor ( n35169 , n30835 , n27833 );
xor ( n35170 , n35169 , n27844 );
not ( n35171 , n35170 );
xor ( n35172 , n32163 , n30139 );
xor ( n35173 , n35172 , n30151 );
and ( n35174 , n35171 , n35173 );
xor ( n35175 , n32045 , n35174 );
xor ( n35176 , n35168 , n35175 );
xor ( n35177 , n35136 , n35176 );
xor ( n35178 , n28863 , n30207 );
xor ( n35179 , n35178 , n30218 );
not ( n35180 , n35179 );
xor ( n35181 , n31088 , n29519 );
xor ( n35182 , n35181 , n29320 );
and ( n35183 , n35180 , n35182 );
xor ( n35184 , n32056 , n35183 );
xor ( n35185 , n27894 , n29399 );
xor ( n35186 , n35185 , n29655 );
not ( n35187 , n35186 );
xor ( n35188 , n28784 , n32043 );
xor ( n35189 , n35188 , n30946 );
and ( n35190 , n35187 , n35189 );
xor ( n35191 , n32065 , n35190 );
xor ( n35192 , n35184 , n35191 );
xor ( n35193 , n29256 , n32120 );
xor ( n35194 , n35193 , n29093 );
not ( n35195 , n35194 );
xor ( n35196 , n31527 , n28107 );
xor ( n35197 , n35196 , n32510 );
and ( n35198 , n35195 , n35197 );
xor ( n35199 , n32075 , n35198 );
xor ( n35200 , n35192 , n35199 );
xor ( n35201 , n32798 , n31100 );
xor ( n35202 , n35201 , n31422 );
not ( n35203 , n35202 );
xor ( n35204 , n31000 , n32256 );
xor ( n35205 , n35204 , n32734 );
and ( n35206 , n35203 , n35205 );
xor ( n35207 , n32095 , n35206 );
xor ( n35208 , n35200 , n35207 );
xor ( n35209 , n27788 , n29306 );
xor ( n35210 , n35209 , n28406 );
not ( n35211 , n35210 );
xor ( n35212 , n31873 , n29964 );
xor ( n35213 , n35212 , n32382 );
and ( n35214 , n35211 , n35213 );
xor ( n35215 , n32105 , n35214 );
xor ( n35216 , n35208 , n35215 );
xor ( n35217 , n35177 , n35216 );
not ( n35218 , n35217 );
xor ( n35219 , n28120 , n30233 );
xor ( n35220 , n35219 , n30243 );
xor ( n35221 , n28580 , n29176 );
xor ( n35222 , n35221 , n29187 );
not ( n35223 , n35222 );
xor ( n35224 , n32008 , n31613 );
xor ( n35225 , n35224 , n28438 );
and ( n35226 , n35223 , n35225 );
xor ( n35227 , n35220 , n35226 );
xor ( n35228 , n29192 , n28212 );
xor ( n35229 , n35228 , n32459 );
xor ( n35230 , n29850 , n29421 );
xor ( n35231 , n35230 , n30643 );
not ( n35232 , n35231 );
xor ( n35233 , n28078 , n31192 );
xor ( n35234 , n35233 , n27700 );
and ( n35235 , n35232 , n35234 );
xor ( n35236 , n35229 , n35235 );
xor ( n35237 , n29525 , n27819 );
xor ( n35238 , n35237 , n30594 );
not ( n35239 , n35220 );
and ( n35240 , n35239 , n35222 );
xor ( n35241 , n35238 , n35240 );
xor ( n35242 , n35236 , n35241 );
xor ( n35243 , n29098 , n28505 );
xor ( n35244 , n35243 , n31038 );
xor ( n35245 , n30301 , n28055 );
xor ( n35246 , n35245 , n28224 );
not ( n35247 , n35246 );
xor ( n35248 , n31694 , n29291 );
xor ( n35249 , n35248 , n31636 );
and ( n35250 , n35247 , n35249 );
xor ( n35251 , n35244 , n35250 );
xor ( n35252 , n35242 , n35251 );
xor ( n35253 , n30171 , n31162 );
xor ( n35254 , n35253 , n29923 );
xor ( n35255 , n31789 , n29148 );
xor ( n35256 , n35255 , n32800 );
not ( n35257 , n35256 );
xor ( n35258 , n32832 , n32510 );
xor ( n35259 , n35258 , n29462 );
and ( n35260 , n35257 , n35259 );
xor ( n35261 , n35254 , n35260 );
xor ( n35262 , n35252 , n35261 );
xor ( n35263 , n33192 , n30321 );
xor ( n35264 , n35263 , n30332 );
xor ( n35265 , n30712 , n28418 );
xor ( n35266 , n35265 , n31969 );
not ( n35267 , n35266 );
xor ( n35268 , n29396 , n32209 );
xor ( n35269 , n35268 , n30389 );
and ( n35270 , n35267 , n35269 );
xor ( n35271 , n35264 , n35270 );
xor ( n35272 , n35262 , n35271 );
xor ( n35273 , n35227 , n35272 );
xor ( n35274 , n35273 , n35009 );
and ( n35275 , n35218 , n35274 );
xor ( n35276 , n35129 , n35275 );
not ( n11876 , n29614 );
and ( n11877 , n11876 , RI173c2cb0_1806);
and ( n11878 , n35276 , n29614 );
or ( n35277 , n11877 , n11878 );
not ( n11879 , RI1754c610_2);
and ( n11880 , n11879 , n35277 );
and ( n11881 , C0 , RI1754c610_2);
or ( n35278 , n11880 , n11881 );
buf ( n35279 , n35278 );
not ( n11882 , n27683 );
and ( n11883 , n11882 , RI19aa3238_2544);
and ( n11884 , RI19aad468_2473 , n27683 );
or ( n35280 , n11883 , n11884 );
not ( n11885 , RI1754c610_2);
and ( n11886 , n11885 , n35280 );
and ( n11887 , C0 , RI1754c610_2);
or ( n35281 , n11886 , n11887 );
buf ( n35282 , n35281 );
xor ( n35283 , n29100 , n28505 );
xor ( n35284 , n35283 , n31038 );
not ( n35285 , n30250 );
and ( n35286 , n35285 , n30253 );
xor ( n35287 , n35284 , n35286 );
xor ( n35288 , n28697 , n32472 );
xor ( n35289 , n35288 , n32323 );
not ( n35290 , n30284 );
and ( n35291 , n35290 , n30307 );
xor ( n35292 , n35289 , n35291 );
xor ( n35293 , n35287 , n35292 );
xor ( n35294 , n30996 , n32256 );
xor ( n35295 , n35294 , n32734 );
not ( n35296 , n30350 );
and ( n35297 , n35296 , n30352 );
xor ( n35298 , n35295 , n35297 );
xor ( n35299 , n35293 , n35298 );
xor ( n35300 , n29918 , n27791 );
xor ( n35301 , n35300 , n30706 );
not ( n35302 , n30391 );
and ( n35303 , n35302 , n30401 );
xor ( n35304 , n35301 , n35303 );
xor ( n35305 , n35299 , n35304 );
xor ( n35306 , n28528 , n27764 );
xor ( n35307 , n35306 , n28125 );
not ( n35308 , n30433 );
and ( n35309 , n35308 , n30445 );
xor ( n35310 , n35307 , n35309 );
xor ( n35311 , n35305 , n35310 );
xor ( n35312 , n30430 , n35311 );
xor ( n35313 , n29408 , n27858 );
xor ( n35314 , n35313 , n27870 );
xor ( n35315 , n30355 , n28684 );
xor ( n35316 , n35315 , n28279 );
not ( n35317 , n35316 );
xor ( n35318 , n28640 , n30271 );
xor ( n35319 , n35318 , n30283 );
and ( n35320 , n35317 , n35319 );
xor ( n35321 , n35314 , n35320 );
xor ( n35322 , n28054 , n29694 );
xor ( n35323 , n35322 , n30457 );
xor ( n35324 , n33227 , n29364 );
xor ( n35325 , n35324 , n29375 );
not ( n35326 , n35325 );
xor ( n35327 , n29882 , n29740 );
xor ( n35328 , n35327 , n29752 );
and ( n35329 , n35326 , n35328 );
xor ( n35330 , n35323 , n35329 );
xor ( n35331 , n35321 , n35330 );
xor ( n35332 , n28556 , n30616 );
xor ( n35333 , n35332 , n30626 );
xor ( n35334 , n28270 , n30443 );
xor ( n35335 , n35334 , n28617 );
not ( n35336 , n35335 );
xor ( n35337 , n28385 , n31921 );
xor ( n35338 , n35337 , n30348 );
and ( n35339 , n35336 , n35338 );
xor ( n35340 , n35333 , n35339 );
xor ( n35341 , n35331 , n35340 );
xor ( n35342 , n27818 , n33390 );
xor ( n35343 , n35342 , n28983 );
xor ( n35344 , n31467 , n33198 );
xor ( n35345 , n35344 , n31714 );
not ( n35346 , n35345 );
xor ( n35347 , n30818 , n28463 );
xor ( n35348 , n35347 , n27752 );
and ( n35349 , n35346 , n35348 );
xor ( n35350 , n35343 , n35349 );
xor ( n35351 , n35341 , n35350 );
xor ( n35352 , n29994 , n28702 );
xor ( n35353 , n35352 , n31065 );
xor ( n35354 , n29114 , n29873 );
xor ( n35355 , n35354 , n32398 );
not ( n35356 , n35355 );
xor ( n35357 , n29030 , n30399 );
xor ( n35358 , n35357 , n29532 );
and ( n35359 , n35356 , n35358 );
xor ( n35360 , n35353 , n35359 );
xor ( n35361 , n35351 , n35360 );
xor ( n35362 , n35312 , n35361 );
xor ( n35363 , n28994 , n29248 );
xor ( n35364 , n35363 , n29438 );
xor ( n35365 , n32603 , n29025 );
xor ( n35366 , n35365 , n29037 );
not ( n35367 , n35366 );
xor ( n35368 , n28962 , n32800 );
xor ( n35369 , n35368 , n32809 );
and ( n35370 , n35367 , n35369 );
xor ( n35371 , n35364 , n35370 );
xor ( n35372 , n28797 , n31978 );
xor ( n35373 , n35372 , n29409 );
xor ( n35374 , n32166 , n30139 );
xor ( n35375 , n35374 , n30151 );
not ( n35376 , n35375 );
xor ( n35377 , n31173 , n29532 );
xor ( n35378 , n35377 , n29544 );
and ( n35379 , n35376 , n35378 );
xor ( n35380 , n35373 , n35379 );
xor ( n35381 , n27749 , n29628 );
xor ( n35382 , n35381 , n29639 );
xor ( n35383 , n30206 , n29561 );
xor ( n35384 , n35383 , n29573 );
not ( n35385 , n35384 );
xor ( n35386 , n29732 , n28304 );
xor ( n35387 , n35386 , n28313 );
and ( n35388 , n35385 , n35387 );
xor ( n35389 , n35382 , n35388 );
xor ( n35390 , n35380 , n35389 );
xor ( n35391 , n28681 , n29711 );
xor ( n35392 , n35391 , n30443 );
xor ( n35393 , n31496 , n28715 );
xor ( n35394 , n35393 , n28727 );
not ( n35395 , n35394 );
xor ( n35396 , n29535 , n30594 );
xor ( n35397 , n35396 , n29224 );
and ( n35398 , n35395 , n35397 );
xor ( n35399 , n35392 , n35398 );
xor ( n35400 , n35390 , n35399 );
xor ( n35401 , n31149 , n31843 );
xor ( n35402 , n35401 , n27779 );
xor ( n35403 , n31421 , n29332 );
xor ( n35404 , n35403 , n29814 );
not ( n35405 , n35404 );
xor ( n35406 , n29716 , n28839 );
xor ( n35407 , n35406 , n28917 );
and ( n35408 , n35405 , n35407 );
xor ( n35409 , n35402 , n35408 );
xor ( n35410 , n35400 , n35409 );
xor ( n35411 , n29836 , n32140 );
xor ( n35412 , n35411 , n31874 );
not ( n35413 , n35364 );
and ( n35414 , n35413 , n35366 );
xor ( n35415 , n35412 , n35414 );
xor ( n35416 , n35410 , n35415 );
xor ( n35417 , n35371 , n35416 );
xor ( n35418 , n35417 , n29843 );
not ( n35419 , n35418 );
not ( n35420 , n32223 );
and ( n35421 , n35420 , n32225 );
xor ( n35422 , n32633 , n35421 );
not ( n35423 , n32633 );
and ( n35424 , n35423 , n32223 );
xor ( n35425 , n32630 , n35424 );
xor ( n35426 , n35425 , n32628 );
not ( n35427 , n32644 );
and ( n35428 , n35427 , n32262 );
xor ( n35429 , n32641 , n35428 );
xor ( n35430 , n35426 , n35429 );
not ( n35431 , n32652 );
and ( n35432 , n35431 , n32281 );
xor ( n35433 , n32649 , n35432 );
xor ( n35434 , n35430 , n35433 );
not ( n35435 , n32660 );
and ( n35436 , n35435 , n32301 );
xor ( n35437 , n32657 , n35436 );
xor ( n35438 , n35434 , n35437 );
xor ( n35439 , n35422 , n35438 );
not ( n35440 , n32673 );
and ( n35441 , n35440 , n32880 );
xor ( n35442 , n32670 , n35441 );
not ( n35443 , n32682 );
and ( n35444 , n35443 , n32895 );
xor ( n35445 , n32679 , n35444 );
xor ( n35446 , n35442 , n35445 );
not ( n35447 , n32692 );
and ( n35448 , n35447 , n32901 );
xor ( n35449 , n32689 , n35448 );
xor ( n35450 , n35446 , n35449 );
not ( n35451 , n32702 );
and ( n35452 , n35451 , n32909 );
xor ( n35453 , n32699 , n35452 );
xor ( n35454 , n35450 , n35453 );
not ( n35455 , n32712 );
and ( n35456 , n35455 , n32917 );
xor ( n35457 , n32709 , n35456 );
xor ( n35458 , n35454 , n35457 );
xor ( n35459 , n35439 , n35458 );
and ( n35460 , n35419 , n35459 );
xor ( n35461 , n35362 , n35460 );
not ( n11888 , n29614 );
and ( n11889 , n11888 , RI1748d540_1047);
and ( n11890 , n35461 , n29614 );
or ( n35462 , n11889 , n11890 );
not ( n11891 , RI1754c610_2);
and ( n11892 , n11891 , n35462 );
and ( n11893 , C0 , RI1754c610_2);
or ( n35463 , n11892 , n11893 );
buf ( n35464 , n35463 );
xor ( n35465 , n30107 , n32778 );
xor ( n35466 , n35465 , n31001 );
not ( n35467 , n30568 );
and ( n35468 , n35467 , n30488 );
xor ( n35469 , n35466 , n35468 );
xor ( n35470 , n29687 , n30972 );
xor ( n35471 , n35470 , n29123 );
not ( n35472 , n35471 );
and ( n35473 , n35472 , n30497 );
xor ( n35474 , n31645 , n35473 );
xor ( n35475 , n30793 , n28771 );
xor ( n35476 , n35475 , n27726 );
not ( n35477 , n35476 );
and ( n35478 , n35477 , n30538 );
xor ( n35479 , n31650 , n35478 );
xor ( n35480 , n35474 , n35479 );
not ( n35481 , n35466 );
and ( n35482 , n35481 , n30568 );
xor ( n35483 , n30493 , n35482 );
xor ( n35484 , n35480 , n35483 );
not ( n35485 , n31640 );
and ( n35486 , n35485 , n30575 );
xor ( n35487 , n31637 , n35486 );
xor ( n35488 , n35484 , n35487 );
xor ( n35489 , n27772 , n31024 );
xor ( n35490 , n35489 , n29306 );
not ( n35491 , n35490 );
and ( n35492 , n35491 , n30595 );
xor ( n35493 , n31661 , n35492 );
xor ( n35494 , n35488 , n35493 );
xor ( n35495 , n35469 , n35494 );
not ( n35496 , n33701 );
and ( n35497 , n35496 , n30607 );
xor ( n35498 , n31668 , n35497 );
not ( n35499 , n33706 );
and ( n35500 , n35499 , n30644 );
xor ( n35501 , n31684 , n35500 );
xor ( n35502 , n35498 , n35501 );
not ( n35503 , n33712 );
and ( n35504 , n35503 , n30675 );
xor ( n35505 , n31698 , n35504 );
xor ( n35506 , n35502 , n35505 );
not ( n35507 , n33718 );
and ( n35508 , n35507 , n30718 );
xor ( n35509 , n31716 , n35508 );
xor ( n35510 , n35506 , n35509 );
not ( n35511 , n33724 );
and ( n35512 , n35511 , n30731 );
xor ( n35513 , n31722 , n35512 );
xor ( n35514 , n35510 , n35513 );
xor ( n35515 , n35495 , n35514 );
xor ( n35516 , n29988 , n28702 );
xor ( n35517 , n35516 , n31065 );
not ( n35518 , n34575 );
and ( n35519 , n35518 , n34577 );
xor ( n35520 , n35517 , n35519 );
xor ( n35521 , n28885 , n30066 );
xor ( n35522 , n35521 , n30007 );
not ( n35523 , n34584 );
and ( n35524 , n35523 , n34586 );
xor ( n35525 , n35522 , n35524 );
xor ( n35526 , n35520 , n35525 );
xor ( n35527 , n29357 , n31763 );
xor ( n35528 , n35527 , n31989 );
not ( n35529 , n34594 );
and ( n35530 , n35529 , n34596 );
xor ( n35531 , n35528 , n35530 );
xor ( n35532 , n35526 , n35531 );
xor ( n35533 , n29241 , n27700 );
xor ( n35534 , n35533 , n27712 );
not ( n35535 , n34604 );
and ( n35536 , n35535 , n34606 );
xor ( n35537 , n35534 , n35536 );
xor ( n35538 , n35532 , n35537 );
xor ( n35539 , n28793 , n31978 );
xor ( n35540 , n35539 , n29409 );
not ( n35541 , n34614 );
and ( n35542 , n35541 , n34616 );
xor ( n35543 , n35540 , n35542 );
xor ( n35544 , n35538 , n35543 );
xor ( n35545 , n34611 , n35544 );
xor ( n35546 , n29288 , n30017 );
xor ( n35547 , n35546 , n30986 );
xor ( n35548 , n30798 , n28771 );
xor ( n35549 , n35548 , n27726 );
not ( n35550 , n35549 );
xor ( n35551 , n32239 , n27844 );
xor ( n35552 , n35551 , n30691 );
and ( n35553 , n35550 , n35552 );
xor ( n35554 , n35547 , n35553 );
xor ( n35555 , n30086 , n28339 );
xor ( n35556 , n35555 , n29910 );
xor ( n35557 , n28303 , n31291 );
xor ( n35558 , n35557 , n27989 );
not ( n35559 , n35558 );
xor ( n35560 , n32357 , n32835 );
xor ( n35561 , n35560 , n31399 );
and ( n35562 , n35559 , n35561 );
xor ( n35563 , n35556 , n35562 );
xor ( n35564 , n35554 , n35563 );
xor ( n35565 , n28352 , n30510 );
xor ( n35566 , n35565 , n30522 );
xor ( n35567 , n29092 , n28493 );
xor ( n35568 , n35567 , n28505 );
not ( n35569 , n35568 );
xor ( n35570 , n30682 , n30869 );
xor ( n35571 , n35570 , n32894 );
and ( n35572 , n35569 , n35571 );
xor ( n35573 , n35566 , n35572 );
xor ( n35574 , n35564 , n35573 );
xor ( n35575 , n29636 , n28148 );
xor ( n35576 , n35575 , n28160 );
xor ( n35577 , n28199 , n29855 );
xor ( n35578 , n35577 , n29079 );
not ( n35579 , n35578 );
xor ( n35580 , n28099 , n31462 );
xor ( n35581 , n35580 , n32275 );
and ( n35582 , n35579 , n35581 );
xor ( n35583 , n35576 , n35582 );
xor ( n35584 , n35574 , n35583 );
xor ( n35585 , n30361 , n28684 );
xor ( n35586 , n35585 , n28279 );
xor ( n35587 , n31113 , n30889 );
xor ( n35588 , n35587 , n30901 );
not ( n35589 , n35588 );
xor ( n35590 , n28920 , n30537 );
xor ( n35591 , n35590 , n30842 );
and ( n35592 , n35589 , n35591 );
xor ( n35593 , n35586 , n35592 );
xor ( n35594 , n35584 , n35593 );
xor ( n35595 , n35545 , n35594 );
not ( n35596 , n35595 );
xor ( n35597 , n30460 , n35311 );
xor ( n35598 , n35597 , n35361 );
and ( n35599 , n35596 , n35598 );
xor ( n35600 , n35515 , n35599 );
not ( n11894 , n29614 );
and ( n11895 , n11894 , RI173e95a8_1618);
and ( n11896 , n35600 , n29614 );
or ( n35601 , n11895 , n11896 );
not ( n11897 , RI1754c610_2);
and ( n11898 , n11897 , n35601 );
and ( n11899 , C0 , RI1754c610_2);
or ( n35602 , n11898 , n11899 );
buf ( n35603 , n35602 );
not ( n35604 , n32406 );
and ( n35605 , n35604 , n32408 );
xor ( n35606 , n32748 , n35605 );
not ( n35607 , n32415 );
and ( n35608 , n35607 , n32428 );
xor ( n35609 , n32755 , n35608 );
xor ( n35610 , n35606 , n35609 );
not ( n35611 , n32436 );
and ( n35612 , n35611 , n32438 );
xor ( n35613 , n32723 , n35612 );
xor ( n35614 , n35610 , n35613 );
not ( n35615 , n32446 );
and ( n35616 , n35615 , n32448 );
xor ( n35617 , n32767 , n35616 );
xor ( n35618 , n35614 , n35617 );
not ( n35619 , n32466 );
and ( n35620 , n35619 , n32474 );
xor ( n35621 , n32783 , n35620 );
xor ( n35622 , n35618 , n35621 );
xor ( n35623 , n32463 , n35622 );
not ( n35624 , n32983 );
and ( n35625 , n35624 , n32997 );
xor ( n35626 , n32810 , n35625 );
not ( n35627 , n33002 );
and ( n35628 , n35627 , n33004 );
xor ( n35629 , n32819 , n35628 );
xor ( n35630 , n35626 , n35629 );
not ( n35631 , n33010 );
and ( n35632 , n35631 , n32978 );
xor ( n35633 , n32840 , n35632 );
xor ( n35634 , n35630 , n35633 );
not ( n35635 , n33016 );
and ( n35636 , n35635 , n33018 );
xor ( n35637 , n32850 , n35636 );
xor ( n35638 , n35634 , n35637 );
xor ( n35639 , n35638 , n34653 );
xor ( n35640 , n35623 , n35639 );
not ( n35641 , n34969 );
and ( n35642 , n35641 , n35011 );
xor ( n35643 , n35640 , n35642 );
not ( n11900 , n29614 );
and ( n11901 , n11900 , RI173f8530_1545);
and ( n11902 , n35643 , n29614 );
or ( n35644 , n11901 , n11902 );
not ( n11903 , RI1754c610_2);
and ( n11904 , n11903 , n35644 );
and ( n11905 , C0 , RI1754c610_2);
or ( n35645 , n11904 , n11905 );
buf ( n35646 , n35645 );
buf ( n35647 , RI174bf130_816);
buf ( n35648 , RI174968e8_1002);
buf ( n35649 , RI17463150_1253);
not ( n35650 , n33953 );
xor ( n35651 , n30203 , n29561 );
xor ( n35652 , n35651 , n29573 );
and ( n35653 , n35650 , n35652 );
xor ( n35654 , n33950 , n35653 );
xor ( n35655 , n35654 , n33991 );
xor ( n35656 , n35655 , n34041 );
xor ( n35657 , n28708 , n29935 );
xor ( n35658 , n35657 , n31279 );
xor ( n35659 , n30590 , n28983 );
xor ( n35660 , n35659 , n28995 );
not ( n35661 , n35660 );
xor ( n35662 , n29487 , n28450 );
xor ( n35663 , n35662 , n30789 );
and ( n35664 , n35661 , n35663 );
xor ( n35665 , n35658 , n35664 );
xor ( n35666 , n28869 , n30218 );
xor ( n35667 , n35666 , n27807 );
xor ( n35668 , n31867 , n29964 );
xor ( n35669 , n35668 , n32382 );
not ( n35670 , n35669 );
xor ( n35671 , n32004 , n31613 );
xor ( n35672 , n35671 , n28438 );
and ( n35673 , n35670 , n35672 );
xor ( n35674 , n35667 , n35673 );
xor ( n35675 , n28586 , n29187 );
xor ( n35676 , n35675 , n29724 );
not ( n35677 , n35658 );
and ( n35678 , n35677 , n35660 );
xor ( n35679 , n35676 , n35678 );
xor ( n35680 , n35674 , n35679 );
xor ( n35681 , n27798 , n30758 );
xor ( n35682 , n35681 , n33390 );
xor ( n35683 , n27914 , n30294 );
xor ( n35684 , n35683 , n30306 );
not ( n35685 , n35684 );
xor ( n35686 , n28195 , n29855 );
xor ( n35687 , n35686 , n29079 );
and ( n35688 , n35685 , n35687 );
xor ( n35689 , n35682 , n35688 );
xor ( n35690 , n35680 , n35689 );
xor ( n35691 , n28177 , n29211 );
xor ( n35692 , n35691 , n28557 );
xor ( n35693 , n30480 , n32991 );
xor ( n35694 , n35693 , n32996 );
not ( n35695 , n35694 );
xor ( n35696 , n27931 , n30364 );
xor ( n35697 , n35696 , n30374 );
and ( n35698 , n35695 , n35697 );
xor ( n35699 , n35692 , n35698 );
xor ( n35700 , n35690 , n35699 );
xor ( n35701 , n31942 , n29346 );
xor ( n35702 , n35701 , n28866 );
xor ( n35703 , n28652 , n30283 );
xor ( n35704 , n35703 , n31089 );
not ( n35705 , n35704 );
xor ( n35706 , n29370 , n31989 );
xor ( n35707 , n35706 , n33898 );
and ( n35708 , n35705 , n35707 );
xor ( n35709 , n35702 , n35708 );
xor ( n35710 , n35700 , n35709 );
xor ( n35711 , n35665 , n35710 );
xor ( n35712 , n32026 , n31874 );
xor ( n35713 , n35712 , n30813 );
xor ( n35714 , n29384 , n33665 );
xor ( n35715 , n35714 , n32209 );
not ( n35716 , n35715 );
xor ( n35717 , n31908 , n30101 );
xor ( n35718 , n35717 , n32426 );
and ( n35719 , n35716 , n35718 );
xor ( n35720 , n35713 , n35719 );
xor ( n35721 , n29243 , n27700 );
xor ( n35722 , n35721 , n27712 );
xor ( n35723 , n28756 , n30823 );
xor ( n35724 , n35723 , n30934 );
not ( n35725 , n35724 );
xor ( n35726 , n31949 , n29346 );
xor ( n35727 , n35726 , n28866 );
and ( n35728 , n35725 , n35727 );
xor ( n35729 , n35722 , n35728 );
xor ( n35730 , n35720 , n35729 );
xor ( n35731 , n30639 , n28174 );
xor ( n35732 , n35731 , n28185 );
xor ( n35733 , n29131 , n32398 );
xor ( n35734 , n35733 , n30364 );
not ( n35735 , n35734 );
xor ( n35736 , n27790 , n29306 );
xor ( n35737 , n35736 , n28406 );
and ( n35738 , n35735 , n35737 );
xor ( n35739 , n35732 , n35738 );
xor ( n35740 , n35730 , n35739 );
xor ( n35741 , n28274 , n30443 );
xor ( n35742 , n35741 , n28617 );
xor ( n35743 , n28389 , n31921 );
xor ( n35744 , n35743 , n30348 );
not ( n35745 , n35744 );
xor ( n35746 , n28968 , n32800 );
xor ( n35747 , n35746 , n32809 );
and ( n35748 , n35745 , n35747 );
xor ( n35749 , n35742 , n35748 );
xor ( n35750 , n35740 , n35749 );
xor ( n35751 , n28010 , n30946 );
xor ( n35752 , n35751 , n30956 );
xor ( n35753 , n30519 , n29062 );
xor ( n35754 , n35753 , n31613 );
not ( n35755 , n35754 );
xor ( n35756 , n29543 , n30594 );
xor ( n35757 , n35756 , n29224 );
and ( n35758 , n35755 , n35757 );
xor ( n35759 , n35752 , n35758 );
xor ( n35760 , n35750 , n35759 );
xor ( n35761 , n35711 , n35760 );
not ( n35762 , n35761 );
xor ( n35763 , n27853 , n29655 );
xor ( n35764 , n35763 , n29601 );
not ( n35765 , n33359 );
and ( n35766 , n35765 , n33361 );
xor ( n35767 , n35764 , n35766 );
xor ( n35768 , n31606 , n29839 );
xor ( n35769 , n35768 , n32031 );
xor ( n35770 , n32127 , n28367 );
xor ( n35771 , n35770 , n29952 );
not ( n35772 , n35771 );
and ( n35773 , n35772 , n33340 );
xor ( n35774 , n35769 , n35773 );
xor ( n35775 , n29299 , n31487 );
xor ( n35776 , n35775 , n31497 );
xor ( n35777 , n31177 , n29532 );
xor ( n35778 , n35777 , n29544 );
not ( n35779 , n35778 );
and ( n35780 , n35779 , n33349 );
xor ( n35781 , n35776 , n35780 );
xor ( n35782 , n35774 , n35781 );
xor ( n35783 , n29431 , n27712 );
xor ( n35784 , n35783 , n30030 );
not ( n35785 , n35764 );
and ( n35786 , n35785 , n33359 );
xor ( n35787 , n35784 , n35786 );
xor ( n35788 , n35782 , n35787 );
xor ( n35789 , n30882 , n32734 );
xor ( n35790 , n35789 , n32744 );
xor ( n35791 , n28231 , n31581 );
xor ( n35792 , n35791 , n28947 );
not ( n35793 , n35792 );
and ( n35794 , n35793 , n33369 );
xor ( n35795 , n35790 , n35794 );
xor ( n35796 , n35788 , n35795 );
xor ( n35797 , n29284 , n30017 );
xor ( n35798 , n35797 , n30986 );
xor ( n35799 , n30327 , n33234 );
xor ( n35800 , n35799 , n31825 );
not ( n35801 , n35800 );
and ( n35802 , n35801 , n33380 );
xor ( n35803 , n35798 , n35802 );
xor ( n35804 , n35796 , n35803 );
xor ( n35805 , n35767 , n35804 );
xor ( n35806 , n28415 , n31247 );
xor ( n35807 , n35806 , n27885 );
xor ( n35808 , n31075 , n32199 );
xor ( n35809 , n35808 , n28380 );
not ( n35810 , n35809 );
and ( n35811 , n35810 , n35667 );
xor ( n35812 , n35807 , n35811 );
xor ( n35813 , n32834 , n32510 );
xor ( n35814 , n35813 , n29462 );
not ( n35815 , n35814 );
and ( n35816 , n35815 , n35676 );
xor ( n35817 , n35663 , n35816 );
xor ( n35818 , n35812 , n35817 );
xor ( n35819 , n28221 , n30457 );
xor ( n35820 , n35819 , n31581 );
xor ( n35821 , n30177 , n31162 );
xor ( n35822 , n35821 , n29923 );
not ( n35823 , n35822 );
and ( n35824 , n35823 , n35682 );
xor ( n35825 , n35820 , n35824 );
xor ( n35826 , n35818 , n35825 );
xor ( n35827 , n29907 , n32091 );
xor ( n35828 , n35827 , n30139 );
xor ( n35829 , n29518 , n30655 );
xor ( n35830 , n35829 , n30665 );
not ( n35831 , n35830 );
and ( n35832 , n35831 , n35692 );
xor ( n35833 , n35828 , n35832 );
xor ( n35834 , n35826 , n35833 );
xor ( n35835 , n30953 , n28355 );
xor ( n35836 , n35835 , n28367 );
xor ( n35837 , n28068 , n31180 );
xor ( n35838 , n35837 , n31192 );
not ( n35839 , n35838 );
and ( n35840 , n35839 , n35702 );
xor ( n35841 , n35836 , n35840 );
xor ( n35842 , n35834 , n35841 );
xor ( n35843 , n35805 , n35842 );
and ( n35844 , n35762 , n35843 );
xor ( n35845 , n35656 , n35844 );
not ( n11906 , n29614 );
and ( n11907 , n11906 , RI17469078_1224);
and ( n11908 , n35845 , n29614 );
or ( n35846 , n11907 , n11908 );
not ( n11909 , RI1754c610_2);
and ( n11910 , n11909 , n35846 );
and ( n11911 , C0 , RI1754c610_2);
or ( n35847 , n11910 , n11911 );
buf ( n35848 , n35847 );
not ( n35849 , n30829 );
xor ( n35850 , n33664 , n31367 );
xor ( n35851 , n35850 , n28800 );
and ( n35852 , n35849 , n35851 );
xor ( n35853 , n30826 , n35852 );
xor ( n35854 , n35853 , n30923 );
xor ( n35855 , n35854 , n31053 );
not ( n35856 , n31622 );
and ( n35857 , n35856 , n31726 );
xor ( n35858 , n35855 , n35857 );
not ( n11912 , n29614 );
and ( n11913 , n11912 , RI17392308_2043);
and ( n11914 , n35858 , n29614 );
or ( n35859 , n11913 , n11914 );
not ( n11915 , RI1754c610_2);
and ( n11916 , n11915 , n35859 );
and ( n11917 , C0 , RI1754c610_2);
or ( n35860 , n11916 , n11917 );
buf ( n35861 , n35860 );
xor ( n35862 , n28936 , n34517 );
xor ( n35863 , n30303 , n28055 );
xor ( n35864 , n35863 , n28224 );
xor ( n35865 , n30217 , n29573 );
xor ( n35866 , n35865 , n30758 );
not ( n35867 , n35866 );
xor ( n35868 , n28241 , n29259 );
xor ( n35869 , n35868 , n29270 );
and ( n35870 , n35867 , n35869 );
xor ( n35871 , n35864 , n35870 );
xor ( n35872 , n30534 , n29752 );
xor ( n35873 , n35872 , n27833 );
xor ( n35874 , n30933 , n27752 );
xor ( n35875 , n35874 , n27764 );
not ( n35876 , n35875 );
xor ( n35877 , n32190 , n29793 );
xor ( n35878 , n35877 , n31909 );
and ( n35879 , n35876 , n35878 );
xor ( n35880 , n35873 , n35879 );
xor ( n35881 , n35871 , n35880 );
xor ( n35882 , n32807 , n31422 );
xor ( n35883 , n35882 , n29011 );
xor ( n35884 , n29247 , n27700 );
xor ( n35885 , n35884 , n27712 );
not ( n35886 , n35885 );
xor ( n35887 , n29262 , n29093 );
xor ( n35888 , n35887 , n29105 );
and ( n35889 , n35886 , n35888 );
xor ( n35890 , n35883 , n35889 );
xor ( n35891 , n35881 , n35890 );
xor ( n35892 , n30397 , n27807 );
xor ( n35893 , n35892 , n27819 );
xor ( n35894 , n29826 , n32130 );
xor ( n35895 , n35894 , n32140 );
not ( n35896 , n35895 );
xor ( n35897 , n28620 , n28327 );
xor ( n35898 , n35897 , n28339 );
and ( n35899 , n35896 , n35898 );
xor ( n35900 , n35893 , n35899 );
xor ( n35901 , n35891 , n35900 );
xor ( n35902 , n29173 , n28185 );
xor ( n35903 , n35902 , n28827 );
xor ( n35904 , n28504 , n30043 );
xor ( n35905 , n35904 , n30053 );
not ( n35906 , n35905 );
xor ( n35907 , n29631 , n28148 );
xor ( n35908 , n35907 , n28160 );
and ( n35909 , n35906 , n35908 );
xor ( n35910 , n35903 , n35909 );
xor ( n35911 , n35901 , n35910 );
xor ( n35912 , n35862 , n35911 );
not ( n35913 , n27898 );
and ( n35914 , n35913 , n27922 );
xor ( n35915 , n29893 , n35914 );
xor ( n35916 , n35915 , n29981 );
xor ( n35917 , n29305 , n31487 );
xor ( n35918 , n35917 , n31497 );
xor ( n35919 , n27900 , n29235 );
xor ( n35920 , n35919 , n30294 );
not ( n35921 , n35920 );
and ( n35922 , n35921 , n28138 );
xor ( n35923 , n35918 , n35922 );
xor ( n35924 , n33389 , n28069 );
xor ( n35925 , n35924 , n28081 );
xor ( n35926 , n30849 , n30114 );
xor ( n35927 , n35926 , n30125 );
not ( n35928 , n35927 );
and ( n35929 , n35928 , n28213 );
xor ( n35930 , n35925 , n35929 );
xor ( n35931 , n35923 , n35930 );
xor ( n35932 , n29398 , n32209 );
xor ( n35933 , n35932 , n30389 );
xor ( n35934 , n30286 , n28043 );
xor ( n35935 , n35934 , n28055 );
not ( n35936 , n35935 );
and ( n35937 , n35936 , n28292 );
xor ( n35938 , n35933 , n35937 );
xor ( n35939 , n35931 , n35938 );
xor ( n35940 , n32365 , n32835 );
xor ( n35941 , n35940 , n31399 );
xor ( n35942 , n29669 , n30842 );
xor ( n35943 , n35942 , n32247 );
not ( n35944 , n35943 );
and ( n35945 , n35944 , n28368 );
xor ( n35946 , n35941 , n35945 );
xor ( n35947 , n35939 , n35946 );
xor ( n35948 , n29693 , n30972 );
xor ( n35949 , n35948 , n29123 );
xor ( n35950 , n31183 , n29544 );
xor ( n35951 , n35950 , n28480 );
not ( n35952 , n35951 );
and ( n35953 , n35952 , n28426 );
xor ( n35954 , n35949 , n35953 );
xor ( n35955 , n35947 , n35954 );
xor ( n35956 , n35916 , n35955 );
not ( n35957 , n35956 );
xor ( n35958 , n30454 , n29123 );
xor ( n35959 , n35958 , n29134 );
not ( n35960 , n32148 );
and ( n35961 , n35960 , n32150 );
xor ( n35962 , n35959 , n35961 );
xor ( n35963 , n31680 , n28001 );
xor ( n35964 , n35963 , n30114 );
not ( n35965 , n32157 );
and ( n35966 , n35965 , n32168 );
xor ( n35967 , n35964 , n35966 );
xor ( n35968 , n35962 , n35967 );
xor ( n35969 , n29811 , n31516 );
xor ( n35970 , n35969 , n31528 );
not ( n35971 , n32176 );
and ( n35972 , n35971 , n32178 );
xor ( n35973 , n35970 , n35972 );
xor ( n35974 , n35968 , n35973 );
xor ( n35975 , n33387 , n28069 );
xor ( n35976 , n35975 , n28081 );
not ( n35977 , n32188 );
and ( n35978 , n35977 , n32201 );
xor ( n35979 , n35976 , n35978 );
xor ( n35980 , n35974 , n35979 );
xor ( n35981 , n28554 , n30616 );
xor ( n35982 , n35981 , n30626 );
not ( n35983 , n32216 );
and ( n35984 , n35983 , n32121 );
xor ( n35985 , n35982 , n35984 );
xor ( n35986 , n35980 , n35985 );
xor ( n35987 , n32213 , n35986 );
not ( n35988 , n32233 );
and ( n35989 , n35988 , n32235 );
xor ( n35990 , n32625 , n35989 );
xor ( n35991 , n35422 , n35990 );
not ( n35992 , n32262 );
and ( n35993 , n35992 , n32264 );
xor ( n35994 , n32644 , n35993 );
xor ( n35995 , n35991 , n35994 );
not ( n35996 , n32281 );
and ( n35997 , n35996 , n32293 );
xor ( n35998 , n32652 , n35997 );
xor ( n35999 , n35995 , n35998 );
not ( n36000 , n32301 );
and ( n36001 , n36000 , n32303 );
xor ( n36002 , n32660 , n36001 );
xor ( n36003 , n35999 , n36002 );
xor ( n36004 , n35987 , n36003 );
and ( n36005 , n35957 , n36004 );
xor ( n36006 , n35912 , n36005 );
not ( n11918 , n29614 );
and ( n11919 , n11918 , RI17397ba0_2016);
and ( n11920 , n36006 , n29614 );
or ( n36007 , n11919 , n11920 );
not ( n11921 , RI1754c610_2);
and ( n11922 , n11921 , n36007 );
and ( n11923 , C0 , RI1754c610_2);
or ( n36008 , n11922 , n11923 );
buf ( n36009 , n36008 );
buf ( n36010 , RI17515908_699);
buf ( n36011 , RI174ba900_830);
not ( n11924 , n27683 );
and ( n11925 , n11924 , RI19a82538_2778);
and ( n11926 , RI19aaa858_2492 , n27683 );
or ( n36012 , n11925 , n11926 );
not ( n11927 , RI1754c610_2);
and ( n11928 , n11927 , n36012 );
and ( n11929 , C0 , RI1754c610_2);
or ( n36013 , n11928 , n11929 );
buf ( n36014 , n36013 );
not ( n11930 , n27683 );
and ( n11931 , n11930 , RI19accea8_2232);
and ( n11932 , RI19a88e38_2732 , n27683 );
or ( n36015 , n11931 , n11932 );
not ( n11933 , RI1754c610_2);
and ( n11934 , n11933 , n36015 );
and ( n11935 , C0 , RI1754c610_2);
or ( n36016 , n11934 , n11935 );
buf ( n36017 , n36016 );
not ( n36018 , n32546 );
xor ( n36019 , n32204 , n28800 );
xor ( n36020 , n36019 , n28812 );
and ( n36021 , n36018 , n36020 );
xor ( n36022 , n32543 , n36021 );
xor ( n36023 , n36022 , n32560 );
xor ( n36024 , n36023 , n32620 );
not ( n36025 , n32707 );
and ( n36026 , n36025 , n32709 );
xor ( n36027 , n32919 , n36026 );
xor ( n36028 , n36027 , n32923 );
xor ( n36029 , n36028 , n32973 );
not ( n36030 , n36029 );
xor ( n36031 , n29916 , n27791 );
xor ( n36032 , n36031 , n30706 );
not ( n36033 , n36032 );
and ( n36034 , n36033 , n33410 );
xor ( n36035 , n34454 , n36034 );
not ( n36036 , n34454 );
and ( n36037 , n36036 , n36032 );
xor ( n36038 , n33415 , n36037 );
not ( n36039 , n34459 );
xor ( n36040 , n29807 , n31516 );
xor ( n36041 , n36040 , n31528 );
and ( n36042 , n36039 , n36041 );
xor ( n36043 , n33424 , n36042 );
xor ( n36044 , n36038 , n36043 );
not ( n36045 , n34465 );
xor ( n36046 , n32376 , n29490 );
xor ( n36047 , n36046 , n29502 );
and ( n36048 , n36045 , n36047 );
xor ( n36049 , n33434 , n36048 );
xor ( n36050 , n36044 , n36049 );
not ( n36051 , n34471 );
xor ( n36052 , n30437 , n28956 );
xor ( n36053 , n36052 , n29995 );
and ( n36054 , n36051 , n36053 );
xor ( n36055 , n33444 , n36054 );
xor ( n36056 , n36050 , n36055 );
not ( n36057 , n33406 );
xor ( n36058 , n29734 , n28304 );
xor ( n36059 , n36058 , n28313 );
and ( n36060 , n36057 , n36059 );
xor ( n36061 , n33403 , n36060 );
xor ( n36062 , n36056 , n36061 );
xor ( n36063 , n36035 , n36062 );
xor ( n36064 , n30185 , n29923 );
xor ( n36065 , n36064 , n29935 );
not ( n36066 , n36065 );
xor ( n36067 , n32363 , n32835 );
xor ( n36068 , n36067 , n31399 );
and ( n36069 , n36066 , n36068 );
xor ( n36070 , n33463 , n36069 );
xor ( n36071 , n29834 , n32140 );
xor ( n36072 , n36071 , n31874 );
not ( n36073 , n36072 );
xor ( n36074 , n28724 , n31279 );
xor ( n36075 , n36074 , n33665 );
and ( n36076 , n36073 , n36075 );
xor ( n36077 , n33472 , n36076 );
xor ( n36078 , n36070 , n36077 );
xor ( n36079 , n29032 , n30399 );
xor ( n36080 , n36079 , n29532 );
not ( n36081 , n36080 );
xor ( n36082 , n28530 , n27764 );
xor ( n36083 , n36082 , n28125 );
and ( n36084 , n36081 , n36083 );
xor ( n36085 , n33482 , n36084 );
xor ( n36086 , n36078 , n36085 );
xor ( n36087 , n30240 , n28250 );
xor ( n36088 , n36087 , n28262 );
not ( n36089 , n36088 );
xor ( n36090 , n30280 , n31309 );
xor ( n36091 , n36090 , n29519 );
and ( n36092 , n36089 , n36091 );
xor ( n36093 , n33492 , n36092 );
xor ( n36094 , n36086 , n36093 );
xor ( n36095 , n31904 , n30101 );
xor ( n36096 , n36095 , n32426 );
not ( n36097 , n36096 );
xor ( n36098 , n30148 , n30918 );
xor ( n36099 , n36098 , n31594 );
and ( n36100 , n36097 , n36099 );
xor ( n36101 , n33502 , n36100 );
xor ( n36102 , n36094 , n36101 );
xor ( n36103 , n36063 , n36102 );
and ( n36104 , n36030 , n36103 );
xor ( n36105 , n36024 , n36104 );
not ( n11936 , n29614 );
and ( n11937 , n11936 , RI17499048_990);
and ( n11938 , n36105 , n29614 );
or ( n36106 , n11937 , n11938 );
not ( n11939 , RI1754c610_2);
and ( n11940 , n11939 , n36106 );
and ( n11941 , C0 , RI1754c610_2);
or ( n36107 , n11940 , n11941 );
buf ( n36108 , n36107 );
buf ( n36109 , RI174aec18_884);
not ( n36110 , n27765 );
and ( n36111 , n36110 , n29857 );
xor ( n36112 , n27739 , n36111 );
not ( n36113 , n29874 );
and ( n36114 , n36113 , n29876 );
xor ( n36115 , n27871 , n36114 );
xor ( n36116 , n36112 , n36115 );
not ( n36117 , n29890 );
and ( n36118 , n36117 , n29893 );
xor ( n36119 , n27949 , n36118 );
xor ( n36120 , n36116 , n36119 );
not ( n36121 , n29911 );
and ( n36122 , n36121 , n29936 );
xor ( n36123 , n28028 , n36122 );
xor ( n36124 , n36120 , n36123 );
not ( n36125 , n29965 );
and ( n36126 , n36125 , n29977 );
xor ( n36127 , n28108 , n36126 );
xor ( n36128 , n36124 , n36127 );
xor ( n36129 , n29980 , n36128 );
not ( n36130 , n35918 );
and ( n36131 , n36130 , n35920 );
xor ( n36132 , n28186 , n36131 );
not ( n36133 , n35925 );
and ( n36134 , n36133 , n35927 );
xor ( n36135 , n28263 , n36134 );
xor ( n36136 , n36132 , n36135 );
not ( n36137 , n35933 );
and ( n36138 , n36137 , n35935 );
xor ( n36139 , n28340 , n36138 );
xor ( n36140 , n36136 , n36139 );
not ( n36141 , n35941 );
and ( n36142 , n36141 , n35943 );
xor ( n36143 , n28419 , n36142 );
xor ( n36144 , n36140 , n36143 );
not ( n36145 , n35949 );
and ( n36146 , n36145 , n35951 );
xor ( n36147 , n28465 , n36146 );
xor ( n36148 , n36144 , n36147 );
xor ( n36149 , n36129 , n36148 );
not ( n36150 , n32411 );
and ( n36151 , n36150 , n32745 );
xor ( n36152 , n32408 , n36151 );
xor ( n36153 , n36152 , n32481 );
xor ( n36154 , n36153 , n33030 );
not ( n36155 , n36154 );
not ( n36156 , n31650 );
and ( n36157 , n36156 , n35476 );
xor ( n36158 , n30553 , n36157 );
xor ( n36159 , n36158 , n31664 );
xor ( n36160 , n36159 , n31725 );
and ( n36161 , n36155 , n36160 );
xor ( n36162 , n36149 , n36161 );
not ( n11942 , n29614 );
and ( n11943 , n11942 , RI17535780_600);
and ( n11944 , n36162 , n29614 );
or ( n36163 , n11943 , n11944 );
not ( n11945 , RI1754c610_2);
and ( n11946 , n11945 , n36163 );
and ( n11947 , C0 , RI1754c610_2);
or ( n36164 , n11946 , n11947 );
buf ( n36165 , n36164 );
not ( n11948 , n27683 );
and ( n11949 , n11948 , RI19a894c8_2729);
and ( n11950 , RI19a936f8_2658 , n27683 );
or ( n36166 , n11949 , n11950 );
not ( n11951 , RI1754c610_2);
and ( n11952 , n11951 , n36166 );
and ( n11953 , C0 , RI1754c610_2);
or ( n36167 , n11952 , n11953 );
buf ( n36168 , n36167 );
buf ( n36169 , RI174a44c0_935);
buf ( n36170 , RI1747fcb0_1113);
buf ( n36171 , RI1747e5b8_1120);
buf ( n36172 , RI17473488_1174);
buf ( n36173 , RI1746cb88_1206);
not ( n11954 , n27683 );
and ( n11955 , n11954 , RI19a8bbb0_2713);
and ( n11956 , RI19a95b88_2642 , n27683 );
or ( n36174 , n11955 , n11956 );
not ( n11957 , RI1754c610_2);
and ( n11958 , n11957 , n36174 );
and ( n11959 , C0 , RI1754c610_2);
or ( n36175 , n11958 , n11959 );
buf ( n36176 , n36175 );
not ( n36177 , n32229 );
and ( n36178 , n36177 , n32630 );
xor ( n36179 , n32225 , n36178 );
not ( n36180 , n32257 );
and ( n36181 , n36180 , n32623 );
xor ( n36182 , n32235 , n36181 );
xor ( n36183 , n36179 , n36182 );
not ( n36184 , n32276 );
and ( n36185 , n36184 , n32641 );
xor ( n36186 , n32264 , n36185 );
xor ( n36187 , n36183 , n36186 );
not ( n36188 , n32296 );
and ( n36189 , n36188 , n32649 );
xor ( n36190 , n32293 , n36189 );
xor ( n36191 , n36187 , n36190 );
not ( n36192 , n32306 );
and ( n36193 , n36192 , n32657 );
xor ( n36194 , n32303 , n36193 );
xor ( n36195 , n36191 , n36194 );
xor ( n36196 , n32638 , n36195 );
not ( n36197 , n32666 );
and ( n36198 , n36197 , n32670 );
xor ( n36199 , n32882 , n36198 );
xor ( n36200 , n36199 , n32878 );
not ( n36201 , n32687 );
and ( n36202 , n36201 , n32689 );
xor ( n36203 , n32903 , n36202 );
xor ( n36204 , n36200 , n36203 );
not ( n36205 , n32697 );
and ( n36206 , n36205 , n32699 );
xor ( n36207 , n32911 , n36206 );
xor ( n36208 , n36204 , n36207 );
xor ( n36209 , n36208 , n36027 );
xor ( n36210 , n36196 , n36209 );
xor ( n36211 , n33013 , n35639 );
not ( n36212 , n31769 );
and ( n36213 , n36212 , n33033 );
xor ( n36214 , n31764 , n36213 );
not ( n36215 , n31779 );
and ( n36216 , n36215 , n33041 );
xor ( n36217 , n31776 , n36216 );
xor ( n36218 , n36214 , n36217 );
not ( n36219 , n31802 );
and ( n36220 , n36219 , n33049 );
xor ( n36221 , n31797 , n36220 );
xor ( n36222 , n36218 , n36221 );
not ( n36223 , n31812 );
and ( n36224 , n36223 , n33057 );
xor ( n36225 , n31809 , n36224 );
xor ( n36226 , n36222 , n36225 );
xor ( n36227 , n36226 , n31739 );
xor ( n36228 , n36211 , n36227 );
not ( n36229 , n36228 );
not ( n36230 , n31886 );
and ( n36231 , n36230 , n31888 );
xor ( n36232 , n34178 , n36231 );
xor ( n36233 , n36232 , n34190 );
not ( n36234 , n33410 );
and ( n36235 , n36234 , n33412 );
xor ( n36236 , n36032 , n36235 );
not ( n36237 , n33419 );
and ( n36238 , n36237 , n33421 );
xor ( n36239 , n36041 , n36238 );
xor ( n36240 , n36236 , n36239 );
not ( n36241 , n33429 );
and ( n36242 , n36241 , n33431 );
xor ( n36243 , n36047 , n36242 );
xor ( n36244 , n36240 , n36243 );
not ( n36245 , n33439 );
and ( n36246 , n36245 , n33441 );
xor ( n36247 , n36053 , n36246 );
xor ( n36248 , n36244 , n36247 );
not ( n36249 , n33449 );
and ( n36250 , n36249 , n33401 );
xor ( n36251 , n36059 , n36250 );
xor ( n36252 , n36248 , n36251 );
xor ( n36253 , n36233 , n36252 );
and ( n36254 , n36229 , n36253 );
xor ( n36255 , n36210 , n36254 );
not ( n11960 , n29614 );
and ( n11961 , n11960 , RI1744dc10_1357);
and ( n11962 , n36255 , n29614 );
or ( n36256 , n11961 , n11962 );
not ( n11963 , RI1754c610_2);
and ( n11964 , n11963 , n36256 );
and ( n11965 , C0 , RI1754c610_2);
or ( n36257 , n11964 , n11965 );
buf ( n36258 , n36257 );
not ( n36259 , n33902 );
and ( n36260 , n36259 , n34097 );
xor ( n36261 , n33899 , n36260 );
xor ( n36262 , n36261 , n33935 );
not ( n36263 , n34194 );
and ( n36264 , n36263 , n33948 );
xor ( n36265 , n35652 , n36264 );
xor ( n36266 , n29394 , n32209 );
xor ( n36267 , n36266 , n30389 );
not ( n36268 , n34199 );
and ( n36269 , n36268 , n33957 );
xor ( n36270 , n36267 , n36269 );
xor ( n36271 , n36265 , n36270 );
xor ( n36272 , n30808 , n32382 );
xor ( n36273 , n36272 , n28463 );
not ( n36274 , n34205 );
and ( n36275 , n36274 , n33967 );
xor ( n36276 , n36273 , n36275 );
xor ( n36277 , n36271 , n36276 );
not ( n36278 , n34211 );
and ( n36279 , n36278 , n33977 );
xor ( n36280 , n33944 , n36279 );
xor ( n36281 , n36277 , n36280 );
xor ( n36282 , n29809 , n31516 );
xor ( n36283 , n36282 , n31528 );
not ( n36284 , n34217 );
and ( n36285 , n36284 , n33983 );
xor ( n36286 , n36283 , n36285 );
xor ( n36287 , n36281 , n36286 );
xor ( n36288 , n36262 , n36287 );
not ( n36289 , n33856 );
and ( n36290 , n36289 , n33828 );
xor ( n36291 , n34067 , n36290 );
xor ( n36292 , n36291 , n34087 );
xor ( n36293 , n36292 , n34127 );
not ( n36294 , n36293 );
and ( n36295 , n36294 , n36024 );
xor ( n36296 , n36288 , n36295 );
not ( n11966 , n29614 );
and ( n11967 , n11966 , RI1747be58_1132);
and ( n11968 , n36296 , n29614 );
or ( n36297 , n11967 , n11968 );
not ( n11969 , RI1754c610_2);
and ( n11970 , n11969 , n36297 );
and ( n11971 , C0 , RI1754c610_2);
or ( n36298 , n11970 , n11971 );
buf ( n36299 , n36298 );
xor ( n36300 , n29206 , n32459 );
xor ( n36301 , n36300 , n30616 );
not ( n36302 , n35392 );
and ( n36303 , n36302 , n35394 );
xor ( n36304 , n36301 , n36303 );
xor ( n36305 , n28752 , n30823 );
xor ( n36306 , n36305 , n30934 );
xor ( n36307 , n32378 , n29490 );
xor ( n36308 , n36307 , n29502 );
not ( n36309 , n36308 );
and ( n36310 , n36309 , n35373 );
xor ( n36311 , n36306 , n36310 );
xor ( n36312 , n27878 , n29387 );
xor ( n36313 , n36312 , n29399 );
xor ( n36314 , n27904 , n29235 );
xor ( n36315 , n36314 , n30294 );
not ( n36316 , n36315 );
and ( n36317 , n36316 , n35382 );
xor ( n36318 , n36313 , n36317 );
xor ( n36319 , n36311 , n36318 );
xor ( n36320 , n29116 , n29873 );
xor ( n36321 , n36320 , n32398 );
not ( n36322 , n36301 );
and ( n36323 , n36322 , n35392 );
xor ( n36324 , n36321 , n36323 );
xor ( n36325 , n36319 , n36324 );
xor ( n36326 , n31707 , n30332 );
xor ( n36327 , n36326 , n32043 );
xor ( n36328 , n29990 , n28702 );
xor ( n36329 , n36328 , n31065 );
not ( n36330 , n36329 );
and ( n36331 , n36330 , n35402 );
xor ( n36332 , n36327 , n36331 );
xor ( n36333 , n36325 , n36332 );
xor ( n36334 , n28350 , n30510 );
xor ( n36335 , n36334 , n30522 );
not ( n36336 , n36335 );
and ( n36337 , n36336 , n35412 );
xor ( n36338 , n35369 , n36337 );
xor ( n36339 , n36333 , n36338 );
xor ( n36340 , n36304 , n36339 );
xor ( n36341 , n30917 , n30348 );
xor ( n36342 , n36341 , n30178 );
not ( n36343 , n36342 );
and ( n36344 , n36343 , n29663 );
xor ( n36345 , n29657 , n36344 );
xor ( n36346 , n28145 , n27726 );
xor ( n36347 , n36346 , n27738 );
xor ( n36348 , n32610 , n29025 );
xor ( n36349 , n36348 , n29037 );
not ( n36350 , n36349 );
and ( n36351 , n36350 , n29678 );
xor ( n36352 , n36347 , n36351 );
xor ( n36353 , n36345 , n36352 );
xor ( n36354 , n28953 , n27948 );
xor ( n36355 , n36354 , n28702 );
xor ( n36356 , n31278 , n30717 );
xor ( n36357 , n36356 , n31367 );
not ( n36358 , n36357 );
and ( n36359 , n36358 , n29700 );
xor ( n36360 , n36355 , n36359 );
xor ( n36361 , n36353 , n36360 );
xor ( n36362 , n31021 , n31594 );
xor ( n36363 , n36362 , n31487 );
xor ( n36364 , n31515 , n28096 );
xor ( n36365 , n36364 , n28107 );
not ( n36366 , n36365 );
and ( n36367 , n36366 , n29753 );
xor ( n36368 , n36363 , n36367 );
xor ( n36369 , n36361 , n36368 );
xor ( n36370 , n29961 , n30164 );
xor ( n36371 , n36370 , n29490 );
xor ( n36372 , n27711 , n27909 );
xor ( n36373 , n36372 , n27921 );
not ( n36374 , n36373 );
and ( n36375 , n36374 , n29801 );
xor ( n36376 , n36371 , n36375 );
xor ( n36377 , n36369 , n36376 );
xor ( n36378 , n36340 , n36377 );
not ( n36379 , n31476 );
and ( n36380 , n36379 , n34286 );
xor ( n36381 , n31463 , n36380 );
xor ( n36382 , n36381 , n31506 );
xor ( n36383 , n36382 , n31621 );
not ( n36384 , n36383 );
xor ( n36385 , n31830 , n34644 );
not ( n36386 , n31834 );
and ( n36387 , n36386 , n31845 );
xor ( n36388 , n34155 , n36387 );
not ( n36389 , n31853 );
and ( n36390 , n36389 , n31855 );
xor ( n36391 , n34162 , n36390 );
xor ( n36392 , n36388 , n36391 );
not ( n36393 , n31876 );
and ( n36394 , n36393 , n31878 );
xor ( n36395 , n34170 , n36394 );
xor ( n36396 , n36392 , n36395 );
xor ( n36397 , n36396 , n36232 );
not ( n36398 , n31896 );
and ( n36399 , n36398 , n31898 );
xor ( n36400 , n34186 , n36399 );
xor ( n36401 , n36397 , n36400 );
xor ( n36402 , n36385 , n36401 );
and ( n36403 , n36384 , n36402 );
xor ( n36404 , n36378 , n36403 );
not ( n11972 , n29614 );
and ( n11973 , n11972 , RI17486c40_1079);
and ( n11974 , n36404 , n29614 );
or ( n36405 , n11973 , n11974 );
not ( n11975 , RI1754c610_2);
and ( n11976 , n11975 , n36405 );
and ( n11977 , C0 , RI1754c610_2);
or ( n36406 , n11976 , n11977 );
buf ( n36407 , n36406 );
not ( n36408 , n29794 );
and ( n36409 , n36408 , n36363 );
xor ( n36410 , n29768 , n36409 );
xor ( n36411 , n36410 , n29843 );
xor ( n36412 , n36411 , n29981 );
not ( n36413 , n34121 );
and ( n36414 , n36413 , n34123 );
xor ( n36415 , n33932 , n36414 );
not ( n36416 , n33888 );
and ( n36417 , n36416 , n34090 );
xor ( n36418 , n33885 , n36417 );
xor ( n36419 , n36418 , n36261 );
not ( n36420 , n33912 );
and ( n36421 , n36420 , n34105 );
xor ( n36422 , n33909 , n36421 );
xor ( n36423 , n36419 , n36422 );
not ( n36424 , n33922 );
and ( n36425 , n36424 , n34113 );
xor ( n36426 , n33919 , n36425 );
xor ( n36427 , n36423 , n36426 );
not ( n36428 , n33932 );
and ( n36429 , n36428 , n34121 );
xor ( n36430 , n33929 , n36429 );
xor ( n36431 , n36427 , n36430 );
xor ( n36432 , n36415 , n36431 );
xor ( n36433 , n36432 , n34221 );
not ( n36434 , n36433 );
xor ( n36435 , n28564 , n30626 );
xor ( n36436 , n36435 , n29740 );
not ( n36437 , n35864 );
and ( n36438 , n36437 , n35866 );
xor ( n36439 , n36436 , n36438 );
xor ( n36440 , n30002 , n30567 );
xor ( n36441 , n36440 , n28647 );
not ( n36442 , n35873 );
and ( n36443 , n36442 , n35875 );
xor ( n36444 , n36441 , n36443 );
xor ( n36445 , n36439 , n36444 );
xor ( n36446 , n27943 , n30374 );
xor ( n36447 , n36446 , n32472 );
not ( n36448 , n35883 );
and ( n36449 , n36448 , n35885 );
xor ( n36450 , n36447 , n36449 );
xor ( n36451 , n36445 , n36450 );
xor ( n36452 , n31126 , n31528 );
xor ( n36453 , n36452 , n32835 );
not ( n36454 , n35893 );
and ( n36455 , n36454 , n35895 );
xor ( n36456 , n36453 , n36455 );
xor ( n36457 , n36451 , n36456 );
xor ( n36458 , n29596 , n28200 );
xor ( n36459 , n36458 , n28212 );
not ( n36460 , n35903 );
and ( n36461 , n36460 , n35905 );
xor ( n36462 , n36459 , n36461 );
xor ( n36463 , n36457 , n36462 );
xor ( n36464 , n35871 , n36463 );
xor ( n36465 , n36464 , n32220 );
and ( n36466 , n36434 , n36465 );
xor ( n36467 , n36412 , n36466 );
not ( n11978 , n29614 );
and ( n11979 , n11978 , RI17524110_654);
and ( n11980 , n36467 , n29614 );
or ( n36468 , n11979 , n11980 );
not ( n11981 , RI1754c610_2);
and ( n11982 , n11981 , n36468 );
and ( n11983 , C0 , RI1754c610_2);
or ( n36469 , n11982 , n11983 );
buf ( n36470 , n36469 );
not ( n11984 , n27683 );
and ( n11985 , n11984 , RI19acc200_2238);
and ( n11986 , RI19a87dd0_2739 , n27683 );
or ( n36471 , n11985 , n11986 );
not ( n11987 , RI1754c610_2);
and ( n11988 , n11987 , n36471 );
and ( n11989 , C0 , RI1754c610_2);
or ( n36472 , n11988 , n11989 );
buf ( n36473 , n36472 );
not ( n11990 , n27683 );
and ( n11991 , n11990 , RI19aa8878_2506);
and ( n11992 , RI19ab29b8_2435 , n27683 );
or ( n36474 , n11991 , n11992 );
not ( n11993 , RI1754c610_2);
and ( n11994 , n11993 , n36474 );
and ( n11995 , C0 , RI1754c610_2);
or ( n36475 , n11994 , n11995 );
buf ( n36476 , n36475 );
xor ( n36477 , n28714 , n29935 );
xor ( n36478 , n36477 , n31279 );
xor ( n36479 , n28034 , n29449 );
xor ( n36480 , n36479 , n29694 );
not ( n36481 , n36480 );
xor ( n36482 , n30238 , n28250 );
xor ( n36483 , n36482 , n28262 );
and ( n36484 , n36481 , n36483 );
xor ( n36485 , n36478 , n36484 );
xor ( n36486 , n29208 , n32459 );
xor ( n36487 , n36486 , n30616 );
not ( n36488 , n36478 );
and ( n36489 , n36488 , n36480 );
xor ( n36490 , n36487 , n36489 );
xor ( n36491 , n29268 , n29093 );
xor ( n36492 , n36491 , n29105 );
xor ( n36493 , n31191 , n29544 );
xor ( n36494 , n36493 , n28480 );
not ( n36495 , n36494 );
xor ( n36496 , n30992 , n32256 );
xor ( n36497 , n36496 , n32734 );
and ( n36498 , n36495 , n36497 );
xor ( n36499 , n36492 , n36498 );
xor ( n36500 , n36490 , n36499 );
xor ( n36501 , n31073 , n32199 );
xor ( n36502 , n36501 , n28380 );
xor ( n36503 , n28811 , n29409 );
xor ( n36504 , n36503 , n29421 );
not ( n36505 , n36504 );
xor ( n36506 , n29685 , n30972 );
xor ( n36507 , n36506 , n29123 );
and ( n36508 , n36505 , n36507 );
xor ( n36509 , n36502 , n36508 );
xor ( n36510 , n36500 , n36509 );
xor ( n36511 , n31244 , n28727 );
xor ( n36512 , n36511 , n29387 );
xor ( n36513 , n29461 , n31950 );
xor ( n36514 , n36513 , n31558 );
not ( n36515 , n36514 );
xor ( n36516 , n27836 , n30857 );
xor ( n36517 , n36516 , n30869 );
and ( n36518 , n36515 , n36517 );
xor ( n36519 , n36512 , n36518 );
xor ( n36520 , n36510 , n36519 );
xor ( n36521 , n29625 , n30799 );
xor ( n36522 , n36521 , n28148 );
xor ( n36523 , n29872 , n30548 );
xor ( n36524 , n36523 , n28673 );
not ( n36525 , n36524 );
xor ( n36526 , n29215 , n28995 );
xor ( n36527 , n36526 , n30780 );
and ( n36528 , n36525 , n36527 );
xor ( n36529 , n36522 , n36528 );
xor ( n36530 , n36520 , n36529 );
xor ( n36531 , n36485 , n36530 );
not ( n36532 , n34678 );
xor ( n36533 , n28132 , n30243 );
xor ( n36534 , n36533 , n31750 );
and ( n36535 , n36532 , n36534 );
xor ( n36536 , n34675 , n36535 );
xor ( n36537 , n28178 , n29211 );
xor ( n36538 , n36537 , n28557 );
not ( n36539 , n36538 );
xor ( n36540 , n30359 , n28684 );
xor ( n36541 , n36540 , n28279 );
and ( n36542 , n36539 , n36541 );
xor ( n36543 , n34692 , n36542 );
xor ( n36544 , n36536 , n36543 );
xor ( n36545 , n31058 , n32323 );
xor ( n36546 , n36545 , n32199 );
not ( n36547 , n36546 );
xor ( n36548 , n30837 , n27833 );
xor ( n36549 , n36548 , n27844 );
and ( n36550 , n36547 , n36549 );
xor ( n36551 , n34702 , n36550 );
xor ( n36552 , n36544 , n36551 );
xor ( n36553 , n29832 , n32140 );
xor ( n36554 , n36553 , n31874 );
not ( n36555 , n36554 );
xor ( n36556 , n31838 , n30151 );
xor ( n36557 , n36556 , n31024 );
and ( n36558 , n36555 , n36557 );
xor ( n36559 , n34712 , n36558 );
xor ( n36560 , n36552 , n36559 );
xor ( n36561 , n29455 , n31950 );
xor ( n36562 , n36561 , n31558 );
not ( n36563 , n36562 );
xor ( n36564 , n28458 , n29502 );
xor ( n36565 , n36564 , n29628 );
and ( n36566 , n36563 , n36565 );
xor ( n36567 , n34722 , n36566 );
xor ( n36568 , n36560 , n36567 );
xor ( n36569 , n36531 , n36568 );
xor ( n36570 , n29943 , n32009 );
xor ( n36571 , n36570 , n30164 );
xor ( n36572 , n32729 , n30475 );
xor ( n36573 , n36572 , n30487 );
not ( n36574 , n36573 );
and ( n36575 , n36574 , n33137 );
xor ( n36576 , n36571 , n36575 );
xor ( n36577 , n28371 , n31909 );
xor ( n36578 , n36577 , n31921 );
not ( n36579 , n36578 );
xor ( n36580 , n31448 , n29011 );
xor ( n36581 , n36580 , n27964 );
and ( n36582 , n36579 , n36581 );
xor ( n36583 , n33133 , n36582 );
not ( n36584 , n36571 );
and ( n36585 , n36584 , n36573 );
xor ( n36586 , n33142 , n36585 );
xor ( n36587 , n36583 , n36586 );
xor ( n36588 , n31912 , n32426 );
xor ( n36589 , n36588 , n31152 );
not ( n36590 , n36589 );
xor ( n36591 , n31240 , n28727 );
xor ( n36592 , n36591 , n29387 );
and ( n36593 , n36590 , n36592 );
xor ( n36594 , n33152 , n36593 );
xor ( n36595 , n36587 , n36594 );
xor ( n36596 , n29054 , n29827 );
xor ( n36597 , n36596 , n29839 );
not ( n36598 , n36597 );
xor ( n36599 , n29087 , n28493 );
xor ( n36600 , n36599 , n28505 );
and ( n36601 , n36598 , n36600 );
xor ( n36602 , n33162 , n36601 );
xor ( n36603 , n36595 , n36602 );
xor ( n36604 , n31056 , n32323 );
xor ( n36605 , n36604 , n32199 );
not ( n36606 , n36605 );
xor ( n36607 , n30024 , n27921 );
xor ( n36608 , n36607 , n28852 );
and ( n36609 , n36606 , n36608 );
xor ( n36610 , n33172 , n36609 );
xor ( n36611 , n36603 , n36610 );
xor ( n36612 , n36576 , n36611 );
xor ( n36613 , n36612 , n33567 );
not ( n36614 , n36613 );
xor ( n36615 , n35449 , n32715 );
xor ( n36616 , n27945 , n30374 );
xor ( n36617 , n36616 , n32472 );
not ( n36618 , n36617 );
xor ( n36619 , n27699 , n28480 );
xor ( n36620 , n36619 , n27909 );
and ( n36621 , n36618 , n36620 );
xor ( n36622 , n32931 , n36621 );
xor ( n36623 , n31111 , n30889 );
xor ( n36624 , n36623 , n30901 );
not ( n36625 , n36624 );
xor ( n36626 , n28261 , n29270 );
xor ( n36627 , n36626 , n30066 );
and ( n36628 , n36625 , n36627 );
xor ( n36629 , n32940 , n36628 );
xor ( n36630 , n36622 , n36629 );
xor ( n36631 , n31397 , n29462 );
xor ( n36632 , n36631 , n29474 );
not ( n36633 , n36632 );
xor ( n36634 , n30547 , n28224 );
xor ( n36635 , n36634 , n28236 );
and ( n36636 , n36633 , n36635 );
xor ( n36637 , n32950 , n36636 );
xor ( n36638 , n36630 , n36637 );
xor ( n36639 , n29435 , n27712 );
xor ( n36640 , n36639 , n30030 );
not ( n36641 , n36640 );
xor ( n36642 , n29501 , n30789 );
xor ( n36643 , n36642 , n30799 );
and ( n36644 , n36641 , n36643 );
xor ( n36645 , n32960 , n36644 );
xor ( n36646 , n36638 , n36645 );
xor ( n36647 , n29749 , n28313 );
xor ( n36648 , n36647 , n31683 );
not ( n36649 , n36648 );
xor ( n36650 , n31793 , n29148 );
xor ( n36651 , n36650 , n32800 );
and ( n36652 , n36649 , n36651 );
xor ( n36653 , n32970 , n36652 );
xor ( n36654 , n36646 , n36653 );
xor ( n36655 , n36615 , n36654 );
and ( n36656 , n36614 , n36655 );
xor ( n36657 , n36569 , n36656 );
not ( n11996 , n29614 );
and ( n11997 , n11996 , RI173d1f98_1732);
and ( n11998 , n36657 , n29614 );
or ( n36658 , n11997 , n11998 );
not ( n11999 , RI1754c610_2);
and ( n12000 , n11999 , n36658 );
and ( n12001 , C0 , RI1754c610_2);
or ( n36659 , n12000 , n12001 );
buf ( n36660 , n36659 );
not ( n12002 , RI1754c610_2);
and ( n12003 , n12002 , RI19a25298_2780);
and ( n12004 , C0 , RI1754c610_2);
or ( n36661 , n12003 , n12004 );
buf ( n36662 , n36661 );
not ( n36663 , n35843 );
not ( n36664 , n31952 );
and ( n36665 , n36664 , n31954 );
xor ( n36666 , n35133 , n36665 );
not ( n36667 , n31979 );
and ( n36668 , n36667 , n31990 );
xor ( n36669 , n35151 , n36668 );
xor ( n36670 , n36666 , n36669 );
not ( n36671 , n31998 );
and ( n36672 , n36671 , n32000 );
xor ( n36673 , n35159 , n36672 );
xor ( n36674 , n36670 , n36673 );
not ( n36675 , n32015 );
and ( n36676 , n36675 , n31933 );
xor ( n36677 , n35165 , n36676 );
xor ( n36678 , n36674 , n36677 );
not ( n36679 , n32021 );
and ( n36680 , n36679 , n32032 );
xor ( n36681 , n35173 , n36680 );
xor ( n36682 , n36678 , n36681 );
xor ( n36683 , n32018 , n36682 );
not ( n36684 , n32051 );
and ( n36685 , n36684 , n32053 );
xor ( n36686 , n35182 , n36685 );
not ( n36687 , n32060 );
and ( n36688 , n36687 , n32062 );
xor ( n36689 , n35189 , n36688 );
xor ( n36690 , n36686 , n36689 );
not ( n36691 , n32070 );
and ( n36692 , n36691 , n32072 );
xor ( n36693 , n35197 , n36692 );
xor ( n36694 , n36690 , n36693 );
not ( n36695 , n32080 );
and ( n36696 , n36695 , n32092 );
xor ( n36697 , n35205 , n36696 );
xor ( n36698 , n36694 , n36697 );
not ( n36699 , n32100 );
and ( n36700 , n36699 , n32102 );
xor ( n36701 , n35213 , n36700 );
xor ( n36702 , n36698 , n36701 );
xor ( n36703 , n36683 , n36702 );
and ( n36704 , n36663 , n36703 );
xor ( n36705 , n35761 , n36704 );
not ( n12005 , n29614 );
and ( n12006 , n12005 , RI17477628_1154);
and ( n12007 , n36705 , n29614 );
or ( n36706 , n12006 , n12007 );
not ( n12008 , RI1754c610_2);
and ( n12009 , n12008 , n36706 );
and ( n12010 , C0 , RI1754c610_2);
or ( n36707 , n12009 , n12010 );
buf ( n36708 , n36707 );
buf ( n36709 , RI174b47f8_856);
buf ( n36710 , RI174a20a8_946);
not ( n12011 , n27683 );
and ( n12012 , n12011 , RI19ab8b38_2390);
and ( n12013 , RI19ac1490_2320 , n27683 );
or ( n36711 , n12012 , n12013 );
not ( n12014 , RI1754c610_2);
and ( n12015 , n12014 , n36711 );
and ( n12016 , C0 , RI1754c610_2);
or ( n36712 , n12015 , n12016 );
buf ( n36713 , n36712 );
buf ( n36714 , RI174686a0_1227);
not ( n36715 , n36534 );
and ( n36716 , n36715 , n34682 );
xor ( n36717 , n34678 , n36716 );
xor ( n36718 , n36717 , n36568 );
not ( n36719 , n30070 );
xor ( n36720 , n27884 , n29387 );
xor ( n36721 , n36720 , n29399 );
and ( n36722 , n36719 , n36721 );
xor ( n36723 , n30067 , n36722 );
xor ( n36724 , n36723 , n30033 );
not ( n36725 , n30152 );
xor ( n36726 , n28211 , n29079 );
xor ( n36727 , n36726 , n28583 );
and ( n36728 , n36725 , n36727 );
xor ( n36729 , n30126 , n36728 );
xor ( n36730 , n36724 , n36729 );
not ( n36731 , n30194 );
xor ( n36732 , n29572 , n32611 );
xor ( n36733 , n36732 , n29161 );
and ( n36734 , n36731 , n36733 );
xor ( n36735 , n30190 , n36734 );
xor ( n36736 , n36730 , n36735 );
not ( n36737 , n30244 );
xor ( n36738 , n27935 , n30364 );
xor ( n36739 , n36738 , n30374 );
and ( n36740 , n36737 , n36739 );
xor ( n36741 , n30222 , n36740 );
xor ( n36742 , n36736 , n36741 );
xor ( n36743 , n36718 , n36742 );
xor ( n36744 , n31787 , n29148 );
xor ( n36745 , n36744 , n32800 );
not ( n36746 , n34875 );
and ( n36747 , n36746 , n34877 );
xor ( n36748 , n36745 , n36747 );
xor ( n36749 , n29670 , n30842 );
xor ( n36750 , n36749 , n32247 );
not ( n36751 , n34884 );
and ( n36752 , n36751 , n34886 );
xor ( n36753 , n36750 , n36752 );
xor ( n36754 , n36748 , n36753 );
xor ( n36755 , n31017 , n31594 );
xor ( n36756 , n36755 , n31487 );
not ( n36757 , n34894 );
and ( n36758 , n36757 , n34896 );
xor ( n36759 , n36756 , n36758 );
xor ( n36760 , n36754 , n36759 );
xor ( n36761 , n27719 , n28533 );
xor ( n36762 , n36761 , n28543 );
not ( n36763 , n34904 );
and ( n36764 , n36763 , n34906 );
xor ( n36765 , n36762 , n36764 );
xor ( n36766 , n36760 , n36765 );
xor ( n36767 , n28074 , n31192 );
xor ( n36768 , n36767 , n27700 );
not ( n36769 , n34914 );
and ( n36770 , n36769 , n34866 );
xor ( n36771 , n36768 , n36770 );
xor ( n36772 , n36766 , n36771 );
xor ( n36773 , n34891 , n36772 );
xor ( n36774 , n30998 , n32256 );
xor ( n36775 , n36774 , n32734 );
not ( n36776 , n34921 );
and ( n36777 , n36776 , n34923 );
xor ( n36778 , n36775 , n36777 );
xor ( n36779 , n31224 , n28741 );
xor ( n36780 , n36779 , n28096 );
not ( n36781 , n34930 );
and ( n36782 , n36781 , n34932 );
xor ( n36783 , n36780 , n36782 );
xor ( n36784 , n36778 , n36783 );
xor ( n36785 , n30714 , n28418 );
xor ( n36786 , n36785 , n31969 );
not ( n36787 , n34940 );
and ( n36788 , n36787 , n34942 );
xor ( n36789 , n36786 , n36788 );
xor ( n36790 , n36784 , n36789 );
xor ( n36791 , n29184 , n28827 );
xor ( n36792 , n36791 , n28839 );
not ( n36793 , n34950 );
and ( n36794 , n36793 , n34952 );
xor ( n36795 , n36792 , n36794 );
xor ( n36796 , n36790 , n36795 );
xor ( n36797 , n30268 , n31697 );
xor ( n36798 , n36797 , n31309 );
not ( n36799 , n34960 );
and ( n36800 , n36799 , n34962 );
xor ( n36801 , n36798 , n36800 );
xor ( n36802 , n36796 , n36801 );
xor ( n36803 , n36773 , n36802 );
not ( n36804 , n36803 );
xor ( n36805 , n29372 , n31989 );
xor ( n36806 , n36805 , n33898 );
xor ( n36807 , n28124 , n30233 );
xor ( n36808 , n36807 , n30243 );
not ( n36809 , n36808 );
and ( n36810 , n36809 , n34544 );
xor ( n36811 , n36806 , n36810 );
not ( n36812 , n34525 );
xor ( n36813 , n29974 , n30813 );
xor ( n36814 , n36813 , n30823 );
and ( n36815 , n36812 , n36814 );
xor ( n36816 , n34522 , n36815 );
xor ( n36817 , n29992 , n28702 );
xor ( n36818 , n36817 , n31065 );
not ( n36819 , n36818 );
xor ( n36820 , n29186 , n28827 );
xor ( n36821 , n36820 , n28839 );
and ( n36822 , n36819 , n36821 );
xor ( n36823 , n34539 , n36822 );
xor ( n36824 , n36816 , n36823 );
not ( n36825 , n36806 );
and ( n36826 , n36825 , n36808 );
xor ( n36827 , n34549 , n36826 );
xor ( n36828 , n36824 , n36827 );
xor ( n36829 , n30787 , n28759 );
xor ( n36830 , n36829 , n28771 );
not ( n36831 , n36830 );
xor ( n36832 , n28799 , n31978 );
xor ( n36833 , n36832 , n29409 );
and ( n36834 , n36831 , n36833 );
xor ( n36835 , n34559 , n36834 );
xor ( n36836 , n36828 , n36835 );
xor ( n36837 , n30545 , n28224 );
xor ( n36838 , n36837 , n28236 );
not ( n36839 , n36838 );
xor ( n36840 , n32777 , n32247 );
xor ( n36841 , n36840 , n32256 );
and ( n36842 , n36839 , n36841 );
xor ( n36843 , n34569 , n36842 );
xor ( n36844 , n36836 , n36843 );
xor ( n36845 , n36811 , n36844 );
xor ( n36846 , n27992 , n29677 );
xor ( n36847 , n36846 , n32778 );
not ( n36848 , n36847 );
and ( n36849 , n36848 , n35517 );
xor ( n36850 , n34580 , n36849 );
xor ( n36851 , n31456 , n27964 );
xor ( n36852 , n36851 , n27975 );
not ( n36853 , n36852 );
and ( n36854 , n36853 , n35522 );
xor ( n36855 , n34589 , n36854 );
xor ( n36856 , n36850 , n36855 );
xor ( n36857 , n32772 , n32247 );
xor ( n36858 , n36857 , n32256 );
not ( n36859 , n36858 );
and ( n36860 , n36859 , n35528 );
xor ( n36861 , n34599 , n36860 );
xor ( n36862 , n36856 , n36861 );
xor ( n36863 , n29806 , n31516 );
xor ( n36864 , n36863 , n31528 );
not ( n36865 , n36864 );
and ( n36866 , n36865 , n35534 );
xor ( n36867 , n34609 , n36866 );
xor ( n36868 , n36862 , n36867 );
xor ( n36869 , n28295 , n31291 );
xor ( n36870 , n36869 , n27989 );
not ( n36871 , n36870 );
and ( n36872 , n36871 , n35540 );
xor ( n36873 , n34619 , n36872 );
xor ( n36874 , n36868 , n36873 );
xor ( n36875 , n36845 , n36874 );
and ( n36876 , n36804 , n36875 );
xor ( n36877 , n36743 , n36876 );
not ( n12017 , n29614 );
and ( n12018 , n12017 , RI17340378_2128);
and ( n12019 , n36877 , n29614 );
or ( n36878 , n12018 , n12019 );
not ( n12020 , RI1754c610_2);
and ( n12021 , n12020 , n36878 );
and ( n12022 , C0 , RI1754c610_2);
or ( n36879 , n12021 , n12022 );
buf ( n36880 , n36879 );
not ( n36881 , n34090 );
and ( n36882 , n36881 , n34092 );
xor ( n36883 , n33888 , n36882 );
xor ( n36884 , n36883 , n36431 );
xor ( n36885 , n36884 , n34221 );
not ( n36886 , n34889 );
xor ( n36887 , n30938 , n29586 );
xor ( n36888 , n36887 , n28355 );
and ( n36889 , n36886 , n36888 );
xor ( n36890 , n34886 , n36889 );
xor ( n36891 , n36890 , n34918 );
xor ( n36892 , n36891 , n34968 );
not ( n36893 , n36892 );
xor ( n36894 , n32501 , n32275 );
xor ( n36895 , n36894 , n31950 );
not ( n36896 , n36895 );
xor ( n36897 , n33383 , n28069 );
xor ( n36898 , n36897 , n28081 );
and ( n36899 , n36896 , n36898 );
xor ( n36900 , n32536 , n36899 );
not ( n36901 , n32526 );
xor ( n36902 , n27849 , n29655 );
xor ( n36903 , n36902 , n29601 );
and ( n36904 , n36901 , n36903 );
xor ( n36905 , n32522 , n36904 );
xor ( n36906 , n32513 , n36905 );
not ( n36907 , n32536 );
and ( n36908 , n36907 , n36895 );
xor ( n36909 , n32533 , n36908 );
xor ( n36910 , n36906 , n36909 );
xor ( n36911 , n36910 , n36022 );
not ( n36912 , n32557 );
xor ( n36913 , n29323 , n31226 );
xor ( n36914 , n36913 , n31516 );
and ( n36915 , n36912 , n36914 );
xor ( n36916 , n32554 , n36915 );
xor ( n36917 , n36911 , n36916 );
xor ( n36918 , n36900 , n36917 );
not ( n36919 , n32568 );
xor ( n36920 , n29581 , n29767 );
xor ( n36921 , n36920 , n30510 );
and ( n36922 , n36919 , n36921 );
xor ( n36923 , n32565 , n36922 );
not ( n36924 , n32577 );
xor ( n36925 , n28873 , n30218 );
xor ( n36926 , n36925 , n27807 );
and ( n36927 , n36924 , n36926 );
xor ( n36928 , n32574 , n36927 );
xor ( n36929 , n36923 , n36928 );
not ( n36930 , n32587 );
xor ( n36931 , n29382 , n33665 );
xor ( n36932 , n36931 , n32209 );
and ( n36933 , n36930 , n36932 );
xor ( n36934 , n32584 , n36933 );
xor ( n36935 , n36929 , n36934 );
not ( n36936 , n32597 );
xor ( n36937 , n29689 , n30972 );
xor ( n36938 , n36937 , n29123 );
and ( n36939 , n36936 , n36938 );
xor ( n36940 , n32594 , n36939 );
xor ( n36941 , n36935 , n36940 );
not ( n36942 , n32617 );
xor ( n36943 , n32986 , n30415 );
xor ( n36944 , n36943 , n30427 );
and ( n36945 , n36942 , n36944 );
xor ( n36946 , n32614 , n36945 );
xor ( n36947 , n36941 , n36946 );
xor ( n36948 , n36918 , n36947 );
and ( n36949 , n36893 , n36948 );
xor ( n36950 , n36885 , n36949 );
not ( n12023 , n29614 );
and ( n12024 , n12023 , RI17444bb0_1401);
and ( n12025 , n36950 , n29614 );
or ( n36951 , n12024 , n12025 );
not ( n12026 , RI1754c610_2);
and ( n12027 , n12026 , n36951 );
and ( n12028 , C0 , RI1754c610_2);
or ( n36952 , n12027 , n12028 );
buf ( n36953 , n36952 );
not ( n12029 , n27683 );
and ( n12030 , n12029 , RI19a8a080_2724);
and ( n12031 , RI19a93fe0_2654 , n27683 );
or ( n36954 , n12030 , n12031 );
not ( n12032 , RI1754c610_2);
and ( n12033 , n12032 , n36954 );
and ( n12034 , C0 , RI1754c610_2);
or ( n36955 , n12033 , n12034 );
buf ( n36956 , n36955 );
xor ( n36957 , n27986 , n28929 );
xor ( n36958 , n36957 , n29677 );
not ( n36959 , n35314 );
and ( n36960 , n36959 , n35316 );
xor ( n36961 , n36958 , n36960 );
xor ( n36962 , n30048 , n28904 );
xor ( n36963 , n36962 , n29291 );
not ( n36964 , n36958 );
and ( n36965 , n36964 , n35314 );
xor ( n36966 , n36963 , n36965 );
xor ( n36967 , n29776 , n28627 );
xor ( n36968 , n36967 , n30089 );
xor ( n36969 , n31306 , n31636 );
xor ( n36970 , n36969 , n30655 );
not ( n36971 , n36970 );
and ( n36972 , n36971 , n35323 );
xor ( n36973 , n36968 , n36972 );
xor ( n36974 , n36966 , n36973 );
xor ( n36975 , n30470 , n32894 );
xor ( n36976 , n36975 , n32991 );
xor ( n36977 , n31160 , n27779 );
xor ( n36978 , n36977 , n27791 );
not ( n36979 , n36978 );
and ( n36980 , n36979 , n35333 );
xor ( n36981 , n36976 , n36980 );
xor ( n36982 , n36974 , n36981 );
xor ( n36983 , n28401 , n31497 );
xor ( n36984 , n36983 , n31247 );
xor ( n36985 , n29852 , n29421 );
xor ( n36986 , n36985 , n30643 );
not ( n36987 , n36986 );
and ( n36988 , n36987 , n35343 );
xor ( n36989 , n36984 , n36988 );
xor ( n36990 , n36982 , n36989 );
xor ( n36991 , n30228 , n28160 );
xor ( n36992 , n36991 , n28250 );
xor ( n36993 , n29090 , n28493 );
xor ( n36994 , n36993 , n28505 );
not ( n36995 , n36994 );
and ( n36996 , n36995 , n35353 );
xor ( n36997 , n36992 , n36996 );
xor ( n36998 , n36990 , n36997 );
xor ( n36999 , n36961 , n36998 );
xor ( n37000 , n29600 , n28200 );
xor ( n37001 , n37000 , n28212 );
xor ( n37002 , n30435 , n28956 );
xor ( n37003 , n37002 , n29995 );
not ( n37004 , n37003 );
xor ( n37005 , n31302 , n31636 );
xor ( n37006 , n37005 , n30655 );
and ( n37007 , n37004 , n37006 );
xor ( n37008 , n37001 , n37007 );
xor ( n37009 , n29122 , n29873 );
xor ( n37010 , n37009 , n32398 );
xor ( n37011 , n31982 , n28785 );
xor ( n37012 , n37011 , n28015 );
not ( n37013 , n37012 );
xor ( n37014 , n28306 , n27989 );
xor ( n37015 , n37014 , n28001 );
and ( n37016 , n37013 , n37015 );
xor ( n37017 , n37010 , n37016 );
xor ( n37018 , n37008 , n37017 );
xor ( n37019 , n28518 , n29724 );
xor ( n37020 , n37019 , n31291 );
xor ( n37021 , n29986 , n28702 );
xor ( n37022 , n37021 , n31065 );
not ( n37023 , n37022 );
xor ( n37024 , n31145 , n31843 );
xor ( n37025 , n37024 , n27779 );
and ( n37026 , n37023 , n37025 );
xor ( n37027 , n37020 , n37026 );
xor ( n37028 , n37018 , n37027 );
xor ( n37029 , n28080 , n31192 );
xor ( n37030 , n37029 , n27700 );
xor ( n37031 , n30324 , n33234 );
xor ( n37032 , n37031 , n31825 );
not ( n37033 , n37032 );
xor ( n37034 , n29621 , n30799 );
xor ( n37035 , n37034 , n28148 );
and ( n37036 , n37033 , n37035 );
xor ( n37037 , n37030 , n37036 );
xor ( n37038 , n37028 , n37037 );
xor ( n37039 , n32322 , n29781 );
xor ( n37040 , n37039 , n29793 );
xor ( n37041 , n28664 , n28236 );
xor ( n37042 , n37041 , n29711 );
not ( n37043 , n37042 );
xor ( n37044 , n27812 , n33390 );
xor ( n37045 , n37044 , n28983 );
and ( n37046 , n37043 , n37045 );
xor ( n37047 , n37040 , n37046 );
xor ( n37048 , n37038 , n37047 );
xor ( n37049 , n36999 , n37048 );
not ( n37050 , n35387 );
and ( n37051 , n37050 , n36313 );
xor ( n37052 , n35384 , n37051 );
xor ( n37053 , n37052 , n35416 );
xor ( n37054 , n37053 , n29843 );
not ( n37055 , n37054 );
not ( n37056 , n31325 );
and ( n37057 , n37056 , n31327 );
xor ( n37058 , n28879 , n37057 );
not ( n37059 , n31337 );
and ( n37060 , n37059 , n31339 );
xor ( n37061 , n28934 , n37060 );
xor ( n37062 , n37058 , n37061 );
not ( n37063 , n31345 );
and ( n37064 , n37063 , n31347 );
xor ( n37065 , n28996 , n37064 );
xor ( n37066 , n37062 , n37065 );
not ( n37067 , n31355 );
and ( n37068 , n37067 , n31368 );
xor ( n37069 , n29063 , n37068 );
xor ( n37070 , n37066 , n37069 );
not ( n37071 , n31374 );
and ( n37072 , n37071 , n31376 );
xor ( n37073 , n29106 , n37072 );
xor ( n37074 , n37070 , n37073 );
xor ( n37075 , n31350 , n37074 );
xor ( n37076 , n31286 , n28917 );
xor ( n37077 , n37076 , n28929 );
not ( n37078 , n36436 );
and ( n37079 , n37078 , n35864 );
xor ( n37080 , n37077 , n37079 );
xor ( n37081 , n29442 , n30030 );
xor ( n37082 , n37081 , n30972 );
not ( n37083 , n36441 );
and ( n37084 , n37083 , n35873 );
xor ( n37085 , n37082 , n37084 );
xor ( n37086 , n37080 , n37085 );
xor ( n37087 , n30648 , n31794 );
xor ( n37088 , n37087 , n28969 );
not ( n37089 , n36447 );
and ( n37090 , n37089 , n35883 );
xor ( n37091 , n37088 , n37090 );
xor ( n37092 , n37086 , n37091 );
xor ( n37093 , n31963 , n27885 );
xor ( n37094 , n37093 , n27897 );
not ( n37095 , n36453 );
and ( n37096 , n37095 , n35893 );
xor ( n37097 , n37094 , n37096 );
xor ( n37098 , n37092 , n37097 );
xor ( n37099 , n30504 , n29051 );
xor ( n37100 , n37099 , n29062 );
not ( n37101 , n36459 );
and ( n37102 , n37101 , n35903 );
xor ( n37103 , n37100 , n37102 );
xor ( n37104 , n37098 , n37103 );
xor ( n37105 , n37075 , n37104 );
and ( n37106 , n37055 , n37105 );
xor ( n37107 , n37049 , n37106 );
not ( n12035 , n29614 );
and ( n12036 , n12035 , RI174b7c78_840);
and ( n12037 , n37107 , n29614 );
or ( n37108 , n12036 , n12037 );
not ( n12038 , RI1754c610_2);
and ( n12039 , n12038 , n37108 );
and ( n12040 , C0 , RI1754c610_2);
or ( n37109 , n12039 , n12040 );
buf ( n37110 , n37109 );
not ( n37111 , n35807 );
and ( n37112 , n37111 , n35809 );
xor ( n37113 , n35672 , n37112 );
not ( n37114 , n35663 );
and ( n37115 , n37114 , n35814 );
xor ( n37116 , n35660 , n37115 );
xor ( n37117 , n37113 , n37116 );
not ( n37118 , n35820 );
and ( n37119 , n37118 , n35822 );
xor ( n37120 , n35687 , n37119 );
xor ( n37121 , n37117 , n37120 );
not ( n37122 , n35828 );
and ( n37123 , n37122 , n35830 );
xor ( n37124 , n35697 , n37123 );
xor ( n37125 , n37121 , n37124 );
not ( n37126 , n35836 );
and ( n37127 , n37126 , n35838 );
xor ( n37128 , n35707 , n37127 );
xor ( n37129 , n37125 , n37128 );
xor ( n37130 , n35841 , n37129 );
xor ( n37131 , n30750 , n29161 );
xor ( n37132 , n37131 , n28069 );
not ( n37133 , n37132 );
xor ( n37134 , n29483 , n28450 );
xor ( n37135 , n37134 , n30789 );
and ( n37136 , n37133 , n37135 );
xor ( n37137 , n35718 , n37136 );
xor ( n37138 , n28830 , n28569 );
xor ( n37139 , n37138 , n29889 );
not ( n37140 , n37139 );
xor ( n37141 , n30710 , n28418 );
xor ( n37142 , n37141 , n31969 );
and ( n37143 , n37140 , n37142 );
xor ( n37144 , n35727 , n37143 );
xor ( n37145 , n37137 , n37144 );
xor ( n37146 , n28060 , n31180 );
xor ( n37147 , n37146 , n31192 );
not ( n37148 , n37147 );
xor ( n37149 , n28048 , n29694 );
xor ( n37150 , n37149 , n30457 );
and ( n37151 , n37148 , n37150 );
xor ( n37152 , n35737 , n37151 );
xor ( n37153 , n37145 , n37152 );
xor ( n37154 , n30609 , n28595 );
xor ( n37155 , n37154 , n28519 );
not ( n37156 , n37155 );
xor ( n37157 , n30420 , n31475 );
xor ( n37158 , n37157 , n31763 );
and ( n37159 , n37156 , n37158 );
xor ( n37160 , n35747 , n37159 );
xor ( n37161 , n37153 , n37160 );
xor ( n37162 , n30199 , n29561 );
xor ( n37163 , n37162 , n29573 );
not ( n37164 , n37163 );
xor ( n37165 , n29512 , n30655 );
xor ( n37166 , n37165 , n30665 );
and ( n37167 , n37164 , n37166 );
xor ( n37168 , n35757 , n37167 );
xor ( n37169 , n37161 , n37168 );
xor ( n37170 , n37130 , n37169 );
not ( n37171 , n32431 );
and ( n37172 , n37171 , n32752 );
xor ( n37173 , n32428 , n37172 );
xor ( n37174 , n36152 , n37173 );
not ( n37175 , n32441 );
and ( n37176 , n37175 , n32721 );
xor ( n37177 , n32438 , n37176 );
xor ( n37178 , n37174 , n37177 );
not ( n37179 , n32461 );
and ( n37180 , n37179 , n32764 );
xor ( n37181 , n32448 , n37180 );
xor ( n37182 , n37178 , n37181 );
not ( n37183 , n32478 );
and ( n37184 , n37183 , n32780 );
xor ( n37185 , n32474 , n37184 );
xor ( n37186 , n37182 , n37185 );
xor ( n37187 , n32750 , n37186 );
not ( n37188 , n32789 );
and ( n37189 , n37188 , n32791 );
xor ( n37190 , n32997 , n37189 );
not ( n37191 , n32814 );
and ( n37192 , n37191 , n32816 );
xor ( n37193 , n33004 , n37192 );
xor ( n37194 , n37190 , n37193 );
xor ( n37195 , n37194 , n32981 );
not ( n37196 , n32845 );
and ( n37197 , n37196 , n32847 );
xor ( n37198 , n33018 , n37197 );
xor ( n37199 , n37195 , n37198 );
not ( n37200 , n32855 );
and ( n37201 , n37200 , n32857 );
xor ( n37202 , n33026 , n37201 );
xor ( n37203 , n37199 , n37202 );
xor ( n37204 , n37187 , n37203 );
not ( n37205 , n37204 );
not ( n37206 , n34277 );
and ( n37207 , n37206 , n31428 );
xor ( n37208 , n34274 , n37207 );
xor ( n37209 , n37208 , n34300 );
xor ( n37210 , n37209 , n34340 );
and ( n37211 , n37205 , n37210 );
xor ( n37212 , n37170 , n37211 );
not ( n12041 , n29614 );
and ( n12042 , n12041 , RI17404380_1487);
and ( n12043 , n37212 , n29614 );
or ( n37213 , n12042 , n12043 );
not ( n12044 , RI1754c610_2);
and ( n12045 , n12044 , n37213 );
and ( n12046 , C0 , RI1754c610_2);
or ( n37214 , n12045 , n12046 );
buf ( n37215 , n37214 );
buf ( n37216 , RI17468358_1228);
not ( n37217 , n33128 );
and ( n37218 , n37217 , n33130 );
xor ( n37219 , n36581 , n37218 );
not ( n37220 , n33137 );
and ( n37221 , n37220 , n33139 );
xor ( n37222 , n36573 , n37221 );
xor ( n37223 , n37219 , n37222 );
not ( n37224 , n33147 );
and ( n37225 , n37224 , n33149 );
xor ( n37226 , n36592 , n37225 );
xor ( n37227 , n37223 , n37226 );
not ( n37228 , n33157 );
and ( n37229 , n37228 , n33159 );
xor ( n37230 , n36600 , n37229 );
xor ( n37231 , n37227 , n37230 );
not ( n37232 , n33167 );
and ( n37233 , n37232 , n33169 );
xor ( n37234 , n36608 , n37233 );
xor ( n37235 , n37231 , n37234 );
xor ( n37236 , n33164 , n37235 );
not ( n37237 , n34764 );
and ( n37238 , n37237 , n34766 );
xor ( n37239 , n33527 , n37238 );
not ( n37240 , n34771 );
and ( n37241 , n37240 , n34759 );
xor ( n37242 , n33536 , n37241 );
xor ( n37243 , n37239 , n37242 );
not ( n37244 , n34777 );
and ( n37245 , n37244 , n34779 );
xor ( n37246 , n33548 , n37245 );
xor ( n37247 , n37243 , n37246 );
not ( n37248 , n33518 );
and ( n37249 , n37248 , n34785 );
xor ( n37250 , n33515 , n37249 );
xor ( n37251 , n37247 , n37250 );
not ( n37252 , n34791 );
and ( n37253 , n37252 , n34793 );
xor ( n37254 , n33564 , n37253 );
xor ( n37255 , n37251 , n37254 );
xor ( n37256 , n37236 , n37255 );
not ( n37257 , n31210 );
and ( n37258 , n37257 , n35046 );
xor ( n37259 , n31206 , n37258 );
xor ( n37260 , n37259 , n31213 );
xor ( n37261 , n37260 , n31317 );
not ( n37262 , n37261 );
not ( n37263 , n31645 );
and ( n37264 , n37263 , n35471 );
xor ( n37265 , n30523 , n37264 );
xor ( n37266 , n37265 , n31664 );
xor ( n37267 , n37266 , n31725 );
and ( n37268 , n37262 , n37267 );
xor ( n37269 , n37256 , n37268 );
not ( n12047 , n29614 );
and ( n12048 , n12047 , RI173f3d00_1567);
and ( n12049 , n37269 , n29614 );
or ( n37270 , n12048 , n12049 );
not ( n12050 , RI1754c610_2);
and ( n12051 , n12050 , n37270 );
and ( n12052 , C0 , RI1754c610_2);
or ( n37271 , n12051 , n12052 );
buf ( n37272 , n37271 );
not ( n37273 , n33883 );
and ( n37274 , n37273 , n33885 );
xor ( n37275 , n34092 , n37274 );
not ( n37276 , n33892 );
and ( n37277 , n37276 , n33899 );
xor ( n37278 , n34099 , n37277 );
xor ( n37279 , n37275 , n37278 );
not ( n37280 , n33907 );
and ( n37281 , n37280 , n33909 );
xor ( n37282 , n34107 , n37281 );
xor ( n37283 , n37279 , n37282 );
not ( n37284 , n33917 );
and ( n37285 , n37284 , n33919 );
xor ( n37286 , n34115 , n37285 );
xor ( n37287 , n37283 , n37286 );
not ( n37288 , n33927 );
and ( n37289 , n37288 , n33929 );
xor ( n37290 , n34123 , n37289 );
xor ( n37291 , n37287 , n37290 );
xor ( n37292 , n33890 , n37291 );
not ( n37293 , n35652 );
and ( n37294 , n37293 , n34194 );
xor ( n37295 , n33953 , n37294 );
not ( n37296 , n36267 );
and ( n37297 , n37296 , n34199 );
xor ( n37298 , n33962 , n37297 );
xor ( n37299 , n37295 , n37298 );
not ( n37300 , n36273 );
and ( n37301 , n37300 , n34205 );
xor ( n37302 , n33972 , n37301 );
xor ( n37303 , n37299 , n37302 );
not ( n37304 , n33944 );
and ( n37305 , n37304 , n34211 );
xor ( n37306 , n33941 , n37305 );
xor ( n37307 , n37303 , n37306 );
not ( n37308 , n36283 );
and ( n37309 , n37308 , n34217 );
xor ( n37310 , n33988 , n37309 );
xor ( n37311 , n37307 , n37310 );
xor ( n37312 , n37292 , n37311 );
not ( n37313 , n35769 );
and ( n37314 , n37313 , n35771 );
xor ( n37315 , n33345 , n37314 );
not ( n37316 , n35776 );
and ( n37317 , n37316 , n35778 );
xor ( n37318 , n33354 , n37317 );
xor ( n37319 , n37315 , n37318 );
not ( n37320 , n35784 );
and ( n37321 , n37320 , n35764 );
xor ( n37322 , n33364 , n37321 );
xor ( n37323 , n37319 , n37322 );
not ( n37324 , n35790 );
and ( n37325 , n37324 , n35792 );
xor ( n37326 , n33374 , n37325 );
xor ( n37327 , n37323 , n37326 );
not ( n37328 , n35798 );
and ( n37329 , n37328 , n35800 );
xor ( n37330 , n33394 , n37329 );
xor ( n37331 , n37327 , n37330 );
xor ( n37332 , n35781 , n37331 );
xor ( n37333 , n37332 , n37129 );
not ( n37334 , n37333 );
not ( n37335 , n33318 );
xor ( n37336 , n32425 , n32167 );
xor ( n37337 , n37336 , n31843 );
and ( n37338 , n37335 , n37337 );
xor ( n37339 , n33315 , n37338 );
xor ( n37340 , n37339 , n33337 );
xor ( n37341 , n37340 , n33397 );
and ( n37342 , n37334 , n37341 );
xor ( n37343 , n37312 , n37342 );
not ( n12053 , n29614 );
and ( n12054 , n12053 , RI17468d30_1225);
and ( n12055 , n37343 , n29614 );
or ( n37344 , n12054 , n12055 );
not ( n12056 , RI1754c610_2);
and ( n12057 , n12056 , n37344 );
and ( n12058 , C0 , RI1754c610_2);
or ( n37345 , n12057 , n12058 );
buf ( n37346 , n37345 );
not ( n37347 , n28056 );
and ( n37348 , n37347 , n28082 );
xor ( n37349 , n29977 , n37348 );
xor ( n37350 , n37349 , n29981 );
xor ( n37351 , n37350 , n35955 );
xor ( n37352 , n36038 , n34475 );
not ( n37353 , n33463 );
and ( n37354 , n37353 , n36065 );
xor ( n37355 , n33460 , n37354 );
not ( n37356 , n33472 );
and ( n37357 , n37356 , n36072 );
xor ( n37358 , n33469 , n37357 );
xor ( n37359 , n37355 , n37358 );
not ( n37360 , n33482 );
and ( n37361 , n37360 , n36080 );
xor ( n37362 , n33479 , n37361 );
xor ( n37363 , n37359 , n37362 );
not ( n37364 , n33492 );
and ( n37365 , n37364 , n36088 );
xor ( n37366 , n33489 , n37365 );
xor ( n37367 , n37363 , n37366 );
not ( n37368 , n33502 );
and ( n37369 , n37368 , n36096 );
xor ( n37370 , n33499 , n37369 );
xor ( n37371 , n37367 , n37370 );
xor ( n37372 , n37352 , n37371 );
not ( n37373 , n37372 );
xor ( n37374 , n28631 , n34497 );
xor ( n37375 , n37374 , n34517 );
and ( n37376 , n37373 , n37375 );
xor ( n37377 , n37351 , n37376 );
not ( n12059 , n29614 );
and ( n12060 , n12059 , RI174053e8_1482);
and ( n12061 , n37377 , n29614 );
or ( n37378 , n12060 , n12061 );
not ( n12062 , RI1754c610_2);
and ( n12063 , n12062 , n37378 );
and ( n12064 , C0 , RI1754c610_2);
or ( n37379 , n12063 , n12064 );
buf ( n37380 , n37379 );
not ( n12065 , n27683 );
and ( n12066 , n12065 , RI19acc9f8_2234);
and ( n12067 , RI19a88a00_2734 , n27683 );
or ( n37381 , n12066 , n12067 );
not ( n12068 , RI1754c610_2);
and ( n12069 , n12068 , n37381 );
and ( n12070 , C0 , RI1754c610_2);
or ( n37382 , n12069 , n12070 );
buf ( n37383 , n37382 );
xor ( n37384 , n35938 , n36148 );
not ( n37385 , n36483 );
xor ( n37386 , n27733 , n28543 );
xor ( n37387 , n37386 , n32120 );
and ( n37388 , n37385 , n37387 );
xor ( n37389 , n36480 , n37388 );
xor ( n37390 , n29072 , n30643 );
xor ( n37391 , n37390 , n29176 );
not ( n37392 , n37391 );
xor ( n37393 , n31576 , n29134 );
xor ( n37394 , n37393 , n27936 );
and ( n37395 , n37392 , n37394 );
xor ( n37396 , n36497 , n37395 );
xor ( n37397 , n37389 , n37396 );
xor ( n37398 , n28610 , n29995 );
xor ( n37399 , n37398 , n28327 );
not ( n37400 , n37399 );
xor ( n37401 , n27984 , n28929 );
xor ( n37402 , n37401 , n29677 );
and ( n37403 , n37400 , n37402 );
xor ( n37404 , n36507 , n37403 );
xor ( n37405 , n37397 , n37404 );
xor ( n37406 , n30515 , n29062 );
xor ( n37407 , n37406 , n31613 );
not ( n37408 , n37407 );
xor ( n37409 , n31916 , n32426 );
xor ( n37410 , n37409 , n31152 );
and ( n37411 , n37408 , n37410 );
xor ( n37412 , n36517 , n37411 );
xor ( n37413 , n37405 , n37412 );
xor ( n37414 , n32359 , n32835 );
xor ( n37415 , n37414 , n31399 );
not ( n37416 , n37415 );
xor ( n37417 , n29970 , n30813 );
xor ( n37418 , n37417 , n30823 );
and ( n37419 , n37416 , n37418 );
xor ( n37420 , n36527 , n37419 );
xor ( n37421 , n37413 , n37420 );
xor ( n37422 , n37384 , n37421 );
not ( n37423 , n34692 );
and ( n37424 , n37423 , n36538 );
xor ( n37425 , n34689 , n37424 );
xor ( n37426 , n34680 , n37425 );
not ( n37427 , n34702 );
and ( n37428 , n37427 , n36546 );
xor ( n37429 , n34699 , n37428 );
xor ( n37430 , n37426 , n37429 );
not ( n37431 , n34712 );
and ( n37432 , n37431 , n36554 );
xor ( n37433 , n34709 , n37432 );
xor ( n37434 , n37430 , n37433 );
not ( n37435 , n34722 );
and ( n37436 , n37435 , n36562 );
xor ( n37437 , n34719 , n37436 );
xor ( n37438 , n37434 , n37437 );
xor ( n37439 , n36559 , n37438 );
xor ( n37440 , n37439 , n30247 );
not ( n37441 , n37440 );
not ( n37442 , n35517 );
and ( n37443 , n37442 , n34575 );
xor ( n37444 , n36847 , n37443 );
not ( n37445 , n35522 );
and ( n37446 , n37445 , n34584 );
xor ( n37447 , n36852 , n37446 );
xor ( n37448 , n37444 , n37447 );
not ( n37449 , n35528 );
and ( n37450 , n37449 , n34594 );
xor ( n37451 , n36858 , n37450 );
xor ( n37452 , n37448 , n37451 );
not ( n37453 , n35534 );
and ( n37454 , n37453 , n34604 );
xor ( n37455 , n36864 , n37454 );
xor ( n37456 , n37452 , n37455 );
not ( n37457 , n35540 );
and ( n37458 , n37457 , n34614 );
xor ( n37459 , n36870 , n37458 );
xor ( n37460 , n37456 , n37459 );
xor ( n37461 , n35543 , n37460 );
xor ( n37462 , n28612 , n29995 );
xor ( n37463 , n37462 , n28327 );
not ( n37464 , n35547 );
and ( n37465 , n37464 , n35549 );
xor ( n37466 , n37463 , n37465 );
xor ( n37467 , n30482 , n32991 );
xor ( n37468 , n37467 , n32996 );
not ( n37469 , n35556 );
and ( n37470 , n37469 , n35558 );
xor ( n37471 , n37468 , n37470 );
xor ( n37472 , n37466 , n37471 );
xor ( n37473 , n31417 , n29332 );
xor ( n37474 , n37473 , n29814 );
not ( n37475 , n35566 );
and ( n37476 , n37475 , n35568 );
xor ( n37477 , n37474 , n37476 );
xor ( n37478 , n37472 , n37477 );
xor ( n37479 , n31608 , n29839 );
xor ( n37480 , n37479 , n32031 );
not ( n37481 , n35576 );
and ( n37482 , n37481 , n35578 );
xor ( n37483 , n37480 , n37482 );
xor ( n37484 , n37478 , n37483 );
xor ( n37485 , n28219 , n30457 );
xor ( n37486 , n37485 , n31581 );
not ( n37487 , n35586 );
and ( n37488 , n37487 , n35588 );
xor ( n37489 , n37486 , n37488 );
xor ( n37490 , n37484 , n37489 );
xor ( n37491 , n37461 , n37490 );
and ( n37492 , n37441 , n37491 );
xor ( n37493 , n37422 , n37492 );
not ( n12071 , n29614 );
and ( n12072 , n12071 , RI1747e900_1119);
and ( n12073 , n37493 , n29614 );
or ( n37494 , n12072 , n12073 );
not ( n12074 , RI1754c610_2);
and ( n12075 , n12074 , n37494 );
and ( n12076 , C0 , RI1754c610_2);
or ( n37495 , n12075 , n12076 );
buf ( n37496 , n37495 );
xor ( n37497 , n34197 , n36287 );
xor ( n37498 , n32733 , n30475 );
xor ( n37499 , n37498 , n30487 );
not ( n37500 , n34224 );
and ( n37501 , n37500 , n33994 );
xor ( n37502 , n37499 , n37501 );
xor ( n37503 , n31023 , n31594 );
xor ( n37504 , n37503 , n31487 );
not ( n37505 , n34229 );
and ( n37506 , n37505 , n34003 );
xor ( n37507 , n37504 , n37506 );
xor ( n37508 , n37502 , n37507 );
xor ( n37509 , n31824 , n29375 );
xor ( n37510 , n37509 , n29767 );
not ( n37511 , n34235 );
and ( n37512 , n37511 , n34013 );
xor ( n37513 , n37510 , n37512 );
xor ( n37514 , n37508 , n37513 );
xor ( n37515 , n28326 , n31065 );
xor ( n37516 , n37515 , n31076 );
not ( n37517 , n34241 );
and ( n37518 , n37517 , n34023 );
xor ( n37519 , n37516 , n37518 );
xor ( n37520 , n37514 , n37519 );
xor ( n37521 , n27896 , n29399 );
xor ( n37522 , n37521 , n29655 );
not ( n37523 , n34247 );
and ( n37524 , n37523 , n34033 );
xor ( n37525 , n37522 , n37524 );
xor ( n37526 , n37520 , n37525 );
xor ( n37527 , n37497 , n37526 );
not ( n37528 , n36888 );
and ( n37529 , n37528 , n36750 );
xor ( n37530 , n34889 , n37529 );
not ( n37531 , n34880 );
xor ( n37532 , n28693 , n32472 );
xor ( n37533 , n37532 , n32323 );
and ( n37534 , n37531 , n37533 );
xor ( n37535 , n34877 , n37534 );
xor ( n37536 , n37535 , n36890 );
not ( n37537 , n34899 );
xor ( n37538 , n32315 , n29781 );
xor ( n37539 , n37538 , n29793 );
and ( n37540 , n37537 , n37539 );
xor ( n37541 , n34896 , n37540 );
xor ( n37542 , n37536 , n37541 );
not ( n37543 , n34909 );
xor ( n37544 , n29367 , n31989 );
xor ( n37545 , n37544 , n33898 );
and ( n37546 , n37543 , n37545 );
xor ( n37547 , n34906 , n37546 );
xor ( n37548 , n37542 , n37547 );
xor ( n37549 , n37548 , n34873 );
xor ( n37550 , n37530 , n37549 );
not ( n37551 , n34926 );
xor ( n37552 , n30650 , n31794 );
xor ( n37553 , n37552 , n28969 );
and ( n37554 , n37551 , n37553 );
xor ( n37555 , n34923 , n37554 );
not ( n37556 , n34935 );
xor ( n37557 , n32421 , n32167 );
xor ( n37558 , n37557 , n31843 );
and ( n37559 , n37556 , n37558 );
xor ( n37560 , n34932 , n37559 );
xor ( n37561 , n37555 , n37560 );
not ( n37562 , n34945 );
xor ( n37563 , n33229 , n29364 );
xor ( n37564 , n37563 , n29375 );
and ( n37565 , n37562 , n37564 );
xor ( n37566 , n34942 , n37565 );
xor ( n37567 , n37561 , n37566 );
not ( n37568 , n34955 );
xor ( n37569 , n27892 , n29399 );
xor ( n37570 , n37569 , n29655 );
and ( n37571 , n37568 , n37570 );
xor ( n37572 , n34952 , n37571 );
xor ( n37573 , n37567 , n37572 );
not ( n37574 , n34965 );
xor ( n37575 , n28887 , n30066 );
xor ( n37576 , n37575 , n30007 );
and ( n37577 , n37574 , n37576 );
xor ( n37578 , n34962 , n37577 );
xor ( n37579 , n37573 , n37578 );
xor ( n37580 , n37550 , n37579 );
not ( n37581 , n37580 );
xor ( n37582 , n31122 , n31528 );
xor ( n37583 , n37582 , n32835 );
not ( n37584 , n35100 );
and ( n37585 , n37584 , n35102 );
xor ( n37586 , n37583 , n37585 );
xor ( n37587 , n29133 , n32398 );
xor ( n37588 , n37587 , n30364 );
xor ( n37589 , n29002 , n29814 );
xor ( n37590 , n37589 , n31131 );
not ( n37591 , n37590 );
and ( n37592 , n37591 , n35081 );
xor ( n37593 , n37588 , n37592 );
xor ( n37594 , n30654 , n31794 );
xor ( n37595 , n37594 , n28969 );
xor ( n37596 , n28791 , n31978 );
xor ( n37597 , n37596 , n29409 );
not ( n37598 , n37597 );
and ( n37599 , n37598 , n35090 );
xor ( n37600 , n37595 , n37599 );
xor ( n37601 , n37593 , n37600 );
xor ( n37602 , n29780 , n28627 );
xor ( n37603 , n37602 , n30089 );
not ( n37604 , n37583 );
and ( n37605 , n37604 , n35100 );
xor ( n37606 , n37603 , n37605 );
xor ( n37607 , n37601 , n37606 );
xor ( n37608 , n31749 , n28262 );
xor ( n37609 , n37608 , n28892 );
xor ( n37610 , n27877 , n29387 );
xor ( n37611 , n37610 , n29399 );
not ( n37612 , n37611 );
and ( n37613 , n37612 , n35110 );
xor ( n37614 , n37609 , n37613 );
xor ( n37615 , n37607 , n37614 );
xor ( n37616 , n32509 , n32275 );
xor ( n37617 , n37616 , n31950 );
xor ( n37618 , n32794 , n31100 );
xor ( n37619 , n37618 , n31422 );
not ( n37620 , n37619 );
and ( n37621 , n37620 , n35120 );
xor ( n37622 , n37617 , n37621 );
xor ( n37623 , n37615 , n37622 );
xor ( n37624 , n37586 , n37623 );
xor ( n37625 , n29760 , n33898 );
xor ( n37626 , n37625 , n29051 );
not ( n37627 , n32515 );
and ( n37628 , n37627 , n32495 );
xor ( n37629 , n37626 , n37628 );
xor ( n37630 , n32161 , n30139 );
xor ( n37631 , n37630 , n30151 );
not ( n37632 , n32520 );
and ( n37633 , n37632 , n32522 );
xor ( n37634 , n37631 , n37633 );
xor ( n37635 , n37629 , n37634 );
not ( n37636 , n32531 );
and ( n37637 , n37636 , n32533 );
xor ( n37638 , n36898 , n37637 );
xor ( n37639 , n37635 , n37638 );
xor ( n37640 , n27994 , n29677 );
xor ( n37641 , n37640 , n32778 );
not ( n37642 , n32541 );
and ( n37643 , n37642 , n32543 );
xor ( n37644 , n37641 , n37643 );
xor ( n37645 , n37639 , n37644 );
xor ( n37646 , n31743 , n28262 );
xor ( n37647 , n37646 , n28892 );
not ( n37648 , n32552 );
and ( n37649 , n37648 , n32554 );
xor ( n37650 , n37647 , n37649 );
xor ( n37651 , n37645 , n37650 );
xor ( n37652 , n37624 , n37651 );
and ( n37653 , n37581 , n37652 );
xor ( n37654 , n37527 , n37653 );
not ( n12077 , n29614 );
and ( n12078 , n12077 , RI174ab798_900);
and ( n12079 , n37654 , n29614 );
or ( n37655 , n12078 , n12079 );
not ( n12080 , RI1754c610_2);
and ( n12081 , n12080 , n37655 );
and ( n12082 , C0 , RI1754c610_2);
or ( n37656 , n12081 , n12082 );
buf ( n37657 , n37656 );
not ( n37658 , n36750 );
and ( n37659 , n37658 , n34884 );
xor ( n37660 , n36888 , n37659 );
not ( n37661 , n37533 );
and ( n37662 , n37661 , n36745 );
xor ( n37663 , n34880 , n37662 );
xor ( n37664 , n37663 , n37530 );
not ( n37665 , n37539 );
and ( n37666 , n37665 , n36756 );
xor ( n37667 , n34899 , n37666 );
xor ( n37668 , n37664 , n37667 );
not ( n37669 , n37545 );
and ( n37670 , n37669 , n36762 );
xor ( n37671 , n34909 , n37670 );
xor ( n37672 , n37668 , n37671 );
not ( n37673 , n34871 );
and ( n37674 , n37673 , n36768 );
xor ( n37675 , n34868 , n37674 );
xor ( n37676 , n37672 , n37675 );
xor ( n37677 , n37660 , n37676 );
not ( n37678 , n37553 );
and ( n37679 , n37678 , n36775 );
xor ( n37680 , n34926 , n37679 );
not ( n37681 , n37558 );
and ( n37682 , n37681 , n36780 );
xor ( n37683 , n34935 , n37682 );
xor ( n37684 , n37680 , n37683 );
not ( n37685 , n37564 );
and ( n37686 , n37685 , n36786 );
xor ( n37687 , n34945 , n37686 );
xor ( n37688 , n37684 , n37687 );
not ( n37689 , n37570 );
and ( n37690 , n37689 , n36792 );
xor ( n37691 , n34955 , n37690 );
xor ( n37692 , n37688 , n37691 );
not ( n37693 , n37576 );
and ( n37694 , n37693 , n36798 );
xor ( n37695 , n34965 , n37694 );
xor ( n37696 , n37692 , n37695 );
xor ( n37697 , n37677 , n37696 );
not ( n37698 , n37077 );
and ( n37699 , n37698 , n36436 );
xor ( n37700 , n35869 , n37699 );
not ( n37701 , n37082 );
and ( n37702 , n37701 , n36441 );
xor ( n37703 , n35878 , n37702 );
xor ( n37704 , n37700 , n37703 );
not ( n37705 , n37088 );
and ( n37706 , n37705 , n36447 );
xor ( n37707 , n35888 , n37706 );
xor ( n37708 , n37704 , n37707 );
not ( n37709 , n37094 );
and ( n37710 , n37709 , n36453 );
xor ( n37711 , n35898 , n37710 );
xor ( n37712 , n37708 , n37711 );
not ( n37713 , n37100 );
and ( n37714 , n37713 , n36459 );
xor ( n37715 , n35908 , n37714 );
xor ( n37716 , n37712 , n37715 );
xor ( n37717 , n37091 , n37716 );
xor ( n37718 , n28299 , n31291 );
xor ( n37719 , n37718 , n27989 );
not ( n37720 , n35959 );
and ( n37721 , n37720 , n32148 );
xor ( n37722 , n37719 , n37721 );
xor ( n37723 , n30266 , n31697 );
xor ( n37724 , n37723 , n31309 );
not ( n37725 , n35964 );
and ( n37726 , n37725 , n32157 );
xor ( n37727 , n37724 , n37726 );
xor ( n37728 , n37722 , n37727 );
xor ( n37729 , n28286 , n28617 );
xor ( n37730 , n37729 , n28627 );
not ( n37731 , n35970 );
and ( n37732 , n37731 , n32176 );
xor ( n37733 , n37730 , n37732 );
xor ( n37734 , n37728 , n37733 );
xor ( n37735 , n32505 , n32275 );
xor ( n37736 , n37735 , n31950 );
not ( n37737 , n35976 );
and ( n37738 , n37737 , n32188 );
xor ( n37739 , n37736 , n37738 );
xor ( n37740 , n37734 , n37739 );
not ( n37741 , n35982 );
and ( n37742 , n37741 , n32216 );
xor ( n37743 , n32144 , n37742 );
xor ( n37744 , n37740 , n37743 );
xor ( n37745 , n37717 , n37744 );
not ( n37746 , n37745 );
xor ( n37747 , n27802 , n30758 );
xor ( n37748 , n37747 , n33390 );
xor ( n37749 , n27918 , n30294 );
xor ( n37750 , n37749 , n30306 );
not ( n37751 , n37750 );
xor ( n37752 , n28770 , n30934 );
xor ( n37753 , n37752 , n28533 );
and ( n37754 , n37751 , n37753 );
xor ( n37755 , n37748 , n37754 );
xor ( n37756 , n31108 , n30889 );
xor ( n37757 , n37756 , n30901 );
xor ( n37758 , n32252 , n30691 );
xor ( n37759 , n37758 , n30475 );
not ( n37760 , n37759 );
xor ( n37761 , n28288 , n28617 );
xor ( n37762 , n37761 , n28627 );
and ( n37763 , n37760 , n37762 );
xor ( n37764 , n37757 , n37763 );
xor ( n37765 , n28949 , n27948 );
xor ( n37766 , n37765 , n28702 );
xor ( n37767 , n28736 , n32809 );
xor ( n37768 , n37767 , n31453 );
not ( n37769 , n37768 );
xor ( n37770 , n32741 , n30487 );
xor ( n37771 , n37770 , n30321 );
and ( n37772 , n37769 , n37771 );
xor ( n37773 , n37766 , n37772 );
xor ( n37774 , n37764 , n37773 );
xor ( n37775 , n32828 , n32510 );
xor ( n37776 , n37775 , n29462 );
xor ( n37777 , n30134 , n28392 );
xor ( n37778 , n37777 , n30918 );
not ( n37779 , n37778 );
xor ( n37780 , n31556 , n28866 );
xor ( n37781 , n37780 , n28878 );
and ( n37782 , n37779 , n37781 );
xor ( n37783 , n37776 , n37782 );
xor ( n37784 , n37774 , n37783 );
xor ( n37785 , n29169 , n28185 );
xor ( n37786 , n37785 , n28827 );
not ( n37787 , n37748 );
and ( n37788 , n37787 , n37750 );
xor ( n37789 , n37786 , n37788 );
xor ( n37790 , n37784 , n37789 );
xor ( n37791 , n29495 , n30789 );
xor ( n37792 , n37791 , n30799 );
xor ( n37793 , n29884 , n29740 );
xor ( n37794 , n37793 , n29752 );
not ( n37795 , n37794 );
xor ( n37796 , n27998 , n29677 );
xor ( n37797 , n37796 , n32778 );
and ( n37798 , n37795 , n37797 );
xor ( n37799 , n37792 , n37798 );
xor ( n37800 , n37790 , n37799 );
xor ( n37801 , n37755 , n37800 );
not ( n37802 , n31138 );
and ( n37803 , n37802 , n35014 );
xor ( n37804 , n31135 , n37803 );
xor ( n37805 , n31103 , n37804 );
not ( n37806 , n31168 );
and ( n37807 , n37806 , n35030 );
xor ( n37808 , n31165 , n37807 );
xor ( n37809 , n37805 , n37808 );
not ( n37810 , n31198 );
and ( n37811 , n37810 , n35038 );
xor ( n37812 , n31195 , n37811 );
xor ( n37813 , n37809 , n37812 );
xor ( n37814 , n37813 , n37259 );
xor ( n37815 , n37801 , n37814 );
and ( n37816 , n37746 , n37815 );
xor ( n37817 , n37697 , n37816 );
not ( n12083 , n29614 );
and ( n12084 , n12083 , RI173dfb70_1665);
and ( n12085 , n37817 , n29614 );
or ( n37818 , n12084 , n12085 );
not ( n12086 , RI1754c610_2);
and ( n12087 , n12086 , n37818 );
and ( n12088 , C0 , RI1754c610_2);
or ( n37819 , n12087 , n12088 );
buf ( n37820 , n37819 );
and ( n37821 , RI1754b788_33 , n34844 );
and ( n37822 , RI1754b788_33 , n34847 );
and ( n37823 , RI1754b788_33 , n34850 );
and ( n37824 , RI1754b788_33 , n34852 );
or ( n37825 , n37821 , n37822 , n37823 , n37824 , C0 , C0 , C0 , C0 );
not ( n12089 , n34859 );
and ( n12090 , n12089 , n37825 );
and ( n12091 , RI1754b788_33 , n34859 );
or ( n37826 , n12090 , n12091 );
not ( n12092 , RI19a22f70_2797);
and ( n12093 , n12092 , n37826 );
and ( n12094 , C0 , RI19a22f70_2797);
or ( n37827 , n12093 , n12094 );
not ( n12095 , n27683 );
and ( n12096 , n12095 , RI19aadb70_2470);
and ( n12097 , n37827 , n27683 );
or ( n37828 , n12096 , n12097 );
not ( n12098 , RI1754c610_2);
and ( n12099 , n12098 , n37828 );
and ( n12100 , C0 , RI1754c610_2);
or ( n37829 , n12099 , n12100 );
buf ( n37830 , n37829 );
not ( n37831 , n33254 );
and ( n37832 , n37831 , n33256 );
xor ( n37833 , n33678 , n37832 );
not ( n37834 , n33654 );
and ( n37835 , n37834 , n33235 );
xor ( n37836 , n33651 , n37835 );
not ( n37837 , n33670 );
and ( n37838 , n37837 , n33244 );
xor ( n37839 , n33667 , n37838 );
xor ( n37840 , n37836 , n37839 );
not ( n37841 , n33678 );
and ( n37842 , n37841 , n33254 );
xor ( n37843 , n33675 , n37842 );
xor ( n37844 , n37840 , n37843 );
not ( n37845 , n33686 );
and ( n37846 , n37845 , n33264 );
xor ( n37847 , n33683 , n37846 );
xor ( n37848 , n37844 , n37847 );
xor ( n37849 , n37848 , n35078 );
xor ( n37850 , n37833 , n37849 );
not ( n37851 , n35086 );
and ( n37852 , n37851 , n37588 );
xor ( n37853 , n35083 , n37852 );
not ( n37854 , n35095 );
and ( n37855 , n37854 , n37595 );
xor ( n37856 , n35092 , n37855 );
xor ( n37857 , n37853 , n37856 );
not ( n37858 , n35105 );
and ( n37859 , n37858 , n37603 );
xor ( n37860 , n35102 , n37859 );
xor ( n37861 , n37857 , n37860 );
not ( n37862 , n35115 );
and ( n37863 , n37862 , n37609 );
xor ( n37864 , n35112 , n37863 );
xor ( n37865 , n37861 , n37864 );
not ( n37866 , n35125 );
and ( n37867 , n37866 , n37617 );
xor ( n37868 , n35122 , n37867 );
xor ( n37869 , n37865 , n37868 );
xor ( n37870 , n37850 , n37869 );
not ( n37871 , n33369 );
and ( n37872 , n37871 , n33371 );
xor ( n37873 , n35792 , n37872 );
xor ( n37874 , n37873 , n35804 );
xor ( n37875 , n37874 , n35842 );
not ( n37876 , n37875 );
not ( n37877 , n33497 );
and ( n37878 , n37877 , n33499 );
xor ( n37879 , n36099 , n37878 );
not ( n37880 , n36068 );
and ( n37881 , n37880 , n33456 );
xor ( n37882 , n36065 , n37881 );
not ( n37883 , n36075 );
and ( n37884 , n37883 , n33467 );
xor ( n37885 , n36072 , n37884 );
xor ( n37886 , n37882 , n37885 );
not ( n37887 , n36083 );
and ( n37888 , n37887 , n33477 );
xor ( n37889 , n36080 , n37888 );
xor ( n37890 , n37886 , n37889 );
not ( n37891 , n36091 );
and ( n37892 , n37891 , n33487 );
xor ( n37893 , n36088 , n37892 );
xor ( n37894 , n37890 , n37893 );
not ( n37895 , n36099 );
and ( n37896 , n37895 , n33497 );
xor ( n37897 , n36096 , n37896 );
xor ( n37898 , n37894 , n37897 );
xor ( n37899 , n37879 , n37898 );
not ( n37900 , n31957 );
and ( n37901 , n37900 , n35131 );
xor ( n37902 , n31954 , n37901 );
not ( n37903 , n31993 );
and ( n37904 , n37903 , n35148 );
xor ( n37905 , n31990 , n37904 );
xor ( n37906 , n37902 , n37905 );
not ( n37907 , n32010 );
and ( n37908 , n37907 , n35156 );
xor ( n37909 , n32000 , n37908 );
xor ( n37910 , n37906 , n37909 );
xor ( n37911 , n37910 , n31940 );
not ( n37912 , n32045 );
and ( n37913 , n37912 , n35170 );
xor ( n37914 , n32032 , n37913 );
xor ( n37915 , n37911 , n37914 );
xor ( n37916 , n37899 , n37915 );
and ( n37917 , n37876 , n37916 );
xor ( n37918 , n37870 , n37917 );
not ( n12101 , n29614 );
and ( n12102 , n12101 , RI173f0538_1584);
and ( n12103 , n37918 , n29614 );
or ( n37919 , n12102 , n12103 );
not ( n12104 , RI1754c610_2);
and ( n12105 , n12104 , n37919 );
and ( n12106 , C0 , RI1754c610_2);
or ( n37920 , n12105 , n12106 );
buf ( n37921 , n37920 );
xor ( n37922 , n34634 , n34150 );
xor ( n37923 , n37922 , n34190 );
not ( n37924 , n37499 );
and ( n37925 , n37924 , n34224 );
xor ( n37926 , n33999 , n37925 );
not ( n37927 , n37504 );
and ( n37928 , n37927 , n34229 );
xor ( n37929 , n34008 , n37928 );
xor ( n37930 , n37926 , n37929 );
not ( n37931 , n37510 );
and ( n37932 , n37931 , n34235 );
xor ( n37933 , n34018 , n37932 );
xor ( n37934 , n37930 , n37933 );
not ( n37935 , n37516 );
and ( n37936 , n37935 , n34241 );
xor ( n37937 , n34028 , n37936 );
xor ( n37938 , n37934 , n37937 );
not ( n37939 , n37522 );
and ( n37940 , n37939 , n34247 );
xor ( n37941 , n34038 , n37940 );
xor ( n37942 , n37938 , n37941 );
xor ( n37943 , n37513 , n37942 );
xor ( n37944 , n37943 , n34395 );
not ( n37945 , n37944 );
xor ( n37946 , n29251 , n32120 );
xor ( n37947 , n37946 , n29093 );
xor ( n37948 , n29004 , n29814 );
xor ( n37949 , n37948 , n31131 );
not ( n37950 , n37949 );
and ( n37951 , n37950 , n34427 );
xor ( n37952 , n37947 , n37951 );
xor ( n37953 , n29390 , n32209 );
xor ( n37954 , n37953 , n30389 );
not ( n37955 , n37954 );
xor ( n37956 , n29537 , n30594 );
xor ( n37957 , n37956 , n29224 );
and ( n37958 , n37955 , n37957 );
xor ( n37959 , n34403 , n37958 );
xor ( n37960 , n31741 , n28262 );
xor ( n37961 , n37960 , n28892 );
not ( n37962 , n37961 );
xor ( n37963 , n32134 , n29952 );
xor ( n37964 , n37963 , n29964 );
and ( n37965 , n37962 , n37964 );
xor ( n37966 , n34412 , n37965 );
xor ( n37967 , n37959 , n37966 );
xor ( n37968 , n30380 , n28812 );
xor ( n37969 , n37968 , n29855 );
not ( n37970 , n37969 );
xor ( n37971 , n28562 , n30626 );
xor ( n37972 , n37971 , n29740 );
and ( n37973 , n37970 , n37972 );
xor ( n37974 , n34422 , n37973 );
xor ( n37975 , n37967 , n37974 );
not ( n37976 , n37947 );
and ( n37977 , n37976 , n37949 );
xor ( n37978 , n34432 , n37977 );
xor ( n37979 , n37975 , n37978 );
xor ( n37980 , n31238 , n28727 );
xor ( n37981 , n37980 , n29387 );
not ( n37982 , n37981 );
xor ( n37983 , n32192 , n29793 );
xor ( n37984 , n37983 , n31909 );
and ( n37985 , n37982 , n37984 );
xor ( n37986 , n34442 , n37985 );
xor ( n37987 , n37979 , n37986 );
xor ( n37988 , n37952 , n37987 );
xor ( n37989 , n28988 , n29248 );
xor ( n37990 , n37989 , n29438 );
xor ( n37991 , n31187 , n29544 );
xor ( n37992 , n37991 , n28480 );
not ( n37993 , n37992 );
xor ( n37994 , n30810 , n32382 );
xor ( n37995 , n37994 , n28463 );
and ( n37996 , n37993 , n37995 );
xor ( n37997 , n37990 , n37996 );
xor ( n37998 , n30158 , n28438 );
xor ( n37999 , n37998 , n28450 );
xor ( n38000 , n29171 , n28185 );
xor ( n38001 , n38000 , n28827 );
not ( n38002 , n38001 );
xor ( n38003 , n27709 , n27909 );
xor ( n38004 , n38003 , n27921 );
and ( n38005 , n38002 , n38004 );
xor ( n38006 , n37999 , n38005 );
xor ( n38007 , n37997 , n38006 );
xor ( n38008 , n28297 , n31291 );
xor ( n38009 , n38008 , n27989 );
xor ( n38010 , n28155 , n27738 );
xor ( n38011 , n38010 , n29259 );
not ( n38012 , n38011 );
xor ( n38013 , n29674 , n30842 );
xor ( n38014 , n38013 , n32247 );
and ( n38015 , n38012 , n38014 );
xor ( n38016 , n38009 , n38015 );
xor ( n38017 , n38007 , n38016 );
xor ( n38018 , n31521 , n28107 );
xor ( n38019 , n38018 , n32510 );
xor ( n38020 , n30686 , n30869 );
xor ( n38021 , n38020 , n32894 );
not ( n38022 , n38021 );
xor ( n38023 , n28782 , n32043 );
xor ( n38024 , n38023 , n30946 );
and ( n38025 , n38022 , n38024 );
xor ( n38026 , n38019 , n38025 );
xor ( n38027 , n38017 , n38026 );
xor ( n38028 , n30094 , n29910 );
xor ( n38029 , n38028 , n32167 );
xor ( n38030 , n31554 , n28866 );
xor ( n38031 , n38030 , n28878 );
not ( n38032 , n38031 );
xor ( n38033 , n30756 , n29161 );
xor ( n38034 , n38033 , n28069 );
and ( n38035 , n38032 , n38034 );
xor ( n38036 , n38029 , n38035 );
xor ( n38037 , n38027 , n38036 );
xor ( n38038 , n37988 , n38037 );
and ( n38039 , n37945 , n38038 );
xor ( n38040 , n37923 , n38039 );
not ( n12107 , n29614 );
and ( n12108 , n12107 , RI17459088_1302);
and ( n12109 , n38040 , n29614 );
or ( n38041 , n12108 , n12109 );
not ( n12110 , RI1754c610_2);
and ( n12111 , n12110 , n38041 );
and ( n12112 , C0 , RI1754c610_2);
or ( n38042 , n12111 , n12112 );
buf ( n38043 , n38042 );
xor ( n38044 , n30521 , n29062 );
xor ( n38045 , n38044 , n31613 );
xor ( n38046 , n29412 , n27870 );
xor ( n38047 , n38046 , n28174 );
not ( n38048 , n38047 );
and ( n38049 , n38048 , n38009 );
xor ( n38050 , n38045 , n38049 );
xor ( n38051 , n30331 , n33234 );
xor ( n38052 , n38051 , n31825 );
not ( n38053 , n38052 );
xor ( n38054 , n28803 , n29409 );
xor ( n38055 , n38054 , n29421 );
and ( n38056 , n38053 , n38055 );
xor ( n38057 , n37995 , n38056 );
xor ( n38058 , n31246 , n28727 );
xor ( n38059 , n38058 , n29387 );
not ( n38060 , n38059 );
xor ( n38061 , n30057 , n29105 );
xor ( n38062 , n38061 , n30567 );
and ( n38063 , n38060 , n38062 );
xor ( n38064 , n38004 , n38063 );
xor ( n38065 , n38057 , n38064 );
not ( n38066 , n38045 );
and ( n38067 , n38066 , n38047 );
xor ( n38068 , n38014 , n38067 );
xor ( n38069 , n38065 , n38068 );
xor ( n38070 , n30138 , n28392 );
xor ( n38071 , n38070 , n30918 );
not ( n38072 , n38071 );
xor ( n38073 , n28485 , n31750 );
xor ( n38074 , n38073 , n30043 );
and ( n38075 , n38072 , n38074 );
xor ( n38076 , n38024 , n38075 );
xor ( n38077 , n38069 , n38076 );
xor ( n38078 , n29198 , n28212 );
xor ( n38079 , n38078 , n32459 );
not ( n38080 , n38079 );
xor ( n38081 , n33658 , n31367 );
xor ( n38082 , n38081 , n28800 );
and ( n38083 , n38080 , n38082 );
xor ( n38084 , n38034 , n38083 );
xor ( n38085 , n38077 , n38084 );
xor ( n38086 , n38050 , n38085 );
xor ( n38087 , n27861 , n29601 );
xor ( n38088 , n38087 , n29199 );
not ( n38089 , n30769 );
and ( n38090 , n38089 , n30781 );
xor ( n38091 , n38088 , n38090 );
xor ( n38092 , n31029 , n30053 );
xor ( n38093 , n38092 , n31697 );
not ( n38094 , n30824 );
and ( n38095 , n38094 , n30826 );
xor ( n38096 , n38093 , n38095 );
xor ( n38097 , n38091 , n38096 );
xor ( n38098 , n29190 , n28212 );
xor ( n38099 , n38098 , n32459 );
not ( n38100 , n30843 );
and ( n38101 , n38100 , n30846 );
xor ( n38102 , n38099 , n38101 );
xor ( n38103 , n38097 , n38102 );
xor ( n38104 , n28884 , n30066 );
xor ( n38105 , n38104 , n30007 );
not ( n38106 , n30877 );
and ( n38107 , n38106 , n30902 );
xor ( n38108 , n38105 , n38107 );
xor ( n38109 , n38103 , n38108 );
xor ( n38110 , n31972 , n27897 );
xor ( n38111 , n38110 , n27858 );
not ( n38112 , n30919 );
and ( n38113 , n38112 , n30759 );
xor ( n38114 , n38111 , n38113 );
xor ( n38115 , n38109 , n38114 );
xor ( n38116 , n38086 , n38115 );
xor ( n38117 , n32285 , n31399 );
xor ( n38118 , n38117 , n29561 );
not ( n38119 , n38118 );
xor ( n38120 , n32739 , n30487 );
xor ( n38121 , n38120 , n30321 );
and ( n38122 , n38119 , n38121 );
xor ( n38123 , n31040 , n38122 );
not ( n38124 , n30960 );
xor ( n38125 , n30288 , n28043 );
xor ( n38126 , n38125 , n28055 );
and ( n38127 , n38124 , n38126 );
xor ( n38128 , n30957 , n38127 );
not ( n38129 , n30987 );
xor ( n38130 , n28456 , n29502 );
xor ( n38131 , n38130 , n29628 );
and ( n38132 , n38129 , n38131 );
xor ( n38133 , n30977 , n38132 );
xor ( n38134 , n38128 , n38133 );
not ( n38135 , n31008 );
xor ( n38136 , n27826 , n31683 );
xor ( n38137 , n38136 , n30857 );
and ( n38138 , n38135 , n38137 );
xor ( n38139 , n31005 , n38138 );
xor ( n38140 , n38134 , n38139 );
not ( n38141 , n31040 );
and ( n38142 , n38141 , n38118 );
xor ( n38143 , n31026 , n38142 );
xor ( n38144 , n38140 , n38143 );
not ( n38145 , n31050 );
xor ( n38146 , n30341 , n31152 );
xor ( n38147 , n38146 , n31162 );
and ( n38148 , n38145 , n38147 );
xor ( n38149 , n31047 , n38148 );
xor ( n38150 , n38144 , n38149 );
xor ( n38151 , n38123 , n38150 );
not ( n38152 , n30497 );
and ( n38153 , n38152 , n30499 );
xor ( n38154 , n35471 , n38153 );
not ( n38155 , n30538 );
and ( n38156 , n38155 , n30550 );
xor ( n38157 , n35476 , n38156 );
xor ( n38158 , n38154 , n38157 );
xor ( n38159 , n38158 , n35469 );
not ( n38160 , n30575 );
and ( n38161 , n38160 , n30578 );
xor ( n38162 , n31640 , n38161 );
xor ( n38163 , n38159 , n38162 );
not ( n38164 , n30595 );
and ( n38165 , n38164 , n30597 );
xor ( n38166 , n35490 , n38165 );
xor ( n38167 , n38163 , n38166 );
xor ( n38168 , n38151 , n38167 );
not ( n38169 , n38168 );
not ( n38170 , n32144 );
and ( n38171 , n38170 , n35982 );
xor ( n38172 , n32141 , n38171 );
not ( n38173 , n32153 );
and ( n38174 , n38173 , n37719 );
xor ( n38175 , n32150 , n38174 );
not ( n38176 , n32171 );
and ( n38177 , n38176 , n37724 );
xor ( n38178 , n32168 , n38177 );
xor ( n38179 , n38175 , n38178 );
not ( n38180 , n32183 );
and ( n38181 , n38180 , n37730 );
xor ( n38182 , n32178 , n38181 );
xor ( n38183 , n38179 , n38182 );
not ( n38184 , n32211 );
and ( n38185 , n38184 , n37736 );
xor ( n38186 , n32201 , n38185 );
xor ( n38187 , n38183 , n38186 );
xor ( n38188 , n38187 , n32146 );
xor ( n38189 , n38172 , n38188 );
xor ( n38190 , n38189 , n36195 );
and ( n38191 , n38169 , n38190 );
xor ( n38192 , n38116 , n38191 );
not ( n12113 , n29614 );
and ( n12114 , n12113 , RI17459a60_1299);
and ( n12115 , n38192 , n29614 );
or ( n38193 , n12114 , n12115 );
not ( n12116 , RI1754c610_2);
and ( n12117 , n12116 , n38193 );
and ( n12118 , C0 , RI1754c610_2);
or ( n38194 , n12117 , n12118 );
buf ( n38195 , n38194 );
not ( n38196 , n36775 );
and ( n38197 , n38196 , n34921 );
xor ( n38198 , n37553 , n38197 );
not ( n38199 , n36780 );
and ( n38200 , n38199 , n34930 );
xor ( n38201 , n37558 , n38200 );
xor ( n38202 , n38198 , n38201 );
not ( n38203 , n36786 );
and ( n38204 , n38203 , n34940 );
xor ( n38205 , n37564 , n38204 );
xor ( n38206 , n38202 , n38205 );
not ( n38207 , n36792 );
and ( n38208 , n38207 , n34950 );
xor ( n38209 , n37570 , n38208 );
xor ( n38210 , n38206 , n38209 );
not ( n38211 , n36798 );
and ( n38212 , n38211 , n34960 );
xor ( n38213 , n37576 , n38212 );
xor ( n38214 , n38210 , n38213 );
xor ( n38215 , n36789 , n38214 );
xor ( n38216 , n30615 , n28595 );
xor ( n38217 , n38216 , n28519 );
not ( n38218 , n33082 );
and ( n38219 , n38218 , n33084 );
xor ( n38220 , n38217 , n38219 );
xor ( n38221 , n30373 , n28279 );
xor ( n38222 , n38221 , n28291 );
not ( n38223 , n33091 );
and ( n38224 , n38223 , n33093 );
xor ( n38225 , n38222 , n38224 );
xor ( n38226 , n38220 , n38225 );
xor ( n38227 , n28000 , n29677 );
xor ( n38228 , n38227 , n32778 );
not ( n38229 , n33101 );
and ( n38230 , n38229 , n33103 );
xor ( n38231 , n38228 , n38230 );
xor ( n38232 , n38226 , n38231 );
xor ( n38233 , n30029 , n27921 );
xor ( n38234 , n38233 , n28852 );
not ( n38235 , n33111 );
and ( n38236 , n38235 , n33073 );
xor ( n38237 , n38234 , n38236 );
xor ( n38238 , n38232 , n38237 );
xor ( n38239 , n31920 , n32426 );
xor ( n38240 , n38239 , n31152 );
not ( n38241 , n33117 );
and ( n38242 , n38241 , n33119 );
xor ( n38243 , n38240 , n38242 );
xor ( n38244 , n38238 , n38243 );
xor ( n38245 , n38215 , n38244 );
not ( n38246 , n36020 );
and ( n38247 , n38246 , n37641 );
xor ( n38248 , n32546 , n38247 );
xor ( n38249 , n38248 , n36917 );
xor ( n38250 , n38249 , n36947 );
not ( n38251 , n38250 );
not ( n38252 , n36497 );
and ( n38253 , n38252 , n37391 );
xor ( n38254 , n36494 , n38253 );
xor ( n38255 , n36485 , n38254 );
not ( n38256 , n36507 );
and ( n38257 , n38256 , n37399 );
xor ( n38258 , n36504 , n38257 );
xor ( n38259 , n38255 , n38258 );
not ( n38260 , n36517 );
and ( n38261 , n38260 , n37407 );
xor ( n38262 , n36514 , n38261 );
xor ( n38263 , n38259 , n38262 );
not ( n38264 , n36527 );
and ( n38265 , n38264 , n37415 );
xor ( n38266 , n36524 , n38265 );
xor ( n38267 , n38263 , n38266 );
xor ( n38268 , n37420 , n38267 );
not ( n38269 , n36541 );
and ( n38270 , n38269 , n34687 );
xor ( n38271 , n36538 , n38270 );
xor ( n38272 , n36717 , n38271 );
not ( n38273 , n36549 );
and ( n38274 , n38273 , n34697 );
xor ( n38275 , n36546 , n38274 );
xor ( n38276 , n38272 , n38275 );
not ( n38277 , n36557 );
and ( n38278 , n38277 , n34707 );
xor ( n38279 , n36554 , n38278 );
xor ( n38280 , n38276 , n38279 );
not ( n38281 , n36565 );
and ( n38282 , n38281 , n34717 );
xor ( n38283 , n36562 , n38282 );
xor ( n38284 , n38280 , n38283 );
xor ( n38285 , n38268 , n38284 );
and ( n38286 , n38251 , n38285 );
xor ( n38287 , n38245 , n38286 );
not ( n12119 , n29614 );
and ( n12120 , n12119 , RI17399c70_2006);
and ( n12121 , n38287 , n29614 );
or ( n38288 , n12120 , n12121 );
not ( n12122 , RI1754c610_2);
and ( n12123 , n12122 , n38288 );
and ( n12124 , C0 , RI1754c610_2);
or ( n38289 , n12123 , n12124 );
buf ( n38290 , n38289 );
not ( n12125 , n27683 );
and ( n12126 , n12125 , RI19acc5c0_2236);
and ( n12127 , RI19a88208_2737 , n27683 );
or ( n38291 , n12126 , n12127 );
not ( n12128 , RI1754c610_2);
and ( n12129 , n12128 , n38291 );
and ( n12130 , C0 , RI1754c610_2);
or ( n38292 , n12129 , n12130 );
buf ( n38293 , n38292 );
xor ( n38294 , n29570 , n32611 );
xor ( n38295 , n38294 , n29161 );
xor ( n38296 , n30664 , n28969 );
xor ( n38297 , n38296 , n28741 );
not ( n38298 , n38297 );
xor ( n38299 , n29830 , n32140 );
xor ( n38300 , n38299 , n31874 );
and ( n38301 , n38298 , n38300 );
xor ( n38302 , n38295 , n38301 );
xor ( n38303 , n33660 , n31367 );
xor ( n38304 , n38303 , n28800 );
not ( n38305 , n38295 );
and ( n38306 , n38305 , n38297 );
xor ( n38307 , n38304 , n38306 );
xor ( n38308 , n30820 , n28463 );
xor ( n38309 , n38308 , n27752 );
xor ( n38310 , n30386 , n28812 );
xor ( n38311 , n38310 , n29855 );
not ( n38312 , n38311 );
xor ( n38313 , n29585 , n29767 );
xor ( n38314 , n38313 , n30510 );
and ( n38315 , n38312 , n38314 );
xor ( n38316 , n38309 , n38315 );
xor ( n38317 , n38307 , n38316 );
xor ( n38318 , n28475 , n29224 );
xor ( n38319 , n38318 , n29235 );
xor ( n38320 , n28490 , n31750 );
xor ( n38321 , n38320 , n30043 );
not ( n38322 , n38321 );
xor ( n38323 , n32274 , n27975 );
xor ( n38324 , n38323 , n29346 );
and ( n38325 , n38322 , n38324 );
xor ( n38326 , n38319 , n38325 );
xor ( n38327 , n38317 , n38326 );
xor ( n38328 , n28899 , n30007 );
xor ( n38329 , n38328 , n30017 );
xor ( n38330 , n29329 , n31226 );
xor ( n38331 , n38330 , n31516 );
not ( n38332 , n38331 );
xor ( n38333 , n30474 , n32894 );
xor ( n38334 , n38333 , n32991 );
and ( n38335 , n38332 , n38334 );
xor ( n38336 , n38329 , n38335 );
xor ( n38337 , n38327 , n38336 );
xor ( n38338 , n31158 , n27779 );
xor ( n38339 , n38338 , n27791 );
xor ( n38340 , n31494 , n28715 );
xor ( n38341 , n38340 , n28727 );
not ( n38342 , n38341 );
xor ( n38343 , n29489 , n28450 );
xor ( n38344 , n38343 , n30789 );
and ( n38345 , n38342 , n38344 );
xor ( n38346 , n38339 , n38345 );
xor ( n38347 , n38337 , n38346 );
xor ( n38348 , n38302 , n38347 );
xor ( n38349 , n38348 , n34300 );
xor ( n38350 , n32757 , n37186 );
xor ( n38351 , n38350 , n37203 );
not ( n38352 , n38351 );
not ( n38353 , n33833 );
and ( n38354 , n38353 , n34067 );
xor ( n38355 , n33830 , n38354 );
not ( n38356 , n33842 );
and ( n38357 , n38356 , n34054 );
xor ( n38358 , n33839 , n38357 );
not ( n38359 , n33851 );
and ( n38360 , n38359 , n34061 );
xor ( n38361 , n33848 , n38360 );
xor ( n38362 , n38358 , n38361 );
xor ( n38363 , n38362 , n33835 );
not ( n38364 , n33867 );
and ( n38365 , n38364 , n34073 );
xor ( n38366 , n33864 , n38365 );
xor ( n38367 , n38363 , n38366 );
not ( n38368 , n33877 );
and ( n38369 , n38368 , n34081 );
xor ( n38370 , n33874 , n38369 );
xor ( n38371 , n38367 , n38370 );
xor ( n38372 , n38355 , n38371 );
xor ( n38373 , n38372 , n36431 );
and ( n38374 , n38352 , n38373 );
xor ( n38375 , n38349 , n38374 );
not ( n12131 , n29614 );
and ( n12132 , n12131 , RI174b0ce8_874);
and ( n12133 , n38375 , n29614 );
or ( n38376 , n12132 , n12133 );
not ( n12134 , RI1754c610_2);
and ( n12135 , n12134 , n38376 );
and ( n12136 , C0 , RI1754c610_2);
or ( n38377 , n12135 , n12136 );
buf ( n38378 , n38377 );
not ( n38379 , n35692 );
and ( n38380 , n38379 , n35694 );
xor ( n38381 , n35830 , n38380 );
xor ( n38382 , n38381 , n35842 );
not ( n38383 , n37135 );
and ( n38384 , n38383 , n35713 );
xor ( n38385 , n37132 , n38384 );
not ( n38386 , n37142 );
and ( n38387 , n38386 , n35722 );
xor ( n38388 , n37139 , n38387 );
xor ( n38389 , n38385 , n38388 );
not ( n38390 , n37150 );
and ( n38391 , n38390 , n35732 );
xor ( n38392 , n37147 , n38391 );
xor ( n38393 , n38389 , n38392 );
not ( n38394 , n37158 );
and ( n38395 , n38394 , n35742 );
xor ( n38396 , n37155 , n38395 );
xor ( n38397 , n38393 , n38396 );
not ( n38398 , n37166 );
and ( n38399 , n38398 , n35752 );
xor ( n38400 , n37163 , n38399 );
xor ( n38401 , n38397 , n38400 );
xor ( n38402 , n38382 , n38401 );
not ( n38403 , n35358 );
and ( n38404 , n38403 , n36992 );
xor ( n38405 , n35355 , n38404 );
xor ( n38406 , n38405 , n35361 );
xor ( n38407 , n30012 , n28647 );
xor ( n38408 , n38407 , n28659 );
not ( n38409 , n38408 );
xor ( n38410 , n30839 , n27833 );
xor ( n38411 , n38410 , n27844 );
and ( n38412 , n38409 , n38411 );
xor ( n38413 , n37006 , n38412 );
xor ( n38414 , n28334 , n31076 );
xor ( n38415 , n38414 , n32091 );
not ( n38416 , n38415 );
xor ( n38417 , n31791 , n29148 );
xor ( n38418 , n38417 , n32800 );
and ( n38419 , n38416 , n38418 );
xor ( n38420 , n37015 , n38419 );
xor ( n38421 , n38413 , n38420 );
xor ( n38422 , n30410 , n30901 );
xor ( n38423 , n38422 , n31475 );
not ( n38424 , n38423 );
xor ( n38425 , n29303 , n31487 );
xor ( n38426 , n38425 , n31497 );
and ( n38427 , n38424 , n38426 );
xor ( n38428 , n37025 , n38427 );
xor ( n38429 , n38421 , n38428 );
xor ( n38430 , n28722 , n31279 );
xor ( n38431 , n38430 , n33665 );
not ( n38432 , n38431 );
xor ( n38433 , n28171 , n29199 );
xor ( n38434 , n38433 , n29211 );
and ( n38435 , n38432 , n38434 );
xor ( n38436 , n37035 , n38435 );
xor ( n38437 , n38429 , n38436 );
xor ( n38438 , n29254 , n32120 );
xor ( n38439 , n38438 , n29093 );
not ( n38440 , n38439 );
xor ( n38441 , n30040 , n28892 );
xor ( n38442 , n38441 , n28904 );
and ( n38443 , n38440 , n38442 );
xor ( n38444 , n37045 , n38443 );
xor ( n38445 , n38437 , n38444 );
xor ( n38446 , n38406 , n38445 );
not ( n38447 , n38446 );
xor ( n38448 , n35056 , n33223 );
xor ( n38449 , n38448 , n33282 );
and ( n38450 , n38447 , n38449 );
xor ( n38451 , n38402 , n38450 );
not ( n12137 , n29614 );
and ( n12138 , n12137 , RI173a9288_1931);
and ( n12139 , n38451 , n29614 );
or ( n38452 , n12138 , n12139 );
not ( n12140 , RI1754c610_2);
and ( n12141 , n12140 , n38452 );
and ( n12142 , C0 , RI1754c610_2);
or ( n38453 , n12141 , n12142 );
buf ( n38454 , n38453 );
not ( n12143 , n27683 );
and ( n12144 , n12143 , RI19ac5978_2287);
and ( n12145 , RI19ace618_2222 , n27683 );
or ( n38455 , n12144 , n12145 );
not ( n12146 , RI1754c610_2);
and ( n12147 , n12146 , n38455 );
and ( n12148 , C0 , RI1754c610_2);
or ( n38456 , n12147 , n12148 );
buf ( n38457 , n38456 );
and ( n38458 , RI1754b878_31 , n34844 );
and ( n38459 , RI1754b878_31 , n34847 );
and ( n38460 , RI1754b878_31 , n34850 );
and ( n38461 , RI1754b878_31 , n34852 );
or ( n38462 , n38458 , n38459 , n38460 , n38461 , C0 , C0 , C0 , C0 );
not ( n12149 , n34859 );
and ( n12150 , n12149 , n38462 );
and ( n12151 , RI1754b878_31 , n34859 );
or ( n38463 , n12150 , n12151 );
not ( n12152 , RI19a22f70_2797);
and ( n12153 , n12152 , n38463 );
and ( n12154 , C0 , RI19a22f70_2797);
or ( n38464 , n12153 , n12154 );
not ( n12155 , n27683 );
and ( n12156 , n12155 , RI19aaa858_2492);
and ( n12157 , n38464 , n27683 );
or ( n38465 , n12156 , n12157 );
not ( n12158 , RI1754c610_2);
and ( n12159 , n12158 , n38465 );
and ( n12160 , C0 , RI1754c610_2);
or ( n38466 , n12159 , n12160 );
buf ( n38467 , n38466 );
xor ( n38468 , n37680 , n37579 );
xor ( n38469 , n30472 , n32894 );
xor ( n38470 , n38469 , n32991 );
not ( n38471 , n38470 );
and ( n38472 , n38471 , n38217 );
xor ( n38473 , n33087 , n38472 );
xor ( n38474 , n31451 , n29011 );
xor ( n38475 , n38474 , n27964 );
not ( n38476 , n38475 );
and ( n38477 , n38476 , n38222 );
xor ( n38478 , n33096 , n38477 );
xor ( n38479 , n38473 , n38478 );
xor ( n38480 , n27882 , n29387 );
xor ( n38481 , n38480 , n29399 );
not ( n38482 , n38481 );
and ( n38483 , n38482 , n38228 );
xor ( n38484 , n33106 , n38483 );
xor ( n38485 , n38479 , n38484 );
not ( n38486 , n33078 );
and ( n38487 , n38486 , n38234 );
xor ( n38488 , n33075 , n38487 );
xor ( n38489 , n38485 , n38488 );
xor ( n38490 , n31633 , n30986 );
xor ( n38491 , n38490 , n31794 );
not ( n38492 , n38491 );
and ( n38493 , n38492 , n38240 );
xor ( n38494 , n33122 , n38493 );
xor ( n38495 , n38489 , n38494 );
xor ( n38496 , n38468 , n38495 );
not ( n38497 , n34128 );
and ( n38498 , n38497 , n34191 );
xor ( n38499 , n38496 , n38498 );
not ( n12161 , n29614 );
and ( n12162 , n12161 , RI17341728_2122);
and ( n12163 , n38499 , n29614 );
or ( n38500 , n12162 , n12163 );
not ( n12164 , RI1754c610_2);
and ( n12165 , n12164 , n38500 );
and ( n12166 , C0 , RI1754c610_2);
or ( n38501 , n12165 , n12166 );
buf ( n38502 , n38501 );
xor ( n38503 , n37265 , n36158 );
not ( n38504 , n30493 );
and ( n38505 , n38504 , n35466 );
xor ( n38506 , n30490 , n38505 );
xor ( n38507 , n38503 , n38506 );
xor ( n38508 , n38507 , n31642 );
not ( n38509 , n31661 );
and ( n38510 , n38509 , n35490 );
xor ( n38511 , n30601 , n38510 );
xor ( n38512 , n38508 , n38511 );
xor ( n38513 , n35487 , n38512 );
not ( n38514 , n31668 );
and ( n38515 , n38514 , n33701 );
xor ( n38516 , n30630 , n38515 );
not ( n38517 , n31684 );
and ( n38518 , n38517 , n33706 );
xor ( n38519 , n30669 , n38518 );
xor ( n38520 , n38516 , n38519 );
not ( n38521 , n31698 );
and ( n38522 , n38521 , n33712 );
xor ( n38523 , n30693 , n38522 );
xor ( n38524 , n38520 , n38523 );
not ( n38525 , n31716 );
and ( n38526 , n38525 , n33718 );
xor ( n38527 , n30725 , n38526 );
xor ( n38528 , n38524 , n38527 );
not ( n38529 , n31722 );
and ( n38530 , n38529 , n33724 );
xor ( n38531 , n30738 , n38530 );
xor ( n38532 , n38528 , n38531 );
xor ( n38533 , n38513 , n38532 );
xor ( n38534 , n32308 , n36003 );
not ( n38535 , n32880 );
and ( n38536 , n38535 , n32882 );
xor ( n38537 , n32673 , n38536 );
not ( n38538 , n32895 );
and ( n38539 , n38538 , n32875 );
xor ( n38540 , n32682 , n38539 );
xor ( n38541 , n38537 , n38540 );
not ( n38542 , n32901 );
and ( n38543 , n38542 , n32903 );
xor ( n38544 , n32692 , n38543 );
xor ( n38545 , n38541 , n38544 );
not ( n38546 , n32909 );
and ( n38547 , n38546 , n32911 );
xor ( n38548 , n32702 , n38547 );
xor ( n38549 , n38545 , n38548 );
not ( n38550 , n32917 );
and ( n38551 , n38550 , n32919 );
xor ( n38552 , n32712 , n38551 );
xor ( n38553 , n38549 , n38552 );
xor ( n38554 , n38534 , n38553 );
not ( n38555 , n38554 );
not ( n38556 , n29450 );
and ( n38557 , n38556 , n29475 );
xor ( n38558 , n28596 , n38557 );
not ( n38559 , n28596 );
and ( n38560 , n38559 , n29450 );
xor ( n38561 , n28570 , n38560 );
xor ( n38562 , n38561 , n28523 );
not ( n38563 , n28685 );
and ( n38564 , n38563 , n29521 );
xor ( n38565 , n28660 , n38564 );
xor ( n38566 , n38562 , n38565 );
not ( n38567 , n28743 );
and ( n38568 , n38567 , n29574 );
xor ( n38569 , n28728 , n38568 );
xor ( n38570 , n38566 , n38569 );
not ( n38571 , n28813 );
and ( n38572 , n38571 , n29603 );
xor ( n38573 , n28787 , n38572 );
xor ( n38574 , n38570 , n38573 );
xor ( n38575 , n38558 , n38574 );
not ( n38576 , n28879 );
and ( n38577 , n38576 , n31325 );
xor ( n38578 , n28853 , n38577 );
not ( n38579 , n28934 );
and ( n38580 , n38579 , n31337 );
xor ( n38581 , n28930 , n38580 );
xor ( n38582 , n38578 , n38581 );
not ( n38583 , n28996 );
and ( n38584 , n38583 , n31345 );
xor ( n38585 , n28971 , n38584 );
xor ( n38586 , n38582 , n38585 );
not ( n38587 , n29063 );
and ( n38588 , n38587 , n31355 );
xor ( n38589 , n29038 , n38588 );
xor ( n38590 , n38586 , n38589 );
not ( n38591 , n29106 );
and ( n38592 , n38591 , n31374 );
xor ( n38593 , n29081 , n38592 );
xor ( n38594 , n38590 , n38593 );
xor ( n38595 , n38575 , n38594 );
and ( n38596 , n38555 , n38595 );
xor ( n38597 , n38533 , n38596 );
not ( n12167 , n29614 );
and ( n12168 , n12167 , RI174ac170_897);
and ( n12169 , n38597 , n29614 );
or ( n38598 , n12168 , n12169 );
not ( n12170 , RI1754c610_2);
and ( n12171 , n12170 , n38598 );
and ( n12172 , C0 , RI1754c610_2);
or ( n38599 , n12171 , n12172 );
buf ( n38600 , n38599 );
xor ( n38601 , n36729 , n30247 );
xor ( n38602 , n38601 , n30461 );
xor ( n38603 , n35900 , n36463 );
xor ( n38604 , n38603 , n32220 );
not ( n38605 , n38604 );
xor ( n38606 , n29042 , n28027 );
xor ( n38607 , n38606 , n29827 );
not ( n38608 , n38607 );
xor ( n38609 , n30994 , n32256 );
xor ( n38610 , n38609 , n32734 );
and ( n38611 , n38608 , n38610 );
xor ( n38612 , n38344 , n38611 );
not ( n38613 , n38314 );
xor ( n38614 , n30297 , n28055 );
xor ( n38615 , n38614 , n28224 );
and ( n38616 , n38613 , n38615 );
xor ( n38617 , n38311 , n38616 );
xor ( n38618 , n38302 , n38617 );
not ( n38619 , n38324 );
xor ( n38620 , n31865 , n29964 );
xor ( n38621 , n38620 , n32382 );
and ( n38622 , n38619 , n38621 );
xor ( n38623 , n38321 , n38622 );
xor ( n38624 , n38618 , n38623 );
not ( n38625 , n38334 );
xor ( n38626 , n29441 , n30030 );
xor ( n38627 , n38626 , n30972 );
and ( n38628 , n38625 , n38627 );
xor ( n38629 , n38331 , n38628 );
xor ( n38630 , n38624 , n38629 );
not ( n38631 , n38344 );
and ( n38632 , n38631 , n38607 );
xor ( n38633 , n38341 , n38632 );
xor ( n38634 , n38630 , n38633 );
xor ( n38635 , n38612 , n38634 );
not ( n38636 , n34270 );
and ( n38637 , n38636 , n31409 );
xor ( n38638 , n34267 , n38637 );
xor ( n38639 , n38638 , n37208 );
xor ( n38640 , n38639 , n34265 );
not ( n38641 , n34289 );
and ( n38642 , n38641 , n31444 );
xor ( n38643 , n34286 , n38642 );
xor ( n38644 , n38640 , n38643 );
not ( n38645 , n34297 );
and ( n38646 , n38645 , n31498 );
xor ( n38647 , n34294 , n38646 );
xor ( n38648 , n38644 , n38647 );
xor ( n38649 , n38635 , n38648 );
and ( n38650 , n38605 , n38649 );
xor ( n38651 , n38602 , n38650 );
not ( n12173 , n29614 );
and ( n12174 , n12173 , RI17488338_1072);
and ( n12175 , n38651 , n29614 );
or ( n38652 , n12174 , n12175 );
not ( n12176 , RI1754c610_2);
and ( n12177 , n12176 , n38652 );
and ( n12178 , C0 , RI1754c610_2);
or ( n38653 , n12177 , n12178 );
buf ( n38654 , n38653 );
not ( n12179 , n27683 );
and ( n12180 , n12179 , RI19aca040_2255);
and ( n12181 , RI19a852b0_2758 , n27683 );
or ( n38655 , n12180 , n12181 );
not ( n12182 , RI1754c610_2);
and ( n12183 , n12182 , n38655 );
and ( n12184 , C0 , RI1754c610_2);
or ( n38656 , n12183 , n12184 );
buf ( n38657 , n38656 );
not ( n38658 , n29657 );
and ( n38659 , n38658 , n36342 );
xor ( n38660 , n29643 , n38659 );
not ( n38661 , n36347 );
and ( n38662 , n38661 , n36349 );
xor ( n38663 , n29695 , n38662 );
xor ( n38664 , n38660 , n38663 );
not ( n38665 , n36355 );
and ( n38666 , n38665 , n36357 );
xor ( n38667 , n29725 , n38666 );
xor ( n38668 , n38664 , n38667 );
not ( n38669 , n36363 );
and ( n38670 , n38669 , n36365 );
xor ( n38671 , n29794 , n38670 );
xor ( n38672 , n38668 , n38671 );
not ( n38673 , n36371 );
and ( n38674 , n38673 , n36373 );
xor ( n38675 , n29840 , n38674 );
xor ( n38676 , n38672 , n38675 );
xor ( n38677 , n36368 , n38676 );
xor ( n38678 , n38677 , n28111 );
not ( n38679 , n36914 );
and ( n38680 , n38679 , n37647 );
xor ( n38681 , n32557 , n38680 );
xor ( n38682 , n38681 , n36917 );
xor ( n38683 , n38682 , n36947 );
not ( n38684 , n38683 );
xor ( n38685 , n30816 , n28463 );
xor ( n38686 , n38685 , n27752 );
not ( n38687 , n35229 );
and ( n38688 , n38687 , n35231 );
xor ( n38689 , n38686 , n38688 );
xor ( n38690 , n28106 , n31462 );
xor ( n38691 , n38690 , n32275 );
not ( n38692 , n38686 );
and ( n38693 , n38692 , n35229 );
xor ( n38694 , n38691 , n38693 );
xor ( n38695 , n29703 , n28947 );
xor ( n38696 , n38695 , n28956 );
not ( n38697 , n38696 );
and ( n38698 , n38697 , n35238 );
xor ( n38699 , n35225 , n38698 );
xor ( n38700 , n38694 , n38699 );
xor ( n38701 , n28877 , n30218 );
xor ( n38702 , n38701 , n27807 );
xor ( n38703 , n27743 , n29628 );
xor ( n38704 , n38703 , n29639 );
not ( n38705 , n38704 );
and ( n38706 , n38705 , n35244 );
xor ( n38707 , n38702 , n38706 );
xor ( n38708 , n38700 , n38707 );
xor ( n38709 , n33233 , n29364 );
xor ( n38710 , n38709 , n29375 );
xor ( n38711 , n29126 , n32398 );
xor ( n38712 , n38711 , n30364 );
not ( n38713 , n38712 );
and ( n38714 , n38713 , n35254 );
xor ( n38715 , n38710 , n38714 );
xor ( n38716 , n38708 , n38715 );
xor ( n38717 , n28147 , n27726 );
xor ( n38718 , n38717 , n27738 );
xor ( n38719 , n32024 , n31874 );
xor ( n38720 , n38719 , n30813 );
not ( n38721 , n38720 );
and ( n38722 , n38721 , n35264 );
xor ( n38723 , n38718 , n38722 );
xor ( n38724 , n38716 , n38723 );
xor ( n38725 , n38689 , n38724 );
xor ( n38726 , n38725 , n29425 );
and ( n38727 , n38684 , n38726 );
xor ( n38728 , n38678 , n38727 );
not ( n12185 , n29614 );
and ( n12186 , n12185 , RI1749aa88_982);
and ( n12187 , n38728 , n29614 );
or ( n38729 , n12186 , n12187 );
not ( n12188 , RI1754c610_2);
and ( n12189 , n12188 , n38729 );
and ( n12190 , C0 , RI1754c610_2);
or ( n38730 , n12189 , n12190 );
buf ( n38731 , n38730 );
not ( n12191 , n27683 );
and ( n12192 , n12191 , RI19abc6c0_2364);
and ( n12193 , RI19ac4dc0_2293 , n27683 );
or ( n38732 , n12192 , n12193 );
not ( n12194 , RI1754c610_2);
and ( n12195 , n12194 , n38732 );
and ( n12196 , C0 , RI1754c610_2);
or ( n38733 , n12195 , n12196 );
buf ( n38734 , n38733 );
not ( n12197 , n27683 );
and ( n12198 , n12197 , RI19a92e10_2662);
and ( n12199 , RI19a9d1a8_2590 , n27683 );
or ( n38735 , n12198 , n12199 );
not ( n12200 , RI1754c610_2);
and ( n12201 , n12200 , n38735 );
and ( n12202 , C0 , RI1754c610_2);
or ( n38736 , n12201 , n12202 );
buf ( n38737 , n38736 );
buf ( n38738 , RI174c9108_785);
not ( n38739 , n33765 );
xor ( n38740 , n32028 , n31874 );
xor ( n38741 , n38740 , n30813 );
and ( n38742 , n38739 , n38741 );
xor ( n38743 , n33762 , n38742 );
xor ( n38744 , n38743 , n33778 );
xor ( n38745 , n28668 , n28236 );
xor ( n38746 , n38745 , n29711 );
xor ( n38747 , n31747 , n28262 );
xor ( n38748 , n38747 , n28892 );
not ( n38749 , n38748 );
xor ( n38750 , n30163 , n28438 );
xor ( n38751 , n38750 , n28450 );
and ( n38752 , n38749 , n38751 );
xor ( n38753 , n38746 , n38752 );
xor ( n38754 , n32243 , n27844 );
xor ( n38755 , n38754 , n30691 );
xor ( n38756 , n28276 , n30443 );
xor ( n38757 , n38756 , n28617 );
not ( n38758 , n38757 );
xor ( n38759 , n32458 , n28583 );
xor ( n38760 , n38759 , n28595 );
and ( n38761 , n38758 , n38760 );
xor ( n38762 , n38755 , n38761 );
xor ( n38763 , n38753 , n38762 );
xor ( n38764 , n28654 , n30283 );
xor ( n38765 , n38764 , n31089 );
xor ( n38766 , n30329 , n33234 );
xor ( n38767 , n38766 , n31825 );
not ( n38768 , n38767 );
xor ( n38769 , n27725 , n28533 );
xor ( n38770 , n38769 , n28543 );
and ( n38771 , n38768 , n38770 );
xor ( n38772 , n38765 , n38771 );
xor ( n38773 , n38763 , n38772 );
xor ( n38774 , n29762 , n33898 );
xor ( n38775 , n38774 , n29051 );
xor ( n38776 , n32380 , n29490 );
xor ( n38777 , n38776 , n29502 );
not ( n38778 , n38777 );
xor ( n38779 , n29386 , n33665 );
xor ( n38780 , n38779 , n32209 );
and ( n38781 , n38778 , n38780 );
xor ( n38782 , n38775 , n38781 );
xor ( n38783 , n38773 , n38782 );
xor ( n38784 , n29230 , n30780 );
xor ( n38785 , n38784 , n28043 );
xor ( n38786 , n30969 , n28852 );
xor ( n38787 , n38786 , n29873 );
not ( n38788 , n38787 );
xor ( n38789 , n31682 , n28001 );
xor ( n38790 , n38789 , n30114 );
and ( n38791 , n38788 , n38790 );
xor ( n38792 , n38785 , n38791 );
xor ( n38793 , n38783 , n38792 );
xor ( n38794 , n38744 , n38793 );
not ( n38795 , n34337 );
and ( n38796 , n38795 , n31600 );
xor ( n38797 , n34334 , n38796 );
xor ( n38798 , n38797 , n34340 );
not ( n38799 , n38691 );
and ( n38800 , n38799 , n38686 );
xor ( n38801 , n35234 , n38800 );
not ( n38802 , n35225 );
and ( n38803 , n38802 , n38696 );
xor ( n38804 , n35222 , n38803 );
xor ( n38805 , n38801 , n38804 );
not ( n38806 , n38702 );
and ( n38807 , n38806 , n38704 );
xor ( n38808 , n35249 , n38807 );
xor ( n38809 , n38805 , n38808 );
not ( n38810 , n38710 );
and ( n38811 , n38810 , n38712 );
xor ( n38812 , n35259 , n38811 );
xor ( n38813 , n38809 , n38812 );
not ( n38814 , n38718 );
and ( n38815 , n38814 , n38720 );
xor ( n38816 , n35269 , n38815 );
xor ( n38817 , n38813 , n38816 );
xor ( n38818 , n38798 , n38817 );
not ( n38819 , n38818 );
xor ( n38820 , n37535 , n34918 );
xor ( n38821 , n38820 , n34968 );
and ( n38822 , n38819 , n38821 );
xor ( n38823 , n38794 , n38822 );
not ( n12203 , n29614 );
and ( n12204 , n12203 , RI1752d698_625);
and ( n12205 , n38823 , n29614 );
or ( n38824 , n12204 , n12205 );
not ( n12206 , RI1754c610_2);
and ( n12207 , n12206 , n38824 );
and ( n12208 , C0 , RI1754c610_2);
or ( n38825 , n12207 , n12208 );
buf ( n38826 , n38825 );
buf ( n38827 , RI17493e40_1015);
buf ( n38828 , RI174693c0_1223);
xor ( n38829 , n38266 , n36530 );
xor ( n38830 , n38829 , n36568 );
not ( n38831 , n35022 );
and ( n38832 , n38831 , n31116 );
xor ( n38833 , n31101 , n38832 );
xor ( n38834 , n38833 , n35052 );
xor ( n38835 , n38834 , n35069 );
not ( n38836 , n38835 );
xor ( n38837 , n32821 , n37203 );
xor ( n38838 , n38837 , n34150 );
and ( n38839 , n38836 , n38838 );
xor ( n38840 , n38830 , n38839 );
not ( n12209 , n29614 );
and ( n12210 , n12209 , RI1749cea0_971);
and ( n12211 , n38840 , n29614 );
or ( n38841 , n12210 , n12211 );
not ( n12212 , RI1754c610_2);
and ( n12213 , n12212 , n38841 );
and ( n12214 , C0 , RI1754c610_2);
or ( n38842 , n12213 , n12214 );
buf ( n38843 , n38842 );
xor ( n38844 , n31883 , n36401 );
xor ( n38845 , n38844 , n33453 );
xor ( n38846 , n27890 , n29399 );
xor ( n38847 , n38846 , n29655 );
not ( n38848 , n38304 );
and ( n38849 , n38848 , n38295 );
xor ( n38850 , n38847 , n38849 );
xor ( n38851 , n31552 , n28866 );
xor ( n38852 , n38851 , n28878 );
not ( n38853 , n38309 );
and ( n38854 , n38853 , n38311 );
xor ( n38855 , n38852 , n38854 );
xor ( n38856 , n38850 , n38855 );
xor ( n38857 , n27731 , n28543 );
xor ( n38858 , n38857 , n32120 );
not ( n38859 , n38319 );
and ( n38860 , n38859 , n38321 );
xor ( n38861 , n38858 , n38860 );
xor ( n38862 , n38856 , n38861 );
xor ( n38863 , n28373 , n31909 );
xor ( n38864 , n38863 , n31921 );
not ( n38865 , n38329 );
and ( n38866 , n38865 , n38331 );
xor ( n38867 , n38864 , n38866 );
xor ( n38868 , n38862 , n38867 );
not ( n38869 , n38339 );
and ( n38870 , n38869 , n38341 );
xor ( n38871 , n38610 , n38870 );
xor ( n38872 , n38868 , n38871 );
xor ( n38873 , n38336 , n38872 );
not ( n38874 , n31424 );
and ( n38875 , n38874 , n34267 );
xor ( n38876 , n31411 , n38875 );
not ( n38877 , n31433 );
and ( n38878 , n38877 , n34274 );
xor ( n38879 , n31430 , n38878 );
xor ( n38880 , n38876 , n38879 );
xor ( n38881 , n38880 , n31406 );
xor ( n38882 , n38881 , n36381 );
not ( n38883 , n31503 );
and ( n38884 , n38883 , n34294 );
xor ( n38885 , n31500 , n38884 );
xor ( n38886 , n38882 , n38885 );
xor ( n38887 , n38873 , n38886 );
not ( n38888 , n38887 );
xor ( n38889 , n34220 , n36287 );
xor ( n38890 , n38889 , n37526 );
and ( n38891 , n38888 , n38890 );
xor ( n38892 , n38845 , n38891 );
not ( n12215 , n29614 );
and ( n12216 , n12215 , RI173ebd08_1606);
and ( n12217 , n38892 , n29614 );
or ( n38893 , n12216 , n12217 );
not ( n12218 , RI1754c610_2);
and ( n12219 , n12218 , n38893 );
and ( n12220 , C0 , RI1754c610_2);
or ( n38894 , n12219 , n12220 );
buf ( n38895 , n38894 );
xor ( n38896 , n35513 , n38532 );
xor ( n38897 , n32117 , n28137 );
xor ( n38898 , n38897 , n28493 );
xor ( n38899 , n32139 , n29952 );
xor ( n38900 , n38899 , n29964 );
not ( n38901 , n38900 );
and ( n38902 , n38901 , n33731 );
xor ( n38903 , n38898 , n38902 );
xor ( n38904 , n27933 , n30364 );
xor ( n38905 , n38904 , n30374 );
xor ( n38906 , n28173 , n29199 );
xor ( n38907 , n38906 , n29211 );
not ( n38908 , n38907 );
and ( n38909 , n38908 , n33740 );
xor ( n38910 , n38905 , n38909 );
xor ( n38911 , n38903 , n38910 );
xor ( n38912 , n31472 , n33198 );
xor ( n38913 , n38912 , n31714 );
xor ( n38914 , n29627 , n30799 );
xor ( n38915 , n38914 , n28148 );
not ( n38916 , n38915 );
and ( n38917 , n38916 , n33750 );
xor ( n38918 , n38913 , n38917 );
xor ( n38919 , n38911 , n38918 );
xor ( n38920 , n28417 , n31247 );
xor ( n38921 , n38920 , n27885 );
not ( n38922 , n38921 );
and ( n38923 , n38922 , n33760 );
xor ( n38924 , n38741 , n38923 );
xor ( n38925 , n38919 , n38924 );
xor ( n38926 , n28040 , n29449 );
xor ( n38927 , n38926 , n29694 );
xor ( n38928 , n30536 , n29752 );
xor ( n38929 , n38928 , n27833 );
not ( n38930 , n38929 );
and ( n38931 , n38930 , n33770 );
xor ( n38932 , n38927 , n38931 );
xor ( n38933 , n38925 , n38932 );
xor ( n38934 , n38896 , n38933 );
not ( n38935 , n37588 );
and ( n38936 , n38935 , n37590 );
xor ( n38937 , n35086 , n38936 );
xor ( n38938 , n38937 , n37869 );
not ( n38939 , n32511 );
and ( n38940 , n38939 , n37626 );
xor ( n38941 , n32497 , n38940 );
not ( n38942 , n36903 );
and ( n38943 , n38942 , n37631 );
xor ( n38944 , n32526 , n38943 );
xor ( n38945 , n38941 , n38944 );
xor ( n38946 , n38945 , n36900 );
xor ( n38947 , n38946 , n38248 );
xor ( n38948 , n38947 , n38681 );
xor ( n38949 , n38938 , n38948 );
not ( n38950 , n38949 );
xor ( n38951 , n32173 , n35986 );
xor ( n38952 , n38951 , n36003 );
and ( n38953 , n38950 , n38952 );
xor ( n38954 , n38934 , n38953 );
not ( n12221 , n29614 );
and ( n12222 , n12221 , RI17337660_2171);
and ( n12223 , n38954 , n29614 );
or ( n38955 , n12222 , n12223 );
not ( n12224 , RI1754c610_2);
and ( n12225 , n12224 , n38955 );
and ( n12226 , C0 , RI1754c610_2);
or ( n38956 , n12225 , n12226 );
buf ( n38957 , n38956 );
not ( n38958 , n34054 );
and ( n38959 , n38958 , n34056 );
xor ( n38960 , n33842 , n38959 );
xor ( n38961 , n38960 , n38371 );
xor ( n38962 , n38961 , n36431 );
xor ( n38963 , n32283 , n31399 );
xor ( n38964 , n38963 , n29561 );
not ( n38965 , n33294 );
and ( n38966 , n38965 , n33296 );
xor ( n38967 , n38964 , n38966 );
xor ( n38968 , n30635 , n28174 );
xor ( n38969 , n38968 , n28185 );
not ( n38970 , n33303 );
and ( n38971 , n38970 , n33305 );
xor ( n38972 , n38969 , n38971 );
xor ( n38973 , n38967 , n38972 );
xor ( n38974 , n29552 , n29474 );
xor ( n38975 , n38974 , n32611 );
not ( n38976 , n33313 );
and ( n38977 , n38976 , n33315 );
xor ( n38978 , n38975 , n38977 );
xor ( n38979 , n38973 , n38978 );
xor ( n38980 , n29594 , n28200 );
xor ( n38981 , n38980 , n28212 );
not ( n38982 , n33323 );
and ( n38983 , n38982 , n33285 );
xor ( n38984 , n38981 , n38983 );
xor ( n38985 , n38979 , n38984 );
xor ( n38986 , n27955 , n31131 );
xor ( n38987 , n38986 , n32366 );
not ( n38988 , n33329 );
and ( n38989 , n38988 , n33331 );
xor ( n38990 , n38987 , n38989 );
xor ( n38991 , n38985 , n38990 );
xor ( n38992 , n33310 , n38991 );
not ( n38993 , n33340 );
and ( n38994 , n38993 , n33342 );
xor ( n38995 , n35771 , n38994 );
not ( n38996 , n33349 );
and ( n38997 , n38996 , n33351 );
xor ( n38998 , n35778 , n38997 );
xor ( n38999 , n38995 , n38998 );
xor ( n39000 , n38999 , n35767 );
xor ( n39001 , n39000 , n37873 );
not ( n39002 , n33380 );
and ( n39003 , n39002 , n33391 );
xor ( n39004 , n35800 , n39003 );
xor ( n39005 , n39001 , n39004 );
xor ( n39006 , n38992 , n39005 );
not ( n39007 , n39006 );
xor ( n39008 , n29232 , n30780 );
xor ( n39009 , n39008 , n28043 );
not ( n39010 , n39009 );
and ( n39011 , n39010 , n32582 );
xor ( n39012 , n36932 , n39011 );
not ( n39013 , n36921 );
xor ( n39014 , n27776 , n31024 );
xor ( n39015 , n39014 , n29306 );
and ( n39016 , n39013 , n39015 );
xor ( n39017 , n32568 , n39016 );
not ( n39018 , n36926 );
xor ( n39019 , n28364 , n30522 );
xor ( n39020 , n39019 , n32009 );
and ( n39021 , n39018 , n39020 );
xor ( n39022 , n32577 , n39021 );
xor ( n39023 , n39017 , n39022 );
not ( n39024 , n36932 );
and ( n39025 , n39024 , n39009 );
xor ( n39026 , n32587 , n39025 );
xor ( n39027 , n39023 , n39026 );
not ( n39028 , n36938 );
xor ( n39029 , n28614 , n29995 );
xor ( n39030 , n39029 , n28327 );
and ( n39031 , n39028 , n39030 );
xor ( n39032 , n32597 , n39031 );
xor ( n39033 , n39027 , n39032 );
not ( n39034 , n36944 );
xor ( n39035 , n31711 , n30332 );
xor ( n39036 , n39035 , n32043 );
and ( n39037 , n39034 , n39036 );
xor ( n39038 , n32617 , n39037 );
xor ( n39039 , n39033 , n39038 );
xor ( n39040 , n39012 , n39039 );
xor ( n39041 , n32471 , n28291 );
xor ( n39042 , n39041 , n29781 );
not ( n39043 , n39042 );
and ( n39044 , n39043 , n38964 );
xor ( n39045 , n33299 , n39044 );
xor ( n39046 , n28095 , n31453 );
xor ( n39047 , n39046 , n31462 );
not ( n39048 , n39047 );
and ( n39049 , n39048 , n38969 );
xor ( n39050 , n33308 , n39049 );
xor ( n39051 , n39045 , n39050 );
not ( n39052 , n37337 );
and ( n39053 , n39052 , n38975 );
xor ( n39054 , n33318 , n39053 );
xor ( n39055 , n39051 , n39054 );
not ( n39056 , n33290 );
and ( n39057 , n39056 , n38981 );
xor ( n39058 , n33287 , n39057 );
xor ( n39059 , n39055 , n39058 );
xor ( n39060 , n29024 , n28878 );
xor ( n39061 , n39060 , n30399 );
not ( n39062 , n39061 );
and ( n39063 , n39062 , n38987 );
xor ( n39064 , n33334 , n39063 );
xor ( n39065 , n39059 , n39064 );
xor ( n39066 , n39040 , n39065 );
and ( n39067 , n39007 , n39066 );
xor ( n39068 , n38962 , n39067 );
not ( n12227 , n29614 );
and ( n12228 , n12227 , RI174689e8_1226);
and ( n12229 , n39068 , n29614 );
or ( n39069 , n12228 , n12229 );
not ( n12230 , RI1754c610_2);
and ( n12231 , n12230 , n39069 );
and ( n12232 , C0 , RI1754c610_2);
or ( n39070 , n12231 , n12232 );
buf ( n39071 , n39070 );
buf ( n39072 , RI1747d208_1126);
not ( n39073 , n29663 );
and ( n39074 , n39073 , n29640 );
xor ( n39075 , n36342 , n39074 );
not ( n39076 , n29678 );
and ( n39077 , n39076 , n29681 );
xor ( n39078 , n36349 , n39077 );
xor ( n39079 , n39075 , n39078 );
not ( n39080 , n29700 );
and ( n39081 , n39080 , n29712 );
xor ( n39082 , n36357 , n39081 );
xor ( n39083 , n39079 , n39082 );
not ( n39084 , n29753 );
and ( n39085 , n39084 , n29768 );
xor ( n39086 , n36365 , n39085 );
xor ( n39087 , n39083 , n39086 );
not ( n39088 , n29801 );
and ( n39089 , n39088 , n29815 );
xor ( n39090 , n36373 , n39089 );
xor ( n39091 , n39087 , n39090 );
xor ( n39092 , n29842 , n39091 );
xor ( n39093 , n39092 , n36128 );
xor ( n39094 , n37080 , n37716 );
xor ( n39095 , n39094 , n37744 );
not ( n39096 , n39095 );
not ( n39097 , n37771 );
xor ( n39098 , n29104 , n28505 );
xor ( n39099 , n39098 , n31038 );
and ( n39100 , n39097 , n39099 );
xor ( n39101 , n37768 , n39100 );
xor ( n39102 , n39101 , n37800 );
xor ( n39103 , n39102 , n37814 );
and ( n39104 , n39096 , n39103 );
xor ( n39105 , n39093 , n39104 );
not ( n12233 , n29614 );
and ( n12234 , n12233 , RI173b6140_1868);
and ( n12235 , n39105 , n29614 );
or ( n39106 , n12234 , n12235 );
not ( n12236 , RI1754c610_2);
and ( n12237 , n12236 , n39106 );
and ( n12238 , C0 , RI1754c610_2);
or ( n39107 , n12237 , n12238 );
buf ( n39108 , n39107 );
not ( n39109 , n38137 );
xor ( n39110 , n31745 , n28262 );
xor ( n39111 , n39110 , n28892 );
and ( n39112 , n39109 , n39111 );
xor ( n39113 , n31008 , n39112 );
xor ( n39114 , n39113 , n38150 );
xor ( n39115 , n39114 , n38167 );
not ( n39116 , n27871 );
and ( n39117 , n39116 , n29874 );
xor ( n39118 , n27845 , n39117 );
xor ( n39119 , n27767 , n39118 );
not ( n39120 , n27949 );
and ( n39121 , n39120 , n29890 );
xor ( n39122 , n27922 , n39121 );
xor ( n39123 , n39119 , n39122 );
not ( n39124 , n28028 );
and ( n39125 , n39124 , n29911 );
xor ( n39126 , n28002 , n39125 );
xor ( n39127 , n39123 , n39126 );
not ( n39128 , n28108 );
and ( n39129 , n39128 , n29965 );
xor ( n39130 , n28082 , n39129 );
xor ( n39131 , n39127 , n39130 );
xor ( n39132 , n36123 , n39131 );
not ( n39133 , n28186 );
and ( n39134 , n39133 , n35918 );
xor ( n39135 , n28161 , n39134 );
not ( n39136 , n28263 );
and ( n39137 , n39136 , n35925 );
xor ( n39138 , n28237 , n39137 );
xor ( n39139 , n39135 , n39138 );
not ( n39140 , n28340 );
and ( n39141 , n39140 , n35933 );
xor ( n39142 , n28314 , n39141 );
xor ( n39143 , n39139 , n39142 );
not ( n39144 , n28419 );
and ( n39145 , n39144 , n35941 );
xor ( n39146 , n28393 , n39145 );
xor ( n39147 , n39143 , n39146 );
not ( n39148 , n28465 );
and ( n39149 , n39148 , n35949 );
xor ( n39150 , n28451 , n39149 );
xor ( n39151 , n39147 , n39150 );
xor ( n39152 , n39132 , n39151 );
not ( n39153 , n39152 );
xor ( n39154 , n36286 , n37311 );
xor ( n39155 , n39154 , n37942 );
and ( n39156 , n39153 , n39155 );
xor ( n39157 , n39115 , n39156 );
not ( n12239 , n29614 );
and ( n12240 , n12239 , RI1750d820_724);
and ( n12241 , n39157 , n29614 );
or ( n39158 , n12240 , n12241 );
not ( n12242 , RI1754c610_2);
and ( n12243 , n12242 , n39158 );
and ( n12244 , C0 , RI1754c610_2);
or ( n39159 , n12243 , n12244 );
buf ( n39160 , n39159 );
xor ( n39161 , n36132 , n39151 );
xor ( n39162 , n39161 , n38267 );
not ( n39163 , n39162 );
not ( n39164 , n32563 );
and ( n39165 , n39164 , n32565 );
xor ( n39166 , n39015 , n39165 );
not ( n39167 , n32572 );
and ( n39168 , n39167 , n32574 );
xor ( n39169 , n39020 , n39168 );
xor ( n39170 , n39166 , n39169 );
not ( n39171 , n32582 );
and ( n39172 , n39171 , n32584 );
xor ( n39173 , n39009 , n39172 );
xor ( n39174 , n39170 , n39173 );
not ( n39175 , n32592 );
and ( n39176 , n39175 , n32594 );
xor ( n39177 , n39030 , n39176 );
xor ( n39178 , n39174 , n39177 );
not ( n39179 , n32612 );
and ( n39180 , n39179 , n32614 );
xor ( n39181 , n39036 , n39180 );
xor ( n39182 , n39178 , n39181 );
xor ( n39183 , n32579 , n39182 );
xor ( n39184 , n39183 , n38991 );
and ( n39185 , n39163 , n39184 );
xor ( n39186 , n34476 , n39185 );
not ( n12245 , n29614 );
and ( n12246 , n12245 , RI17339a78_2160);
and ( n12247 , n39186 , n29614 );
or ( n39187 , n12246 , n12247 );
not ( n12248 , RI1754c610_2);
and ( n12249 , n12248 , n39187 );
and ( n12250 , C0 , RI1754c610_2);
or ( n39188 , n12249 , n12250 );
buf ( n39189 , n39188 );
not ( n12251 , n27683 );
and ( n12252 , n12251 , RI19aa17f8_2556);
and ( n12253 , RI19aab938_2485 , n27683 );
or ( n39190 , n12252 , n12253 );
not ( n12254 , RI1754c610_2);
and ( n12255 , n12254 , n39190 );
and ( n12256 , C0 , RI1754c610_2);
or ( n39191 , n12255 , n12256 );
buf ( n39192 , n39191 );
not ( n39193 , n36745 );
and ( n39194 , n39193 , n34875 );
xor ( n39195 , n37533 , n39194 );
xor ( n39196 , n39195 , n37660 );
not ( n39197 , n36756 );
and ( n39198 , n39197 , n34894 );
xor ( n39199 , n37539 , n39198 );
xor ( n39200 , n39196 , n39199 );
not ( n39201 , n36762 );
and ( n39202 , n39201 , n34904 );
xor ( n39203 , n37545 , n39202 );
xor ( n39204 , n39200 , n39203 );
not ( n39205 , n36768 );
and ( n39206 , n39205 , n34914 );
xor ( n39207 , n34871 , n39206 );
xor ( n39208 , n39204 , n39207 );
xor ( n39209 , n36759 , n39208 );
xor ( n39210 , n39209 , n38214 );
not ( n39211 , n33599 );
and ( n39212 , n39211 , n33601 );
xor ( n39213 , n34825 , n39212 );
xor ( n39214 , n39213 , n34837 );
xor ( n39215 , n39214 , n33880 );
not ( n39216 , n39215 );
not ( n39217 , n33279 );
and ( n39218 , n39217 , n33691 );
xor ( n39219 , n33276 , n39218 );
xor ( n39220 , n39219 , n33282 );
xor ( n39221 , n39220 , n37623 );
and ( n39222 , n39216 , n39221 );
xor ( n39223 , n39210 , n39222 );
not ( n12257 , n29614 );
and ( n12258 , n12257 , RI173e5de0_1635);
and ( n12259 , n39223 , n29614 );
or ( n39224 , n12258 , n12259 );
not ( n12260 , RI1754c610_2);
and ( n12261 , n12260 , n39224 );
and ( n12262 , C0 , RI1754c610_2);
or ( n39225 , n12261 , n12262 );
buf ( n39226 , n39225 );
and ( n39227 , RI1754c430_6 , n34844 );
and ( n39228 , RI1754c430_6 , n34847 );
and ( n39229 , RI1754c430_6 , n34850 );
and ( n39230 , RI1754c430_6 , n34852 );
and ( n39231 , RI1754c430_6 , n34854 );
and ( n39232 , RI1754c430_6 , n34856 );
nor ( n39233 , n34846 , RI1754a630_70 , RI1754a6a8_69);
and ( n39234 , RI1754c430_6 , n39233 );
or ( n39235 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39234 , C0 );
not ( n12263 , n34859 );
and ( n12264 , n12263 , n39235 );
and ( n12265 , RI1754c430_6 , n34859 );
or ( n39236 , n12264 , n12265 );
not ( n12266 , RI19a22f70_2797);
and ( n12267 , n12266 , n39236 );
and ( n12268 , C0 , RI19a22f70_2797);
or ( n39237 , n12267 , n12268 );
not ( n12269 , n27683 );
and ( n12270 , n12269 , RI19a88460_2736);
and ( n12271 , n39237 , n27683 );
or ( n39238 , n12270 , n12271 );
not ( n12272 , RI1754c610_2);
and ( n12273 , n12272 , n39238 );
and ( n12274 , C0 , RI1754c610_2);
or ( n39239 , n12273 , n12274 );
buf ( n39240 , n39239 );
not ( n12275 , n27683 );
and ( n12276 , n12275 , RI19a97820_2629);
and ( n12277 , RI19aa1438_2558 , n27683 );
or ( n39241 , n12276 , n12277 );
not ( n12278 , RI1754c610_2);
and ( n12279 , n12278 , n39241 );
and ( n12280 , C0 , RI1754c610_2);
or ( n39242 , n12279 , n12280 );
buf ( n39243 , n39242 );
not ( n39244 , n36963 );
and ( n39245 , n39244 , n36958 );
xor ( n39246 , n35319 , n39245 );
not ( n39247 , n35319 );
and ( n39248 , n39247 , n36963 );
xor ( n39249 , n35316 , n39248 );
not ( n39250 , n35328 );
and ( n39251 , n39250 , n36968 );
xor ( n39252 , n35325 , n39251 );
xor ( n39253 , n39249 , n39252 );
not ( n39254 , n35338 );
and ( n39255 , n39254 , n36976 );
xor ( n39256 , n35335 , n39255 );
xor ( n39257 , n39253 , n39256 );
not ( n39258 , n35348 );
and ( n39259 , n39258 , n36984 );
xor ( n39260 , n35345 , n39259 );
xor ( n39261 , n39257 , n39260 );
xor ( n39262 , n39261 , n38405 );
xor ( n39263 , n39246 , n39262 );
not ( n39264 , n38411 );
and ( n39265 , n39264 , n37001 );
xor ( n39266 , n38408 , n39265 );
not ( n39267 , n38418 );
and ( n39268 , n39267 , n37010 );
xor ( n39269 , n38415 , n39268 );
xor ( n39270 , n39266 , n39269 );
not ( n39271 , n38426 );
and ( n39272 , n39271 , n37020 );
xor ( n39273 , n38423 , n39272 );
xor ( n39274 , n39270 , n39273 );
not ( n39275 , n38434 );
and ( n39276 , n39275 , n37030 );
xor ( n39277 , n38431 , n39276 );
xor ( n39278 , n39274 , n39277 );
not ( n39279 , n38442 );
and ( n39280 , n39279 , n37040 );
xor ( n39281 , n38439 , n39280 );
xor ( n39282 , n39278 , n39281 );
xor ( n39283 , n39263 , n39282 );
xor ( n39284 , n33144 , n37235 );
xor ( n39285 , n39284 , n37255 );
not ( n39286 , n39285 );
not ( n39287 , n33805 );
and ( n39288 , n39287 , n32347 );
xor ( n39289 , n33802 , n39288 );
xor ( n39290 , n39289 , n33824 );
xor ( n39291 , n39290 , n32786 );
and ( n39292 , n39286 , n39291 );
xor ( n39293 , n39283 , n39292 );
not ( n12281 , n29614 );
and ( n12282 , n12281 , RI17340d50_2125);
and ( n12283 , n39293 , n29614 );
or ( n39294 , n12282 , n12283 );
not ( n12284 , RI1754c610_2);
and ( n12285 , n12284 , n39294 );
and ( n12286 , C0 , RI1754c610_2);
or ( n39295 , n12285 , n12286 );
buf ( n39296 , n39295 );
buf ( n39297 , RI17482758_1100);
buf ( n39298 , RI1748a750_1061);
buf ( n39299 , RI175085a0_740);
buf ( n39300 , RI1750f1e8_719);
xor ( n39301 , n38623 , n38347 );
xor ( n39302 , n39301 , n34300 );
xor ( n39303 , n38143 , n31053 );
xor ( n39304 , n39303 , n35494 );
not ( n39305 , n39304 );
xor ( n39306 , n37202 , n33030 );
xor ( n39307 , n39306 , n33069 );
and ( n39308 , n39305 , n39307 );
xor ( n39309 , n39302 , n39308 );
not ( n12287 , n29614 );
and ( n12288 , n12287 , RI173a0c00_1972);
and ( n12289 , n39309 , n29614 );
or ( n39310 , n12288 , n12289 );
not ( n12290 , RI1754c610_2);
and ( n12291 , n12290 , n39310 );
and ( n12292 , C0 , RI1754c610_2);
or ( n39311 , n12291 , n12292 );
buf ( n39312 , n39311 );
xor ( n39313 , n30377 , n35311 );
xor ( n39314 , n39313 , n35361 );
xor ( n39315 , n35043 , n37814 );
xor ( n39316 , n39315 , n33223 );
not ( n39317 , n39316 );
not ( n39318 , n35369 );
and ( n39319 , n39318 , n36335 );
xor ( n39320 , n35366 , n39319 );
not ( n39321 , n35378 );
and ( n39322 , n39321 , n36306 );
xor ( n39323 , n35375 , n39322 );
xor ( n39324 , n39323 , n37052 );
not ( n39325 , n35397 );
and ( n39326 , n39325 , n36321 );
xor ( n39327 , n35394 , n39326 );
xor ( n39328 , n39324 , n39327 );
not ( n39329 , n35407 );
and ( n39330 , n39329 , n36327 );
xor ( n39331 , n35404 , n39330 );
xor ( n39332 , n39328 , n39331 );
xor ( n39333 , n39332 , n35371 );
xor ( n39334 , n39320 , n39333 );
not ( n39335 , n29695 );
and ( n39336 , n39335 , n36347 );
xor ( n39337 , n29681 , n39336 );
xor ( n39338 , n29659 , n39337 );
not ( n39339 , n29725 );
and ( n39340 , n39339 , n36355 );
xor ( n39341 , n29712 , n39340 );
xor ( n39342 , n39338 , n39341 );
xor ( n39343 , n39342 , n36410 );
not ( n39344 , n29840 );
and ( n39345 , n39344 , n36371 );
xor ( n39346 , n29815 , n39345 );
xor ( n39347 , n39343 , n39346 );
xor ( n39348 , n39334 , n39347 );
and ( n39349 , n39317 , n39348 );
xor ( n39350 , n39314 , n39349 );
not ( n12293 , n29614 );
and ( n12294 , n12293 , RI173a7848_1939);
and ( n12295 , n39350 , n29614 );
or ( n39351 , n12294 , n12295 );
not ( n12296 , RI1754c610_2);
and ( n12297 , n12296 , n39351 );
and ( n12298 , C0 , RI1754c610_2);
or ( n39352 , n12297 , n12298 );
buf ( n39353 , n39352 );
not ( n12299 , RI1754c610_2);
and ( n12300 , n12299 , RI175373a0_595);
and ( n12301 , C0 , RI1754c610_2);
or ( n39354 , n12300 , n12301 );
buf ( n39355 , n39354 );
not ( n12302 , n27683 );
and ( n12303 , n12302 , RI19ab5d48_2410);
and ( n12304 , RI19abf0f0_2340 , n27683 );
or ( n39356 , n12303 , n12304 );
not ( n12305 , RI1754c610_2);
and ( n12306 , n12305 , n39356 );
and ( n12307 , C0 , RI1754c610_2);
or ( n39357 , n12306 , n12307 );
buf ( n39358 , n39357 );
xor ( n39359 , n32317 , n29781 );
xor ( n39360 , n39359 , n29793 );
not ( n39361 , n39360 );
and ( n39362 , n39361 , n37463 );
xor ( n39363 , n35552 , n39362 );
or ( n39364 , n35141 , RI175385e8_592);
or ( n39365 , n39364 , RI17537fd0_593);
or ( n39366 , n39365 , RI175379b8_594);
or ( n39367 , n39366 , RI175373a0_595);
or ( n39368 , n39367 , RI17536d88_596);
or ( n39369 , n39368 , RI17536770_597);
xor ( n39370 , n39363 , n39369 );
not ( n39371 , n35552 );
and ( n39372 , n39371 , n39360 );
xor ( n39373 , n35549 , n39372 );
not ( n39374 , n35561 );
xor ( n39375 , n30560 , n31038 );
xor ( n39376 , n39375 , n30271 );
and ( n39377 , n39374 , n39376 );
xor ( n39378 , n35558 , n39377 );
xor ( n39379 , n39373 , n39378 );
not ( n39380 , n35571 );
xor ( n39381 , n28778 , n32043 );
xor ( n39382 , n39381 , n30946 );
and ( n39383 , n39380 , n39382 );
xor ( n39384 , n35568 , n39383 );
xor ( n39385 , n39379 , n39384 );
not ( n39386 , n35581 );
xor ( n39387 , n27902 , n29235 );
xor ( n39388 , n39387 , n30294 );
and ( n39389 , n39386 , n39388 );
xor ( n39390 , n35578 , n39389 );
xor ( n39391 , n39385 , n39390 );
not ( n39392 , n35591 );
xor ( n39393 , n27851 , n29655 );
xor ( n39394 , n39393 , n29601 );
and ( n39395 , n39392 , n39394 );
xor ( n39396 , n35588 , n39395 );
xor ( n39397 , n39391 , n39396 );
xor ( n39398 , n39370 , n39397 );
not ( n39399 , n32342 );
and ( n39400 , n39399 , n33786 );
xor ( n39401 , n32339 , n39400 );
xor ( n39402 , n32330 , n39401 );
not ( n39403 , n32352 );
and ( n39404 , n39403 , n33802 );
xor ( n39405 , n32349 , n39404 );
xor ( n39406 , n39402 , n39405 );
not ( n39407 , n32383 );
and ( n39408 , n39407 , n33810 );
xor ( n39409 , n32370 , n39408 );
xor ( n39410 , n39406 , n39409 );
not ( n39411 , n32400 );
and ( n39412 , n39411 , n33818 );
xor ( n39413 , n32390 , n39412 );
xor ( n39414 , n39410 , n39413 );
xor ( n39415 , n39398 , n39414 );
xor ( n39416 , n37683 , n37579 );
xor ( n39417 , n39416 , n38495 );
not ( n39418 , n39417 );
xor ( n39419 , n34901 , n36772 );
xor ( n39420 , n39419 , n36802 );
and ( n39421 , n39418 , n39420 );
xor ( n39422 , n39415 , n39421 );
or ( n39423 , n27689 , RI1753a460_587);
or ( n39424 , n39423 , RI17539218_590);
or ( n39425 , n39424 , RI175379b8_594);
or ( n39426 , n39425 , RI17536770_597);
or ( n39427 , n39426 , RI17539e48_588);
xor ( n39428 , n39422 , n39427 );
not ( n12308 , n29614 );
and ( n12309 , n12308 , RI1746be68_1210);
and ( n12310 , n39428 , n29614 );
or ( n39429 , n12309 , n12310 );
not ( n12311 , RI1754c610_2);
and ( n12312 , n12311 , n39429 );
and ( n12313 , C0 , RI1754c610_2);
or ( n39430 , n12312 , n12313 );
buf ( n39431 , n39430 );
not ( n39432 , n38217 );
and ( n39433 , n39432 , n33082 );
xor ( n39434 , n38470 , n39433 );
not ( n39435 , n38222 );
and ( n39436 , n39435 , n33091 );
xor ( n39437 , n38475 , n39436 );
xor ( n39438 , n39434 , n39437 );
not ( n39439 , n38228 );
and ( n39440 , n39439 , n33101 );
xor ( n39441 , n38481 , n39440 );
xor ( n39442 , n39438 , n39441 );
not ( n39443 , n38234 );
and ( n39444 , n39443 , n33111 );
xor ( n39445 , n33078 , n39444 );
xor ( n39446 , n39442 , n39445 );
not ( n39447 , n38240 );
and ( n39448 , n39447 , n33117 );
xor ( n39449 , n38491 , n39448 );
xor ( n39450 , n39446 , n39449 );
xor ( n39451 , n38231 , n39450 );
not ( n39452 , n36581 );
and ( n39453 , n39452 , n33128 );
xor ( n39454 , n36578 , n39453 );
xor ( n39455 , n39454 , n36576 );
not ( n39456 , n36592 );
and ( n39457 , n39456 , n33147 );
xor ( n39458 , n36589 , n39457 );
xor ( n39459 , n39455 , n39458 );
not ( n39460 , n36600 );
and ( n39461 , n39460 , n33157 );
xor ( n39462 , n36597 , n39461 );
xor ( n39463 , n39459 , n39462 );
not ( n39464 , n36608 );
and ( n39465 , n39464 , n33167 );
xor ( n39466 , n36605 , n39465 );
xor ( n39467 , n39463 , n39466 );
xor ( n39468 , n39451 , n39467 );
not ( n39469 , n33553 );
and ( n39470 , n39469 , n33513 );
xor ( n39471 , n34785 , n39470 );
xor ( n39472 , n39471 , n34797 );
xor ( n39473 , n39472 , n34837 );
not ( n39474 , n39473 );
not ( n39475 , n35173 );
and ( n39476 , n39475 , n32021 );
xor ( n39477 , n35170 , n39476 );
xor ( n39478 , n39477 , n35176 );
xor ( n39479 , n39478 , n35216 );
and ( n39480 , n39474 , n39479 );
xor ( n39481 , n39468 , n39480 );
not ( n12314 , n29614 );
and ( n12315 , n12314 , RI17493120_1019);
and ( n12316 , n39481 , n29614 );
or ( n39482 , n12315 , n12316 );
not ( n12317 , RI1754c610_2);
and ( n12318 , n12317 , n39482 );
and ( n12319 , C0 , RI1754c610_2);
or ( n39483 , n12318 , n12319 );
buf ( n39484 , n39483 );
xor ( n39485 , n29374 , n31989 );
xor ( n39486 , n39485 , n33898 );
not ( n39487 , n39486 );
and ( n39488 , n39487 , n38088 );
xor ( n39489 , n30800 , n39488 );
not ( n39490 , n30800 );
and ( n39491 , n39490 , n39486 );
xor ( n39492 , n30781 , n39491 );
xor ( n39493 , n39492 , n35853 );
not ( n39494 , n30870 );
xor ( n39495 , n29838 , n32140 );
xor ( n39496 , n39495 , n31874 );
and ( n39497 , n39494 , n39496 );
xor ( n39498 , n30846 , n39497 );
xor ( n39499 , n39493 , n39498 );
not ( n39500 , n30905 );
xor ( n39501 , n30347 , n31152 );
xor ( n39502 , n39501 , n31162 );
and ( n39503 , n39500 , n39502 );
xor ( n39504 , n30902 , n39503 );
xor ( n39505 , n39499 , n39504 );
xor ( n39506 , n39505 , n30767 );
xor ( n39507 , n39489 , n39506 );
xor ( n39508 , n39507 , n38150 );
not ( n39509 , n33584 );
and ( n39510 , n39509 , n34807 );
xor ( n39511 , n33581 , n39510 );
xor ( n39512 , n39511 , n33617 );
not ( n39513 , n34061 );
and ( n39514 , n39513 , n34049 );
xor ( n39515 , n33851 , n39514 );
xor ( n39516 , n38960 , n39515 );
xor ( n39517 , n39516 , n38355 );
not ( n39518 , n34073 );
and ( n39519 , n39518 , n34075 );
xor ( n39520 , n33867 , n39519 );
xor ( n39521 , n39517 , n39520 );
not ( n39522 , n34081 );
and ( n39523 , n39522 , n34083 );
xor ( n39524 , n33877 , n39523 );
xor ( n39525 , n39521 , n39524 );
xor ( n39526 , n39512 , n39525 );
not ( n39527 , n39526 );
not ( n39528 , n35667 );
and ( n39529 , n39528 , n35669 );
xor ( n39530 , n35809 , n39529 );
not ( n39531 , n35676 );
and ( n39532 , n39531 , n35658 );
xor ( n39533 , n35814 , n39532 );
xor ( n39534 , n39530 , n39533 );
not ( n39535 , n35682 );
and ( n39536 , n39535 , n35684 );
xor ( n39537 , n35822 , n39536 );
xor ( n39538 , n39534 , n39537 );
xor ( n39539 , n39538 , n38381 );
not ( n39540 , n35702 );
and ( n39541 , n39540 , n35704 );
xor ( n39542 , n35838 , n39541 );
xor ( n39543 , n39539 , n39542 );
xor ( n39544 , n35689 , n39543 );
not ( n39545 , n35713 );
and ( n39546 , n39545 , n35715 );
xor ( n39547 , n37135 , n39546 );
not ( n39548 , n35722 );
and ( n39549 , n39548 , n35724 );
xor ( n39550 , n37142 , n39549 );
xor ( n39551 , n39547 , n39550 );
not ( n39552 , n35732 );
and ( n39553 , n39552 , n35734 );
xor ( n39554 , n37150 , n39553 );
xor ( n39555 , n39551 , n39554 );
not ( n39556 , n35742 );
and ( n39557 , n39556 , n35744 );
xor ( n39558 , n37158 , n39557 );
xor ( n39559 , n39555 , n39558 );
not ( n39560 , n35752 );
and ( n39561 , n39560 , n35754 );
xor ( n39562 , n37166 , n39561 );
xor ( n39563 , n39559 , n39562 );
xor ( n39564 , n39544 , n39563 );
and ( n39565 , n39527 , n39564 );
xor ( n39566 , n39508 , n39565 );
not ( n12320 , n29614 );
and ( n12321 , n12320 , RI174acb48_894);
and ( n12322 , n39566 , n29614 );
or ( n39567 , n12321 , n12322 );
not ( n12323 , RI1754c610_2);
and ( n12324 , n12323 , n39567 );
and ( n12325 , C0 , RI1754c610_2);
or ( n39568 , n12324 , n12325 );
buf ( n39569 , n39568 );
and ( n39570 , RI1754b800_32 , n34844 );
and ( n39571 , RI1754b800_32 , n34847 );
and ( n39572 , RI1754b800_32 , n34850 );
and ( n39573 , RI1754b800_32 , n34852 );
or ( n39574 , n39570 , n39571 , n39572 , n39573 , C0 , C0 , C0 , C0 );
not ( n12326 , n34859 );
and ( n12327 , n12326 , n39574 );
and ( n12328 , RI1754b800_32 , n34859 );
or ( n39575 , n12327 , n12328 );
not ( n12329 , RI19a22f70_2797);
and ( n12330 , n12329 , n39575 );
and ( n12331 , C0 , RI19a22f70_2797);
or ( n39576 , n12330 , n12331 );
not ( n12332 , n27683 );
and ( n12333 , n12332 , RI19aac388_2481);
and ( n12334 , n39576 , n27683 );
or ( n39577 , n12333 , n12334 );
not ( n12335 , RI1754c610_2);
and ( n12336 , n12335 , n39577 );
and ( n12337 , C0 , RI1754c610_2);
or ( n39578 , n12336 , n12337 );
buf ( n39579 , n39578 );
not ( n39580 , n31534 );
and ( n39581 , n39580 , n34303 );
xor ( n39582 , n31531 , n39581 );
or ( n39583 , n35140 , RI17538c00_591);
or ( n39584 , n39583 , RI175385e8_592);
or ( n39585 , n39584 , RI17537fd0_593);
or ( n39586 , n39585 , RI175379b8_594);
or ( n39587 , n39586 , RI17536d88_596);
xor ( n39588 , n39582 , n39587 );
not ( n39589 , n31546 );
and ( n39590 , n39589 , n34310 );
xor ( n39591 , n31543 , n39590 );
xor ( n39592 , n39588 , n39591 );
not ( n39593 , n31565 );
and ( n39594 , n39593 , n34318 );
xor ( n39595 , n31562 , n39594 );
xor ( n39596 , n39592 , n39595 );
not ( n39597 , n31595 );
and ( n39598 , n39597 , n34326 );
xor ( n39599 , n31582 , n39598 );
xor ( n39600 , n39596 , n39599 );
not ( n39601 , n31618 );
and ( n39602 , n39601 , n34334 );
xor ( n39603 , n31615 , n39602 );
xor ( n39604 , n39600 , n39603 );
xor ( n39605 , n34339 , n39604 );
not ( n39606 , n35234 );
and ( n39607 , n39606 , n38691 );
xor ( n39608 , n35231 , n39607 );
xor ( n39609 , n39608 , n35227 );
not ( n39610 , n35249 );
and ( n39611 , n39610 , n38702 );
xor ( n39612 , n35246 , n39611 );
xor ( n39613 , n39609 , n39612 );
not ( n39614 , n35259 );
and ( n39615 , n39614 , n38710 );
xor ( n39616 , n35256 , n39615 );
xor ( n39617 , n39613 , n39616 );
not ( n39618 , n35269 );
and ( n39619 , n39618 , n38718 );
xor ( n39620 , n35266 , n39619 );
xor ( n39621 , n39617 , n39620 );
xor ( n39622 , n39605 , n39621 );
not ( n39623 , n35151 );
and ( n39624 , n39623 , n31979 );
xor ( n39625 , n35148 , n39624 );
xor ( n39626 , n35136 , n39625 );
not ( n39627 , n35159 );
and ( n39628 , n39627 , n31998 );
xor ( n39629 , n35156 , n39628 );
xor ( n39630 , n39626 , n39629 );
not ( n39631 , n35165 );
and ( n39632 , n39631 , n32015 );
xor ( n39633 , n31938 , n39632 );
xor ( n39634 , n39630 , n39633 );
xor ( n39635 , n39634 , n39477 );
xor ( n39636 , n36666 , n39635 );
not ( n39637 , n35182 );
and ( n39638 , n39637 , n32051 );
xor ( n39639 , n35179 , n39638 );
not ( n39640 , n35189 );
and ( n39641 , n39640 , n32060 );
xor ( n39642 , n35186 , n39641 );
xor ( n39643 , n39639 , n39642 );
not ( n39644 , n35197 );
and ( n39645 , n39644 , n32070 );
xor ( n39646 , n35194 , n39645 );
xor ( n39647 , n39643 , n39646 );
not ( n39648 , n35205 );
and ( n39649 , n39648 , n32080 );
xor ( n39650 , n35202 , n39649 );
xor ( n39651 , n39647 , n39650 );
not ( n39652 , n35213 );
and ( n39653 , n39652 , n32100 );
xor ( n39654 , n35210 , n39653 );
xor ( n39655 , n39651 , n39654 );
xor ( n39656 , n39636 , n39655 );
not ( n39657 , n39656 );
and ( n39658 , n39657 , n33826 );
xor ( n39659 , n39622 , n39658 );
not ( n12338 , n29614 );
and ( n12339 , n12338 , RI173cda98_1753);
and ( n12340 , n39659 , n29614 );
or ( n39660 , n12339 , n12340 );
not ( n12341 , RI1754c610_2);
and ( n12342 , n12341 , n39660 );
and ( n12343 , C0 , RI1754c610_2);
or ( n39661 , n12342 , n12343 );
buf ( n39662 , n39661 );
not ( n39663 , n34800 );
and ( n39664 , n39663 , n34802 );
xor ( n39665 , n33575 , n39664 );
or ( n39666 , RI17539218_590 , RI175385e8_592);
or ( n39667 , n39666 , RI17537fd0_593);
or ( n39668 , n39667 , RI17536770_597);
or ( n39669 , n39668 , RI17539e48_588);
xor ( n39670 , n39665 , n39669 );
not ( n39671 , n33575 );
and ( n39672 , n39671 , n34800 );
xor ( n39673 , n33572 , n39672 );
xor ( n39674 , n39673 , n39511 );
not ( n39675 , n33594 );
and ( n39676 , n39675 , n34815 );
xor ( n39677 , n33591 , n39676 );
xor ( n39678 , n39674 , n39677 );
not ( n39679 , n33604 );
and ( n39680 , n39679 , n34823 );
xor ( n39681 , n33601 , n39680 );
xor ( n39682 , n39678 , n39681 );
not ( n39683 , n33614 );
and ( n39684 , n39683 , n34831 );
xor ( n39685 , n33611 , n39684 );
xor ( n39686 , n39682 , n39685 );
xor ( n39687 , n39670 , n39686 );
xor ( n39688 , n39687 , n34087 );
xor ( n39689 , n39022 , n36947 );
not ( n39690 , n33299 );
and ( n39691 , n39690 , n39042 );
xor ( n39692 , n33296 , n39691 );
not ( n39693 , n33308 );
and ( n39694 , n39693 , n39047 );
xor ( n39695 , n33305 , n39694 );
xor ( n39696 , n39692 , n39695 );
xor ( n39697 , n39696 , n37339 );
xor ( n39698 , n39697 , n33292 );
not ( n39699 , n33334 );
and ( n39700 , n39699 , n39061 );
xor ( n39701 , n33331 , n39700 );
xor ( n39702 , n39698 , n39701 );
xor ( n39703 , n39689 , n39702 );
not ( n39704 , n39703 );
xor ( n39705 , n32538 , n37651 );
xor ( n39706 , n39705 , n39182 );
and ( n39707 , n39704 , n39706 );
xor ( n39708 , n39688 , n39707 );
or ( n39709 , n35140 , RI175385e8_592);
or ( n39710 , n39709 , RI17536d88_596);
or ( n39711 , n39710 , RI17539e48_588);
xor ( n39712 , n39708 , n39711 );
not ( n12344 , n29614 );
and ( n12345 , n12344 , RI174686a0_1227);
and ( n12346 , n39712 , n29614 );
or ( n39713 , n12345 , n12346 );
not ( n12347 , RI1754c610_2);
and ( n12348 , n12347 , n39713 );
and ( n12349 , C0 , RI1754c610_2);
or ( n39714 , n12348 , n12349 );
buf ( n39715 , n39714 );
not ( n12350 , n27683 );
and ( n12351 , n12350 , RI19aa0358_2567);
and ( n12352 , RI19aa9f70_2496 , n27683 );
or ( n39716 , n12351 , n12352 );
not ( n12353 , RI1754c610_2);
and ( n12354 , n12353 , n39716 );
and ( n12355 , C0 , RI1754c610_2);
or ( n39717 , n12354 , n12355 );
buf ( n39718 , n39717 );
xor ( n39719 , n36422 , n33935 );
xor ( n39720 , n39719 , n36287 );
not ( n39721 , n38024 );
and ( n39722 , n39721 , n38071 );
xor ( n39723 , n38021 , n39722 );
xor ( n39724 , n39723 , n38037 );
not ( n39725 , n35851 );
and ( n39726 , n39725 , n38093 );
xor ( n39727 , n30829 , n39726 );
xor ( n39728 , n39489 , n39727 );
not ( n39729 , n39496 );
and ( n39730 , n39729 , n38099 );
xor ( n39731 , n30870 , n39730 );
xor ( n39732 , n39728 , n39731 );
not ( n39733 , n39502 );
and ( n39734 , n39733 , n38105 );
xor ( n39735 , n30905 , n39734 );
xor ( n39736 , n39732 , n39735 );
not ( n39737 , n30765 );
and ( n39738 , n39737 , n38111 );
xor ( n39739 , n30762 , n39738 );
xor ( n39740 , n39736 , n39739 );
xor ( n39741 , n39724 , n39740 );
not ( n39742 , n39741 );
not ( n39743 , n35757 );
and ( n39744 , n39743 , n37163 );
xor ( n39745 , n35754 , n39744 );
xor ( n39746 , n39745 , n35760 );
xor ( n39747 , n39746 , n39333 );
and ( n39748 , n39742 , n39747 );
xor ( n39749 , n39720 , n39748 );
not ( n12356 , n29614 );
and ( n12357 , n12356 , RI173e7820_1627);
and ( n12358 , n39749 , n29614 );
or ( n39750 , n12357 , n12358 );
not ( n12359 , RI1754c610_2);
and ( n12360 , n12359 , n39750 );
and ( n12361 , C0 , RI1754c610_2);
or ( n39751 , n12360 , n12361 );
buf ( n39752 , n39751 );
not ( n12362 , n27683 );
and ( n12363 , n12362 , RI19aa9bb0_2498);
and ( n12364 , RI19ab36d8_2428 , n27683 );
or ( n39753 , n12363 , n12364 );
not ( n12365 , RI1754c610_2);
and ( n12366 , n12365 , n39753 );
and ( n12367 , C0 , RI1754c610_2);
or ( n39754 , n12366 , n12367 );
buf ( n39755 , n39754 );
not ( n39756 , n33087 );
and ( n39757 , n39756 , n38470 );
xor ( n39758 , n33084 , n39757 );
not ( n39759 , n33096 );
and ( n39760 , n39759 , n38475 );
xor ( n39761 , n33093 , n39760 );
xor ( n39762 , n39758 , n39761 );
not ( n39763 , n33106 );
and ( n39764 , n39763 , n38481 );
xor ( n39765 , n33103 , n39764 );
xor ( n39766 , n39762 , n39765 );
xor ( n39767 , n39766 , n33080 );
not ( n39768 , n33122 );
and ( n39769 , n39768 , n38491 );
xor ( n39770 , n33119 , n39769 );
xor ( n39771 , n39767 , n39770 );
xor ( n39772 , n38488 , n39771 );
not ( n39773 , n33133 );
and ( n39774 , n39773 , n36578 );
xor ( n39775 , n33130 , n39774 );
not ( n39776 , n33142 );
and ( n39777 , n39776 , n36571 );
xor ( n39778 , n33139 , n39777 );
xor ( n39779 , n39775 , n39778 );
not ( n39780 , n33152 );
and ( n39781 , n39780 , n36589 );
xor ( n39782 , n33149 , n39781 );
xor ( n39783 , n39779 , n39782 );
not ( n39784 , n33162 );
and ( n39785 , n39784 , n36597 );
xor ( n39786 , n33159 , n39785 );
xor ( n39787 , n39783 , n39786 );
not ( n39788 , n33172 );
and ( n39789 , n39788 , n36605 );
xor ( n39790 , n33169 , n39789 );
xor ( n39791 , n39787 , n39790 );
xor ( n39792 , n39772 , n39791 );
xor ( n39793 , n31099 , n29320 );
xor ( n39794 , n39793 , n29332 );
not ( n39795 , n39794 );
xor ( n39796 , n30046 , n28904 );
xor ( n39797 , n39796 , n29291 );
and ( n39798 , n39795 , n39797 );
xor ( n39799 , n37797 , n39798 );
not ( n39800 , n37762 );
xor ( n39801 , n29234 , n30780 );
xor ( n39802 , n39801 , n28043 );
and ( n39803 , n39800 , n39802 );
xor ( n39804 , n37759 , n39803 );
xor ( n39805 , n39804 , n39101 );
not ( n39806 , n37781 );
xor ( n39807 , n31580 , n29134 );
xor ( n39808 , n39807 , n27936 );
and ( n39809 , n39806 , n39808 );
xor ( n39810 , n37778 , n39809 );
xor ( n39811 , n39805 , n39810 );
xor ( n39812 , n39811 , n37755 );
not ( n39813 , n37797 );
and ( n39814 , n39813 , n39794 );
xor ( n39815 , n37794 , n39814 );
xor ( n39816 , n39812 , n39815 );
xor ( n39817 , n39799 , n39816 );
xor ( n39818 , n39817 , n35052 );
not ( n39819 , n39818 );
xor ( n39820 , n38128 , n31053 );
xor ( n39821 , n39820 , n35494 );
and ( n39822 , n39819 , n39821 );
xor ( n39823 , n39792 , n39822 );
not ( n12368 , n29614 );
and ( n12369 , n12368 , RI173f39b8_1568);
and ( n12370 , n39823 , n29614 );
or ( n39824 , n12369 , n12370 );
not ( n12371 , RI1754c610_2);
and ( n12372 , n12371 , n39824 );
and ( n12373 , C0 , RI1754c610_2);
or ( n39825 , n12372 , n12373 );
buf ( n39826 , n39825 );
not ( n12374 , n27683 );
and ( n12375 , n12374 , RI19a99440_2617);
and ( n12376 , RI19aa2e78_2546 , n27683 );
or ( n39827 , n12375 , n12376 );
not ( n12377 , RI1754c610_2);
and ( n12378 , n12377 , n39827 );
and ( n12379 , C0 , RI1754c610_2);
or ( n39828 , n12378 , n12379 );
buf ( n39829 , n39828 );
xor ( n39830 , n32548 , n37651 );
xor ( n39831 , n39830 , n39182 );
xor ( n39832 , n34643 , n34150 );
xor ( n39833 , n39832 , n34190 );
not ( n39834 , n39833 );
not ( n39835 , n34728 );
and ( n39836 , n39835 , n30054 );
xor ( n39837 , n36721 , n39836 );
not ( n39838 , n36721 );
and ( n39839 , n39838 , n34728 );
xor ( n39840 , n30070 , n39839 );
not ( n39841 , n30031 );
and ( n39842 , n39841 , n34733 );
xor ( n39843 , n30018 , n39842 );
xor ( n39844 , n39840 , n39843 );
not ( n39845 , n36727 );
and ( n39846 , n39845 , n34739 );
xor ( n39847 , n30152 , n39846 );
xor ( n39848 , n39844 , n39847 );
not ( n39849 , n36733 );
and ( n39850 , n39849 , n34745 );
xor ( n39851 , n30194 , n39850 );
xor ( n39852 , n39848 , n39851 );
not ( n39853 , n36739 );
and ( n39854 , n39853 , n34751 );
xor ( n39855 , n30244 , n39854 );
xor ( n39856 , n39852 , n39855 );
xor ( n39857 , n39837 , n39856 );
xor ( n39858 , n28897 , n30007 );
xor ( n39859 , n39858 , n30017 );
not ( n39860 , n39859 );
and ( n39861 , n39860 , n35284 );
xor ( n39862 , n30258 , n39861 );
xor ( n39863 , n29717 , n28839 );
xor ( n39864 , n39863 , n28917 );
not ( n39865 , n39864 );
and ( n39866 , n39865 , n35289 );
xor ( n39867 , n30333 , n39866 );
xor ( n39868 , n39862 , n39867 );
xor ( n39869 , n29903 , n32091 );
xor ( n39870 , n39869 , n30139 );
not ( n39871 , n39870 );
and ( n39872 , n39871 , n35295 );
xor ( n39873 , n30375 , n39872 );
xor ( n39874 , n39868 , n39873 );
xor ( n39875 , n28443 , n29975 );
xor ( n39876 , n39875 , n28759 );
not ( n39877 , n39876 );
and ( n39878 , n39877 , n35301 );
xor ( n39879 , n30428 , n39878 );
xor ( n39880 , n39874 , n39879 );
xor ( n39881 , n29566 , n32611 );
xor ( n39882 , n39881 , n29161 );
not ( n39883 , n39882 );
and ( n39884 , n39883 , n35307 );
xor ( n39885 , n30458 , n39884 );
xor ( n39886 , n39880 , n39885 );
xor ( n39887 , n39857 , n39886 );
and ( n39888 , n39834 , n39887 );
xor ( n39889 , n39831 , n39888 );
not ( n12380 , n29614 );
and ( n12381 , n12380 , RI173fe458_1516);
and ( n12382 , n39889 , n29614 );
or ( n39890 , n12381 , n12382 );
not ( n12383 , RI1754c610_2);
and ( n12384 , n12383 , n39890 );
and ( n12385 , C0 , RI1754c610_2);
or ( n39891 , n12384 , n12385 );
buf ( n39892 , n39891 );
xor ( n39893 , n38316 , n38872 );
xor ( n39894 , n39893 , n38886 );
xor ( n39895 , n39054 , n39702 );
not ( n39896 , n33345 );
and ( n39897 , n39896 , n35769 );
xor ( n39898 , n33342 , n39897 );
not ( n39899 , n33354 );
and ( n39900 , n39899 , n35776 );
xor ( n39901 , n33351 , n39900 );
xor ( n39902 , n39898 , n39901 );
not ( n39903 , n33364 );
and ( n39904 , n39903 , n35784 );
xor ( n39905 , n33361 , n39904 );
xor ( n39906 , n39902 , n39905 );
not ( n39907 , n33374 );
and ( n39908 , n39907 , n35790 );
xor ( n39909 , n33371 , n39908 );
xor ( n39910 , n39906 , n39909 );
not ( n39911 , n33394 );
and ( n39912 , n39911 , n35798 );
xor ( n39913 , n33391 , n39912 );
xor ( n39914 , n39910 , n39913 );
xor ( n39915 , n39895 , n39914 );
not ( n39916 , n39915 );
not ( n39917 , n31529 );
and ( n39918 , n39917 , n31531 );
xor ( n39919 , n34306 , n39918 );
not ( n39920 , n31539 );
and ( n39921 , n39920 , n31543 );
xor ( n39922 , n34313 , n39921 );
xor ( n39923 , n39919 , n39922 );
not ( n39924 , n31560 );
and ( n39925 , n39924 , n31562 );
xor ( n39926 , n34321 , n39925 );
xor ( n39927 , n39923 , n39926 );
not ( n39928 , n31571 );
and ( n39929 , n39928 , n31582 );
xor ( n39930 , n34329 , n39929 );
xor ( n39931 , n39927 , n39930 );
not ( n39932 , n31600 );
and ( n39933 , n39932 , n31615 );
xor ( n39934 , n34337 , n39933 );
xor ( n39935 , n39931 , n39934 );
xor ( n39936 , n31597 , n39935 );
not ( n39937 , n35238 );
and ( n39938 , n39937 , n35220 );
xor ( n39939 , n38696 , n39938 );
xor ( n39940 , n38689 , n39939 );
not ( n39941 , n35244 );
and ( n39942 , n39941 , n35246 );
xor ( n39943 , n38704 , n39942 );
xor ( n39944 , n39940 , n39943 );
not ( n39945 , n35254 );
and ( n39946 , n39945 , n35256 );
xor ( n39947 , n38712 , n39946 );
xor ( n39948 , n39944 , n39947 );
not ( n39949 , n35264 );
and ( n39950 , n39949 , n35266 );
xor ( n39951 , n38720 , n39950 );
xor ( n39952 , n39948 , n39951 );
xor ( n39953 , n39936 , n39952 );
and ( n39954 , n39916 , n39953 );
xor ( n39955 , n39894 , n39954 );
not ( n12386 , n29614 );
and ( n12387 , n12386 , RI173964a8_2023);
and ( n12388 , n39955 , n29614 );
or ( n39956 , n12387 , n12388 );
not ( n12389 , RI1754c610_2);
and ( n12390 , n12389 , n39956 );
and ( n12391 , C0 , RI1754c610_2);
or ( n39957 , n12390 , n12391 );
buf ( n39958 , n39957 );
xor ( n39959 , n33974 , n34221 );
xor ( n39960 , n39959 , n34251 );
xor ( n39961 , n32990 , n30415 );
xor ( n39962 , n39961 , n30427 );
not ( n39963 , n34352 );
and ( n39964 , n39963 , n34354 );
xor ( n39965 , n39962 , n39964 );
xor ( n39966 , n30188 , n29923 );
xor ( n39967 , n39966 , n29935 );
not ( n39968 , n34361 );
and ( n39969 , n39968 , n34363 );
xor ( n39970 , n39967 , n39969 );
xor ( n39971 , n39965 , n39970 );
xor ( n39972 , n33897 , n28015 );
xor ( n39973 , n39972 , n28027 );
not ( n39974 , n34371 );
and ( n39975 , n39974 , n34373 );
xor ( n39976 , n39973 , n39975 );
xor ( n39977 , n39971 , n39976 );
xor ( n39978 , n32198 , n29793 );
xor ( n39979 , n39978 , n31909 );
not ( n39980 , n34381 );
and ( n39981 , n39980 , n34343 );
xor ( n39982 , n39979 , n39981 );
xor ( n39983 , n39977 , n39982 );
xor ( n39984 , n30388 , n28812 );
xor ( n39985 , n39984 , n29855 );
not ( n39986 , n34387 );
and ( n39987 , n39986 , n34389 );
xor ( n39988 , n39985 , n39987 );
xor ( n39989 , n39983 , n39988 );
xor ( n39990 , n34384 , n39989 );
not ( n39991 , n34398 );
and ( n39992 , n39991 , n34400 );
xor ( n39993 , n37957 , n39992 );
not ( n39994 , n34407 );
and ( n39995 , n39994 , n34409 );
xor ( n39996 , n37964 , n39995 );
xor ( n39997 , n39993 , n39996 );
not ( n39998 , n34417 );
and ( n39999 , n39998 , n34419 );
xor ( n40000 , n37972 , n39999 );
xor ( n40001 , n39997 , n40000 );
not ( n40002 , n34427 );
and ( n40003 , n40002 , n34429 );
xor ( n40004 , n37949 , n40003 );
xor ( n40005 , n40001 , n40004 );
not ( n40006 , n34437 );
and ( n40007 , n40006 , n34439 );
xor ( n40008 , n37984 , n40007 );
xor ( n40009 , n40005 , n40008 );
xor ( n40010 , n39990 , n40009 );
not ( n40011 , n40010 );
not ( n40012 , n29188 );
and ( n40013 , n40012 , n29212 );
xor ( n40014 , n34973 , n40013 );
or ( n40015 , n39583 , RI17537fd0_593);
or ( n40016 , n40015 , RI175373a0_595);
or ( n40017 , n40016 , RI17536d88_596);
xor ( n40018 , n40014 , n40017 );
not ( n40019 , n29249 );
and ( n40020 , n40019 , n29271 );
xor ( n40021 , n34984 , n40020 );
xor ( n40022 , n40018 , n40021 );
not ( n40023 , n29292 );
and ( n40024 , n40023 , n29135 );
xor ( n40025 , n34990 , n40024 );
xor ( n40026 , n40022 , n40025 );
not ( n40027 , n29308 );
and ( n40028 , n40027 , n29333 );
xor ( n40029 , n34998 , n40028 );
xor ( n40030 , n40026 , n40029 );
not ( n40031 , n29376 );
and ( n40032 , n40031 , n29400 );
xor ( n40033 , n35006 , n40032 );
xor ( n40034 , n40030 , n40033 );
xor ( n40035 , n29424 , n40034 );
not ( n40036 , n28521 );
and ( n40037 , n40036 , n29503 );
xor ( n40038 , n28506 , n40037 );
xor ( n40039 , n38558 , n40038 );
not ( n40040 , n29521 );
and ( n40041 , n40040 , n29545 );
xor ( n40042 , n28685 , n40041 );
xor ( n40043 , n40039 , n40042 );
not ( n40044 , n29574 );
and ( n40045 , n40044 , n29588 );
xor ( n40046 , n28743 , n40045 );
xor ( n40047 , n40043 , n40046 );
not ( n40048 , n29603 );
and ( n40049 , n40048 , n29606 );
xor ( n40050 , n28813 , n40049 );
xor ( n40051 , n40047 , n40050 );
xor ( n40052 , n40035 , n40051 );
and ( n40053 , n40011 , n40052 );
xor ( n40054 , n39960 , n40053 );
not ( n12392 , n29614 );
and ( n12393 , n12392 , RI174a09b0_953);
and ( n12394 , n40054 , n29614 );
or ( n40055 , n12393 , n12394 );
not ( n12395 , RI1754c610_2);
and ( n12396 , n12395 , n40055 );
and ( n12397 , C0 , RI1754c610_2);
or ( n40056 , n12396 , n12397 );
buf ( n40057 , n40056 );
not ( n12398 , n27683 );
and ( n12399 , n12398 , RI19a9ca28_2593);
and ( n12400 , RI19aa62f8_2521 , n27683 );
or ( n40058 , n12399 , n12400 );
not ( n12401 , RI1754c610_2);
and ( n12402 , n12401 , n40058 );
and ( n12403 , C0 , RI1754c610_2);
or ( n40059 , n12402 , n12403 );
buf ( n40060 , n40059 );
xor ( n40061 , n36043 , n34475 );
xor ( n40062 , n40061 , n37371 );
xor ( n40063 , n34378 , n39989 );
xor ( n40064 , n40063 , n40009 );
not ( n40065 , n40064 );
not ( n40066 , n35697 );
and ( n40067 , n40066 , n35828 );
xor ( n40068 , n35694 , n40067 );
xor ( n40069 , n40068 , n35710 );
xor ( n40070 , n40069 , n35760 );
and ( n40071 , n40065 , n40070 );
xor ( n40072 , n40062 , n40071 );
not ( n12404 , n29614 );
and ( n12405 , n12404 , RI174c48d8_799);
and ( n12406 , n40072 , n29614 );
or ( n40073 , n12405 , n12406 );
not ( n12407 , RI1754c610_2);
and ( n12408 , n12407 , n40073 );
and ( n12409 , C0 , RI1754c610_2);
or ( n40074 , n12408 , n12409 );
buf ( n40075 , n40074 );
not ( n40076 , n37995 );
and ( n40077 , n40076 , n38052 );
xor ( n40078 , n37992 , n40077 );
not ( n40079 , n38004 );
and ( n40080 , n40079 , n38059 );
xor ( n40081 , n38001 , n40080 );
xor ( n40082 , n40078 , n40081 );
not ( n40083 , n38014 );
and ( n40084 , n40083 , n38045 );
xor ( n40085 , n38011 , n40084 );
xor ( n40086 , n40082 , n40085 );
xor ( n40087 , n40086 , n39723 );
not ( n40088 , n38034 );
and ( n40089 , n40088 , n38079 );
xor ( n40090 , n38031 , n40089 );
xor ( n40091 , n40087 , n40090 );
xor ( n40092 , n38064 , n40091 );
not ( n40093 , n38088 );
and ( n40094 , n40093 , n30769 );
xor ( n40095 , n39486 , n40094 );
not ( n40096 , n38093 );
and ( n40097 , n40096 , n30824 );
xor ( n40098 , n35851 , n40097 );
xor ( n40099 , n40095 , n40098 );
not ( n40100 , n38099 );
and ( n40101 , n40100 , n30843 );
xor ( n40102 , n39496 , n40101 );
xor ( n40103 , n40099 , n40102 );
not ( n40104 , n38105 );
and ( n40105 , n40104 , n30877 );
xor ( n40106 , n39502 , n40105 );
xor ( n40107 , n40103 , n40106 );
not ( n40108 , n38111 );
and ( n40109 , n40108 , n30919 );
xor ( n40110 , n30765 , n40109 );
xor ( n40111 , n40107 , n40110 );
xor ( n40112 , n40092 , n40111 );
not ( n40113 , n34739 );
and ( n40114 , n40113 , n30102 );
xor ( n40115 , n36727 , n40114 );
xor ( n40116 , n40115 , n39856 );
xor ( n40117 , n40116 , n39886 );
not ( n40118 , n40117 );
xor ( n40119 , n39260 , n35361 );
xor ( n40120 , n40119 , n38445 );
and ( n40121 , n40118 , n40120 );
xor ( n40122 , n40112 , n40121 );
not ( n12410 , n29614 );
and ( n12411 , n12410 , RI17455f50_1317);
and ( n12412 , n40122 , n29614 );
or ( n40123 , n12411 , n12412 );
not ( n12413 , RI1754c610_2);
and ( n12414 , n12413 , n40123 );
and ( n12415 , C0 , RI1754c610_2);
or ( n40124 , n12414 , n12415 );
buf ( n40125 , n40124 );
not ( n40126 , n33522 );
and ( n40127 , n40126 , n33524 );
xor ( n40128 , n34766 , n40127 );
xor ( n40129 , n40128 , n34797 );
xor ( n40130 , n40129 , n34837 );
not ( n40131 , n37626 );
and ( n40132 , n40131 , n32515 );
xor ( n40133 , n32511 , n40132 );
not ( n40134 , n37631 );
and ( n40135 , n40134 , n32520 );
xor ( n40136 , n36903 , n40135 );
xor ( n40137 , n40133 , n40136 );
not ( n40138 , n36898 );
and ( n40139 , n40138 , n32531 );
xor ( n40140 , n36895 , n40139 );
xor ( n40141 , n40137 , n40140 );
not ( n40142 , n37641 );
and ( n40143 , n40142 , n32541 );
xor ( n40144 , n36020 , n40143 );
xor ( n40145 , n40141 , n40144 );
not ( n40146 , n37647 );
and ( n40147 , n40146 , n32552 );
xor ( n40148 , n36914 , n40147 );
xor ( n40149 , n40145 , n40148 );
xor ( n40150 , n37634 , n40149 );
not ( n40151 , n39015 );
and ( n40152 , n40151 , n32563 );
xor ( n40153 , n36921 , n40152 );
not ( n40154 , n39020 );
and ( n40155 , n40154 , n32572 );
xor ( n40156 , n36926 , n40155 );
xor ( n40157 , n40153 , n40156 );
xor ( n40158 , n40157 , n39012 );
not ( n40159 , n39030 );
and ( n40160 , n40159 , n32592 );
xor ( n40161 , n36938 , n40160 );
xor ( n40162 , n40158 , n40161 );
not ( n40163 , n39036 );
and ( n40164 , n40163 , n32612 );
xor ( n40165 , n36944 , n40164 );
xor ( n40166 , n40162 , n40165 );
xor ( n40167 , n40150 , n40166 );
not ( n40168 , n40167 );
xor ( n40169 , n37860 , n35128 );
xor ( n40170 , n40169 , n36917 );
and ( n40171 , n40168 , n40170 );
xor ( n40172 , n40130 , n40171 );
not ( n12416 , n29614 );
and ( n12417 , n12416 , RI17468358_1228);
and ( n12418 , n40172 , n29614 );
or ( n40173 , n12417 , n12418 );
not ( n12419 , RI1754c610_2);
and ( n12420 , n12419 , n40173 );
and ( n12421 , C0 , RI1754c610_2);
or ( n40174 , n12420 , n12421 );
buf ( n40175 , n40174 );
xor ( n40176 , n37355 , n33505 );
xor ( n40177 , n40176 , n39635 );
not ( n40178 , n33962 );
and ( n40179 , n40178 , n36267 );
xor ( n40180 , n33959 , n40179 );
xor ( n40181 , n35654 , n40180 );
not ( n40182 , n33972 );
and ( n40183 , n40182 , n36273 );
xor ( n40184 , n33969 , n40183 );
xor ( n40185 , n40181 , n40184 );
xor ( n40186 , n40185 , n33946 );
not ( n40187 , n33988 );
and ( n40188 , n40187 , n36283 );
xor ( n40189 , n33985 , n40188 );
xor ( n40190 , n40186 , n40189 );
xor ( n40191 , n37298 , n40190 );
not ( n40192 , n33999 );
and ( n40193 , n40192 , n37499 );
xor ( n40194 , n33996 , n40193 );
not ( n40195 , n34008 );
and ( n40196 , n40195 , n37504 );
xor ( n40197 , n34005 , n40196 );
xor ( n40198 , n40194 , n40197 );
not ( n40199 , n34018 );
and ( n40200 , n40199 , n37510 );
xor ( n40201 , n34015 , n40200 );
xor ( n40202 , n40198 , n40201 );
not ( n40203 , n34028 );
and ( n40204 , n40203 , n37516 );
xor ( n40205 , n34025 , n40204 );
xor ( n40206 , n40202 , n40205 );
not ( n40207 , n34038 );
and ( n40208 , n40207 , n37522 );
xor ( n40209 , n34035 , n40208 );
xor ( n40210 , n40206 , n40209 );
xor ( n40211 , n40191 , n40210 );
not ( n40212 , n40211 );
not ( n40213 , n34105 );
and ( n40214 , n40213 , n34107 );
xor ( n40215 , n33912 , n40214 );
xor ( n40216 , n40215 , n36431 );
xor ( n40217 , n40216 , n34221 );
and ( n40218 , n40212 , n40217 );
xor ( n40219 , n40177 , n40218 );
not ( n12422 , n29614 );
and ( n12423 , n12422 , RI1746d8a8_1202);
and ( n12424 , n40219 , n29614 );
or ( n40220 , n12423 , n12424 );
not ( n12425 , RI1754c610_2);
and ( n12426 , n12425 , n40220 );
and ( n12427 , C0 , RI1754c610_2);
or ( n40221 , n12426 , n12427 );
buf ( n40222 , n40221 );
buf ( n40223 , RI174ace90_893);
buf ( n40224 , RI174a6590_925);
not ( n40225 , n35672 );
and ( n40226 , n40225 , n35807 );
xor ( n40227 , n35669 , n40226 );
xor ( n40228 , n40227 , n35665 );
not ( n40229 , n35687 );
and ( n40230 , n40229 , n35820 );
xor ( n40231 , n35684 , n40230 );
xor ( n40232 , n40228 , n40231 );
xor ( n40233 , n40232 , n40068 );
not ( n40234 , n35707 );
and ( n40235 , n40234 , n35836 );
xor ( n40236 , n35704 , n40235 );
xor ( n40237 , n40233 , n40236 );
xor ( n40238 , n37124 , n40237 );
not ( n40239 , n35718 );
and ( n40240 , n40239 , n37132 );
xor ( n40241 , n35715 , n40240 );
not ( n40242 , n35727 );
and ( n40243 , n40242 , n37139 );
xor ( n40244 , n35724 , n40243 );
xor ( n40245 , n40241 , n40244 );
not ( n40246 , n35737 );
and ( n40247 , n40246 , n37147 );
xor ( n40248 , n35734 , n40247 );
xor ( n40249 , n40245 , n40248 );
not ( n40250 , n35747 );
and ( n40251 , n40250 , n37155 );
xor ( n40252 , n35744 , n40251 );
xor ( n40253 , n40249 , n40252 );
xor ( n40254 , n40253 , n39745 );
xor ( n40255 , n40238 , n40254 );
xor ( n40256 , n32047 , n36682 );
xor ( n40257 , n40256 , n36702 );
not ( n40258 , n40257 );
xor ( n40259 , n37663 , n37549 );
xor ( n40260 , n40259 , n37579 );
and ( n40261 , n40258 , n40260 );
xor ( n40262 , n40255 , n40261 );
not ( n12428 , n29614 );
and ( n12429 , n12428 , RI173f0880_1583);
and ( n12430 , n40262 , n29614 );
or ( n40263 , n12429 , n12430 );
not ( n12431 , RI1754c610_2);
and ( n12432 , n12431 , n40263 );
and ( n12433 , C0 , RI1754c610_2);
or ( n40264 , n12432 , n12433 );
buf ( n40265 , n40264 );
xor ( n40266 , n39454 , n36611 );
xor ( n40267 , n40266 , n33567 );
not ( n40268 , n35081 );
and ( n40269 , n40268 , n35083 );
xor ( n40270 , n37590 , n40269 );
not ( n40271 , n35090 );
and ( n40272 , n40271 , n35092 );
xor ( n40273 , n37597 , n40272 );
xor ( n40274 , n40270 , n40273 );
xor ( n40275 , n40274 , n37586 );
not ( n40276 , n35110 );
and ( n40277 , n40276 , n35112 );
xor ( n40278 , n37611 , n40277 );
xor ( n40279 , n40275 , n40278 );
not ( n40280 , n35120 );
and ( n40281 , n40280 , n35122 );
xor ( n40282 , n37619 , n40281 );
xor ( n40283 , n40279 , n40282 );
xor ( n40284 , n35097 , n40283 );
xor ( n40285 , n40284 , n32560 );
not ( n40286 , n40285 );
not ( n40287 , n33235 );
and ( n40288 , n40287 , n33237 );
xor ( n40289 , n33654 , n40288 );
not ( n40290 , n33244 );
and ( n40291 , n40290 , n33246 );
xor ( n40292 , n33670 , n40291 );
xor ( n40293 , n40289 , n40292 );
xor ( n40294 , n40293 , n37833 );
not ( n40295 , n33264 );
and ( n40296 , n40295 , n33266 );
xor ( n40297 , n33686 , n40296 );
xor ( n40298 , n40294 , n40297 );
not ( n40299 , n33274 );
and ( n40300 , n40299 , n33276 );
xor ( n40301 , n33694 , n40300 );
xor ( n40302 , n40298 , n40301 );
xor ( n40303 , n33261 , n40302 );
not ( n40304 , n37595 );
and ( n40305 , n40304 , n37597 );
xor ( n40306 , n35095 , n40305 );
xor ( n40307 , n38937 , n40306 );
not ( n40308 , n37603 );
and ( n40309 , n40308 , n37583 );
xor ( n40310 , n35105 , n40309 );
xor ( n40311 , n40307 , n40310 );
not ( n40312 , n37609 );
and ( n40313 , n40312 , n37611 );
xor ( n40314 , n35115 , n40313 );
xor ( n40315 , n40311 , n40314 );
not ( n40316 , n37617 );
and ( n40317 , n40316 , n37619 );
xor ( n40318 , n35125 , n40317 );
xor ( n40319 , n40315 , n40318 );
xor ( n40320 , n40303 , n40319 );
and ( n40321 , n40286 , n40320 );
xor ( n40322 , n40267 , n40321 );
not ( n12434 , n29614 );
and ( n12435 , n12434 , RI17468010_1229);
and ( n12436 , n40322 , n29614 );
or ( n40323 , n12435 , n12436 );
not ( n12437 , RI1754c610_2);
and ( n12438 , n12437 , n40323 );
and ( n12439 , C0 , RI1754c610_2);
or ( n40324 , n12438 , n12439 );
buf ( n40325 , n40324 );
not ( n40326 , n37957 );
and ( n40327 , n40326 , n34398 );
xor ( n40328 , n37954 , n40327 );
not ( n40329 , n37964 );
and ( n40330 , n40329 , n34407 );
xor ( n40331 , n37961 , n40330 );
xor ( n40332 , n40328 , n40331 );
not ( n40333 , n37972 );
and ( n40334 , n40333 , n34417 );
xor ( n40335 , n37969 , n40334 );
xor ( n40336 , n40332 , n40335 );
xor ( n40337 , n40336 , n37952 );
not ( n40338 , n37984 );
and ( n40339 , n40338 , n34437 );
xor ( n40340 , n37981 , n40339 );
xor ( n40341 , n40337 , n40340 );
xor ( n40342 , n40004 , n40341 );
xor ( n40343 , n40342 , n40091 );
xor ( n40344 , n33452 , n36252 );
not ( n40345 , n33456 );
and ( n40346 , n40345 , n33460 );
xor ( n40347 , n36068 , n40346 );
not ( n40348 , n33467 );
and ( n40349 , n40348 , n33469 );
xor ( n40350 , n36075 , n40349 );
xor ( n40351 , n40347 , n40350 );
not ( n40352 , n33477 );
and ( n40353 , n40352 , n33479 );
xor ( n40354 , n36083 , n40353 );
xor ( n40355 , n40351 , n40354 );
not ( n40356 , n33487 );
and ( n40357 , n40356 , n33489 );
xor ( n40358 , n36091 , n40357 );
xor ( n40359 , n40355 , n40358 );
xor ( n40360 , n40359 , n37879 );
xor ( n40361 , n40344 , n40360 );
not ( n40362 , n40361 );
not ( n40363 , n36487 );
and ( n40364 , n40363 , n36478 );
xor ( n40365 , n37387 , n40364 );
not ( n40366 , n36492 );
and ( n40367 , n40366 , n36494 );
xor ( n40368 , n37394 , n40367 );
xor ( n40369 , n40365 , n40368 );
not ( n40370 , n36502 );
and ( n40371 , n40370 , n36504 );
xor ( n40372 , n37402 , n40371 );
xor ( n40373 , n40369 , n40372 );
not ( n40374 , n36512 );
and ( n40375 , n40374 , n36514 );
xor ( n40376 , n37410 , n40375 );
xor ( n40377 , n40373 , n40376 );
not ( n40378 , n36522 );
and ( n40379 , n40378 , n36524 );
xor ( n40380 , n37418 , n40379 );
xor ( n40381 , n40377 , n40380 );
xor ( n40382 , n36490 , n40381 );
xor ( n40383 , n40382 , n37438 );
and ( n40384 , n40362 , n40383 );
xor ( n40385 , n40343 , n40384 );
not ( n12440 , n29614 );
and ( n12441 , n12440 , RI1752b280_632);
and ( n12442 , n40385 , n29614 );
or ( n40386 , n12441 , n12442 );
not ( n12443 , RI1754c610_2);
and ( n12444 , n12443 , n40386 );
and ( n12445 , C0 , RI1754c610_2);
or ( n40387 , n12444 , n12445 );
buf ( n40388 , n40387 );
xor ( n40389 , n40140 , n38948 );
xor ( n40390 , n40389 , n39039 );
xor ( n40391 , n31893 , n36401 );
xor ( n40392 , n40391 , n33453 );
not ( n40393 , n40392 );
not ( n40394 , n32931 );
and ( n40395 , n40394 , n36617 );
xor ( n40396 , n32928 , n40395 );
not ( n40397 , n32940 );
and ( n40398 , n40397 , n36624 );
xor ( n40399 , n32937 , n40398 );
xor ( n40400 , n40396 , n40399 );
not ( n40401 , n32950 );
and ( n40402 , n40401 , n36632 );
xor ( n40403 , n32947 , n40402 );
xor ( n40404 , n40400 , n40403 );
not ( n40405 , n32960 );
and ( n40406 , n40405 , n36640 );
xor ( n40407 , n32957 , n40406 );
xor ( n40408 , n40404 , n40407 );
not ( n40409 , n32970 );
and ( n40410 , n40409 , n36648 );
xor ( n40411 , n32967 , n40410 );
xor ( n40412 , n40408 , n40411 );
xor ( n40413 , n36653 , n40412 );
not ( n40414 , n39802 );
xor ( n40415 , n31627 , n30986 );
xor ( n40416 , n40415 , n31794 );
and ( n40417 , n40414 , n40416 );
xor ( n40418 , n37762 , n40417 );
not ( n40419 , n39099 );
xor ( n40420 , n31481 , n30189 );
xor ( n40421 , n40420 , n28715 );
and ( n40422 , n40419 , n40421 );
xor ( n40423 , n37771 , n40422 );
xor ( n40424 , n40418 , n40423 );
not ( n40425 , n39808 );
xor ( n40426 , n31785 , n29148 );
xor ( n40427 , n40426 , n32800 );
and ( n40428 , n40425 , n40427 );
xor ( n40429 , n37781 , n40428 );
xor ( n40430 , n40424 , n40429 );
not ( n40431 , n37753 );
xor ( n40432 , n31155 , n27779 );
xor ( n40433 , n40432 , n27791 );
and ( n40434 , n40431 , n40433 );
xor ( n40435 , n37750 , n40434 );
xor ( n40436 , n40430 , n40435 );
xor ( n40437 , n40436 , n39799 );
xor ( n40438 , n40413 , n40437 );
and ( n40439 , n40393 , n40438 );
xor ( n40440 , n40390 , n40439 );
not ( n12446 , n29614 );
and ( n12447 , n12446 , RI17500f80_757);
and ( n12448 , n40440 , n29614 );
or ( n40441 , n12447 , n12448 );
not ( n12449 , RI1754c610_2);
and ( n12450 , n12449 , n40441 );
and ( n12451 , C0 , RI1754c610_2);
or ( n40442 , n12450 , n12451 );
buf ( n40443 , n40442 );
xor ( n40444 , n38593 , n29109 );
not ( n40445 , n35869 );
and ( n40446 , n40445 , n37077 );
xor ( n40447 , n35866 , n40446 );
not ( n40448 , n35878 );
and ( n40449 , n40448 , n37082 );
xor ( n40450 , n35875 , n40449 );
xor ( n40451 , n40447 , n40450 );
not ( n40452 , n35888 );
and ( n40453 , n40452 , n37088 );
xor ( n40454 , n35885 , n40453 );
xor ( n40455 , n40451 , n40454 );
not ( n40456 , n35898 );
and ( n40457 , n40456 , n37094 );
xor ( n40458 , n35895 , n40457 );
xor ( n40459 , n40455 , n40458 );
not ( n40460 , n35908 );
and ( n40461 , n40460 , n37100 );
xor ( n40462 , n35905 , n40461 );
xor ( n40463 , n40459 , n40462 );
xor ( n40464 , n40444 , n40463 );
xor ( n40465 , n33955 , n34221 );
xor ( n40466 , n40465 , n34251 );
not ( n40467 , n40466 );
not ( n40468 , n33731 );
and ( n40469 , n40468 , n33733 );
xor ( n40470 , n38900 , n40469 );
not ( n40471 , n33740 );
and ( n40472 , n40471 , n33742 );
xor ( n40473 , n38907 , n40472 );
xor ( n40474 , n40470 , n40473 );
not ( n40475 , n33750 );
and ( n40476 , n40475 , n33752 );
xor ( n40477 , n38915 , n40476 );
xor ( n40478 , n40474 , n40477 );
not ( n40479 , n33760 );
and ( n40480 , n40479 , n33762 );
xor ( n40481 , n38921 , n40480 );
xor ( n40482 , n40478 , n40481 );
not ( n40483 , n33770 );
and ( n40484 , n40483 , n33772 );
xor ( n40485 , n38929 , n40484 );
xor ( n40486 , n40482 , n40485 );
xor ( n40487 , n33747 , n40486 );
xor ( n40488 , n27929 , n30364 );
xor ( n40489 , n40488 , n30374 );
not ( n40490 , n38746 );
and ( n40491 , n40490 , n38748 );
xor ( n40492 , n40489 , n40491 );
xor ( n40493 , n29252 , n32120 );
xor ( n40494 , n40493 , n29093 );
not ( n40495 , n38755 );
and ( n40496 , n40495 , n38757 );
xor ( n40497 , n40494 , n40496 );
xor ( n40498 , n40492 , n40497 );
xor ( n40499 , n30894 , n32744 );
xor ( n40500 , n40499 , n33198 );
not ( n40501 , n38765 );
and ( n40502 , n40501 , n38767 );
xor ( n40503 , n40500 , n40502 );
xor ( n40504 , n40498 , n40503 );
xor ( n40505 , n31175 , n29532 );
xor ( n40506 , n40505 , n29544 );
not ( n40507 , n38775 );
and ( n40508 , n40507 , n38777 );
xor ( n40509 , n40506 , n40508 );
xor ( n40510 , n40504 , n40509 );
xor ( n40511 , n28411 , n31247 );
xor ( n40512 , n40511 , n27885 );
not ( n40513 , n38785 );
and ( n40514 , n40513 , n38787 );
xor ( n40515 , n40512 , n40514 );
xor ( n40516 , n40510 , n40515 );
xor ( n40517 , n40487 , n40516 );
and ( n40518 , n40467 , n40517 );
xor ( n40519 , n40464 , n40518 );
not ( n12452 , n29614 );
and ( n12453 , n12452 , RI17400f00_1503);
and ( n12454 , n40519 , n29614 );
or ( n40520 , n12453 , n12454 );
not ( n12455 , RI1754c610_2);
and ( n12456 , n12455 , n40520 );
and ( n12457 , C0 , RI1754c610_2);
or ( n40521 , n12456 , n12457 );
buf ( n40522 , n40521 );
xor ( n40523 , n32646 , n36195 );
xor ( n40524 , n40523 , n36209 );
xor ( n40525 , n32769 , n37186 );
xor ( n40526 , n40525 , n37203 );
not ( n40527 , n40526 );
xor ( n40528 , n39603 , n31621 );
xor ( n40529 , n40528 , n35272 );
and ( n40530 , n40527 , n40529 );
xor ( n40531 , n40524 , n40530 );
not ( n12458 , n29614 );
and ( n12459 , n12458 , RI173a2cd0_1962);
and ( n12460 , n40531 , n29614 );
or ( n40532 , n12459 , n12460 );
not ( n12461 , RI1754c610_2);
and ( n12462 , n12461 , n40532 );
and ( n12463 , C0 , RI1754c610_2);
or ( n40533 , n12462 , n12463 );
buf ( n40534 , n40533 );
buf ( n40535 , RI174b9460_834);
not ( n12464 , n27683 );
and ( n12465 , n12464 , RI19aaeb60_2463);
and ( n12466 , RI19ab8958_2391 , n27683 );
or ( n40536 , n12465 , n12466 );
not ( n12467 , RI1754c610_2);
and ( n12468 , n12467 , n40536 );
and ( n12469 , C0 , RI1754c610_2);
or ( n40537 , n12468 , n12469 );
buf ( n40538 , n40537 );
not ( n12470 , n27683 );
and ( n12471 , n12470 , RI19aaad80_2489);
and ( n12472 , RI19ab4bf0_2418 , n27683 );
or ( n40539 , n12471 , n12472 );
not ( n12473 , RI1754c610_2);
and ( n12474 , n12473 , n40539 );
and ( n12475 , C0 , RI1754c610_2);
or ( n40540 , n12474 , n12475 );
buf ( n40541 , n40540 );
buf ( n40542 , RI174b0310_877);
xor ( n40543 , n31620 , n39935 );
xor ( n40544 , n40543 , n39952 );
not ( n40545 , n34529 );
and ( n40546 , n40545 , n34520 );
xor ( n40547 , n36814 , n40546 );
not ( n40548 , n34534 );
and ( n40549 , n40548 , n34536 );
xor ( n40550 , n36821 , n40549 );
xor ( n40551 , n40547 , n40550 );
not ( n40552 , n34544 );
and ( n40553 , n40552 , n34546 );
xor ( n40554 , n36808 , n40553 );
xor ( n40555 , n40551 , n40554 );
not ( n40556 , n34554 );
and ( n40557 , n40556 , n34556 );
xor ( n40558 , n36833 , n40557 );
xor ( n40559 , n40555 , n40558 );
not ( n40560 , n34564 );
and ( n40561 , n40560 , n34566 );
xor ( n40562 , n36841 , n40561 );
xor ( n40563 , n40559 , n40562 );
xor ( n40564 , n34532 , n40563 );
xor ( n40565 , n40564 , n35544 );
not ( n40566 , n40565 );
not ( n40567 , n37006 );
and ( n40568 , n40567 , n38408 );
xor ( n40569 , n37003 , n40568 );
not ( n40570 , n37015 );
and ( n40571 , n40570 , n38415 );
xor ( n40572 , n37012 , n40571 );
xor ( n40573 , n40569 , n40572 );
not ( n40574 , n37025 );
and ( n40575 , n40574 , n38423 );
xor ( n40576 , n37022 , n40575 );
xor ( n40577 , n40573 , n40576 );
not ( n40578 , n37035 );
and ( n40579 , n40578 , n38431 );
xor ( n40580 , n37032 , n40579 );
xor ( n40581 , n40577 , n40580 );
not ( n40582 , n37045 );
and ( n40583 , n40582 , n38439 );
xor ( n40584 , n37042 , n40583 );
xor ( n40585 , n40581 , n40584 );
xor ( n40586 , n38420 , n40585 );
xor ( n40587 , n40586 , n34918 );
and ( n40588 , n40566 , n40587 );
xor ( n40589 , n40544 , n40588 );
not ( n12476 , n29614 );
and ( n12477 , n12476 , RI174a5f00_927);
and ( n12478 , n40589 , n29614 );
or ( n40590 , n12477 , n12478 );
not ( n12479 , RI1754c610_2);
and ( n12480 , n12479 , n40590 );
and ( n12481 , C0 , RI1754c610_2);
or ( n40591 , n12480 , n12481 );
buf ( n40592 , n40591 );
buf ( n40593 , RI174a2a80_943);
xor ( n40594 , n35962 , n37744 );
xor ( n40595 , n40594 , n35438 );
not ( n40596 , n38615 );
and ( n40597 , n40596 , n38852 );
xor ( n40598 , n38314 , n40597 );
xor ( n40599 , n40598 , n38634 );
xor ( n40600 , n40599 , n38648 );
not ( n40601 , n40600 );
and ( n40602 , n40601 , n39115 );
xor ( n40603 , n40595 , n40602 );
not ( n12482 , n29614 );
and ( n12483 , n12482 , RI174b2728_866);
and ( n12484 , n40603 , n29614 );
or ( n40604 , n12483 , n12484 );
not ( n12485 , RI1754c610_2);
and ( n12486 , n12485 , n40604 );
and ( n12487 , C0 , RI1754c610_2);
or ( n40605 , n12486 , n12487 );
buf ( n40606 , n40605 );
buf ( n40607 , RI1749a0b0_985);
buf ( n40608 , RI174816f0_1105);
not ( n12488 , n27683 );
and ( n12489 , n12488 , RI19ab7530_2399);
and ( n12490 , RI19ac04a0_2329 , n27683 );
or ( n40609 , n12489 , n12490 );
not ( n12491 , RI1754c610_2);
and ( n12492 , n12491 , n40609 );
and ( n12493 , C0 , RI1754c610_2);
or ( n40610 , n12492 , n12493 );
buf ( n40611 , n40610 );
buf ( n40612 , RI174789d8_1148);
buf ( n40613 , RI1746b148_1214);
buf ( n40614 , RI17516da8_695);
not ( n40615 , n34392 );
xor ( n40616 , n29471 , n31558 );
xor ( n40617 , n40616 , n29025 );
and ( n40618 , n40615 , n40617 );
xor ( n40619 , n34389 , n40618 );
xor ( n40620 , n40619 , n34395 );
xor ( n40621 , n40620 , n34445 );
not ( n40622 , n33837 );
and ( n40623 , n40622 , n33839 );
xor ( n40624 , n34056 , n40623 );
xor ( n40625 , n40624 , n34087 );
xor ( n40626 , n40625 , n34127 );
not ( n40627 , n40626 );
not ( n40628 , n37010 );
and ( n40629 , n40628 , n37012 );
xor ( n40630 , n38418 , n40629 );
xor ( n40631 , n40630 , n39282 );
xor ( n40632 , n40631 , n37676 );
and ( n40633 , n40627 , n40632 );
xor ( n40634 , n40621 , n40633 );
not ( n12494 , n29614 );
and ( n12495 , n12494 , RI174146b8_1408);
and ( n12496 , n40634 , n29614 );
or ( n40635 , n12495 , n12496 );
not ( n12497 , RI1754c610_2);
and ( n12498 , n12497 , n40635 );
and ( n12499 , C0 , RI1754c610_2);
or ( n40636 , n12498 , n12499 );
buf ( n40637 , n40636 );
and ( n40638 , RI1754b530_38 , n34844 );
and ( n40639 , RI1754b530_38 , n34847 );
and ( n40640 , RI1754b530_38 , n34850 );
or ( n40641 , n40638 , n40639 , n40640 , C0 , C0 , C0 , C0 , C0 );
not ( n12500 , n34859 );
and ( n12501 , n12500 , n40641 );
and ( n12502 , RI1754b530_38 , n34859 );
or ( n40642 , n12501 , n12502 );
not ( n12503 , RI19a22f70_2797);
and ( n12504 , n12503 , n40642 );
and ( n12505 , C0 , RI19a22f70_2797);
or ( n40643 , n12504 , n12505 );
not ( n12506 , n27683 );
and ( n12507 , n12506 , RI19ab54d8_2414);
and ( n12508 , n40643 , n27683 );
or ( n40644 , n12507 , n12508 );
not ( n12509 , RI1754c610_2);
and ( n12510 , n12509 , n40644 );
and ( n12511 , C0 , RI1754c610_2);
or ( n40645 , n12510 , n12511 );
buf ( n40646 , n40645 );
not ( n40647 , n37001 );
and ( n40648 , n40647 , n37003 );
xor ( n40649 , n38411 , n40648 );
xor ( n40650 , n40649 , n40630 );
not ( n40651 , n37020 );
and ( n40652 , n40651 , n37022 );
xor ( n40653 , n38426 , n40652 );
xor ( n40654 , n40650 , n40653 );
not ( n40655 , n37030 );
and ( n40656 , n40655 , n37032 );
xor ( n40657 , n38434 , n40656 );
xor ( n40658 , n40654 , n40657 );
not ( n40659 , n37040 );
and ( n40660 , n40659 , n37042 );
xor ( n40661 , n38442 , n40660 );
xor ( n40662 , n40658 , n40661 );
xor ( n40663 , n37008 , n40662 );
xor ( n40664 , n40663 , n39208 );
xor ( n40665 , n40180 , n33991 );
xor ( n40666 , n40665 , n34041 );
not ( n40667 , n40666 );
and ( n40668 , n40667 , n37870 );
xor ( n40669 , n40664 , n40668 );
not ( n12512 , n29614 );
and ( n12513 , n12512 , RI173d3348_1726);
and ( n12514 , n40669 , n29614 );
or ( n40670 , n12513 , n12514 );
not ( n12515 , RI1754c610_2);
and ( n12516 , n12515 , n40670 );
and ( n12517 , C0 , RI1754c610_2);
or ( n40671 , n12516 , n12517 );
buf ( n40672 , n40671 );
xor ( n40673 , n38548 , n35458 );
not ( n40674 , n36620 );
and ( n40675 , n40674 , n32926 );
xor ( n40676 , n36617 , n40675 );
not ( n40677 , n36627 );
and ( n40678 , n40677 , n32935 );
xor ( n40679 , n36624 , n40678 );
xor ( n40680 , n40676 , n40679 );
not ( n40681 , n36635 );
and ( n40682 , n40681 , n32945 );
xor ( n40683 , n36632 , n40682 );
xor ( n40684 , n40680 , n40683 );
not ( n40685 , n36643 );
and ( n40686 , n40685 , n32955 );
xor ( n40687 , n36640 , n40686 );
xor ( n40688 , n40684 , n40687 );
not ( n40689 , n36651 );
and ( n40690 , n40689 , n32965 );
xor ( n40691 , n36648 , n40690 );
xor ( n40692 , n40688 , n40691 );
xor ( n40693 , n40673 , n40692 );
not ( n40694 , n38790 );
xor ( n40695 , n29179 , n28827 );
xor ( n40696 , n40695 , n28839 );
and ( n40697 , n40694 , n40696 );
xor ( n40698 , n38787 , n40697 );
xor ( n40699 , n40698 , n38793 );
xor ( n40700 , n40699 , n40563 );
not ( n40701 , n40700 );
xor ( n40702 , n37137 , n40254 );
not ( n40703 , n36306 );
and ( n40704 , n40703 , n36308 );
xor ( n40705 , n35378 , n40704 );
not ( n40706 , n36313 );
and ( n40707 , n40706 , n36315 );
xor ( n40708 , n35387 , n40707 );
xor ( n40709 , n40705 , n40708 );
not ( n40710 , n36321 );
and ( n40711 , n40710 , n36301 );
xor ( n40712 , n35397 , n40711 );
xor ( n40713 , n40709 , n40712 );
not ( n40714 , n36327 );
and ( n40715 , n40714 , n36329 );
xor ( n40716 , n35407 , n40715 );
xor ( n40717 , n40713 , n40716 );
xor ( n40718 , n40717 , n39320 );
xor ( n40719 , n40702 , n40718 );
and ( n40720 , n40701 , n40719 );
xor ( n40721 , n40693 , n40720 );
not ( n12518 , n29614 );
and ( n12519 , n12518 , RI173fca18_1524);
and ( n12520 , n40721 , n29614 );
or ( n40722 , n12519 , n12520 );
not ( n12521 , RI1754c610_2);
and ( n12522 , n12521 , n40722 );
and ( n12523 , C0 , RI1754c610_2);
or ( n40723 , n12522 , n12523 );
buf ( n40724 , n40723 );
xor ( n40725 , n33201 , n31317 );
xor ( n40726 , n40725 , n40302 );
xor ( n40727 , n33046 , n36227 );
not ( n40728 , n31848 );
and ( n40729 , n40728 , n34153 );
xor ( n40730 , n31845 , n40729 );
not ( n40731 , n31858 );
and ( n40732 , n40731 , n34160 );
xor ( n40733 , n31855 , n40732 );
xor ( n40734 , n40730 , n40733 );
not ( n40735 , n31881 );
and ( n40736 , n40735 , n34168 );
xor ( n40737 , n31878 , n40736 );
xor ( n40738 , n40734 , n40737 );
not ( n40739 , n31891 );
and ( n40740 , n40739 , n34176 );
xor ( n40741 , n31888 , n40740 );
xor ( n40742 , n40738 , n40741 );
xor ( n40743 , n40742 , n34450 );
xor ( n40744 , n40727 , n40743 );
not ( n40745 , n40744 );
xor ( n40746 , n34660 , n32863 );
xor ( n40747 , n40746 , n34644 );
and ( n40748 , n40745 , n40747 );
xor ( n40749 , n40726 , n40748 );
not ( n12524 , n29614 );
and ( n12525 , n12524 , RI17462e08_1254);
and ( n12526 , n40749 , n29614 );
or ( n40750 , n12525 , n12526 );
not ( n12527 , RI1754c610_2);
and ( n12528 , n12527 , n40750 );
and ( n12529 , C0 , RI1754c610_2);
or ( n40751 , n12528 , n12529 );
buf ( n40752 , n40751 );
xor ( n40753 , n31686 , n30741 );
not ( n40754 , n33736 );
and ( n40755 , n40754 , n38898 );
xor ( n40756 , n33733 , n40755 );
not ( n40757 , n33745 );
and ( n40758 , n40757 , n38905 );
xor ( n40759 , n33742 , n40758 );
xor ( n40760 , n40756 , n40759 );
not ( n40761 , n33755 );
and ( n40762 , n40761 , n38913 );
xor ( n40763 , n33752 , n40762 );
xor ( n40764 , n40760 , n40763 );
xor ( n40765 , n40764 , n38743 );
not ( n40766 , n33775 );
and ( n40767 , n40766 , n38927 );
xor ( n40768 , n33772 , n40767 );
xor ( n40769 , n40765 , n40768 );
xor ( n40770 , n40753 , n40769 );
xor ( n40771 , n36324 , n40718 );
xor ( n40772 , n40771 , n38676 );
not ( n40773 , n40772 );
not ( n40774 , n34707 );
and ( n40775 , n40774 , n34709 );
xor ( n40776 , n36557 , n40775 );
xor ( n40777 , n40776 , n38284 );
xor ( n40778 , n40777 , n39856 );
and ( n40779 , n40773 , n40778 );
xor ( n40780 , n40770 , n40779 );
not ( n12530 , n29614 );
and ( n12531 , n12530 , RI173d50d0_1717);
and ( n12532 , n40780 , n29614 );
or ( n40781 , n12531 , n12532 );
not ( n12533 , RI1754c610_2);
and ( n12534 , n12533 , n40781 );
and ( n12535 , C0 , RI1754c610_2);
or ( n40782 , n12534 , n12535 );
buf ( n40783 , n40782 );
not ( n12536 , n27683 );
and ( n12537 , n12536 , RI19ac25e8_2311);
and ( n12538 , RI19acb648_2244 , n27683 );
or ( n40784 , n12537 , n12538 );
not ( n12539 , RI1754c610_2);
and ( n12540 , n12539 , n40784 );
and ( n12541 , C0 , RI1754c610_2);
or ( n40785 , n12540 , n12541 );
buf ( n40786 , n40785 );
not ( n40787 , n37792 );
and ( n40788 , n40787 , n37794 );
xor ( n40789 , n39797 , n40788 );
not ( n40790 , n40416 );
and ( n40791 , n40790 , n37757 );
xor ( n40792 , n39802 , n40791 );
not ( n40793 , n40421 );
and ( n40794 , n40793 , n37766 );
xor ( n40795 , n39099 , n40794 );
xor ( n40796 , n40792 , n40795 );
not ( n40797 , n40427 );
and ( n40798 , n40797 , n37776 );
xor ( n40799 , n39808 , n40798 );
xor ( n40800 , n40796 , n40799 );
not ( n40801 , n40433 );
and ( n40802 , n40801 , n37786 );
xor ( n40803 , n37753 , n40802 );
xor ( n40804 , n40800 , n40803 );
not ( n40805 , n39797 );
and ( n40806 , n40805 , n37792 );
xor ( n40807 , n39794 , n40806 );
xor ( n40808 , n40804 , n40807 );
xor ( n40809 , n40789 , n40808 );
not ( n40810 , n31116 );
and ( n40811 , n40810 , n31077 );
xor ( n40812 , n35022 , n40811 );
not ( n40813 , n31132 );
and ( n40814 , n40813 , n31135 );
xor ( n40815 , n35016 , n40814 );
xor ( n40816 , n40812 , n40815 );
not ( n40817 , n31163 );
and ( n40818 , n40817 , n31165 );
xor ( n40819 , n35033 , n40818 );
xor ( n40820 , n40816 , n40819 );
not ( n40821 , n31193 );
and ( n40822 , n40821 , n31195 );
xor ( n40823 , n35041 , n40822 );
xor ( n40824 , n40820 , n40823 );
not ( n40825 , n31203 );
and ( n40826 , n40825 , n31206 );
xor ( n40827 , n35049 , n40826 );
xor ( n40828 , n40824 , n40827 );
xor ( n40829 , n40809 , n40828 );
xor ( n40830 , n31850 , n36401 );
xor ( n40831 , n40830 , n33453 );
not ( n40832 , n40831 );
and ( n40833 , n40832 , n39894 );
xor ( n40834 , n40829 , n40833 );
not ( n12542 , n29614 );
and ( n12543 , n12542 , RI173c1f90_1810);
and ( n12544 , n40834 , n29614 );
or ( n40835 , n12543 , n12544 );
not ( n12545 , RI1754c610_2);
and ( n12546 , n12545 , n40835 );
and ( n12547 , C0 , RI1754c610_2);
or ( n40836 , n12546 , n12547 );
buf ( n40837 , n40836 );
xor ( n40838 , n32619 , n39182 );
xor ( n40839 , n40838 , n38991 );
not ( n40840 , n34984 );
and ( n40841 , n40840 , n29249 );
xor ( n40842 , n34981 , n40841 );
xor ( n40843 , n34976 , n40842 );
not ( n40844 , n34990 );
and ( n40845 , n40844 , n29292 );
xor ( n40846 , n29163 , n40845 );
xor ( n40847 , n40843 , n40846 );
not ( n40848 , n34998 );
and ( n40849 , n40848 , n29308 );
xor ( n40850 , n34995 , n40849 );
xor ( n40851 , n40847 , n40850 );
not ( n40852 , n35006 );
and ( n40853 , n40852 , n29376 );
xor ( n40854 , n35003 , n40853 );
xor ( n40855 , n40851 , n40854 );
xor ( n40856 , n40018 , n40855 );
xor ( n40857 , n40856 , n38574 );
not ( n40858 , n40857 );
xor ( n40859 , n38157 , n35494 );
xor ( n40860 , n40859 , n35514 );
and ( n40861 , n40858 , n40860 );
xor ( n40862 , n40839 , n40861 );
not ( n12548 , n29614 );
and ( n12549 , n12548 , RI174a96c8_910);
and ( n12550 , n40862 , n29614 );
or ( n40863 , n12549 , n12550 );
not ( n12551 , RI1754c610_2);
and ( n12552 , n12551 , n40863 );
and ( n12553 , C0 , RI1754c610_2);
or ( n40864 , n12552 , n12553 );
buf ( n40865 , n40864 );
xor ( n40866 , n38243 , n39450 );
xor ( n40867 , n40866 , n39467 );
xor ( n40868 , n35674 , n39543 );
xor ( n40869 , n40868 , n39563 );
not ( n40870 , n40869 );
not ( n40871 , n31428 );
and ( n40872 , n40871 , n31430 );
xor ( n40873 , n34277 , n40872 );
xor ( n40874 , n40873 , n38648 );
not ( n40875 , n34306 );
and ( n40876 , n40875 , n31529 );
xor ( n40877 , n34303 , n40876 );
not ( n40878 , n34313 );
and ( n40879 , n40878 , n31539 );
xor ( n40880 , n34310 , n40879 );
xor ( n40881 , n40877 , n40880 );
not ( n40882 , n34321 );
and ( n40883 , n40882 , n31560 );
xor ( n40884 , n34318 , n40883 );
xor ( n40885 , n40881 , n40884 );
not ( n40886 , n34329 );
and ( n40887 , n40886 , n31571 );
xor ( n40888 , n34326 , n40887 );
xor ( n40889 , n40885 , n40888 );
xor ( n40890 , n40889 , n38797 );
xor ( n40891 , n40874 , n40890 );
and ( n40892 , n40870 , n40891 );
xor ( n40893 , n40867 , n40892 );
not ( n12554 , n29614 );
and ( n12555 , n12554 , RI1749ec28_962);
and ( n12556 , n40893 , n29614 );
or ( n40894 , n12555 , n12556 );
not ( n12557 , RI1754c610_2);
and ( n12558 , n12557 , n40894 );
and ( n12559 , C0 , RI1754c610_2);
or ( n40895 , n12558 , n12559 );
buf ( n40896 , n40895 );
xor ( n40897 , n40730 , n31925 );
xor ( n40898 , n40897 , n34475 );
not ( n40899 , n36821 );
and ( n40900 , n40899 , n34534 );
xor ( n40901 , n36818 , n40900 );
xor ( n40902 , n40901 , n36844 );
xor ( n40903 , n40902 , n36874 );
not ( n40904 , n40903 );
xor ( n40905 , n36594 , n39791 );
xor ( n40906 , n40128 , n34762 );
not ( n40907 , n33543 );
and ( n40908 , n40907 , n33545 );
xor ( n40909 , n34779 , n40908 );
xor ( n40910 , n40906 , n40909 );
xor ( n40911 , n40910 , n39471 );
not ( n40912 , n33559 );
and ( n40913 , n40912 , n33561 );
xor ( n40914 , n34793 , n40913 );
xor ( n40915 , n40911 , n40914 );
xor ( n40916 , n40905 , n40915 );
and ( n40917 , n40904 , n40916 );
xor ( n40918 , n40898 , n40917 );
not ( n12560 , n29614 );
and ( n12561 , n12560 , RI17449098_1380);
and ( n12562 , n40918 , n29614 );
or ( n40919 , n12561 , n12562 );
not ( n12563 , RI1754c610_2);
and ( n12564 , n12563 , n40919 );
and ( n12565 , C0 , RI1754c610_2);
or ( n40920 , n12564 , n12565 );
buf ( n40921 , n40920 );
not ( n40922 , n38905 );
and ( n40923 , n40922 , n38907 );
xor ( n40924 , n33745 , n40923 );
xor ( n40925 , n40924 , n40769 );
not ( n40926 , n38751 );
xor ( n40927 , n28908 , n29889 );
xor ( n40928 , n40927 , n30537 );
and ( n40929 , n40926 , n40928 );
xor ( n40930 , n38748 , n40929 );
not ( n40931 , n38760 );
xor ( n40932 , n31415 , n29332 );
xor ( n40933 , n40932 , n29814 );
and ( n40934 , n40931 , n40933 );
xor ( n40935 , n38757 , n40934 );
xor ( n40936 , n40930 , n40935 );
not ( n40937 , n38770 );
xor ( n40938 , n30528 , n29752 );
xor ( n40939 , n40938 , n27833 );
and ( n40940 , n40937 , n40939 );
xor ( n40941 , n38767 , n40940 );
xor ( n40942 , n40936 , n40941 );
not ( n40943 , n38780 );
xor ( n40944 , n30658 , n28969 );
xor ( n40945 , n40944 , n28741 );
and ( n40946 , n40943 , n40945 );
xor ( n40947 , n38777 , n40946 );
xor ( n40948 , n40942 , n40947 );
xor ( n40949 , n40948 , n40698 );
xor ( n40950 , n40925 , n40949 );
xor ( n40951 , n29548 , n40051 );
xor ( n40952 , n40951 , n37074 );
not ( n40953 , n40952 );
not ( n40954 , n36814 );
and ( n40955 , n40954 , n34529 );
xor ( n40956 , n34525 , n40955 );
xor ( n40957 , n40956 , n40901 );
xor ( n40958 , n40957 , n36811 );
not ( n40959 , n36833 );
and ( n40960 , n40959 , n34554 );
xor ( n40961 , n36830 , n40960 );
xor ( n40962 , n40958 , n40961 );
not ( n40963 , n36841 );
and ( n40964 , n40963 , n34564 );
xor ( n40965 , n36838 , n40964 );
xor ( n40966 , n40962 , n40965 );
xor ( n40967 , n40558 , n40966 );
xor ( n40968 , n40967 , n37460 );
and ( n40969 , n40953 , n40968 );
xor ( n40970 , n40950 , n40969 );
not ( n12566 , n29614 );
and ( n12567 , n12566 , RI17393370_2038);
and ( n12568 , n40970 , n29614 );
or ( n40971 , n12567 , n12568 );
not ( n12569 , RI1754c610_2);
and ( n12570 , n12569 , n40971 );
and ( n12571 , C0 , RI1754c610_2);
or ( n40972 , n12570 , n12571 );
buf ( n40973 , n40972 );
not ( n40974 , n38969 );
and ( n40975 , n40974 , n33303 );
xor ( n40976 , n39047 , n40975 );
xor ( n40977 , n40976 , n39065 );
xor ( n40978 , n40977 , n37331 );
xor ( n40979 , n39595 , n31621 );
xor ( n40980 , n40979 , n35272 );
not ( n40981 , n40980 );
and ( n40982 , n40981 , n40343 );
xor ( n40983 , n40978 , n40982 );
not ( n12572 , n29614 );
and ( n12573 , n12572 , RI174ccee8_773);
and ( n12574 , n40983 , n29614 );
or ( n40984 , n12573 , n12574 );
not ( n12575 , RI1754c610_2);
and ( n12576 , n12575 , n40984 );
and ( n12577 , C0 , RI1754c610_2);
or ( n40985 , n12576 , n12577 );
buf ( n40986 , n40985 );
not ( n12578 , n27683 );
and ( n12579 , n12578 , RI19a90cc8_2677);
and ( n12580 , RI19a9ad18_2606 , n27683 );
or ( n40987 , n12579 , n12580 );
not ( n12581 , RI1754c610_2);
and ( n12582 , n12581 , n40987 );
and ( n12583 , C0 , RI1754c610_2);
or ( n40988 , n12582 , n12583 );
buf ( n40989 , n40988 );
not ( n40990 , n35323 );
and ( n40991 , n40990 , n35325 );
xor ( n40992 , n36970 , n40991 );
xor ( n40993 , n36961 , n40992 );
not ( n40994 , n35333 );
and ( n40995 , n40994 , n35335 );
xor ( n40996 , n36978 , n40995 );
xor ( n40997 , n40993 , n40996 );
not ( n40998 , n35343 );
and ( n40999 , n40998 , n35345 );
xor ( n41000 , n36986 , n40999 );
xor ( n41001 , n40997 , n41000 );
not ( n41002 , n35353 );
and ( n41003 , n41002 , n35355 );
xor ( n41004 , n36994 , n41003 );
xor ( n41005 , n41001 , n41004 );
xor ( n41006 , n35321 , n41005 );
xor ( n41007 , n41006 , n40585 );
not ( n41008 , n41007 );
xor ( n41009 , n33904 , n37291 );
xor ( n41010 , n41009 , n37311 );
and ( n41011 , n41008 , n41010 );
xor ( n41012 , n33506 , n41011 );
not ( n12584 , n29614 );
and ( n12585 , n12584 , RI1740d098_1444);
and ( n12586 , n41012 , n29614 );
or ( n41013 , n12585 , n12586 );
not ( n12587 , RI1754c610_2);
and ( n12588 , n12587 , n41013 );
and ( n12589 , C0 , RI1754c610_2);
or ( n41014 , n12588 , n12589 );
buf ( n41015 , n41014 );
xor ( n41016 , n34601 , n35544 );
xor ( n41017 , n41016 , n35594 );
xor ( n41018 , n41000 , n36998 );
xor ( n41019 , n41018 , n37048 );
not ( n41020 , n41019 );
xor ( n41021 , n39090 , n36377 );
xor ( n41022 , n41021 , n39131 );
and ( n41023 , n41020 , n41022 );
xor ( n41024 , n41017 , n41023 );
not ( n12590 , n29614 );
and ( n12591 , n12590 , RI1747f2d8_1116);
and ( n12592 , n41024 , n29614 );
or ( n41025 , n12591 , n12592 );
not ( n12593 , RI1754c610_2);
and ( n12594 , n12593 , n41025 );
and ( n12595 , C0 , RI1754c610_2);
or ( n41026 , n12594 , n12595 );
buf ( n41027 , n41026 );
xor ( n41028 , n32785 , n37186 );
xor ( n41029 , n41028 , n37203 );
xor ( n41030 , n34227 , n37526 );
not ( n41031 , n34357 );
xor ( n41032 , n29949 , n32009 );
xor ( n41033 , n41032 , n30164 );
and ( n41034 , n41031 , n41033 );
xor ( n41035 , n34354 , n41034 );
not ( n41036 , n34366 );
xor ( n41037 , n29541 , n30594 );
xor ( n41038 , n41037 , n29224 );
and ( n41039 , n41036 , n41038 );
xor ( n41040 , n34363 , n41039 );
xor ( n41041 , n41035 , n41040 );
not ( n41042 , n34376 );
xor ( n41043 , n29886 , n29740 );
xor ( n41044 , n41043 , n29752 );
and ( n41045 , n41042 , n41044 );
xor ( n41046 , n34373 , n41045 );
xor ( n41047 , n41041 , n41046 );
xor ( n41048 , n41047 , n34350 );
xor ( n41049 , n41048 , n40619 );
xor ( n41050 , n41030 , n41049 );
not ( n41051 , n41050 );
xor ( n41052 , n39550 , n38401 );
not ( n41053 , n35373 );
and ( n41054 , n41053 , n35375 );
xor ( n41055 , n36308 , n41054 );
not ( n41056 , n35382 );
and ( n41057 , n41056 , n35384 );
xor ( n41058 , n36315 , n41057 );
xor ( n41059 , n41055 , n41058 );
xor ( n41060 , n41059 , n36304 );
not ( n41061 , n35402 );
and ( n41062 , n41061 , n35404 );
xor ( n41063 , n36329 , n41062 );
xor ( n41064 , n41060 , n41063 );
not ( n41065 , n35412 );
and ( n41066 , n41065 , n35364 );
xor ( n41067 , n36335 , n41066 );
xor ( n41068 , n41064 , n41067 );
xor ( n41069 , n41052 , n41068 );
and ( n41070 , n41051 , n41069 );
xor ( n41071 , n41029 , n41070 );
not ( n12596 , n29614 );
and ( n12597 , n12596 , RI174a37a0_939);
and ( n12598 , n41071 , n29614 );
or ( n41072 , n12597 , n12598 );
not ( n12599 , RI1754c610_2);
and ( n12600 , n12599 , n41072 );
and ( n12601 , C0 , RI1754c610_2);
or ( n41073 , n12600 , n12601 );
buf ( n41074 , n41073 );
xor ( n41075 , n38209 , n37696 );
xor ( n41076 , n41075 , n39450 );
xor ( n41077 , n40691 , n36654 );
xor ( n41078 , n41077 , n40808 );
not ( n41079 , n41078 );
xor ( n41080 , n40095 , n39740 );
not ( n41081 , n38126 );
xor ( n41082 , n29433 , n27712 );
xor ( n41083 , n41082 , n30030 );
and ( n41084 , n41081 , n41083 );
xor ( n41085 , n30960 , n41084 );
not ( n41086 , n38131 );
xor ( n41087 , n28514 , n29724 );
xor ( n41088 , n41087 , n31291 );
and ( n41089 , n41086 , n41088 );
xor ( n41090 , n30987 , n41089 );
xor ( n41091 , n41085 , n41090 );
xor ( n41092 , n41091 , n39113 );
xor ( n41093 , n41092 , n38123 );
not ( n41094 , n38147 );
xor ( n41095 , n29156 , n29037 );
xor ( n41096 , n41095 , n31180 );
and ( n41097 , n41094 , n41096 );
xor ( n41098 , n31050 , n41097 );
xor ( n41099 , n41093 , n41098 );
xor ( n41100 , n41080 , n41099 );
and ( n41101 , n41079 , n41100 );
xor ( n41102 , n41076 , n41101 );
not ( n12602 , n29614 );
and ( n12603 , n12602 , RI173f3670_1569);
and ( n12604 , n41102 , n29614 );
or ( n41103 , n12603 , n12604 );
not ( n12605 , RI1754c610_2);
and ( n12606 , n12605 , n41103 );
and ( n12607 , C0 , RI1754c610_2);
or ( n41104 , n12606 , n12607 );
buf ( n41105 , n41104 );
xor ( n41106 , n36701 , n39655 );
not ( n41107 , n38847 );
and ( n41108 , n41107 , n38304 );
xor ( n41109 , n38300 , n41108 );
not ( n41110 , n38852 );
and ( n41111 , n41110 , n38309 );
xor ( n41112 , n38615 , n41111 );
xor ( n41113 , n41109 , n41112 );
not ( n41114 , n38858 );
and ( n41115 , n41114 , n38319 );
xor ( n41116 , n38621 , n41115 );
xor ( n41117 , n41113 , n41116 );
not ( n41118 , n38864 );
and ( n41119 , n41118 , n38329 );
xor ( n41120 , n38627 , n41119 );
xor ( n41121 , n41117 , n41120 );
not ( n41122 , n38610 );
and ( n41123 , n41122 , n38339 );
xor ( n41124 , n38607 , n41123 );
xor ( n41125 , n41121 , n41124 );
xor ( n41126 , n41106 , n41125 );
xor ( n41127 , n31670 , n30741 );
xor ( n41128 , n41127 , n40769 );
not ( n41129 , n41128 );
xor ( n41130 , n30078 , n34755 );
xor ( n41131 , n41130 , n35311 );
and ( n41132 , n41129 , n41131 );
xor ( n41133 , n41126 , n41132 );
not ( n12608 , n29614 );
and ( n12609 , n12608 , RI174a4e98_932);
and ( n12610 , n41133 , n29614 );
or ( n41134 , n12609 , n12610 );
not ( n12611 , RI1754c610_2);
and ( n12612 , n12611 , n41134 );
and ( n12613 , C0 , RI1754c610_2);
or ( n41135 , n12612 , n12613 );
buf ( n41136 , n41135 );
xor ( n41137 , n40624 , n34052 );
xor ( n41138 , n41137 , n36291 );
not ( n41139 , n33862 );
and ( n41140 , n41139 , n33864 );
xor ( n41141 , n34075 , n41140 );
xor ( n41142 , n41138 , n41141 );
not ( n41143 , n33872 );
and ( n41144 , n41143 , n33874 );
xor ( n41145 , n34083 , n41144 );
xor ( n41146 , n41142 , n41145 );
xor ( n41147 , n33853 , n41146 );
xor ( n41148 , n41147 , n37291 );
xor ( n41149 , n39327 , n35416 );
xor ( n41150 , n41149 , n29843 );
not ( n41151 , n41150 );
xor ( n41152 , n39126 , n28111 );
xor ( n41153 , n41152 , n28468 );
and ( n41154 , n41151 , n41153 );
xor ( n41155 , n41148 , n41154 );
not ( n12614 , n29614 );
and ( n12615 , n12614 , RI17454858_1324);
and ( n12616 , n41155 , n29614 );
or ( n41156 , n12615 , n12616 );
not ( n12617 , RI1754c610_2);
and ( n12618 , n12617 , n41156 );
and ( n12619 , C0 , RI1754c610_2);
or ( n41157 , n12618 , n12619 );
buf ( n41158 , n41157 );
xor ( n41159 , n40318 , n37869 );
xor ( n41160 , n41159 , n38948 );
not ( n41161 , n40928 );
and ( n41162 , n41161 , n40489 );
xor ( n41163 , n38751 , n41162 );
xor ( n41164 , n41163 , n40949 );
xor ( n41165 , n41164 , n34572 );
not ( n41166 , n41165 );
not ( n41167 , n36041 );
and ( n41168 , n41167 , n33419 );
xor ( n41169 , n34459 , n41168 );
xor ( n41170 , n41169 , n36062 );
xor ( n41171 , n41170 , n36102 );
and ( n41172 , n41166 , n41171 );
xor ( n41173 , n41160 , n41172 );
not ( n12620 , n29614 );
and ( n12621 , n12620 , RI17403318_1492);
and ( n12622 , n41173 , n29614 );
or ( n41174 , n12621 , n12622 );
not ( n12623 , RI1754c610_2);
and ( n12624 , n12623 , n41174 );
and ( n12625 , C0 , RI1754c610_2);
or ( n41175 , n12624 , n12625 );
buf ( n41176 , n41175 );
not ( n12626 , n27683 );
and ( n12627 , n12626 , RI19aaca18_2478);
and ( n12628 , RI19ab63d8_2407 , n27683 );
or ( n41177 , n12627 , n12628 );
not ( n12629 , RI1754c610_2);
and ( n12630 , n12629 , n41177 );
and ( n12631 , C0 , RI1754c610_2);
or ( n41178 , n12630 , n12631 );
buf ( n41179 , n41178 );
not ( n41180 , n34580 );
and ( n41181 , n41180 , n36847 );
xor ( n41182 , n34577 , n41181 );
not ( n41183 , n34589 );
and ( n41184 , n41183 , n36852 );
xor ( n41185 , n34586 , n41184 );
xor ( n41186 , n41182 , n41185 );
not ( n41187 , n34599 );
and ( n41188 , n41187 , n36858 );
xor ( n41189 , n34596 , n41188 );
xor ( n41190 , n41186 , n41189 );
not ( n41191 , n34609 );
and ( n41192 , n41191 , n36864 );
xor ( n41193 , n34606 , n41192 );
xor ( n41194 , n41190 , n41193 );
not ( n41195 , n34619 );
and ( n41196 , n41195 , n36870 );
xor ( n41197 , n34616 , n41196 );
xor ( n41198 , n41194 , n41197 );
xor ( n41199 , n36873 , n41198 );
not ( n41200 , n39376 );
and ( n41201 , n41200 , n37468 );
xor ( n41202 , n35561 , n41201 );
xor ( n41203 , n39370 , n41202 );
not ( n41204 , n39382 );
and ( n41205 , n41204 , n37474 );
xor ( n41206 , n35571 , n41205 );
xor ( n41207 , n41203 , n41206 );
not ( n41208 , n39388 );
and ( n41209 , n41208 , n37480 );
xor ( n41210 , n35581 , n41209 );
xor ( n41211 , n41207 , n41210 );
not ( n41212 , n39394 );
and ( n41213 , n41212 , n37486 );
xor ( n41214 , n35591 , n41213 );
xor ( n41215 , n41211 , n41214 );
xor ( n41216 , n41199 , n41215 );
not ( n41217 , n38962 );
and ( n41218 , n41217 , n39006 );
xor ( n41219 , n41216 , n41218 );
not ( n12632 , n29614 );
and ( n12633 , n12632 , RI174a2a80_943);
and ( n12634 , n41219 , n29614 );
or ( n41220 , n12633 , n12634 );
not ( n12635 , RI1754c610_2);
and ( n12636 , n12635 , n41220 );
and ( n12637 , C0 , RI1754c610_2);
or ( n41221 , n12636 , n12637 );
buf ( n41222 , n41221 );
not ( n12638 , n27683 );
and ( n12639 , n12638 , RI19a9fae8_2571);
and ( n12640 , RI19aa9868_2499 , n27683 );
or ( n41223 , n12639 , n12640 );
not ( n12641 , RI1754c610_2);
and ( n12642 , n12641 , n41223 );
and ( n12643 , C0 , RI1754c610_2);
or ( n41224 , n12642 , n12643 );
buf ( n41225 , n41224 );
xor ( n41226 , n35749 , n39563 );
xor ( n41227 , n41226 , n35416 );
xor ( n41228 , n39654 , n35216 );
not ( n41229 , n38300 );
and ( n41230 , n41229 , n38847 );
xor ( n41231 , n38297 , n41230 );
xor ( n41232 , n41231 , n40598 );
not ( n41233 , n38621 );
and ( n41234 , n41233 , n38858 );
xor ( n41235 , n38324 , n41234 );
xor ( n41236 , n41232 , n41235 );
not ( n41237 , n38627 );
and ( n41238 , n41237 , n38864 );
xor ( n41239 , n38334 , n41238 );
xor ( n41240 , n41236 , n41239 );
xor ( n41241 , n41240 , n38612 );
xor ( n41242 , n41228 , n41241 );
not ( n41243 , n41242 );
xor ( n41244 , n34928 , n36802 );
xor ( n41245 , n41244 , n33125 );
and ( n41246 , n41243 , n41245 );
xor ( n41247 , n41227 , n41246 );
not ( n12644 , n29614 );
and ( n12645 , n12644 , RI173f0bc8_1582);
and ( n12646 , n41247 , n29614 );
or ( n41248 , n12645 , n12646 );
not ( n12647 , RI1754c610_2);
and ( n12648 , n12647 , n41248 );
and ( n12649 , C0 , RI1754c610_2);
or ( n41249 , n12648 , n12649 );
buf ( n41250 , n41249 );
xor ( n41251 , n39462 , n36611 );
xor ( n41252 , n41251 , n33567 );
xor ( n41253 , n36101 , n37371 );
xor ( n41254 , n41253 , n36682 );
not ( n41255 , n41254 );
xor ( n41256 , n34656 , n32863 );
xor ( n41257 , n41256 , n34644 );
and ( n41258 , n41255 , n41257 );
xor ( n41259 , n41252 , n41258 );
not ( n12650 , n29614 );
and ( n12651 , n12650 , RI173ab9e8_1919);
and ( n12652 , n41259 , n29614 );
or ( n41260 , n12651 , n12652 );
not ( n12653 , RI1754c610_2);
and ( n12654 , n12653 , n41260 );
and ( n12655 , C0 , RI1754c610_2);
or ( n41261 , n12654 , n12655 );
buf ( n41262 , n41261 );
not ( n41263 , n31236 );
and ( n41264 , n41263 , n31249 );
xor ( n41265 , n33630 , n41264 );
xor ( n41266 , n41265 , n33648 );
xor ( n41267 , n41266 , n33697 );
xor ( n41268 , n37909 , n32048 );
xor ( n41269 , n41268 , n32108 );
not ( n41270 , n41269 );
xor ( n41271 , n41120 , n41241 );
not ( n41272 , n31409 );
and ( n41273 , n41272 , n31411 );
xor ( n41274 , n34270 , n41273 );
xor ( n41275 , n41274 , n40873 );
not ( n41276 , n31438 );
and ( n41277 , n41276 , n31389 );
xor ( n41278 , n34262 , n41277 );
xor ( n41279 , n41275 , n41278 );
not ( n41280 , n31444 );
and ( n41281 , n41280 , n31463 );
xor ( n41282 , n34289 , n41281 );
xor ( n41283 , n41279 , n41282 );
not ( n41284 , n31498 );
and ( n41285 , n41284 , n31500 );
xor ( n41286 , n34297 , n41285 );
xor ( n41287 , n41283 , n41286 );
xor ( n41288 , n41271 , n41287 );
and ( n41289 , n41270 , n41288 );
xor ( n41290 , n41267 , n41289 );
not ( n12656 , n29614 );
and ( n12657 , n12656 , RI1744efc0_1351);
and ( n12658 , n41290 , n29614 );
or ( n41291 , n12657 , n12658 );
not ( n12659 , RI1754c610_2);
and ( n12660 , n12659 , n41291 );
and ( n12661 , C0 , RI1754c610_2);
or ( n41292 , n12660 , n12661 );
buf ( n41293 , n41292 );
buf ( n41294 , RI17470350_1189);
xor ( n41295 , n41067 , n36339 );
xor ( n41296 , n41295 , n36377 );
xor ( n41297 , n35554 , n37490 );
not ( n41298 , n32332 );
and ( n41299 , n41298 , n32313 );
xor ( n41300 , n33794 , n41299 );
not ( n41301 , n32337 );
and ( n41302 , n41301 , n32339 );
xor ( n41303 , n33788 , n41302 );
xor ( n41304 , n41300 , n41303 );
not ( n41305 , n32347 );
and ( n41306 , n41305 , n32349 );
xor ( n41307 , n33805 , n41306 );
xor ( n41308 , n41304 , n41307 );
not ( n41309 , n32368 );
and ( n41310 , n41309 , n32370 );
xor ( n41311 , n33813 , n41310 );
xor ( n41312 , n41308 , n41311 );
not ( n41313 , n32388 );
and ( n41314 , n41313 , n32390 );
xor ( n41315 , n33821 , n41314 );
xor ( n41316 , n41312 , n41315 );
xor ( n41317 , n41297 , n41316 );
not ( n41318 , n41317 );
xor ( n41319 , n40098 , n39740 );
xor ( n41320 , n41319 , n41099 );
and ( n41321 , n41318 , n41320 );
xor ( n41322 , n41296 , n41321 );
not ( n12662 , n29614 );
and ( n12663 , n12662 , RI17534d30_602);
and ( n12664 , n41322 , n29614 );
or ( n41323 , n12663 , n12664 );
not ( n12665 , RI1754c610_2);
and ( n12666 , n12665 , n41323 );
and ( n12667 , C0 , RI1754c610_2);
or ( n41324 , n12666 , n12667 );
buf ( n41325 , n41324 );
xor ( n41326 , n38307 , n38872 );
xor ( n41327 , n41326 , n38886 );
not ( n41328 , n41327 );
xor ( n41329 , n35629 , n34669 );
xor ( n41330 , n41329 , n31831 );
and ( n41331 , n41328 , n41330 );
xor ( n41332 , n40052 , n41331 );
not ( n12668 , n29614 );
and ( n12669 , n12668 , RI173fb320_1531);
and ( n12670 , n41332 , n29614 );
or ( n41333 , n12669 , n12670 );
not ( n12671 , RI1754c610_2);
and ( n12672 , n12671 , n41333 );
and ( n12673 , C0 , RI1754c610_2);
or ( n41334 , n12672 , n12673 );
buf ( n41335 , n41334 );
xor ( n41336 , n36135 , n39151 );
xor ( n41337 , n41336 , n38267 );
xor ( n41338 , n36203 , n32923 );
xor ( n41339 , n41338 , n32973 );
not ( n41340 , n41339 );
not ( n41341 , n37786 );
and ( n41342 , n41341 , n37748 );
xor ( n41343 , n40433 , n41342 );
xor ( n41344 , n41343 , n40808 );
xor ( n41345 , n41344 , n40828 );
and ( n41346 , n41340 , n41345 );
xor ( n41347 , n41337 , n41346 );
not ( n12674 , n29614 );
and ( n12675 , n12674 , RI17451a68_1338);
and ( n12676 , n41347 , n29614 );
or ( n41348 , n12675 , n12676 );
not ( n12677 , RI1754c610_2);
and ( n12678 , n12677 , n41348 );
and ( n12679 , C0 , RI1754c610_2);
or ( n41349 , n12678 , n12679 );
buf ( n41350 , n41349 );
and ( n41351 , RI19a822e0_2779 , n27689 );
not ( n12680 , RI1754c610_2);
and ( n12681 , n12680 , n41351 );
and ( n12682 , C0 , RI1754c610_2);
or ( n41352 , n12681 , n12682 );
buf ( n41353 , n41352 );
not ( n12683 , n27683 );
and ( n12684 , n12683 , RI19abd890_2354);
and ( n12685 , RI19ac63c8_2283 , n27683 );
or ( n41354 , n12684 , n12685 );
not ( n12686 , RI1754c610_2);
and ( n12687 , n12686 , n41354 );
and ( n12688 , C0 , RI1754c610_2);
or ( n41355 , n12687 , n12688 );
buf ( n41356 , n41355 );
buf ( n41357 , RI1746fcc0_1191);
xor ( n41358 , n36035 , n41169 );
not ( n41359 , n36047 );
and ( n41360 , n41359 , n33429 );
xor ( n41361 , n34465 , n41360 );
xor ( n41362 , n41358 , n41361 );
not ( n41363 , n36053 );
and ( n41364 , n41363 , n33439 );
xor ( n41365 , n34471 , n41364 );
xor ( n41366 , n41362 , n41365 );
not ( n41367 , n36059 );
and ( n41368 , n41367 , n33449 );
xor ( n41369 , n33406 , n41368 );
xor ( n41370 , n41366 , n41369 );
xor ( n41371 , n36239 , n41370 );
xor ( n41372 , n41371 , n37898 );
xor ( n41373 , n40737 , n31925 );
xor ( n41374 , n41373 , n34475 );
not ( n41375 , n41374 );
not ( n41376 , n33527 );
and ( n41377 , n41376 , n34764 );
xor ( n41378 , n33524 , n41377 );
not ( n41379 , n33536 );
and ( n41380 , n41379 , n34771 );
xor ( n41381 , n33533 , n41380 );
xor ( n41382 , n41378 , n41381 );
not ( n41383 , n33548 );
and ( n41384 , n41383 , n34777 );
xor ( n41385 , n33545 , n41384 );
xor ( n41386 , n41382 , n41385 );
xor ( n41387 , n41386 , n33520 );
not ( n41388 , n33564 );
and ( n41389 , n41388 , n34791 );
xor ( n41390 , n33561 , n41389 );
xor ( n41391 , n41387 , n41390 );
xor ( n41392 , n37250 , n41391 );
xor ( n41393 , n41392 , n39686 );
and ( n41394 , n41375 , n41393 );
xor ( n41395 , n41372 , n41394 );
not ( n12689 , n29614 );
and ( n12690 , n12689 , RI17471d90_1181);
and ( n12691 , n41395 , n29614 );
or ( n41396 , n12690 , n12691 );
not ( n12692 , RI1754c610_2);
and ( n12693 , n12692 , n41396 );
and ( n12694 , C0 , RI1754c610_2);
or ( n41397 , n12693 , n12694 );
buf ( n41398 , n41397 );
xor ( n41399 , n37889 , n36102 );
xor ( n41400 , n41399 , n32048 );
xor ( n41401 , n33869 , n41146 );
xor ( n41402 , n41401 , n37291 );
not ( n41403 , n41402 );
xor ( n41404 , n37047 , n40662 );
xor ( n41405 , n41404 , n39208 );
and ( n41406 , n41403 , n41405 );
xor ( n41407 , n41400 , n41406 );
not ( n12695 , n29614 );
and ( n12696 , n12695 , RI17481060_1107);
and ( n12697 , n41407 , n29614 );
or ( n41408 , n12696 , n12697 );
not ( n12698 , RI1754c610_2);
and ( n12699 , n12698 , n41408 );
and ( n12700 , C0 , RI1754c610_2);
or ( n41409 , n12699 , n12700 );
buf ( n41410 , n41409 );
xor ( n41411 , n40481 , n38933 );
not ( n41412 , n40489 );
and ( n41413 , n41412 , n38746 );
xor ( n41414 , n40928 , n41413 );
not ( n41415 , n40494 );
and ( n41416 , n41415 , n38755 );
xor ( n41417 , n40933 , n41416 );
xor ( n41418 , n41414 , n41417 );
not ( n41419 , n40500 );
and ( n41420 , n41419 , n38765 );
xor ( n41421 , n40939 , n41420 );
xor ( n41422 , n41418 , n41421 );
not ( n41423 , n40506 );
and ( n41424 , n41423 , n38775 );
xor ( n41425 , n40945 , n41424 );
xor ( n41426 , n41422 , n41425 );
not ( n41427 , n40512 );
and ( n41428 , n41427 , n38785 );
xor ( n41429 , n40696 , n41428 );
xor ( n41430 , n41426 , n41429 );
xor ( n41431 , n41411 , n41430 );
xor ( n41432 , n41369 , n36062 );
xor ( n41433 , n41432 , n36102 );
not ( n41434 , n41433 );
xor ( n41435 , n41035 , n34395 );
xor ( n41436 , n41435 , n34445 );
and ( n41437 , n41434 , n41436 );
xor ( n41438 , n41431 , n41437 );
not ( n12701 , n29614 );
and ( n12702 , n12701 , RI173afb88_1899);
and ( n12703 , n41438 , n29614 );
or ( n41439 , n12702 , n12703 );
not ( n12704 , RI1754c610_2);
and ( n12705 , n12704 , n41439 );
and ( n12706 , C0 , RI1754c610_2);
or ( n41440 , n12705 , n12706 );
buf ( n41441 , n41440 );
xor ( n41442 , n34571 , n40563 );
xor ( n41443 , n41442 , n35544 );
xor ( n41444 , n39758 , n33125 );
xor ( n41445 , n41444 , n33175 );
not ( n41446 , n41445 );
not ( n41447 , n34097 );
and ( n41448 , n41447 , n34099 );
xor ( n41449 , n33902 , n41448 );
xor ( n41450 , n41449 , n36431 );
xor ( n41451 , n41450 , n34221 );
and ( n41452 , n41446 , n41451 );
xor ( n41453 , n41443 , n41452 );
not ( n12707 , n29614 );
and ( n12708 , n12707 , RI173bca40_1836);
and ( n12709 , n41453 , n29614 );
or ( n41454 , n12708 , n12709 );
not ( n12710 , RI1754c610_2);
and ( n12711 , n12710 , n41454 );
and ( n12712 , C0 , RI1754c610_2);
or ( n41455 , n12711 , n12712 );
buf ( n41456 , n41455 );
buf ( n41457 , RI174cd410_772);
not ( n12713 , n27683 );
and ( n12714 , n12713 , RI19aa5218_2529);
and ( n12715 , RI19aaf628_2458 , n27683 );
or ( n41458 , n12714 , n12715 );
not ( n12716 , RI1754c610_2);
and ( n12717 , n12716 , n41458 );
and ( n12718 , C0 , RI1754c610_2);
or ( n41459 , n12717 , n12718 );
buf ( n41460 , n41459 );
xor ( n41461 , n41112 , n41241 );
xor ( n41462 , n41461 , n41287 );
not ( n41463 , n34807 );
and ( n41464 , n41463 , n34809 );
xor ( n41465 , n33584 , n41464 );
xor ( n41466 , n39670 , n41465 );
not ( n41467 , n34815 );
and ( n41468 , n41467 , n34817 );
xor ( n41469 , n33594 , n41468 );
xor ( n41470 , n41466 , n41469 );
not ( n41471 , n34823 );
and ( n41472 , n41471 , n34825 );
xor ( n41473 , n33604 , n41472 );
xor ( n41474 , n41470 , n41473 );
not ( n41475 , n34831 );
and ( n41476 , n41475 , n34833 );
xor ( n41477 , n33614 , n41476 );
xor ( n41478 , n41474 , n41477 );
xor ( n41479 , n34820 , n41478 );
xor ( n41480 , n41479 , n41146 );
not ( n41481 , n41480 );
not ( n41482 , n34348 );
and ( n41483 , n41482 , n39979 );
xor ( n41484 , n34345 , n41483 );
xor ( n41485 , n41484 , n41049 );
not ( n41486 , n34403 );
and ( n41487 , n41486 , n37954 );
xor ( n41488 , n34400 , n41487 );
not ( n41489 , n34412 );
and ( n41490 , n41489 , n37961 );
xor ( n41491 , n34409 , n41490 );
xor ( n41492 , n41488 , n41491 );
not ( n41493 , n34422 );
and ( n41494 , n41493 , n37969 );
xor ( n41495 , n34419 , n41494 );
xor ( n41496 , n41492 , n41495 );
not ( n41497 , n34432 );
and ( n41498 , n41497 , n37947 );
xor ( n41499 , n34429 , n41498 );
xor ( n41500 , n41496 , n41499 );
not ( n41501 , n34442 );
and ( n41502 , n41501 , n37981 );
xor ( n41503 , n34439 , n41502 );
xor ( n41504 , n41500 , n41503 );
xor ( n41505 , n41485 , n41504 );
and ( n41506 , n41481 , n41505 );
xor ( n41507 , n41462 , n41506 );
not ( n12719 , n29614 );
and ( n12720 , n12719 , RI173d8550_1701);
and ( n12721 , n41507 , n29614 );
or ( n41508 , n12720 , n12721 );
not ( n12722 , RI1754c610_2);
and ( n12723 , n12722 , n41508 );
and ( n12724 , C0 , RI1754c610_2);
or ( n41509 , n12723 , n12724 );
buf ( n41510 , n41509 );
buf ( n41511 , RI1748d540_1047);
xor ( n41512 , n35880 , n36463 );
xor ( n41513 , n41512 , n32220 );
not ( n41514 , n33794 );
and ( n41515 , n41514 , n32332 );
xor ( n41516 , n32328 , n41515 );
xor ( n41517 , n41516 , n33791 );
xor ( n41518 , n41517 , n39289 );
not ( n41519 , n33813 );
and ( n41520 , n41519 , n32368 );
xor ( n41521 , n33810 , n41520 );
xor ( n41522 , n41518 , n41521 );
not ( n41523 , n33821 );
and ( n41524 , n41523 , n32388 );
xor ( n41525 , n33818 , n41524 );
xor ( n41526 , n41522 , n41525 );
xor ( n41527 , n41307 , n41526 );
not ( n41528 , n32748 );
and ( n41529 , n41528 , n32406 );
xor ( n41530 , n32745 , n41529 );
not ( n41531 , n32755 );
and ( n41532 , n41531 , n32415 );
xor ( n41533 , n32752 , n41532 );
xor ( n41534 , n41530 , n41533 );
xor ( n41535 , n41534 , n32726 );
not ( n41536 , n32767 );
and ( n41537 , n41536 , n32446 );
xor ( n41538 , n32764 , n41537 );
xor ( n41539 , n41535 , n41538 );
not ( n41540 , n32783 );
and ( n41541 , n41540 , n32466 );
xor ( n41542 , n32780 , n41541 );
xor ( n41543 , n41539 , n41542 );
xor ( n41544 , n41527 , n41543 );
not ( n41545 , n41544 );
xor ( n41546 , n37198 , n33030 );
xor ( n41547 , n41546 , n33069 );
and ( n41548 , n41545 , n41547 );
xor ( n41549 , n41513 , n41548 );
not ( n12725 , n29614 );
and ( n12726 , n12725 , RI1744d580_1359);
and ( n12727 , n41549 , n29614 );
or ( n41550 , n12726 , n12727 );
not ( n12728 , RI1754c610_2);
and ( n12729 , n12728 , n41550 );
and ( n12730 , C0 , RI1754c610_2);
or ( n41551 , n12729 , n12730 );
buf ( n41552 , n41551 );
not ( n12731 , n27683 );
and ( n12732 , n12731 , RI19abaa28_2376);
and ( n12733 , RI19ac3290_2305 , n27683 );
or ( n41553 , n12732 , n12733 );
not ( n12734 , RI1754c610_2);
and ( n12735 , n12734 , n41553 );
and ( n12736 , C0 , RI1754c610_2);
or ( n41554 , n12735 , n12736 );
buf ( n41555 , n41554 );
buf ( n41556 , RI174709e0_1187);
buf ( n41557 , RI19ad0700_2208);
xor ( n41558 , n39441 , n38495 );
xor ( n41559 , n41558 , n36611 );
xor ( n41560 , n32599 , n39182 );
xor ( n41561 , n41560 , n38991 );
not ( n41562 , n41561 );
xor ( n41563 , n36567 , n37438 );
xor ( n41564 , n41563 , n30247 );
and ( n41565 , n41562 , n41564 );
xor ( n41566 , n41559 , n41565 );
not ( n12737 , n29614 );
and ( n12738 , n12737 , RI17399fb8_2005);
and ( n12739 , n41566 , n29614 );
or ( n41567 , n12738 , n12739 );
not ( n12740 , RI1754c610_2);
and ( n12741 , n12740 , n41567 );
and ( n12742 , C0 , RI1754c610_2);
or ( n41568 , n12741 , n12742 );
buf ( n41569 , n41568 );
xor ( n41570 , n36139 , n39151 );
xor ( n41571 , n41570 , n38267 );
xor ( n41572 , n35433 , n32663 );
xor ( n41573 , n41572 , n32715 );
not ( n41574 , n41573 );
not ( n41575 , n38964 );
and ( n41576 , n41575 , n33294 );
xor ( n41577 , n39042 , n41576 );
xor ( n41578 , n41577 , n40976 );
not ( n41579 , n38975 );
and ( n41580 , n41579 , n33313 );
xor ( n41581 , n37337 , n41580 );
xor ( n41582 , n41578 , n41581 );
not ( n41583 , n38981 );
and ( n41584 , n41583 , n33323 );
xor ( n41585 , n33290 , n41584 );
xor ( n41586 , n41582 , n41585 );
not ( n41587 , n38987 );
and ( n41588 , n41587 , n33329 );
xor ( n41589 , n39061 , n41588 );
xor ( n41590 , n41586 , n41589 );
xor ( n41591 , n38990 , n41590 );
xor ( n41592 , n41591 , n35804 );
and ( n41593 , n41574 , n41592 );
xor ( n41594 , n41571 , n41593 );
not ( n12743 , n29614 );
and ( n12744 , n12743 , RI173a67e0_1944);
and ( n12745 , n41594 , n29614 );
or ( n41595 , n12744 , n12745 );
not ( n12746 , RI1754c610_2);
and ( n12747 , n12746 , n41595 );
and ( n12748 , C0 , RI1754c610_2);
or ( n41596 , n12747 , n12748 );
buf ( n41597 , n41596 );
not ( n12749 , n27683 );
and ( n12750 , n12749 , RI19ac81c8_2269);
and ( n12751 , RI19a82f88_2773 , n27683 );
or ( n41598 , n12750 , n12751 );
not ( n12752 , RI1754c610_2);
and ( n12753 , n12752 , n41598 );
and ( n12754 , C0 , RI1754c610_2);
or ( n41599 , n12753 , n12754 );
buf ( n41600 , n41599 );
xor ( n41601 , n39588 , n31621 );
xor ( n41602 , n41601 , n35272 );
xor ( n41603 , n30831 , n38115 );
not ( n41604 , n30936 );
and ( n41605 , n41604 , n30957 );
xor ( n41606 , n41083 , n41605 );
not ( n41607 , n30974 );
and ( n41608 , n41607 , n30977 );
xor ( n41609 , n41088 , n41608 );
xor ( n41610 , n41606 , n41609 );
not ( n41611 , n31003 );
and ( n41612 , n41611 , n31005 );
xor ( n41613 , n39111 , n41612 );
xor ( n41614 , n41610 , n41613 );
not ( n41615 , n31013 );
and ( n41616 , n41615 , n31026 );
xor ( n41617 , n38121 , n41616 );
xor ( n41618 , n41614 , n41617 );
not ( n41619 , n31045 );
and ( n41620 , n41619 , n31047 );
xor ( n41621 , n41096 , n41620 );
xor ( n41622 , n41618 , n41621 );
xor ( n41623 , n41603 , n41622 );
not ( n41624 , n41623 );
xor ( n41625 , n40085 , n38037 );
xor ( n41626 , n41625 , n39740 );
and ( n41627 , n41624 , n41626 );
xor ( n41628 , n41602 , n41627 );
or ( n41629 , RI17539218_590 , RI17538c00_591);
or ( n41630 , n41629 , RI175385e8_592);
or ( n41631 , n41630 , RI17537fd0_593);
or ( n41632 , n41631 , RI17536d88_596);
or ( n41633 , n41632 , RI17539e48_588);
xor ( n41634 , n41628 , n41633 );
not ( n12755 , n29614 );
and ( n12756 , n12755 , RI1746ec58_1196);
and ( n12757 , n41634 , n29614 );
or ( n41635 , n12756 , n12757 );
not ( n12758 , RI1754c610_2);
and ( n12759 , n12758 , n41635 );
and ( n12760 , C0 , RI1754c610_2);
or ( n41636 , n12759 , n12760 );
buf ( n41637 , n41636 );
xor ( n41638 , n34911 , n36772 );
xor ( n41639 , n41638 , n36802 );
xor ( n41640 , n32922 , n38553 );
not ( n41641 , n32926 );
and ( n41642 , n41641 , n32928 );
xor ( n41643 , n36620 , n41642 );
not ( n41644 , n32935 );
and ( n41645 , n41644 , n32937 );
xor ( n41646 , n36627 , n41645 );
xor ( n41647 , n41643 , n41646 );
not ( n41648 , n32945 );
and ( n41649 , n41648 , n32947 );
xor ( n41650 , n36635 , n41649 );
xor ( n41651 , n41647 , n41650 );
not ( n41652 , n32955 );
and ( n41653 , n41652 , n32957 );
xor ( n41654 , n36643 , n41653 );
xor ( n41655 , n41651 , n41654 );
not ( n41656 , n32965 );
and ( n41657 , n41656 , n32967 );
xor ( n41658 , n36651 , n41657 );
xor ( n41659 , n41655 , n41658 );
xor ( n41660 , n41640 , n41659 );
not ( n41661 , n41660 );
not ( n41662 , n38055 );
and ( n41663 , n41662 , n37990 );
xor ( n41664 , n38052 , n41663 );
xor ( n41665 , n41664 , n38085 );
xor ( n41666 , n41665 , n38115 );
and ( n41667 , n41661 , n41666 );
xor ( n41668 , n41639 , n41667 );
not ( n12761 , n29614 );
and ( n12762 , n12761 , RI173f3328_1570);
and ( n12763 , n41668 , n29614 );
or ( n41669 , n12762 , n12763 );
not ( n12764 , RI1754c610_2);
and ( n12765 , n12764 , n41669 );
and ( n12766 , C0 , RI1754c610_2);
or ( n41670 , n12765 , n12766 );
buf ( n41671 , n41670 );
not ( n41672 , n37990 );
and ( n41673 , n41672 , n37992 );
xor ( n41674 , n38055 , n41673 );
not ( n41675 , n37999 );
and ( n41676 , n41675 , n38001 );
xor ( n41677 , n38062 , n41676 );
xor ( n41678 , n41674 , n41677 );
not ( n41679 , n38009 );
and ( n41680 , n41679 , n38011 );
xor ( n41681 , n38047 , n41680 );
xor ( n41682 , n41678 , n41681 );
not ( n41683 , n38019 );
and ( n41684 , n41683 , n38021 );
xor ( n41685 , n38074 , n41684 );
xor ( n41686 , n41682 , n41685 );
not ( n41687 , n38029 );
and ( n41688 , n41687 , n38031 );
xor ( n41689 , n38082 , n41688 );
xor ( n41690 , n41686 , n41689 );
xor ( n41691 , n37997 , n41690 );
xor ( n41692 , n41691 , n39506 );
not ( n41693 , n40950 );
and ( n41694 , n41693 , n40952 );
xor ( n41695 , n41692 , n41694 );
not ( n12767 , n29614 );
and ( n12768 , n12767 , RI17343e88_2110);
and ( n12769 , n41695 , n29614 );
or ( n41696 , n12768 , n12769 );
not ( n12770 , RI1754c610_2);
and ( n12771 , n12770 , n41696 );
and ( n12772 , C0 , RI1754c610_2);
or ( n41697 , n12771 , n12772 );
buf ( n41698 , n41697 );
xor ( n41699 , n40289 , n37849 );
xor ( n41700 , n41699 , n37869 );
xor ( n41701 , n38998 , n35804 );
xor ( n41702 , n41701 , n35842 );
not ( n41703 , n41702 );
xor ( n41704 , n33859 , n41146 );
xor ( n41705 , n41704 , n37291 );
and ( n41706 , n41703 , n41705 );
xor ( n41707 , n41700 , n41706 );
not ( n12773 , n29614 );
and ( n12774 , n12773 , RI1733d240_2143);
and ( n12775 , n41707 , n29614 );
or ( n41708 , n12774 , n12775 );
not ( n12776 , RI1754c610_2);
and ( n12777 , n12776 , n41708 );
and ( n12778 , C0 , RI1754c610_2);
or ( n41709 , n12777 , n12778 );
buf ( n41710 , n41709 );
xor ( n41711 , n39646 , n35216 );
xor ( n41712 , n41711 , n41241 );
xor ( n41713 , n40106 , n39740 );
xor ( n41714 , n41713 , n41099 );
not ( n41715 , n41714 );
xor ( n41716 , n41542 , n32786 );
xor ( n41717 , n41716 , n32863 );
and ( n41718 , n41715 , n41717 );
xor ( n41719 , n41712 , n41718 );
not ( n12779 , n29614 );
and ( n12780 , n12779 , RI173a08b8_1973);
and ( n12781 , n41719 , n29614 );
or ( n41720 , n12780 , n12781 );
not ( n12782 , RI1754c610_2);
and ( n12783 , n12782 , n41720 );
and ( n12784 , C0 , RI1754c610_2);
or ( n41721 , n12783 , n12784 );
buf ( n41722 , n41721 );
xor ( n41723 , n33436 , n36252 );
xor ( n41724 , n41723 , n40360 );
not ( n41725 , n33570 );
and ( n41726 , n41725 , n33572 );
xor ( n41727 , n34802 , n41726 );
not ( n41728 , n33579 );
and ( n41729 , n41728 , n33581 );
xor ( n41730 , n34809 , n41729 );
xor ( n41731 , n41727 , n41730 );
not ( n41732 , n33589 );
and ( n41733 , n41732 , n33591 );
xor ( n41734 , n34817 , n41733 );
xor ( n41735 , n41731 , n41734 );
xor ( n41736 , n41735 , n39213 );
not ( n41737 , n33609 );
and ( n41738 , n41737 , n33611 );
xor ( n41739 , n34833 , n41738 );
xor ( n41740 , n41736 , n41739 );
xor ( n41741 , n33606 , n41740 );
xor ( n41742 , n41741 , n38371 );
not ( n41743 , n41742 );
xor ( n41744 , n35360 , n41005 );
xor ( n41745 , n41744 , n40585 );
and ( n41746 , n41743 , n41745 );
xor ( n41747 , n41724 , n41746 );
not ( n12785 , n29614 );
and ( n12786 , n12785 , RI174809d0_1109);
and ( n12787 , n41747 , n29614 );
or ( n41748 , n12786 , n12787 );
not ( n12788 , RI1754c610_2);
and ( n12789 , n12788 , n41748 );
and ( n12790 , C0 , RI1754c610_2);
or ( n41749 , n12789 , n12790 );
buf ( n41750 , n41749 );
xor ( n41751 , n40649 , n39282 );
xor ( n41752 , n41751 , n37676 );
xor ( n41753 , n39078 , n36377 );
xor ( n41754 , n41753 , n39131 );
not ( n41755 , n41754 );
xor ( n41756 , n37707 , n40463 );
not ( n41757 , n37719 );
and ( n41758 , n41757 , n35959 );
xor ( n41759 , n32153 , n41758 );
not ( n41760 , n37724 );
and ( n41761 , n41760 , n35964 );
xor ( n41762 , n32171 , n41761 );
xor ( n41763 , n41759 , n41762 );
not ( n41764 , n37730 );
and ( n41765 , n41764 , n35970 );
xor ( n41766 , n32183 , n41765 );
xor ( n41767 , n41763 , n41766 );
not ( n41768 , n37736 );
and ( n41769 , n41768 , n35976 );
xor ( n41770 , n32211 , n41769 );
xor ( n41771 , n41767 , n41770 );
xor ( n41772 , n41771 , n38172 );
xor ( n41773 , n41756 , n41772 );
and ( n41774 , n41755 , n41773 );
xor ( n41775 , n41752 , n41774 );
not ( n12791 , n29614 );
and ( n12792 , n12791 , RI174b7fc0_839);
and ( n12793 , n41775 , n29614 );
or ( n41776 , n12792 , n12793 );
not ( n12794 , RI1754c610_2);
and ( n12795 , n12794 , n41776 );
and ( n12796 , C0 , RI1754c610_2);
or ( n41777 , n12795 , n12796 );
buf ( n41778 , n41777 );
xor ( n41779 , n34541 , n40563 );
xor ( n41780 , n41779 , n35544 );
not ( n41781 , n28138 );
and ( n41782 , n41781 , n28161 );
xor ( n41783 , n35920 , n41782 );
not ( n41784 , n28213 );
and ( n41785 , n41784 , n28237 );
xor ( n41786 , n35927 , n41785 );
xor ( n41787 , n41783 , n41786 );
not ( n41788 , n28292 );
and ( n41789 , n41788 , n28314 );
xor ( n41790 , n35935 , n41789 );
xor ( n41791 , n41787 , n41790 );
not ( n41792 , n28368 );
and ( n41793 , n41792 , n28393 );
xor ( n41794 , n35943 , n41793 );
xor ( n41795 , n41791 , n41794 );
not ( n41796 , n28426 );
and ( n41797 , n41796 , n28451 );
xor ( n41798 , n35951 , n41797 );
xor ( n41799 , n41795 , n41798 );
xor ( n41800 , n28342 , n41799 );
xor ( n41801 , n41800 , n40381 );
not ( n41802 , n41801 );
not ( n41803 , n36968 );
and ( n41804 , n41803 , n36970 );
xor ( n41805 , n35328 , n41804 );
xor ( n41806 , n39246 , n41805 );
not ( n41807 , n36976 );
and ( n41808 , n41807 , n36978 );
xor ( n41809 , n35338 , n41808 );
xor ( n41810 , n41806 , n41809 );
not ( n41811 , n36984 );
and ( n41812 , n41811 , n36986 );
xor ( n41813 , n35348 , n41812 );
xor ( n41814 , n41810 , n41813 );
not ( n41815 , n36992 );
and ( n41816 , n41815 , n36994 );
xor ( n41817 , n35358 , n41816 );
xor ( n41818 , n41814 , n41817 );
xor ( n41819 , n36989 , n41818 );
xor ( n41820 , n41819 , n40662 );
and ( n41821 , n41802 , n41820 );
xor ( n41822 , n41780 , n41821 );
not ( n12797 , n29614 );
and ( n12798 , n12797 , RI173d5aa8_1714);
and ( n12799 , n41822 , n29614 );
or ( n41823 , n12798 , n12799 );
not ( n12800 , RI1754c610_2);
and ( n12801 , n12800 , n41823 );
and ( n12802 , C0 , RI1754c610_2);
or ( n41824 , n12801 , n12802 );
buf ( n41825 , n41824 );
xor ( n41826 , n32344 , n41316 );
xor ( n41827 , n41826 , n35622 );
xor ( n41828 , n30154 , n34755 );
xor ( n41829 , n41828 , n35311 );
not ( n41830 , n41829 );
and ( n41831 , n41830 , n41076 );
xor ( n41832 , n41827 , n41831 );
not ( n12803 , n29614 );
and ( n12804 , n12803 , RI173d6480_1711);
and ( n12805 , n41832 , n29614 );
or ( n41833 , n12804 , n12805 );
not ( n12806 , RI1754c610_2);
and ( n12807 , n12806 , n41833 );
and ( n12808 , C0 , RI1754c610_2);
or ( n41834 , n12807 , n12808 );
buf ( n41835 , n41834 );
xor ( n41836 , n40292 , n37849 );
xor ( n41837 , n41836 , n37869 );
xor ( n41838 , n33637 , n35069 );
not ( n41839 , n33240 );
and ( n41840 , n41839 , n33651 );
xor ( n41841 , n33237 , n41840 );
not ( n41842 , n33249 );
and ( n41843 , n41842 , n33667 );
xor ( n41844 , n33246 , n41843 );
xor ( n41845 , n41841 , n41844 );
not ( n41846 , n33259 );
and ( n41847 , n41846 , n33675 );
xor ( n41848 , n33256 , n41847 );
xor ( n41849 , n41845 , n41848 );
not ( n41850 , n33269 );
and ( n41851 , n41850 , n33683 );
xor ( n41852 , n33266 , n41851 );
xor ( n41853 , n41849 , n41852 );
xor ( n41854 , n41853 , n39219 );
xor ( n41855 , n41838 , n41854 );
not ( n41856 , n41855 );
xor ( n41857 , n37181 , n32481 );
xor ( n41858 , n41857 , n33030 );
and ( n41859 , n41856 , n41858 );
xor ( n41860 , n41837 , n41859 );
not ( n12809 , n29614 );
and ( n12810 , n12809 , RI17476278_1160);
and ( n12811 , n41860 , n29614 );
or ( n41861 , n12810 , n12811 );
not ( n12812 , RI1754c610_2);
and ( n12813 , n12812 , n41861 );
and ( n12814 , C0 , RI1754c610_2);
or ( n41862 , n12813 , n12814 );
buf ( n41863 , n41862 );
not ( n12815 , n27683 );
and ( n12816 , n12815 , RI19a83438_2771);
and ( n12817 , RI19ab54d8_2414 , n27683 );
or ( n41864 , n12816 , n12817 );
not ( n12818 , RI1754c610_2);
and ( n12819 , n12818 , n41864 );
and ( n12820 , C0 , RI1754c610_2);
or ( n41865 , n12819 , n12820 );
buf ( n41866 , n41865 );
xor ( n41867 , n39413 , n32403 );
xor ( n41868 , n41867 , n32481 );
xor ( n41869 , n38753 , n40516 );
xor ( n41870 , n41869 , n40966 );
not ( n41871 , n41870 );
xor ( n41872 , n41491 , n34445 );
not ( n41873 , n38062 );
and ( n41874 , n41873 , n37999 );
xor ( n41875 , n38059 , n41874 );
xor ( n41876 , n41664 , n41875 );
xor ( n41877 , n41876 , n38050 );
not ( n41878 , n38074 );
and ( n41879 , n41878 , n38019 );
xor ( n41880 , n38071 , n41879 );
xor ( n41881 , n41877 , n41880 );
not ( n41882 , n38082 );
and ( n41883 , n41882 , n38029 );
xor ( n41884 , n38079 , n41883 );
xor ( n41885 , n41881 , n41884 );
xor ( n41886 , n41872 , n41885 );
and ( n41887 , n41871 , n41886 );
xor ( n41888 , n41868 , n41887 );
not ( n12821 , n29614 );
and ( n12822 , n12821 , RI1745e920_1275);
and ( n12823 , n41888 , n29614 );
or ( n41889 , n12822 , n12823 );
not ( n12824 , RI1754c610_2);
and ( n12825 , n12824 , n41889 );
and ( n12826 , C0 , RI1754c610_2);
or ( n41890 , n12825 , n12826 );
buf ( n41891 , n41890 );
xor ( n41892 , n41685 , n41885 );
xor ( n41893 , n41892 , n30923 );
xor ( n41894 , n34516 , n31380 );
xor ( n41895 , n41894 , n36463 );
not ( n41896 , n41895 );
xor ( n41897 , n40877 , n34340 );
xor ( n41898 , n41897 , n38817 );
and ( n41899 , n41896 , n41898 );
xor ( n41900 , n41893 , n41899 );
not ( n12827 , n29614 );
and ( n12828 , n12827 , RI173c0208_1819);
and ( n12829 , n41900 , n29614 );
or ( n41901 , n12828 , n12829 );
not ( n12830 , RI1754c610_2);
and ( n12831 , n12830 , n41901 );
and ( n12832 , C0 , RI1754c610_2);
or ( n41902 , n12831 , n12832 );
buf ( n41903 , n41902 );
xor ( n41904 , n41063 , n36339 );
xor ( n41905 , n41904 , n36377 );
xor ( n41906 , n38633 , n38347 );
xor ( n41907 , n41906 , n34300 );
not ( n41908 , n41907 );
xor ( n41909 , n38220 , n39450 );
xor ( n41910 , n41909 , n39467 );
and ( n41911 , n41908 , n41910 );
xor ( n41912 , n41905 , n41911 );
not ( n12833 , n29614 );
and ( n12834 , n12833 , RI173f0f10_1581);
and ( n12835 , n41912 , n29614 );
or ( n41913 , n12834 , n12835 );
not ( n12836 , RI1754c610_2);
and ( n12837 , n12836 , n41913 );
and ( n12838 , C0 , RI1754c610_2);
or ( n41914 , n12837 , n12838 );
buf ( n41915 , n41914 );
not ( n41916 , n39962 );
and ( n41917 , n41916 , n34352 );
xor ( n41918 , n41033 , n41917 );
not ( n41919 , n39967 );
and ( n41920 , n41919 , n34361 );
xor ( n41921 , n41038 , n41920 );
xor ( n41922 , n41918 , n41921 );
not ( n41923 , n39973 );
and ( n41924 , n41923 , n34371 );
xor ( n41925 , n41044 , n41924 );
xor ( n41926 , n41922 , n41925 );
not ( n41927 , n39979 );
and ( n41928 , n41927 , n34381 );
xor ( n41929 , n34348 , n41928 );
xor ( n41930 , n41926 , n41929 );
not ( n41931 , n39985 );
and ( n41932 , n41931 , n34387 );
xor ( n41933 , n40617 , n41932 );
xor ( n41934 , n41930 , n41933 );
xor ( n41935 , n39976 , n41934 );
xor ( n41936 , n41935 , n40341 );
not ( n41937 , n41893 );
and ( n41938 , n41937 , n41895 );
xor ( n41939 , n41936 , n41938 );
not ( n12839 , n29614 );
and ( n12840 , n12839 , RI174a5528_930);
and ( n12841 , n41939 , n29614 );
or ( n41940 , n12840 , n12841 );
not ( n12842 , RI1754c610_2);
and ( n12843 , n12842 , n41940 );
and ( n12844 , C0 , RI1754c610_2);
or ( n41941 , n12843 , n12844 );
buf ( n41942 , n41941 );
not ( n41943 , n30428 );
and ( n41944 , n41943 , n39876 );
xor ( n41945 , n30401 , n41944 );
xor ( n41946 , n41945 , n30461 );
xor ( n41947 , n41946 , n39262 );
xor ( n41948 , n33934 , n37291 );
xor ( n41949 , n41948 , n37311 );
not ( n41950 , n41949 );
xor ( n41951 , n36311 , n40718 );
xor ( n41952 , n41951 , n38676 );
and ( n41953 , n41950 , n41952 );
xor ( n41954 , n41947 , n41953 );
not ( n12845 , n29614 );
and ( n12846 , n12845 , RI173ab358_1921);
and ( n12847 , n41954 , n29614 );
or ( n41955 , n12846 , n12847 );
not ( n12848 , RI1754c610_2);
and ( n12849 , n12848 , n41955 );
and ( n12850 , C0 , RI1754c610_2);
or ( n41956 , n12849 , n12850 );
buf ( n41957 , n41956 );
xor ( n41958 , n40201 , n34041 );
xor ( n41959 , n41958 , n41934 );
xor ( n41960 , n33376 , n39005 );
xor ( n41961 , n41960 , n39543 );
not ( n41962 , n41961 );
xor ( n41963 , n35051 , n37814 );
xor ( n41964 , n41963 , n33223 );
and ( n41965 , n41962 , n41964 );
xor ( n41966 , n41959 , n41965 );
not ( n12851 , n29614 );
and ( n12852 , n12851 , RI1748b128_1058);
and ( n12853 , n41966 , n29614 );
or ( n41967 , n12852 , n12853 );
not ( n12854 , RI1754c610_2);
and ( n12855 , n12854 , n41967 );
and ( n12856 , C0 , RI1754c610_2);
or ( n41968 , n12855 , n12856 );
buf ( n41969 , n41968 );
xor ( n41970 , n35064 , n33223 );
xor ( n41971 , n41970 , n33282 );
not ( n41972 , n35284 );
and ( n41973 , n41972 , n30250 );
xor ( n41974 , n39859 , n41973 );
not ( n41975 , n35289 );
and ( n41976 , n41975 , n30284 );
xor ( n41977 , n39864 , n41976 );
xor ( n41978 , n41974 , n41977 );
not ( n41979 , n35295 );
and ( n41980 , n41979 , n30350 );
xor ( n41981 , n39870 , n41980 );
xor ( n41982 , n41978 , n41981 );
not ( n41983 , n35301 );
and ( n41984 , n41983 , n30391 );
xor ( n41985 , n39876 , n41984 );
xor ( n41986 , n41982 , n41985 );
not ( n41987 , n35307 );
and ( n41988 , n41987 , n30433 );
xor ( n41989 , n39882 , n41988 );
xor ( n41990 , n41986 , n41989 );
xor ( n41991 , n35310 , n41990 );
xor ( n41992 , n41991 , n41005 );
not ( n41993 , n41992 );
xor ( n41994 , n40347 , n37898 );
xor ( n41995 , n41994 , n37915 );
and ( n41996 , n41993 , n41995 );
xor ( n41997 , n41971 , n41996 );
not ( n12857 , n29614 );
and ( n12858 , n12857 , RI17520858_665);
and ( n12859 , n41997 , n29614 );
or ( n41998 , n12858 , n12859 );
not ( n12860 , RI1754c610_2);
and ( n12861 , n12860 , n41998 );
and ( n12862 , C0 , RI1754c610_2);
or ( n41999 , n12861 , n12862 );
buf ( n42000 , n41999 );
xor ( n42001 , n34582 , n35544 );
xor ( n42002 , n42001 , n35594 );
xor ( n42003 , n39727 , n39506 );
xor ( n42004 , n42003 , n38150 );
not ( n42005 , n42004 );
not ( n42006 , n30375 );
and ( n42007 , n42006 , n39870 );
xor ( n42008 , n30352 , n42007 );
xor ( n42009 , n42008 , n30461 );
xor ( n42010 , n42009 , n39262 );
and ( n42011 , n42005 , n42010 );
xor ( n42012 , n42002 , n42011 );
not ( n12863 , n29614 );
and ( n12864 , n12863 , RI174479a0_1387);
and ( n12865 , n42012 , n29614 );
or ( n42013 , n12864 , n12865 );
not ( n12866 , RI1754c610_2);
and ( n12867 , n12866 , n42013 );
and ( n12868 , C0 , RI1754c610_2);
or ( n42014 , n12867 , n12868 );
buf ( n42015 , n42014 );
xor ( n42016 , n40888 , n34340 );
xor ( n42017 , n42016 , n38817 );
not ( n42018 , n41033 );
and ( n42019 , n42018 , n39962 );
xor ( n42020 , n34357 , n42019 );
not ( n42021 , n41038 );
and ( n42022 , n42021 , n39967 );
xor ( n42023 , n34366 , n42022 );
xor ( n42024 , n42020 , n42023 );
not ( n42025 , n41044 );
and ( n42026 , n42025 , n39973 );
xor ( n42027 , n34376 , n42026 );
xor ( n42028 , n42024 , n42027 );
xor ( n42029 , n42028 , n41484 );
not ( n42030 , n40617 );
and ( n42031 , n42030 , n39985 );
xor ( n42032 , n34392 , n42031 );
xor ( n42033 , n42029 , n42032 );
xor ( n42034 , n41933 , n42033 );
xor ( n42035 , n42034 , n37987 );
not ( n42036 , n42035 );
not ( n42037 , n31216 );
and ( n42038 , n42037 , n31227 );
xor ( n42039 , n33625 , n42038 );
xor ( n42040 , n42039 , n41265 );
not ( n42041 , n31257 );
and ( n42042 , n42041 , n31259 );
xor ( n42043 , n33186 , n42042 );
xor ( n42044 , n42040 , n42043 );
not ( n42045 , n31267 );
and ( n42046 , n42045 , n31280 );
xor ( n42047 , n33640 , n42046 );
xor ( n42048 , n42044 , n42047 );
xor ( n42049 , n42048 , n33623 );
xor ( n42050 , n31234 , n42049 );
xor ( n42051 , n42050 , n37849 );
and ( n42052 , n42036 , n42051 );
xor ( n42053 , n42017 , n42052 );
not ( n12869 , n29614 );
and ( n12870 , n12869 , RI173fa948_1534);
and ( n12871 , n42053 , n29614 );
or ( n42054 , n12870 , n12871 );
not ( n12872 , RI1754c610_2);
and ( n12873 , n12872 , n42054 );
and ( n12874 , C0 , RI1754c610_2);
or ( n42055 , n12873 , n12874 );
buf ( n42056 , n42055 );
xor ( n42057 , n38589 , n29109 );
xor ( n42058 , n42057 , n40463 );
not ( n42059 , n41126 );
and ( n42060 , n42059 , n41128 );
xor ( n42061 , n42058 , n42060 );
not ( n12875 , n29614 );
and ( n12876 , n12875 , RI174968e8_1002);
and ( n12877 , n42061 , n29614 );
or ( n42062 , n12876 , n12877 );
not ( n12878 , RI1754c610_2);
and ( n12879 , n12878 , n42062 );
and ( n12880 , C0 , RI1754c610_2);
or ( n42063 , n12879 , n12880 );
buf ( n42064 , n42063 );
buf ( n42065 , RI174aadc0_903);
not ( n12881 , n27683 );
and ( n12882 , n12881 , RI19ac6bc0_2279);
and ( n12883 , RI19acf680_2215 , n27683 );
or ( n42066 , n12882 , n12883 );
not ( n12884 , RI1754c610_2);
and ( n12885 , n12884 , n42066 );
and ( n12886 , C0 , RI1754c610_2);
or ( n42067 , n12885 , n12886 );
buf ( n42068 , n42067 );
buf ( n42069 , RI174b1378_872);
xor ( n42070 , n33656 , n41854 );
xor ( n42071 , n42070 , n40283 );
xor ( n42072 , n29697 , n39091 );
xor ( n42073 , n42072 , n36128 );
not ( n42074 , n42073 );
xor ( n42075 , n39629 , n35176 );
xor ( n42076 , n42075 , n35216 );
and ( n42077 , n42074 , n42076 );
xor ( n42078 , n42071 , n42077 );
not ( n12887 , n29614 );
and ( n12888 , n12887 , RI173cf4d8_1745);
and ( n12889 , n42078 , n29614 );
or ( n42079 , n12888 , n12889 );
not ( n12890 , RI1754c610_2);
and ( n12891 , n12890 , n42079 );
and ( n12892 , C0 , RI1754c610_2);
or ( n42080 , n12891 , n12892 );
buf ( n42081 , n42080 );
xor ( n42082 , n39252 , n35361 );
xor ( n42083 , n42082 , n38445 );
not ( n42084 , n42083 );
xor ( n42085 , n38565 , n28816 );
xor ( n42086 , n42085 , n29109 );
and ( n42087 , n42084 , n42086 );
xor ( n42088 , n40719 , n42087 );
not ( n12893 , n29614 );
and ( n12894 , n12893 , RI173d0f18_1737);
and ( n12895 , n42088 , n29614 );
or ( n42089 , n12894 , n12895 );
not ( n12896 , RI1754c610_2);
and ( n12897 , n12896 , n42089 );
and ( n12898 , C0 , RI1754c610_2);
or ( n42090 , n12897 , n12898 );
buf ( n42091 , n42090 );
buf ( n42092 , RI174a1d60_947);
buf ( n42093 , RI174a8660_915);
xor ( n42094 , n36783 , n38214 );
xor ( n42095 , n42094 , n38244 );
xor ( n42096 , n32589 , n39182 );
xor ( n42097 , n42096 , n38991 );
not ( n42098 , n42097 );
xor ( n42099 , n37326 , n39914 );
xor ( n42100 , n42099 , n40237 );
and ( n42101 , n42098 , n42100 );
xor ( n42102 , n42095 , n42101 );
not ( n12899 , n29614 );
and ( n12900 , n12899 , RI174537f0_1329);
and ( n12901 , n42102 , n29614 );
or ( n42103 , n12900 , n12901 );
not ( n12902 , RI1754c610_2);
and ( n12903 , n12902 , n42103 );
and ( n12904 , C0 , RI1754c610_2);
or ( n42104 , n12903 , n12904 );
buf ( n42105 , n42104 );
not ( n12905 , n27683 );
and ( n12906 , n12905 , RI19a9a610_2609);
and ( n12907 , RI19aa3c88_2539 , n27683 );
or ( n42106 , n12906 , n12907 );
not ( n12908 , RI1754c610_2);
and ( n12909 , n12908 , n42106 );
and ( n12910 , C0 , RI1754c610_2);
or ( n42107 , n12909 , n12910 );
buf ( n42108 , n42107 );
buf ( n42109 , RI17472df8_1176);
buf ( n42110 , RI174796f8_1144);
xor ( n42111 , n33815 , n39414 );
xor ( n42112 , n42111 , n37186 );
xor ( n42113 , n40661 , n39282 );
xor ( n42114 , n42113 , n37676 );
not ( n42115 , n42114 );
xor ( n42116 , n38694 , n38817 );
xor ( n42117 , n42116 , n40034 );
and ( n42118 , n42115 , n42117 );
xor ( n42119 , n42112 , n42118 );
not ( n12911 , n29614 );
and ( n12912 , n12911 , RI173f81e8_1546);
and ( n12913 , n42119 , n29614 );
or ( n42120 , n12912 , n12913 );
not ( n12914 , RI1754c610_2);
and ( n12915 , n12914 , n42120 );
and ( n12916 , C0 , RI1754c610_2);
or ( n42121 , n12915 , n12916 );
buf ( n42122 , n42121 );
buf ( n42123 , RI17466918_1236);
xor ( n42124 , n36444 , n37104 );
xor ( n42125 , n42124 , n35986 );
not ( n42126 , n41571 );
and ( n42127 , n42126 , n41573 );
xor ( n42128 , n42125 , n42127 );
not ( n12917 , n29614 );
and ( n12918 , n12917 , RI17397ee8_2015);
and ( n12919 , n42128 , n29614 );
or ( n42129 , n12918 , n12919 );
not ( n12920 , RI1754c610_2);
and ( n12921 , n12920 , n42129 );
and ( n12922 , C0 , RI1754c610_2);
or ( n42130 , n12921 , n12922 );
buf ( n42131 , n42130 );
xor ( n42132 , n37902 , n32048 );
xor ( n42133 , n42132 , n32108 );
xor ( n42134 , n37703 , n40463 );
xor ( n42135 , n42134 , n41772 );
not ( n42136 , n42135 );
xor ( n42137 , n38016 , n41690 );
xor ( n42138 , n42137 , n39506 );
and ( n42139 , n42136 , n42138 );
xor ( n42140 , n42133 , n42139 );
not ( n12923 , n29614 );
and ( n12924 , n12923 , RI173cb338_1765);
and ( n12925 , n42140 , n29614 );
or ( n42141 , n12924 , n12925 );
not ( n12926 , RI1754c610_2);
and ( n12927 , n12926 , n42141 );
and ( n12928 , C0 , RI1754c610_2);
or ( n42142 , n12927 , n12928 );
buf ( n42143 , n42142 );
not ( n12929 , n27683 );
and ( n12930 , n12929 , RI19ac1850_2318);
and ( n12931 , RI19acadd8_2249 , n27683 );
or ( n42144 , n12930 , n12931 );
not ( n12932 , RI1754c610_2);
and ( n12933 , n12932 , n42144 );
and ( n12934 , C0 , RI1754c610_2);
or ( n42145 , n12933 , n12934 );
buf ( n42146 , n42145 );
not ( n42147 , n32864 );
xor ( n42148 , n37691 , n37579 );
xor ( n42149 , n42148 , n38495 );
and ( n42150 , n42147 , n42149 );
xor ( n42151 , n32716 , n42150 );
not ( n12935 , n29614 );
and ( n12936 , n12935 , RI174c9630_784);
and ( n12937 , n42151 , n29614 );
or ( n42152 , n12936 , n12937 );
not ( n12938 , RI1754c610_2);
and ( n12939 , n12938 , n42152 );
and ( n12940 , C0 , RI1754c610_2);
or ( n42153 , n12939 , n12940 );
buf ( n42154 , n42153 );
buf ( n42155 , RI17488d10_1069);
buf ( n42156 , RI1750a9b8_733);
xor ( n42157 , n39277 , n38445 );
xor ( n42158 , n42157 , n37549 );
xor ( n42159 , n32662 , n36195 );
xor ( n42160 , n42159 , n36209 );
not ( n42161 , n42160 );
xor ( n42162 , n37959 , n41504 );
xor ( n42163 , n42162 , n41690 );
and ( n42164 , n42161 , n42163 );
xor ( n42165 , n42158 , n42164 );
not ( n12941 , n29614 );
and ( n12942 , n12941 , RI173f2fe0_1571);
and ( n12943 , n42165 , n29614 );
or ( n42166 , n12942 , n12943 );
not ( n12944 , RI1754c610_2);
and ( n12945 , n12944 , n42166 );
and ( n12946 , C0 , RI1754c610_2);
or ( n42167 , n12945 , n12946 );
buf ( n42168 , n42167 );
xor ( n42169 , n37444 , n36874 );
not ( n42170 , n37463 );
and ( n42171 , n42170 , n35547 );
xor ( n42172 , n39360 , n42171 );
not ( n42173 , n37468 );
and ( n42174 , n42173 , n35556 );
xor ( n42175 , n39376 , n42174 );
xor ( n42176 , n42172 , n42175 );
not ( n42177 , n37474 );
and ( n42178 , n42177 , n35566 );
xor ( n42179 , n39382 , n42178 );
xor ( n42180 , n42176 , n42179 );
not ( n42181 , n37480 );
and ( n42182 , n42181 , n35576 );
xor ( n42183 , n39388 , n42182 );
xor ( n42184 , n42180 , n42183 );
not ( n42185 , n37486 );
and ( n42186 , n42185 , n35586 );
xor ( n42187 , n39394 , n42186 );
xor ( n42188 , n42184 , n42187 );
xor ( n42189 , n42169 , n42188 );
xor ( n42190 , n36753 , n39208 );
xor ( n42191 , n42190 , n38214 );
not ( n42192 , n42191 );
xor ( n42193 , n39273 , n38445 );
xor ( n42194 , n42193 , n37549 );
and ( n42195 , n42192 , n42194 );
xor ( n42196 , n42189 , n42195 );
not ( n12947 , n29614 );
and ( n12948 , n12947 , RI1746bb20_1211);
and ( n12949 , n42196 , n29614 );
or ( n42197 , n12948 , n12949 );
not ( n12950 , RI1754c610_2);
and ( n12951 , n12950 , n42197 );
and ( n12952 , C0 , RI1754c610_2);
or ( n42198 , n12951 , n12952 );
buf ( n42199 , n42198 );
xor ( n42200 , n34444 , n40009 );
xor ( n42201 , n42200 , n38085 );
xor ( n42202 , n40676 , n36654 );
xor ( n42203 , n42202 , n40808 );
not ( n42204 , n42203 );
xor ( n42205 , n38699 , n38817 );
xor ( n42206 , n42205 , n40034 );
and ( n42207 , n42204 , n42206 );
xor ( n42208 , n42201 , n42207 );
not ( n12953 , n29614 );
and ( n12954 , n12953 , RI173362b0_2177);
and ( n12955 , n42208 , n29614 );
or ( n42209 , n12954 , n12955 );
not ( n12956 , RI1754c610_2);
and ( n12957 , n12956 , n42209 );
and ( n12958 , C0 , RI1754c610_2);
or ( n42210 , n12957 , n12958 );
buf ( n42211 , n42210 );
not ( n12959 , n27683 );
and ( n12960 , n12959 , RI19a8a878_2721);
and ( n12961 , RI19a946e8_2651 , n27683 );
or ( n42212 , n12960 , n12961 );
not ( n12962 , RI1754c610_2);
and ( n12963 , n12962 , n42212 );
and ( n12964 , C0 , RI1754c610_2);
or ( n42213 , n12963 , n12964 );
buf ( n42214 , n42213 );
not ( n12965 , n27683 );
and ( n12966 , n12965 , RI19ac0ba8_2325);
and ( n12967 , RI19ac9de8_2256 , n27683 );
or ( n42215 , n12966 , n12967 );
not ( n12968 , RI1754c610_2);
and ( n12969 , n12968 , n42215 );
and ( n12970 , C0 , RI1754c610_2);
or ( n42216 , n12969 , n12970 );
buf ( n42217 , n42216 );
not ( n12971 , n27683 );
and ( n12972 , n12971 , RI19a9e8a0_2580);
and ( n12973 , RI19aa8080_2509 , n27683 );
or ( n42218 , n12972 , n12973 );
not ( n12974 , RI1754c610_2);
and ( n12975 , n12974 , n42218 );
and ( n12976 , C0 , RI1754c610_2);
or ( n42219 , n12975 , n12976 );
buf ( n42220 , n42219 );
not ( n12977 , n27683 );
and ( n12978 , n12977 , RI19a85058_2759);
and ( n12979 , RI19ac4f28_2292 , n27683 );
or ( n42221 , n12978 , n12979 );
not ( n12980 , RI1754c610_2);
and ( n12981 , n12980 , n42221 );
and ( n12982 , C0 , RI1754c610_2);
or ( n42222 , n12981 , n12982 );
buf ( n42223 , n42222 );
xor ( n42224 , n39681 , n33617 );
xor ( n42225 , n42224 , n39525 );
xor ( n42226 , n35493 , n38512 );
xor ( n42227 , n42226 , n38532 );
not ( n42228 , n42227 );
and ( n42229 , n42228 , n39283 );
xor ( n42230 , n42225 , n42229 );
not ( n12983 , n29614 );
and ( n12984 , n12983 , RI173ad0e0_1912);
and ( n12985 , n42230 , n29614 );
or ( n42231 , n12984 , n12985 );
not ( n12986 , RI1754c610_2);
and ( n12987 , n12986 , n42231 );
and ( n12988 , C0 , RI1754c610_2);
or ( n42232 , n12987 , n12988 );
buf ( n42233 , n42232 );
xor ( n42234 , n38205 , n37696 );
xor ( n42235 , n42234 , n39450 );
xor ( n42236 , n40435 , n39816 );
xor ( n42237 , n42236 , n35052 );
not ( n42238 , n42237 );
xor ( n42239 , n34496 , n29610 );
xor ( n42240 , n42239 , n31380 );
and ( n42241 , n42238 , n42240 );
xor ( n42242 , n42235 , n42241 );
not ( n12989 , n29614 );
and ( n12990 , n12989 , RI174893a0_1067);
and ( n12991 , n42242 , n29614 );
or ( n42243 , n12990 , n12991 );
not ( n12992 , RI1754c610_2);
and ( n12993 , n12992 , n42243 );
and ( n12994 , C0 , RI1754c610_2);
or ( n42244 , n12993 , n12994 );
buf ( n42245 , n42244 );
not ( n42246 , n34153 );
and ( n42247 , n42246 , n34155 );
xor ( n42248 , n31848 , n42247 );
not ( n42249 , n34160 );
and ( n42250 , n42249 , n34162 );
xor ( n42251 , n31858 , n42250 );
xor ( n42252 , n42248 , n42251 );
not ( n42253 , n34168 );
and ( n42254 , n42253 , n34170 );
xor ( n42255 , n31881 , n42254 );
xor ( n42256 , n42252 , n42255 );
not ( n42257 , n34176 );
and ( n42258 , n42257 , n34178 );
xor ( n42259 , n31891 , n42258 );
xor ( n42260 , n42256 , n42259 );
not ( n42261 , n34184 );
and ( n42262 , n42261 , n34186 );
xor ( n42263 , n31922 , n42262 );
xor ( n42264 , n42260 , n42263 );
xor ( n42265 , n34165 , n42264 );
xor ( n42266 , n42265 , n41370 );
xor ( n42267 , n34238 , n37526 );
xor ( n42268 , n42267 , n41049 );
not ( n42269 , n42268 );
xor ( n42270 , n35795 , n37331 );
xor ( n42271 , n42270 , n37129 );
and ( n42272 , n42269 , n42271 );
xor ( n42273 , n42266 , n42272 );
not ( n12995 , n29614 );
and ( n12996 , n12995 , RI174c43b0_800);
and ( n12997 , n42273 , n29614 );
or ( n42274 , n12996 , n12997 );
not ( n12998 , RI1754c610_2);
and ( n12999 , n12998 , n42274 );
and ( n13000 , C0 , RI1754c610_2);
or ( n42275 , n12999 , n13000 );
buf ( n42276 , n42275 );
xor ( n42277 , n37650 , n40149 );
xor ( n42278 , n42277 , n40166 );
xor ( n42279 , n31119 , n40828 );
xor ( n42280 , n42279 , n42049 );
not ( n42281 , n42280 );
xor ( n42282 , n38581 , n29109 );
xor ( n42283 , n42282 , n40463 );
and ( n42284 , n42281 , n42283 );
xor ( n42285 , n42278 , n42284 );
not ( n13001 , n29614 );
and ( n13002 , n13001 , RI173d9270_1697);
and ( n13003 , n42285 , n29614 );
or ( n42286 , n13002 , n13003 );
not ( n13004 , RI1754c610_2);
and ( n13005 , n13004 , n42286 );
and ( n13006 , C0 , RI1754c610_2);
or ( n42287 , n13005 , n13006 );
buf ( n42288 , n42287 );
buf ( n42289 , RI174713b8_1184);
buf ( n42290 , RI17500530_759);
buf ( n42291 , RI17466288_1238);
not ( n42292 , n40529 );
xor ( n42293 , n38516 , n31725 );
not ( n42294 , n38898 );
and ( n42295 , n42294 , n38900 );
xor ( n42296 , n33736 , n42295 );
xor ( n42297 , n42296 , n40924 );
not ( n42298 , n38913 );
and ( n42299 , n42298 , n38915 );
xor ( n42300 , n33755 , n42299 );
xor ( n42301 , n42297 , n42300 );
not ( n42302 , n38741 );
and ( n42303 , n42302 , n38921 );
xor ( n42304 , n33765 , n42303 );
xor ( n42305 , n42301 , n42304 );
not ( n42306 , n38927 );
and ( n42307 , n42306 , n38929 );
xor ( n42308 , n33775 , n42307 );
xor ( n42309 , n42305 , n42308 );
xor ( n42310 , n42293 , n42309 );
and ( n42311 , n42292 , n42310 );
xor ( n42312 , n40526 , n42311 );
not ( n13007 , n29614 );
and ( n13008 , n13007 , RI173b1280_1892);
and ( n13009 , n42312 , n29614 );
or ( n42313 , n13008 , n13009 );
not ( n13010 , RI1754c610_2);
and ( n13011 , n13010 , n42313 );
and ( n13012 , C0 , RI1754c610_2);
or ( n42314 , n13011 , n13012 );
buf ( n42315 , n42314 );
not ( n42316 , n29422 );
and ( n42317 , n42316 , n35003 );
xor ( n42318 , n29400 , n42317 );
xor ( n42319 , n42318 , n29425 );
xor ( n42320 , n42319 , n29610 );
xor ( n42321 , n39434 , n38495 );
xor ( n42322 , n42321 , n36611 );
not ( n42323 , n42322 );
xor ( n42324 , n38254 , n36530 );
xor ( n42325 , n42324 , n36568 );
and ( n42326 , n42323 , n42325 );
xor ( n42327 , n42320 , n42326 );
not ( n13013 , n29614 );
and ( n13014 , n13013 , RI1752e0e8_623);
and ( n13015 , n42327 , n29614 );
or ( n42328 , n13014 , n13015 );
not ( n13016 , RI1754c610_2);
and ( n13017 , n13016 , n42328 );
and ( n13018 , C0 , RI1754c610_2);
or ( n42329 , n13017 , n13018 );
buf ( n42330 , n42329 );
xor ( n42331 , n38671 , n39347 );
not ( n42332 , n27792 );
and ( n42333 , n42332 , n27713 );
xor ( n42334 , n29857 , n42333 );
not ( n42335 , n27820 );
and ( n42336 , n42335 , n27845 );
xor ( n42337 , n29876 , n42336 );
xor ( n42338 , n42334 , n42337 );
xor ( n42339 , n42338 , n35915 );
not ( n42340 , n27976 );
and ( n42341 , n42340 , n28002 );
xor ( n42342 , n29936 , n42341 );
xor ( n42343 , n42339 , n42342 );
xor ( n42344 , n42343 , n37349 );
xor ( n42345 , n42331 , n42344 );
xor ( n42346 , n38885 , n31506 );
xor ( n42347 , n42346 , n31621 );
not ( n42348 , n42347 );
xor ( n42349 , n36583 , n39791 );
xor ( n42350 , n42349 , n40915 );
and ( n42351 , n42348 , n42350 );
xor ( n42352 , n42345 , n42351 );
not ( n13019 , n29614 );
and ( n13020 , n13019 , RI173f1258_1580);
and ( n13021 , n42352 , n29614 );
or ( n42353 , n13020 , n13021 );
not ( n13022 , RI1754c610_2);
and ( n13023 , n13022 , n42353 );
and ( n13024 , C0 , RI1754c610_2);
or ( n42354 , n13023 , n13024 );
buf ( n42355 , n42354 );
xor ( n42356 , n34405 , n40009 );
xor ( n42357 , n42356 , n38085 );
xor ( n42358 , n37242 , n41391 );
xor ( n42359 , n42358 , n39686 );
not ( n42360 , n42359 );
xor ( n42361 , n39537 , n35842 );
xor ( n42362 , n42361 , n38401 );
and ( n42363 , n42360 , n42362 );
xor ( n42364 , n42357 , n42363 );
not ( n13025 , n29614 );
and ( n13026 , n13025 , RI17445c18_1396);
and ( n13027 , n42364 , n29614 );
or ( n42365 , n13026 , n13027 );
not ( n13028 , RI1754c610_2);
and ( n13029 , n13028 , n42365 );
and ( n13030 , C0 , RI1754c610_2);
or ( n42366 , n13029 , n13030 );
buf ( n42367 , n42366 );
xor ( n42368 , n37362 , n33505 );
xor ( n42369 , n42368 , n39635 );
xor ( n42370 , n34078 , n39525 );
xor ( n42371 , n36883 , n41449 );
xor ( n42372 , n42371 , n40215 );
not ( n42373 , n34113 );
and ( n42374 , n42373 , n34115 );
xor ( n42375 , n33922 , n42374 );
xor ( n42376 , n42372 , n42375 );
xor ( n42377 , n42376 , n36415 );
xor ( n42378 , n42370 , n42377 );
not ( n42379 , n42378 );
xor ( n42380 , n33823 , n39414 );
xor ( n42381 , n42380 , n37186 );
and ( n42382 , n42379 , n42381 );
xor ( n42383 , n42369 , n42382 );
not ( n13031 , n29614 );
and ( n13032 , n13031 , RI17512fc8_707);
and ( n13033 , n42383 , n29614 );
or ( n42384 , n13032 , n13033 );
not ( n13034 , RI1754c610_2);
and ( n13035 , n13034 , n42384 );
and ( n13036 , C0 , RI1754c610_2);
or ( n42385 , n13035 , n13036 );
buf ( n42386 , n42385 );
xor ( n42387 , n39166 , n40166 );
xor ( n42388 , n42387 , n41590 );
not ( n42389 , n32974 );
and ( n42390 , n42389 , n33070 );
xor ( n42391 , n42388 , n42390 );
not ( n13037 , n29614 );
and ( n13038 , n13037 , RI174b4b40_855);
and ( n13039 , n42391 , n29614 );
or ( n42392 , n13038 , n13039 );
not ( n13040 , RI1754c610_2);
and ( n13041 , n13040 , n42392 );
and ( n13042 , C0 , RI1754c610_2);
or ( n42393 , n13041 , n13042 );
buf ( n42394 , n42393 );
not ( n13043 , n27683 );
and ( n13044 , n13043 , RI19a9f548_2574);
and ( n13045 , RI19aa90e8_2502 , n27683 );
or ( n42395 , n13044 , n13045 );
not ( n13046 , RI1754c610_2);
and ( n13047 , n13046 , n42395 );
and ( n13048 , C0 , RI1754c610_2);
or ( n42396 , n13047 , n13048 );
buf ( n42397 , n42396 );
xor ( n42398 , n35985 , n37744 );
xor ( n42399 , n42398 , n35438 );
not ( n42400 , n42399 );
xor ( n42401 , n39965 , n41934 );
xor ( n42402 , n42401 , n40341 );
and ( n42403 , n42400 , n42402 );
xor ( n42404 , n41820 , n42403 );
not ( n13049 , n29614 );
and ( n13050 , n13049 , RI173f2c98_1572);
and ( n13051 , n42404 , n29614 );
or ( n42405 , n13050 , n13051 );
not ( n13052 , RI1754c610_2);
and ( n13053 , n13052 , n42405 );
and ( n13054 , C0 , RI1754c610_2);
or ( n42406 , n13053 , n13054 );
buf ( n42407 , n42406 );
xor ( n42408 , n38519 , n31725 );
xor ( n42409 , n42408 , n42309 );
xor ( n42410 , n30571 , n38167 );
xor ( n42411 , n42410 , n33728 );
not ( n42412 , n42411 );
xor ( n42413 , n36143 , n39151 );
xor ( n42414 , n42413 , n38267 );
and ( n42415 , n42412 , n42414 );
xor ( n42416 , n42409 , n42415 );
not ( n13055 , n29614 );
and ( n13056 , n13055 , RI1747df28_1122);
and ( n13057 , n42416 , n29614 );
or ( n42417 , n13056 , n13057 );
not ( n13058 , RI1754c610_2);
and ( n13059 , n13058 , n42417 );
and ( n13060 , C0 , RI1754c610_2);
or ( n42418 , n13059 , n13060 );
buf ( n42419 , n42418 );
xor ( n42420 , n36765 , n39208 );
xor ( n42421 , n42420 , n38214 );
not ( n42422 , n38934 );
and ( n42423 , n42422 , n38949 );
xor ( n42424 , n42421 , n42423 );
not ( n13061 , n29614 );
and ( n13062 , n13061 , RI175274a0_644);
and ( n13063 , n42424 , n29614 );
or ( n42425 , n13062 , n13063 );
not ( n13064 , RI1754c610_2);
and ( n13065 , n13064 , n42425 );
and ( n13066 , C0 , RI1754c610_2);
or ( n42426 , n13065 , n13066 );
buf ( n42427 , n42426 );
xor ( n42428 , n37073 , n38594 );
xor ( n42429 , n42428 , n37716 );
xor ( n42430 , n41530 , n32786 );
xor ( n42431 , n42430 , n32863 );
not ( n42432 , n42431 );
xor ( n42433 , n37222 , n39467 );
xor ( n42434 , n42433 , n41391 );
and ( n42435 , n42432 , n42434 );
xor ( n42436 , n42429 , n42435 );
not ( n13067 , n29614 );
and ( n13068 , n13067 , RI174a6c20_923);
and ( n13069 , n42436 , n29614 );
or ( n42437 , n13068 , n13069 );
not ( n13070 , RI1754c610_2);
and ( n13071 , n13070 , n42437 );
and ( n13072 , C0 , RI1754c610_2);
or ( n42438 , n13071 , n13072 );
buf ( n42439 , n42438 );
not ( n13073 , n27683 );
and ( n13074 , n13073 , RI19a83d20_2767);
and ( n13075 , RI19ab9df8_2381 , n27683 );
or ( n42440 , n13074 , n13075 );
not ( n13076 , RI1754c610_2);
and ( n13077 , n13076 , n42440 );
and ( n13078 , C0 , RI1754c610_2);
or ( n42441 , n13077 , n13078 );
buf ( n42442 , n42441 );
xor ( n42443 , n39685 , n33617 );
xor ( n42444 , n42443 , n39525 );
xor ( n42445 , n29666 , n39091 );
xor ( n42446 , n42445 , n36128 );
not ( n42447 , n42446 );
xor ( n42448 , n29276 , n40034 );
xor ( n42449 , n42448 , n40051 );
and ( n42450 , n42447 , n42449 );
xor ( n42451 , n42444 , n42450 );
not ( n13079 , n29614 );
and ( n13080 , n13079 , RI1749f600_959);
and ( n13081 , n42451 , n29614 );
or ( n42452 , n13080 , n13081 );
not ( n13082 , RI1754c610_2);
and ( n13083 , n13082 , n42452 );
and ( n13084 , C0 , RI1754c610_2);
or ( n42453 , n13083 , n13084 );
buf ( n42454 , n42453 );
xor ( n42455 , n40156 , n39039 );
xor ( n42456 , n42455 , n39065 );
xor ( n42457 , n37246 , n41391 );
xor ( n42458 , n42457 , n39686 );
not ( n42459 , n42458 );
xor ( n42460 , n39909 , n33397 );
xor ( n42461 , n42460 , n35710 );
and ( n42462 , n42459 , n42461 );
xor ( n42463 , n42456 , n42462 );
not ( n13085 , n29614 );
and ( n13086 , n13085 , RI1738c098_2073);
and ( n13087 , n42463 , n29614 );
or ( n42464 , n13086 , n13087 );
not ( n13088 , RI1754c610_2);
and ( n13089 , n13088 , n42464 );
and ( n13090 , C0 , RI1754c610_2);
or ( n42465 , n13089 , n13090 );
buf ( n42466 , n42465 );
xor ( n42467 , n32480 , n35622 );
xor ( n42468 , n42467 , n35639 );
xor ( n42469 , n35380 , n41068 );
xor ( n42470 , n42469 , n39091 );
not ( n42471 , n42470 );
xor ( n42472 , n33672 , n41854 );
xor ( n42473 , n42472 , n40283 );
and ( n42474 , n42471 , n42473 );
xor ( n42475 , n42468 , n42474 );
not ( n13091 , n29614 );
and ( n13092 , n13091 , RI17338d58_2164);
and ( n13093 , n42475 , n29614 );
or ( n42476 , n13092 , n13093 );
not ( n13094 , RI1754c610_2);
and ( n13095 , n13094 , n42476 );
and ( n13096 , C0 , RI1754c610_2);
or ( n42477 , n13095 , n13096 );
buf ( n42478 , n42477 );
xor ( n42479 , n35304 , n41990 );
xor ( n42480 , n42479 , n41005 );
xor ( n42481 , n35910 , n36463 );
xor ( n42482 , n42481 , n32220 );
not ( n42483 , n42482 );
xor ( n42484 , n37502 , n37942 );
xor ( n42485 , n42484 , n34395 );
and ( n42486 , n42483 , n42485 );
xor ( n42487 , n42480 , n42486 );
not ( n13097 , n29614 );
and ( n13098 , n13097 , RI173f2950_1573);
and ( n13099 , n42487 , n29614 );
or ( n42488 , n13098 , n13099 );
not ( n13100 , RI1754c610_2);
and ( n13101 , n13100 , n42488 );
and ( n13102 , C0 , RI1754c610_2);
or ( n42489 , n13101 , n13102 );
buf ( n42490 , n42489 );
xor ( n42491 , n39855 , n36742 );
not ( n42492 , n30258 );
and ( n42493 , n42492 , n39859 );
xor ( n42494 , n30253 , n42493 );
not ( n42495 , n30333 );
and ( n42496 , n42495 , n39864 );
xor ( n42497 , n30307 , n42496 );
xor ( n42498 , n42494 , n42497 );
xor ( n42499 , n42498 , n42008 );
xor ( n42500 , n42499 , n41945 );
not ( n42501 , n30458 );
and ( n42502 , n42501 , n39882 );
xor ( n42503 , n30445 , n42502 );
xor ( n42504 , n42500 , n42503 );
xor ( n42505 , n42491 , n42504 );
xor ( n42506 , n41231 , n38634 );
xor ( n42507 , n42506 , n38648 );
not ( n42508 , n42507 );
xor ( n42509 , n35990 , n35438 );
xor ( n42510 , n42509 , n35458 );
and ( n42511 , n42508 , n42510 );
xor ( n42512 , n42505 , n42511 );
not ( n13103 , n29614 );
and ( n13104 , n13103 , RI17406108_1478);
and ( n13105 , n42512 , n29614 );
or ( n42513 , n13104 , n13105 );
not ( n13106 , RI1754c610_2);
and ( n13107 , n13106 , n42513 );
and ( n13108 , C0 , RI1754c610_2);
or ( n42514 , n13107 , n13108 );
buf ( n42515 , n42514 );
not ( n13109 , n27683 );
and ( n13110 , n13109 , RI19a9efa8_2577);
and ( n13111 , RI19aa8878_2506 , n27683 );
or ( n42516 , n13110 , n13111 );
not ( n13112 , RI1754c610_2);
and ( n13113 , n13112 , n42516 );
and ( n13114 , C0 , RI1754c610_2);
or ( n42517 , n13113 , n13114 );
buf ( n42518 , n42517 );
xor ( n42519 , n29939 , n36128 );
xor ( n42520 , n42519 , n36148 );
xor ( n42521 , n39934 , n40890 );
xor ( n42522 , n42521 , n38724 );
not ( n42523 , n42522 );
xor ( n42524 , n34769 , n37255 );
xor ( n42525 , n42524 , n41478 );
and ( n42526 , n42523 , n42525 );
xor ( n42527 , n42520 , n42526 );
not ( n13115 , n29614 );
and ( n13116 , n13115 , RI173f15a0_1579);
and ( n13117 , n42527 , n29614 );
or ( n42528 , n13116 , n13117 );
not ( n13118 , RI1754c610_2);
and ( n13119 , n13118 , n42528 );
and ( n13120 , C0 , RI1754c610_2);
or ( n42529 , n13119 , n13120 );
buf ( n42530 , n42529 );
xor ( n42531 , n39199 , n37676 );
xor ( n42532 , n42531 , n37696 );
xor ( n42533 , n40407 , n32973 );
xor ( n42534 , n42533 , n39816 );
not ( n42535 , n42534 );
not ( n42536 , n37387 );
and ( n42537 , n42536 , n36487 );
xor ( n42538 , n36483 , n42537 );
not ( n42539 , n37394 );
and ( n42540 , n42539 , n36492 );
xor ( n42541 , n37391 , n42540 );
xor ( n42542 , n42538 , n42541 );
not ( n42543 , n37402 );
and ( n42544 , n42543 , n36502 );
xor ( n42545 , n37399 , n42544 );
xor ( n42546 , n42542 , n42545 );
not ( n42547 , n37410 );
and ( n42548 , n42547 , n36512 );
xor ( n42549 , n37407 , n42548 );
xor ( n42550 , n42546 , n42549 );
not ( n42551 , n37418 );
and ( n42552 , n42551 , n36522 );
xor ( n42553 , n37415 , n42552 );
xor ( n42554 , n42550 , n42553 );
xor ( n42555 , n40380 , n42554 );
xor ( n42556 , n42555 , n34725 );
and ( n42557 , n42535 , n42556 );
xor ( n42558 , n42532 , n42557 );
not ( n13121 , n29614 );
and ( n13122 , n13121 , RI17508ac8_739);
and ( n13123 , n42558 , n29614 );
or ( n42559 , n13122 , n13123 );
not ( n13124 , RI1754c610_2);
and ( n13125 , n13124 , n42559 );
and ( n13126 , C0 , RI1754c610_2);
or ( n42560 , n13125 , n13126 );
buf ( n42561 , n42560 );
not ( n42562 , n36703 );
xor ( n42563 , n41315 , n41526 );
xor ( n42564 , n42563 , n41543 );
and ( n42565 , n42562 , n42564 );
xor ( n42566 , n35843 , n42565 );
not ( n13127 , n29614 );
and ( n13128 , n13127 , RI17486268_1082);
and ( n13129 , n42566 , n29614 );
or ( n42567 , n13128 , n13129 );
not ( n13130 , RI1754c610_2);
and ( n13131 , n13130 , n42567 );
and ( n13132 , C0 , RI1754c610_2);
or ( n42568 , n13131 , n13132 );
buf ( n42569 , n42568 );
not ( n13133 , n27683 );
and ( n13134 , n13133 , RI19acf1d0_2217);
and ( n13135 , RI19a9fcc8_2570 , n27683 );
or ( n42570 , n13134 , n13135 );
not ( n13136 , RI1754c610_2);
and ( n13137 , n13136 , n42570 );
and ( n13138 , C0 , RI1754c610_2);
or ( n42571 , n13137 , n13138 );
buf ( n42572 , n42571 );
xor ( n42573 , n31536 , n39935 );
xor ( n42574 , n42573 , n39952 );
xor ( n42575 , n32942 , n41659 );
xor ( n42576 , n42575 , n37800 );
not ( n42577 , n42576 );
xor ( n42578 , n38523 , n31725 );
xor ( n42579 , n42578 , n42309 );
and ( n42580 , n42577 , n42579 );
xor ( n42581 , n42574 , n42580 );
not ( n13139 , n29614 );
and ( n13140 , n13139 , RI173cc3a0_1760);
and ( n13141 , n42581 , n29614 );
or ( n42582 , n13140 , n13141 );
not ( n13142 , RI1754c610_2);
and ( n13143 , n13142 , n42582 );
and ( n13144 , C0 , RI1754c610_2);
or ( n42583 , n13143 , n13144 );
buf ( n42584 , n42583 );
not ( n13145 , n27683 );
and ( n13146 , n13145 , RI19aa6b68_2518);
and ( n13147 , RI19ab0e10_2447 , n27683 );
or ( n42585 , n13146 , n13147 );
not ( n13148 , RI1754c610_2);
and ( n13149 , n13148 , n42585 );
and ( n13150 , C0 , RI1754c610_2);
or ( n42586 , n13149 , n13150 );
buf ( n42587 , n42586 );
xor ( n42588 , n38473 , n39771 );
xor ( n42589 , n42588 , n39791 );
not ( n42590 , n34682 );
and ( n42591 , n42590 , n34673 );
xor ( n42592 , n36534 , n42591 );
not ( n42593 , n34687 );
and ( n42594 , n42593 , n34689 );
xor ( n42595 , n36541 , n42594 );
xor ( n42596 , n42592 , n42595 );
not ( n42597 , n34697 );
and ( n42598 , n42597 , n34699 );
xor ( n42599 , n36549 , n42598 );
xor ( n42600 , n42596 , n42599 );
xor ( n42601 , n42600 , n40776 );
not ( n42602 , n34717 );
and ( n42603 , n42602 , n34719 );
xor ( n42604 , n36565 , n42603 );
xor ( n42605 , n42601 , n42604 );
xor ( n42606 , n34694 , n42605 );
not ( n42607 , n34733 );
and ( n42608 , n42607 , n30075 );
xor ( n42609 , n30031 , n42608 );
xor ( n42610 , n39837 , n42609 );
xor ( n42611 , n42610 , n40115 );
not ( n42612 , n34745 );
and ( n42613 , n42612 , n30166 );
xor ( n42614 , n36733 , n42613 );
xor ( n42615 , n42611 , n42614 );
not ( n42616 , n34751 );
and ( n42617 , n42616 , n30219 );
xor ( n42618 , n36739 , n42617 );
xor ( n42619 , n42615 , n42618 );
xor ( n42620 , n42606 , n42619 );
not ( n42621 , n42620 );
xor ( n42622 , n40799 , n40437 );
xor ( n42623 , n38833 , n35019 );
not ( n42624 , n35033 );
and ( n42625 , n42624 , n31163 );
xor ( n42626 , n35030 , n42625 );
xor ( n42627 , n42623 , n42626 );
not ( n42628 , n35041 );
and ( n42629 , n42628 , n31193 );
xor ( n42630 , n35038 , n42629 );
xor ( n42631 , n42627 , n42630 );
not ( n42632 , n35049 );
and ( n42633 , n42632 , n31203 );
xor ( n42634 , n35046 , n42633 );
xor ( n42635 , n42631 , n42634 );
xor ( n42636 , n42622 , n42635 );
and ( n42637 , n42621 , n42636 );
xor ( n42638 , n42589 , n42637 );
not ( n13151 , n29614 );
and ( n13152 , n13151 , RI17414d48_1406);
and ( n13153 , n42638 , n29614 );
or ( n42639 , n13152 , n13153 );
not ( n13154 , RI1754c610_2);
and ( n13155 , n13154 , n42639 );
and ( n13156 , C0 , RI1754c610_2);
or ( n42640 , n13155 , n13156 );
buf ( n42641 , n42640 );
xor ( n42642 , n37882 , n36102 );
xor ( n42643 , n42642 , n32048 );
xor ( n42644 , n35563 , n37490 );
xor ( n42645 , n42644 , n41316 );
not ( n42646 , n42645 );
xor ( n42647 , n39677 , n33617 );
xor ( n42648 , n42647 , n39525 );
and ( n42649 , n42646 , n42648 );
xor ( n42650 , n42643 , n42649 );
not ( n13157 , n29614 );
and ( n13158 , n13157 , RI17449728_1378);
and ( n13159 , n42650 , n29614 );
or ( n42651 , n13158 , n13159 );
not ( n13160 , RI1754c610_2);
and ( n13161 , n13160 , n42651 );
and ( n13162 , C0 , RI1754c610_2);
or ( n42652 , n13161 , n13162 );
buf ( n42653 , n42652 );
xor ( n42654 , n36735 , n30247 );
xor ( n42655 , n42654 , n30461 );
not ( n42656 , n40464 );
and ( n42657 , n42656 , n40466 );
xor ( n42658 , n42655 , n42657 );
not ( n13163 , n29614 );
and ( n13164 , n13163 , RI173f2608_1574);
and ( n13165 , n42658 , n29614 );
or ( n42659 , n13164 , n13165 );
not ( n13166 , RI1754c610_2);
and ( n13167 , n13166 , n42659 );
and ( n13168 , C0 , RI1754c610_2);
or ( n42660 , n13167 , n13168 );
buf ( n42661 , n42660 );
not ( n13169 , n27683 );
and ( n13170 , n13169 , RI19aaeea8_2462);
and ( n13171 , RI19ab8b38_2390 , n27683 );
or ( n42662 , n13170 , n13171 );
not ( n13172 , RI1754c610_2);
and ( n13173 , n13172 , n42662 );
and ( n13174 , C0 , RI1754c610_2);
or ( n42663 , n13173 , n13174 );
buf ( n42664 , n42663 );
and ( n42665 , RI1754bcb0_22 , n34844 );
and ( n42666 , RI1754bcb0_22 , n34847 );
and ( n42667 , RI1754bcb0_22 , n34850 );
and ( n42668 , RI1754bcb0_22 , n34852 );
and ( n42669 , RI1754bcb0_22 , n34854 );
or ( n42670 , n42665 , n42666 , n42667 , n42668 , n42669 , C0 , C0 , C0 );
not ( n13175 , n34859 );
and ( n13176 , n13175 , n42670 );
and ( n13177 , RI1754bcb0_22 , n34859 );
or ( n42671 , n13176 , n13177 );
not ( n13178 , RI19a22f70_2797);
and ( n13179 , n13178 , n42671 );
and ( n13180 , C0 , RI19a22f70_2797);
or ( n42672 , n13179 , n13180 );
not ( n13181 , n27683 );
and ( n13182 , n13181 , RI19a9cc08_2592);
and ( n13183 , n42672 , n27683 );
or ( n42673 , n13182 , n13183 );
not ( n13184 , RI1754c610_2);
and ( n13185 , n13184 , n42673 );
and ( n13186 , C0 , RI1754c610_2);
or ( n42674 , n13185 , n13186 );
buf ( n42675 , n42674 );
buf ( n42676 , RI1749aa88_982);
xor ( n42677 , n36243 , n41370 );
xor ( n42678 , n42677 , n37898 );
xor ( n42679 , n31478 , n41287 );
xor ( n42680 , n42679 , n39935 );
not ( n42681 , n42680 );
xor ( n42682 , n37941 , n40210 );
xor ( n42683 , n42682 , n39989 );
and ( n42684 , n42681 , n42683 );
xor ( n42685 , n42678 , n42684 );
not ( n13187 , n29614 );
and ( n13188 , n13187 , RI173ec050_1605);
and ( n13189 , n42685 , n29614 );
or ( n42686 , n13188 , n13189 );
not ( n13190 , RI1754c610_2);
and ( n13191 , n13190 , n42686 );
and ( n13192 , C0 , RI1754c610_2);
or ( n42687 , n13191 , n13192 );
buf ( n42688 , n42687 );
buf ( n42689 , RI174809d0_1109);
not ( n42690 , n36253 );
xor ( n42691 , n35803 , n37331 );
xor ( n42692 , n42691 , n37129 );
and ( n42693 , n42690 , n42692 );
xor ( n42694 , n36228 , n42693 );
not ( n13193 , n29614 );
and ( n13194 , n13193 , RI1745c850_1285);
and ( n13195 , n42694 , n29614 );
or ( n42695 , n13194 , n13195 );
not ( n13196 , RI1754c610_2);
and ( n13197 , n13196 , n42695 );
and ( n13198 , C0 , RI1754c610_2);
or ( n42696 , n13197 , n13198 );
buf ( n42697 , n42696 );
not ( n13199 , n27683 );
and ( n13200 , n13199 , RI19a85c10_2754);
and ( n13201 , RI19a23678_2793 , n27683 );
or ( n42698 , n13200 , n13201 );
not ( n13202 , RI1754c610_2);
and ( n13203 , n13202 , n42698 );
and ( n13204 , C0 , RI1754c610_2);
or ( n42699 , n13203 , n13204 );
buf ( n42700 , n42699 );
xor ( n42701 , n38346 , n38872 );
xor ( n42702 , n42701 , n38886 );
not ( n42703 , n37049 );
and ( n42704 , n42703 , n37054 );
xor ( n42705 , n42702 , n42704 );
not ( n13205 , n29614 );
and ( n13206 , n13205 , RI1733aae0_2155);
and ( n13207 , n42705 , n29614 );
or ( n42706 , n13206 , n13207 );
not ( n13208 , RI1754c610_2);
and ( n13209 , n13208 , n42706 );
and ( n13210 , C0 , RI1754c610_2);
or ( n42707 , n13209 , n13210 );
buf ( n42708 , n42707 );
buf ( n42709 , RI17511b28_711);
not ( n13211 , n27683 );
and ( n13212 , n13211 , RI19a932c0_2660);
and ( n13213 , RI19a9d658_2588 , n27683 );
or ( n42710 , n13212 , n13213 );
not ( n13214 , RI1754c610_2);
and ( n13215 , n13214 , n42710 );
and ( n13216 , C0 , RI1754c610_2);
or ( n42711 , n13215 , n13216 );
buf ( n42712 , n42711 );
buf ( n42713 , RI174b8650_837);
xor ( n42714 , n37295 , n40190 );
xor ( n42715 , n42714 , n40210 );
not ( n42716 , n42715 );
and ( n42717 , n42716 , n35855 );
xor ( n42718 , n31926 , n42717 );
not ( n13217 , n29614 );
and ( n13218 , n13217 , RI173be138_1829);
and ( n13219 , n42718 , n29614 );
or ( n42719 , n13218 , n13219 );
not ( n13220 , RI1754c610_2);
and ( n13221 , n13220 , n42719 );
and ( n13222 , C0 , RI1754c610_2);
or ( n42720 , n13221 , n13222 );
buf ( n42721 , n42720 );
xor ( n42722 , n42592 , n38284 );
xor ( n42723 , n42722 , n39856 );
xor ( n42724 , n35817 , n37129 );
xor ( n42725 , n42724 , n37169 );
not ( n42726 , n42725 );
xor ( n42727 , n34488 , n29610 );
xor ( n42728 , n42727 , n31380 );
and ( n42729 , n42726 , n42728 );
xor ( n42730 , n42723 , n42729 );
not ( n13223 , n29614 );
and ( n13224 , n13223 , RI17413308_1414);
and ( n13225 , n42730 , n29614 );
or ( n42731 , n13224 , n13225 );
not ( n13226 , RI1754c610_2);
and ( n13227 , n13226 , n42731 );
and ( n13228 , C0 , RI1754c610_2);
or ( n42732 , n13227 , n13228 );
buf ( n42733 , n42732 );
xor ( n42734 , n35068 , n33223 );
xor ( n42735 , n42734 , n33282 );
xor ( n42736 , n38537 , n35458 );
xor ( n42737 , n42736 , n40692 );
not ( n42738 , n42737 );
xor ( n42739 , n38804 , n39621 );
xor ( n42740 , n42739 , n40855 );
and ( n42741 , n42738 , n42740 );
xor ( n42742 , n42735 , n42741 );
not ( n13229 , n29614 );
and ( n13230 , n13229 , RI173d2628_1730);
and ( n13231 , n42742 , n29614 );
or ( n42743 , n13230 , n13231 );
not ( n13232 , RI1754c610_2);
and ( n13233 , n13232 , n42743 );
and ( n13234 , C0 , RI1754c610_2);
or ( n42744 , n13233 , n13234 );
buf ( n42745 , n42744 );
buf ( n42746 , RI17472768_1178);
buf ( n42747 , RI17476c50_1157);
xor ( n42748 , n37128 , n40237 );
xor ( n42749 , n42748 , n40254 );
xor ( n42750 , n40956 , n36844 );
xor ( n42751 , n42750 , n36874 );
not ( n42752 , n42751 );
xor ( n42753 , n37966 , n41504 );
xor ( n42754 , n42753 , n41690 );
and ( n42755 , n42752 , n42754 );
xor ( n42756 , n42749 , n42755 );
not ( n13235 , n29614 );
and ( n13236 , n13235 , RI175342e0_604);
and ( n13237 , n42756 , n29614 );
or ( n42757 , n13236 , n13237 );
not ( n13238 , RI1754c610_2);
and ( n13239 , n13238 , n42757 );
and ( n13240 , C0 , RI1754c610_2);
or ( n42758 , n13239 , n13240 );
buf ( n42759 , n42758 );
xor ( n42760 , n40580 , n37048 );
xor ( n42761 , n42760 , n36772 );
xor ( n42762 , n32862 , n37203 );
xor ( n42763 , n42762 , n34150 );
not ( n42764 , n42763 );
and ( n42765 , n42764 , n42002 );
xor ( n42766 , n42761 , n42765 );
not ( n13241 , n29614 );
and ( n13242 , n13241 , RI173a2988_1963);
and ( n13243 , n42766 , n29614 );
or ( n42767 , n13242 , n13243 );
not ( n13244 , RI1754c610_2);
and ( n13245 , n13244 , n42767 );
and ( n13246 , C0 , RI1754c610_2);
or ( n42768 , n13245 , n13246 );
buf ( n42769 , n42768 );
not ( n13247 , n27683 );
and ( n13248 , n13247 , RI19abe808_2345);
and ( n13249 , RI19ac7700_2274 , n27683 );
or ( n42770 , n13248 , n13249 );
not ( n13250 , RI1754c610_2);
and ( n13251 , n13250 , n42770 );
and ( n13252 , C0 , RI1754c610_2);
or ( n42771 , n13251 , n13252 );
buf ( n42772 , n42771 );
not ( n13253 , n27683 );
and ( n13254 , n13253 , RI19ab5a00_2411);
and ( n13255 , RI19abef88_2341 , n27683 );
or ( n42773 , n13254 , n13255 );
not ( n13256 , RI1754c610_2);
and ( n13257 , n13256 , n42773 );
and ( n13258 , C0 , RI1754c610_2);
or ( n42774 , n13257 , n13258 );
buf ( n42775 , n42774 );
xor ( n42776 , n34947 , n36802 );
xor ( n42777 , n42776 , n33125 );
not ( n42778 , n41252 );
and ( n42779 , n42778 , n41254 );
xor ( n42780 , n42777 , n42779 );
not ( n13259 , n29614 );
and ( n13260 , n13259 , RI17490d08_1030);
and ( n13261 , n42780 , n29614 );
or ( n42781 , n13260 , n13261 );
not ( n13262 , RI1754c610_2);
and ( n13263 , n13262 , n42781 );
and ( n13264 , C0 , RI1754c610_2);
or ( n42782 , n13263 , n13264 );
buf ( n42783 , n42782 );
not ( n13265 , n27683 );
and ( n13266 , n13265 , RI19ac7700_2274);
and ( n13267 , RI19a82538_2778 , n27683 );
or ( n42784 , n13266 , n13267 );
not ( n13268 , RI1754c610_2);
and ( n13269 , n13268 , n42784 );
and ( n13270 , C0 , RI1754c610_2);
or ( n42785 , n13269 , n13270 );
buf ( n42786 , n42785 );
xor ( n42787 , n39146 , n28468 );
xor ( n42788 , n42787 , n36530 );
xor ( n42789 , n38816 , n39621 );
xor ( n42790 , n42789 , n40855 );
not ( n42791 , n42790 );
xor ( n42792 , n39673 , n33617 );
xor ( n42793 , n42792 , n39525 );
and ( n42794 , n42791 , n42793 );
xor ( n42795 , n42788 , n42794 );
not ( n13271 , n29614 );
and ( n13272 , n13271 , RI173f18e8_1578);
and ( n13273 , n42795 , n29614 );
or ( n42796 , n13272 , n13273 );
not ( n13274 , RI1754c610_2);
and ( n13275 , n13274 , n42796 );
and ( n13276 , C0 , RI1754c610_2);
or ( n42797 , n13275 , n13276 );
buf ( n42798 , n42797 );
not ( n13277 , n27683 );
and ( n13278 , n13277 , RI19a97460_2631);
and ( n13279 , RI19aa0f10_2561 , n27683 );
or ( n42799 , n13278 , n13279 );
not ( n13280 , RI1754c610_2);
and ( n13281 , n13280 , n42799 );
and ( n13282 , C0 , RI1754c610_2);
or ( n42800 , n13281 , n13282 );
buf ( n42801 , n42800 );
xor ( n42802 , n37856 , n35128 );
xor ( n42803 , n42802 , n36917 );
not ( n42804 , n41559 );
and ( n42805 , n42804 , n41561 );
xor ( n42806 , n42803 , n42805 );
not ( n13283 , n29614 );
and ( n13284 , n13283 , RI1738b6c0_2076);
and ( n13285 , n42806 , n29614 );
or ( n42807 , n13284 , n13285 );
not ( n13286 , RI1754c610_2);
and ( n13287 , n13286 , n42807 );
and ( n13288 , C0 , RI1754c610_2);
or ( n42808 , n13287 , n13288 );
buf ( n42809 , n42808 );
not ( n42810 , n36288 );
and ( n42811 , n42810 , n36293 );
xor ( n42812 , n36103 , n42811 );
not ( n13289 , n29614 );
and ( n13290 , n13289 , RI1746d560_1203);
and ( n13291 , n42812 , n29614 );
or ( n42813 , n13290 , n13291 );
not ( n13292 , RI1754c610_2);
and ( n13293 , n13292 , n42813 );
and ( n13294 , C0 , RI1754c610_2);
or ( n42814 , n13293 , n13294 );
buf ( n42815 , n42814 );
not ( n13295 , n27683 );
and ( n13296 , n13295 , RI19ac2cf0_2308);
and ( n13297 , RI19acbc60_2241 , n27683 );
or ( n42816 , n13296 , n13297 );
not ( n13298 , RI1754c610_2);
and ( n13299 , n13298 , n42816 );
and ( n13300 , C0 , RI1754c610_2);
or ( n42817 , n13299 , n13300 );
buf ( n42818 , n42817 );
xor ( n42819 , n37836 , n33697 );
xor ( n42820 , n42819 , n35128 );
xor ( n42821 , n31860 , n36401 );
xor ( n42822 , n42821 , n33453 );
not ( n42823 , n42822 );
xor ( n42824 , n34141 , n33069 );
xor ( n42825 , n42824 , n42264 );
and ( n42826 , n42823 , n42825 );
xor ( n42827 , n42820 , n42826 );
not ( n13301 , n29614 );
and ( n13302 , n13301 , RI17463150_1253);
and ( n13303 , n42827 , n29614 );
or ( n42828 , n13302 , n13303 );
not ( n13304 , RI1754c610_2);
and ( n13305 , n13304 , n42828 );
and ( n13306 , C0 , RI1754c610_2);
or ( n42829 , n13305 , n13306 );
buf ( n42830 , n42829 );
xor ( n42831 , n41880 , n38085 );
xor ( n42832 , n42831 , n38115 );
xor ( n42833 , n32402 , n41316 );
xor ( n42834 , n42833 , n35622 );
not ( n42835 , n42834 );
xor ( n42836 , n34805 , n41478 );
xor ( n42837 , n42836 , n41146 );
and ( n42838 , n42835 , n42837 );
xor ( n42839 , n42832 , n42838 );
not ( n13307 , n29614 );
and ( n13308 , n13307 , RI173aeb20_1904);
and ( n13309 , n42839 , n29614 );
or ( n42840 , n13308 , n13309 );
not ( n13310 , RI1754c610_2);
and ( n13311 , n13310 , n42840 );
and ( n13312 , C0 , RI1754c610_2);
or ( n42841 , n13311 , n13312 );
buf ( n42842 , n42841 );
xor ( n42843 , n35117 , n40283 );
xor ( n42844 , n42843 , n32560 );
xor ( n42845 , n39281 , n38445 );
xor ( n42846 , n42845 , n37549 );
not ( n42847 , n42846 );
xor ( n42848 , n39639 , n35216 );
xor ( n42849 , n42848 , n41241 );
and ( n42850 , n42847 , n42849 );
xor ( n42851 , n42844 , n42850 );
not ( n13313 , n29614 );
and ( n13314 , n13313 , RI175217d0_662);
and ( n13315 , n42851 , n29614 );
or ( n42852 , n13314 , n13315 );
not ( n13316 , RI1754c610_2);
and ( n13317 , n13316 , n42852 );
and ( n13318 , C0 , RI1754c610_2);
or ( n42853 , n13317 , n13318 );
buf ( n42854 , n42853 );
not ( n13319 , n27683 );
and ( n13320 , n13319 , RI19ac90c8_2262);
and ( n13321 , RI19a841d0_2765 , n27683 );
or ( n42855 , n13320 , n13321 );
not ( n13322 , RI1754c610_2);
and ( n13323 , n13322 , n42855 );
and ( n13324 , C0 , RI1754c610_2);
or ( n42856 , n13323 , n13324 );
buf ( n42857 , n42856 );
not ( n13325 , n27683 );
and ( n13326 , n13325 , RI19aa5fb0_2523);
and ( n13327 , RI19ab01e0_2453 , n27683 );
or ( n42858 , n13326 , n13327 );
not ( n13328 , RI1754c610_2);
and ( n13329 , n13328 , n42858 );
and ( n13330 , C0 , RI1754c610_2);
or ( n42859 , n13329 , n13330 );
buf ( n42860 , n42859 );
not ( n13331 , n27683 );
and ( n13332 , n13331 , RI19a89bd0_2726);
and ( n13333 , RI19a93d88_2655 , n27683 );
or ( n42861 , n13332 , n13333 );
not ( n13334 , RI1754c610_2);
and ( n13335 , n13334 , n42861 );
and ( n13336 , C0 , RI1754c610_2);
or ( n42862 , n13335 , n13336 );
buf ( n42863 , n42862 );
not ( n42864 , n42754 );
xor ( n42865 , n37404 , n38267 );
xor ( n42866 , n42865 , n38284 );
and ( n42867 , n42864 , n42866 );
xor ( n42868 , n42751 , n42867 );
not ( n13337 , n29614 );
and ( n13338 , n13337 , RI174adef8_888);
and ( n13339 , n42868 , n29614 );
or ( n42869 , n13338 , n13339 );
not ( n13340 , RI1754c610_2);
and ( n13341 , n13340 , n42869 );
and ( n13342 , C0 , RI1754c610_2);
or ( n42870 , n13341 , n13342 );
buf ( n42871 , n42870 );
xor ( n42872 , n40136 , n38948 );
xor ( n42873 , n42872 , n39039 );
xor ( n42874 , n39405 , n32403 );
xor ( n42875 , n42874 , n32481 );
not ( n42876 , n42875 );
xor ( n42877 , n33446 , n36252 );
xor ( n42878 , n42877 , n40360 );
and ( n42879 , n42876 , n42878 );
xor ( n42880 , n42873 , n42879 );
not ( n13343 , n29614 );
and ( n13344 , n13343 , RI173dc3a8_1682);
and ( n13345 , n42880 , n29614 );
or ( n42881 , n13344 , n13345 );
not ( n13346 , RI1754c610_2);
and ( n13347 , n13346 , n42881 );
and ( n13348 , C0 , RI1754c610_2);
or ( n42882 , n13347 , n13348 );
buf ( n42883 , n42882 );
xor ( n42884 , n37483 , n42188 );
xor ( n42885 , n42884 , n41526 );
not ( n42886 , n42885 );
xor ( n42887 , n41004 , n36998 );
xor ( n42888 , n42887 , n37048 );
and ( n42889 , n42886 , n42888 );
xor ( n42890 , n42579 , n42889 );
not ( n13349 , n29614 );
and ( n13350 , n13349 , RI173e98f0_1617);
and ( n13351 , n42890 , n29614 );
or ( n42891 , n13350 , n13351 );
not ( n13352 , RI1754c610_2);
and ( n13353 , n13352 , n42891 );
and ( n13354 , C0 , RI1754c610_2);
or ( n42892 , n13353 , n13354 );
buf ( n42893 , n42892 );
not ( n13355 , n27683 );
and ( n13356 , n13355 , RI19a9b1c8_2604);
and ( n13357 , RI19aa4a98_2532 , n27683 );
or ( n42894 , n13356 , n13357 );
not ( n13358 , RI1754c610_2);
and ( n13359 , n13358 , n42894 );
and ( n13360 , C0 , RI1754c610_2);
or ( n42895 , n13359 , n13360 );
buf ( n42896 , n42895 );
xor ( n42897 , n41058 , n36339 );
xor ( n42898 , n42897 , n36377 );
xor ( n42899 , n37933 , n40210 );
xor ( n42900 , n42899 , n39989 );
not ( n42901 , n42900 );
xor ( n42902 , n28030 , n42344 );
xor ( n42903 , n42902 , n41799 );
and ( n42904 , n42901 , n42903 );
xor ( n42905 , n42898 , n42904 );
not ( n13361 , n29614 );
and ( n13362 , n13361 , RI1738d100_2068);
and ( n13363 , n42905 , n29614 );
or ( n42906 , n13362 , n13363 );
not ( n13364 , RI1754c610_2);
and ( n13365 , n13364 , n42906 );
and ( n13366 , C0 , RI1754c610_2);
or ( n42907 , n13365 , n13366 );
buf ( n42908 , n42907 );
xor ( n42909 , n39782 , n33175 );
xor ( n42910 , n42909 , n34797 );
xor ( n42911 , n41585 , n39065 );
xor ( n42912 , n42911 , n37331 );
not ( n42913 , n42912 );
xor ( n42914 , n34754 , n42619 );
xor ( n42915 , n42914 , n41990 );
and ( n42916 , n42913 , n42915 );
xor ( n42917 , n42910 , n42916 );
not ( n13367 , n29614 );
and ( n13368 , n13367 , RI1739a300_2004);
and ( n13369 , n42917 , n29614 );
or ( n42918 , n13368 , n13369 );
not ( n13370 , RI1754c610_2);
and ( n13371 , n13370 , n42918 );
and ( n13372 , C0 , RI1754c610_2);
or ( n42919 , n13371 , n13372 );
buf ( n42920 , n42919 );
xor ( n42921 , n38527 , n31725 );
xor ( n42922 , n42921 , n42309 );
not ( n42923 , n42922 );
xor ( n42924 , n31505 , n41287 );
xor ( n42925 , n42924 , n39935 );
and ( n42926 , n42923 , n42925 );
xor ( n42927 , n41773 , n42926 );
not ( n13373 , n29614 );
and ( n13374 , n13373 , RI17516880_696);
and ( n13375 , n42927 , n29614 );
or ( n42928 , n13374 , n13375 );
not ( n13376 , RI1754c610_2);
and ( n13377 , n13376 , n42928 );
and ( n13378 , C0 , RI1754c610_2);
or ( n42929 , n13377 , n13378 );
buf ( n42930 , n42929 );
xor ( n42931 , n40376 , n42554 );
xor ( n42932 , n42931 , n34725 );
not ( n42933 , n29236 );
and ( n42934 , n42933 , n34971 );
xor ( n42935 , n29212 , n42934 );
not ( n42936 , n29274 );
and ( n42937 , n42936 , n34981 );
xor ( n42938 , n29271 , n42937 );
xor ( n42939 , n42935 , n42938 );
xor ( n42940 , n42939 , n29165 );
not ( n42941 , n29348 );
and ( n42942 , n42941 , n34995 );
xor ( n42943 , n29333 , n42942 );
xor ( n42944 , n42940 , n42943 );
xor ( n42945 , n42944 , n42318 );
xor ( n42946 , n35008 , n42945 );
xor ( n42947 , n42946 , n34497 );
not ( n42948 , n42947 );
xor ( n42949 , n38358 , n33880 );
xor ( n42950 , n42949 , n33935 );
and ( n42951 , n42948 , n42950 );
xor ( n42952 , n42932 , n42951 );
not ( n13379 , n29614 );
and ( n13380 , n13379 , RI173f1c30_1577);
and ( n13381 , n42952 , n29614 );
or ( n42953 , n13380 , n13381 );
not ( n13382 , RI1754c610_2);
and ( n13383 , n13382 , n42953 );
and ( n13384 , C0 , RI1754c610_2);
or ( n42954 , n13383 , n13384 );
buf ( n42955 , n42954 );
buf ( n42956 , RI1748b128_1058);
buf ( n42957 , RI174d0cc8_761);
buf ( n42958 , RI174765c0_1159);
xor ( n42959 , n32684 , n36209 );
xor ( n42960 , n42959 , n40412 );
not ( n42961 , n35515 );
and ( n42962 , n42961 , n35595 );
xor ( n42963 , n42960 , n42962 );
not ( n13385 , n29614 );
and ( n13386 , n13385 , RI173da968_1690);
and ( n13387 , n42963 , n29614 );
or ( n42964 , n13386 , n13387 );
not ( n13388 , RI1754c610_2);
and ( n13389 , n13388 , n42964 );
and ( n13390 , C0 , RI1754c610_2);
or ( n42965 , n13389 , n13390 );
buf ( n42966 , n42965 );
xor ( n42967 , n29506 , n40051 );
xor ( n42968 , n42967 , n37074 );
xor ( n42969 , n36861 , n41198 );
xor ( n42970 , n42969 , n41215 );
not ( n42971 , n42970 );
xor ( n42972 , n32385 , n41316 );
xor ( n42973 , n42972 , n35622 );
and ( n42974 , n42971 , n42973 );
xor ( n42975 , n42968 , n42974 );
not ( n13391 , n29614 );
and ( n13392 , n13391 , RI1744cef0_1361);
and ( n13393 , n42975 , n29614 );
or ( n42976 , n13392 , n13393 );
not ( n13394 , RI1754c610_2);
and ( n13395 , n13394 , n42976 );
and ( n13396 , C0 , RI1754c610_2);
or ( n42977 , n13395 , n13396 );
buf ( n42978 , n42977 );
xor ( n42979 , n38006 , n41690 );
xor ( n42980 , n42979 , n39506 );
xor ( n42981 , n34424 , n40009 );
xor ( n42982 , n42981 , n38085 );
not ( n42983 , n42982 );
xor ( n42984 , n40252 , n35760 );
xor ( n42985 , n42984 , n39333 );
and ( n42986 , n42983 , n42985 );
xor ( n42987 , n42980 , n42986 );
not ( n13397 , n29614 );
and ( n13398 , n13397 , RI1747d208_1126);
and ( n13399 , n42987 , n29614 );
or ( n42988 , n13398 , n13399 );
not ( n13400 , RI1754c610_2);
and ( n13401 , n13400 , n42988 );
and ( n13402 , C0 , RI1754c610_2);
or ( n42989 , n13401 , n13402 );
buf ( n42990 , n42989 );
xor ( n42991 , n33990 , n34221 );
xor ( n42992 , n42991 , n34251 );
xor ( n42993 , n37389 , n38267 );
xor ( n42994 , n42993 , n38284 );
not ( n42995 , n42994 );
xor ( n42996 , n37085 , n37716 );
xor ( n42997 , n42996 , n37744 );
and ( n42998 , n42995 , n42997 );
xor ( n42999 , n42992 , n42998 );
not ( n13403 , n29614 );
and ( n13404 , n13403 , RI1749ffd8_956);
and ( n13405 , n42999 , n29614 );
or ( n43000 , n13404 , n13405 );
not ( n13406 , RI1754c610_2);
and ( n13407 , n13406 , n43000 );
and ( n13408 , C0 , RI1754c610_2);
or ( n43001 , n13407 , n13408 );
buf ( n43002 , n43001 );
xor ( n43003 , n38166 , n35494 );
xor ( n43004 , n43003 , n35514 );
not ( n43005 , n42357 );
and ( n43006 , n43005 , n42359 );
xor ( n43007 , n43004 , n43006 );
not ( n13409 , n29614 );
and ( n13410 , n13409 , RI1744e930_1353);
and ( n13411 , n43007 , n29614 );
or ( n43008 , n13410 , n13411 );
not ( n13412 , RI1754c610_2);
and ( n13413 , n13412 , n43008 );
and ( n13414 , C0 , RI1754c610_2);
or ( n43009 , n13413 , n13414 );
buf ( n43010 , n43009 );
xor ( n43011 , n29609 , n40051 );
xor ( n43012 , n43011 , n37074 );
not ( n43013 , n43012 );
xor ( n43014 , n37275 , n34127 );
xor ( n43015 , n43014 , n40190 );
and ( n43016 , n43013 , n43015 );
xor ( n43017 , n40778 , n43016 );
not ( n13415 , n29614 );
and ( n13416 , n13415 , RI173f1f78_1576);
and ( n13417 , n43017 , n29614 );
or ( n43018 , n13416 , n13417 );
not ( n13418 , RI1754c610_2);
and ( n13419 , n13418 , n43018 );
and ( n13420 , C0 , RI1754c610_2);
or ( n43019 , n13419 , n13420 );
buf ( n43020 , n43019 );
xor ( n43021 , n32694 , n36209 );
xor ( n43022 , n43021 , n40412 );
not ( n43023 , n34559 );
and ( n43024 , n43023 , n36830 );
xor ( n43025 , n34556 , n43024 );
xor ( n43026 , n43025 , n34572 );
xor ( n43027 , n43026 , n34622 );
not ( n43028 , n43027 );
and ( n43029 , n43028 , n42320 );
xor ( n43030 , n43022 , n43029 );
not ( n13421 , n29614 );
and ( n13422 , n13421 , RI174cf828_765);
and ( n13423 , n43030 , n29614 );
or ( n43031 , n13422 , n13423 );
not ( n13424 , RI1754c610_2);
and ( n13425 , n13424 , n43031 );
and ( n13426 , C0 , RI1754c610_2);
or ( n43032 , n13425 , n13426 );
buf ( n43033 , n43032 );
xor ( n43034 , n41235 , n38634 );
xor ( n43035 , n43034 , n38648 );
xor ( n43036 , n39599 , n31621 );
xor ( n43037 , n43036 , n35272 );
not ( n43038 , n43037 );
xor ( n43039 , n42553 , n37421 );
xor ( n43040 , n43039 , n42605 );
and ( n43041 , n43038 , n43040 );
xor ( n43042 , n43035 , n43041 );
not ( n13427 , n29614 );
and ( n13428 , n13427 , RI1745df48_1278);
and ( n13429 , n43042 , n29614 );
or ( n43043 , n13428 , n13429 );
not ( n13430 , RI1754c610_2);
and ( n13431 , n13430 , n43043 );
and ( n13432 , C0 , RI1754c610_2);
or ( n43044 , n13431 , n13432 );
buf ( n43045 , n43044 );
xor ( n43046 , n37711 , n40463 );
xor ( n43047 , n43046 , n41772 );
not ( n43048 , n43047 );
xor ( n43049 , n38444 , n40585 );
xor ( n43050 , n43049 , n34918 );
and ( n43051 , n43048 , n43050 );
xor ( n43052 , n42728 , n43051 );
not ( n13433 , n29614 );
and ( n13434 , n13433 , RI1745f2f8_1272);
and ( n13435 , n43052 , n29614 );
or ( n43053 , n13434 , n13435 );
not ( n13436 , RI1754c610_2);
and ( n13437 , n13436 , n43053 );
and ( n13438 , C0 , RI1754c610_2);
or ( n43054 , n13437 , n13438 );
buf ( n43055 , n43054 );
xor ( n43056 , n40657 , n39282 );
xor ( n43057 , n43056 , n37676 );
xor ( n43058 , n28110 , n42344 );
xor ( n43059 , n43058 , n41799 );
not ( n43060 , n43059 );
xor ( n43061 , n32933 , n41659 );
xor ( n43062 , n43061 , n37800 );
and ( n43063 , n43060 , n43062 );
xor ( n43064 , n43057 , n43063 );
not ( n13439 , n29614 );
and ( n13440 , n13439 , RI1748dbd0_1045);
and ( n13441 , n43064 , n29614 );
or ( n43065 , n13440 , n13441 );
not ( n13442 , RI1754c610_2);
and ( n13443 , n13442 , n43065 );
and ( n13444 , C0 , RI1754c610_2);
or ( n43066 , n13443 , n13444 );
buf ( n43067 , n43066 );
buf ( n43068 , RI1747dbe0_1123);
buf ( n43069 , RI1746a428_1218);
xor ( n43070 , n41469 , n39686 );
xor ( n43071 , n43070 , n34087 );
not ( n43072 , n42844 );
and ( n43073 , n43072 , n42846 );
xor ( n43074 , n43071 , n43073 );
not ( n13445 , n29614 );
and ( n13446 , n13445 , RI1750a490_734);
and ( n13447 , n43074 , n29614 );
or ( n43075 , n13446 , n13447 );
not ( n13448 , RI1754c610_2);
and ( n13449 , n13448 , n43075 );
and ( n13450 , C0 , RI1754c610_2);
or ( n43076 , n13449 , n13450 );
buf ( n43077 , n43076 );
xor ( n43078 , n34882 , n36772 );
xor ( n43079 , n43078 , n36802 );
not ( n43080 , n41337 );
and ( n43081 , n43080 , n41339 );
xor ( n43082 , n43079 , n43081 );
not ( n13451 , n29614 );
and ( n13452 , n13451 , RI17414370_1409);
and ( n13453 , n43082 , n29614 );
or ( n43083 , n13452 , n13453 );
not ( n13454 , RI1754c610_2);
and ( n13455 , n13454 , n43083 );
and ( n13456 , C0 , RI1754c610_2);
or ( n43084 , n13455 , n13456 );
buf ( n43085 , n43084 );
not ( n43086 , n27689 );
and ( n43087 , RI19a250b8_2781 , n43086 );
or ( n43088 , n27689 , n27683 );
not ( n13457 , n43088 );
and ( n13458 , n13457 , RI19a24ed8_2782);
and ( n13459 , n43087 , n43088 );
or ( n43089 , n13458 , n13459 );
not ( n13460 , RI1754c610_2);
and ( n13461 , n13460 , n43089 );
and ( n13462 , C0 , RI1754c610_2);
or ( n43090 , n13461 , n13462 );
buf ( n43091 , n43090 );
buf ( n43092 , RI174cb520_778);
xor ( n43093 , n40148 , n38948 );
xor ( n43094 , n43093 , n39039 );
xor ( n43095 , n38850 , n41125 );
xor ( n43096 , n43095 , n31506 );
not ( n43097 , n43096 );
xor ( n43098 , n40038 , n38574 );
xor ( n43099 , n43098 , n38594 );
and ( n43100 , n43097 , n43099 );
xor ( n43101 , n43094 , n43100 );
not ( n13463 , n29614 );
and ( n13464 , n13463 , RI173c3340_1804);
and ( n13465 , n43101 , n29614 );
or ( n43102 , n13464 , n13465 );
not ( n13466 , RI1754c610_2);
and ( n13467 , n13466 , n43102 );
and ( n13468 , C0 , RI1754c610_2);
or ( n43103 , n13467 , n13468 );
buf ( n43104 , n43103 );
buf ( n43105 , RI1748ec38_1040);
buf ( n43106 , RI1747be58_1132);
not ( n13469 , n27683 );
and ( n13470 , n13469 , RI19ac52e8_2290);
and ( n13471 , RI19acdf10_2225 , n27683 );
or ( n43107 , n13470 , n13471 );
not ( n13472 , RI1754c610_2);
and ( n13473 , n13472 , n43107 );
and ( n13474 , C0 , RI1754c610_2);
or ( n43108 , n13473 , n13474 );
buf ( n43109 , n43108 );
xor ( n43110 , n34631 , n34150 );
xor ( n43111 , n43110 , n34190 );
xor ( n43112 , n40473 , n38933 );
xor ( n43113 , n43112 , n41430 );
not ( n43114 , n43113 );
and ( n43115 , n43114 , n42532 );
xor ( n43116 , n43111 , n43115 );
not ( n13475 , n29614 );
and ( n13476 , n13475 , RI174af5f0_881);
and ( n13477 , n43116 , n29614 );
or ( n43117 , n13476 , n13477 );
not ( n13478 , RI1754c610_2);
and ( n13479 , n13478 , n43117 );
and ( n13480 , C0 , RI1754c610_2);
or ( n43118 , n13479 , n13480 );
buf ( n43119 , n43118 );
not ( n43120 , n42100 );
xor ( n43121 , n38036 , n41690 );
xor ( n43122 , n43121 , n39506 );
and ( n43123 , n43120 , n43122 );
xor ( n43124 , n42097 , n43123 );
not ( n13481 , n29614 );
and ( n13482 , n13481 , RI1746c4f8_1208);
and ( n13483 , n43124 , n29614 );
or ( n43125 , n13482 , n13483 );
not ( n13484 , RI1754c610_2);
and ( n13485 , n13484 , n43125 );
and ( n13486 , C0 , RI1754c610_2);
or ( n43126 , n13485 , n13486 );
buf ( n43127 , n43126 );
not ( n13487 , n27683 );
and ( n13488 , n13487 , RI19aca4f0_2253);
and ( n13489 , RI19a859b8_2755 , n27683 );
or ( n43128 , n13488 , n13489 );
not ( n13490 , RI1754c610_2);
and ( n13491 , n13490 , n43128 );
and ( n13492 , C0 , RI1754c610_2);
or ( n43129 , n13491 , n13492 );
buf ( n43130 , n43129 );
not ( n13493 , n27683 );
and ( n13494 , n13493 , RI19ac4dc0_2293);
and ( n13495 , RI19acda60_2227 , n27683 );
or ( n43131 , n13494 , n13495 );
not ( n13496 , RI1754c610_2);
and ( n13497 , n13496 , n43131 );
and ( n13498 , C0 , RI1754c610_2);
or ( n43132 , n13497 , n13498 );
buf ( n43133 , n43132 );
not ( n13499 , n27683 );
and ( n13500 , n13499 , RI19ab9a38_2383);
and ( n13501 , RI19ac25e8_2311 , n27683 );
or ( n43134 , n13500 , n13501 );
not ( n13502 , RI1754c610_2);
and ( n13503 , n13502 , n43134 );
and ( n13504 , C0 , RI1754c610_2);
or ( n43135 , n13503 , n13504 );
buf ( n43136 , n43135 );
xor ( n43137 , n27873 , n42344 );
xor ( n43138 , n43137 , n41799 );
not ( n43139 , n43138 );
xor ( n43140 , n38182 , n32220 );
xor ( n43141 , n43140 , n32309 );
and ( n43142 , n43139 , n43141 );
xor ( n43143 , n38821 , n43142 );
not ( n13505 , n29614 );
and ( n13506 , n13505 , RI174b8308_838);
and ( n13507 , n43143 , n29614 );
or ( n43144 , n13506 , n13507 );
not ( n13508 , RI1754c610_2);
and ( n13509 , n13508 , n43144 );
and ( n13510 , C0 , RI1754c610_2);
or ( n43145 , n13509 , n13510 );
buf ( n43146 , n43145 );
xor ( n43147 , n40756 , n33778 );
xor ( n43148 , n43147 , n38793 );
xor ( n43149 , n33799 , n39414 );
xor ( n43150 , n43149 , n37186 );
not ( n43151 , n43150 );
xor ( n43152 , n32906 , n38553 );
xor ( n43153 , n43152 , n41659 );
and ( n43154 , n43151 , n43153 );
xor ( n43155 , n43148 , n43154 );
not ( n13511 , n29614 );
and ( n13512 , n13511 , RI17345238_2104);
and ( n13513 , n43155 , n29614 );
or ( n43156 , n13512 , n13513 );
not ( n13514 , RI1754c610_2);
and ( n13515 , n13514 , n43156 );
and ( n13516 , C0 , RI1754c610_2);
or ( n43157 , n13515 , n13516 );
buf ( n43158 , n43157 );
xor ( n43159 , n37366 , n33505 );
xor ( n43160 , n43159 , n39635 );
xor ( n43161 , n39562 , n38401 );
xor ( n43162 , n43161 , n41068 );
not ( n43163 , n43162 );
xor ( n43164 , n40153 , n39039 );
xor ( n43165 , n43164 , n39065 );
and ( n43166 , n43163 , n43165 );
xor ( n43167 , n43160 , n43166 );
not ( n13517 , n29614 );
and ( n13518 , n13517 , RI17502420_753);
and ( n13519 , n43167 , n29614 );
or ( n43168 , n13518 , n13519 );
not ( n13520 , RI1754c610_2);
and ( n13521 , n13520 , n43168 );
and ( n13522 , C0 , RI1754c610_2);
or ( n43169 , n13521 , n13522 );
buf ( n43170 , n43169 );
not ( n13523 , n27683 );
and ( n13524 , n13523 , RI19a8af08_2718);
and ( n13525 , RI19a952a0_2646 , n27683 );
or ( n43171 , n13524 , n13525 );
not ( n13526 , RI1754c610_2);
and ( n13527 , n13526 , n43171 );
and ( n13528 , C0 , RI1754c610_2);
or ( n43172 , n13527 , n13528 );
buf ( n43173 , n43172 );
xor ( n43174 , n31781 , n34644 );
xor ( n43175 , n43174 , n36401 );
xor ( n43176 , n40184 , n33991 );
xor ( n43177 , n43176 , n34041 );
not ( n43178 , n43177 );
xor ( n43179 , n33326 , n38991 );
xor ( n43180 , n43179 , n39005 );
and ( n43181 , n43178 , n43180 );
xor ( n43182 , n43175 , n43181 );
not ( n13529 , n29614 );
and ( n13530 , n13529 , RI174c3e88_801);
and ( n13531 , n43182 , n29614 );
or ( n43183 , n13530 , n13531 );
not ( n13532 , RI1754c610_2);
and ( n13533 , n13532 , n43183 );
and ( n13534 , C0 , RI1754c610_2);
or ( n43184 , n13533 , n13534 );
buf ( n43185 , n43184 );
not ( n43186 , n40587 );
xor ( n43187 , n36981 , n41818 );
xor ( n43188 , n43187 , n40662 );
and ( n43189 , n43186 , n43188 );
xor ( n43190 , n40565 , n43189 );
not ( n13535 , n29614 );
and ( n13536 , n13535 , RI1746b7d8_1212);
and ( n13537 , n43190 , n29614 );
or ( n43191 , n13536 , n13537 );
not ( n13538 , RI1754c610_2);
and ( n13539 , n13538 , n43191 );
and ( n13540 , C0 , RI1754c610_2);
or ( n43192 , n13539 , n13540 );
buf ( n43193 , n43192 );
xor ( n43194 , n31435 , n41287 );
xor ( n43195 , n43194 , n39935 );
xor ( n43196 , n33366 , n39005 );
xor ( n43197 , n43196 , n39543 );
not ( n43198 , n43197 );
xor ( n43199 , n38715 , n38817 );
xor ( n43200 , n43199 , n40034 );
and ( n43201 , n43198 , n43200 );
xor ( n43202 , n43195 , n43201 );
not ( n13541 , n29614 );
and ( n13542 , n13541 , RI173967f0_2022);
and ( n13543 , n43202 , n29614 );
or ( n43203 , n13542 , n13543 );
not ( n13544 , RI1754c610_2);
and ( n13545 , n13544 , n43203 );
and ( n13546 , C0 , RI1754c610_2);
or ( n43204 , n13545 , n13546 );
buf ( n43205 , n43204 );
xor ( n43206 , n34504 , n31380 );
xor ( n43207 , n43206 , n36463 );
xor ( n43208 , n40042 , n38574 );
xor ( n43209 , n43208 , n38594 );
not ( n43210 , n43209 );
xor ( n43211 , n31042 , n41622 );
xor ( n43212 , n43211 , n38512 );
and ( n43213 , n43210 , n43212 );
xor ( n43214 , n43207 , n43213 );
not ( n13547 , n29614 );
and ( n13548 , n13547 , RI174741a8_1170);
and ( n13549 , n43214 , n29614 );
or ( n43215 , n13548 , n13549 );
not ( n13550 , RI1754c610_2);
and ( n13551 , n13550 , n43215 );
and ( n13552 , C0 , RI1754c610_2);
or ( n43216 , n13551 , n13552 );
buf ( n43217 , n43216 );
xor ( n43218 , n35679 , n39543 );
xor ( n43219 , n43218 , n39563 );
not ( n43220 , n38845 );
and ( n43221 , n43220 , n38887 );
xor ( n43222 , n43219 , n43221 );
not ( n13553 , n29614 );
and ( n13554 , n13553 , RI173dd0c8_1678);
and ( n13555 , n43222 , n29614 );
or ( n43223 , n13554 , n13555 );
not ( n13556 , RI1754c610_2);
and ( n13557 , n13556 , n43223 );
and ( n13558 , C0 , RI1754c610_2);
or ( n43224 , n13557 , n13558 );
buf ( n43225 , n43224 );
buf ( n43226 , RI17499390_989);
xor ( n43227 , n42599 , n38284 );
xor ( n43228 , n43227 , n39856 );
not ( n43229 , n43228 );
and ( n43230 , n43229 , n42058 );
xor ( n43231 , n41131 , n43230 );
not ( n13559 , n29614 );
and ( n13560 , n13559 , RI174796f8_1144);
and ( n13561 , n43231 , n29614 );
or ( n43232 , n13560 , n13561 );
not ( n13562 , RI1754c610_2);
and ( n13563 , n13562 , n43232 );
and ( n13564 , C0 , RI1754c610_2);
or ( n43233 , n13563 , n13564 );
buf ( n43234 , n43233 );
buf ( n43235 , RI174c05d0_812);
xor ( n43236 , n41385 , n33567 );
xor ( n43237 , n43236 , n33617 );
xor ( n43238 , n41852 , n33282 );
xor ( n43239 , n43238 , n37623 );
not ( n43240 , n43239 );
xor ( n43241 , n32219 , n35986 );
xor ( n43242 , n43241 , n36003 );
and ( n43243 , n43240 , n43242 );
xor ( n43244 , n43237 , n43243 );
not ( n13565 , n29614 );
and ( n13566 , n13565 , RI1748a0c0_1063);
and ( n13567 , n43244 , n29614 );
or ( n43245 , n13566 , n13567 );
not ( n13568 , RI1754c610_2);
and ( n13569 , n13568 , n43245 );
and ( n13570 , C0 , RI1754c610_2);
or ( n43246 , n13569 , n13570 );
buf ( n43247 , n43246 );
xor ( n43248 , n39337 , n29843 );
xor ( n43249 , n43248 , n29981 );
not ( n43250 , n36378 );
and ( n43251 , n43250 , n36383 );
xor ( n43252 , n43249 , n43251 );
not ( n13571 , n29614 );
and ( n13572 , n13571 , RI17478690_1149);
and ( n13573 , n43252 , n29614 );
or ( n43253 , n13572 , n13573 );
not ( n13574 , RI1754c610_2);
and ( n13575 , n13574 , n43253 );
and ( n13576 , C0 , RI1754c610_2);
or ( n43254 , n13575 , n13576 );
buf ( n43255 , n43254 );
buf ( n43256 , RI174aef60_883);
buf ( n43257 , RI174a7fd0_917);
buf ( n43258 , RI174844e0_1091);
buf ( n43259 , RI1750c380_728);
not ( n43260 , n41083 );
and ( n43261 , n43260 , n30936 );
xor ( n43262 , n38126 , n43261 );
not ( n43263 , n41088 );
and ( n43264 , n43263 , n30974 );
xor ( n43265 , n38131 , n43264 );
xor ( n43266 , n43262 , n43265 );
not ( n43267 , n39111 );
and ( n43268 , n43267 , n31003 );
xor ( n43269 , n38137 , n43268 );
xor ( n43270 , n43266 , n43269 );
not ( n43271 , n38121 );
and ( n43272 , n43271 , n31013 );
xor ( n43273 , n38118 , n43272 );
xor ( n43274 , n43270 , n43273 );
not ( n43275 , n41096 );
and ( n43276 , n43275 , n31045 );
xor ( n43277 , n38147 , n43276 );
xor ( n43278 , n43274 , n43277 );
xor ( n43279 , n41621 , n43278 );
xor ( n43280 , n43279 , n31664 );
xor ( n43281 , n42039 , n33648 );
xor ( n43282 , n43281 , n33697 );
not ( n43283 , n43282 );
xor ( n43284 , n37061 , n38594 );
xor ( n43285 , n43284 , n37716 );
and ( n43286 , n43283 , n43285 );
xor ( n43287 , n43280 , n43286 );
not ( n13577 , n29614 );
and ( n13578 , n13577 , RI17336fd0_2173);
and ( n13579 , n43287 , n29614 );
or ( n43288 , n13578 , n13579 );
not ( n13580 , RI1754c610_2);
and ( n13581 , n13580 , n43288 );
and ( n13582 , C0 , RI1754c610_2);
or ( n43289 , n13581 , n13582 );
buf ( n43290 , n43289 );
xor ( n43291 , n31316 , n42049 );
xor ( n43292 , n43291 , n37849 );
xor ( n43293 , n41109 , n41241 );
xor ( n43294 , n43293 , n41287 );
not ( n43295 , n43294 );
xor ( n43296 , n39996 , n40341 );
xor ( n43297 , n43296 , n40091 );
and ( n43298 , n43295 , n43297 );
xor ( n43299 , n43292 , n43298 );
not ( n13583 , n29614 );
and ( n13584 , n13583 , RI174a89a8_914);
and ( n13585 , n43299 , n29614 );
or ( n43300 , n13584 , n13585 );
not ( n13586 , RI1754c610_2);
and ( n13587 , n13586 , n43300 );
and ( n13588 , C0 , RI1754c610_2);
or ( n43301 , n13587 , n13588 );
buf ( n43302 , n43301 );
xor ( n43303 , n36940 , n32620 );
xor ( n43304 , n43303 , n33337 );
not ( n43305 , n40621 );
and ( n43306 , n43305 , n40626 );
xor ( n43307 , n43304 , n43306 );
not ( n13589 , n29614 );
and ( n13590 , n13589 , RI17342100_2119);
and ( n13591 , n43307 , n29614 );
or ( n43308 , n13590 , n13591 );
not ( n13592 , RI1754c610_2);
and ( n13593 , n13592 , n43308 );
and ( n13594 , C0 , RI1754c610_2);
or ( n43309 , n13593 , n13594 );
buf ( n43310 , n43309 );
xor ( n43311 , n34736 , n42619 );
xor ( n43312 , n43311 , n41990 );
xor ( n43313 , n35251 , n39952 );
xor ( n43314 , n43313 , n42945 );
not ( n43315 , n43314 );
xor ( n43316 , n37739 , n41772 );
xor ( n43317 , n43316 , n32663 );
and ( n43318 , n43315 , n43317 );
xor ( n43319 , n43312 , n43318 );
not ( n13595 , n29614 );
and ( n13596 , n13595 , RI173dee50_1669);
and ( n13597 , n43319 , n29614 );
or ( n43320 , n13596 , n13597 );
not ( n13598 , RI1754c610_2);
and ( n13599 , n13598 , n43320 );
and ( n13600 , C0 , RI1754c610_2);
or ( n43321 , n13599 , n13600 );
buf ( n43322 , n43321 );
xor ( n43323 , n38573 , n28816 );
xor ( n43324 , n43323 , n29109 );
not ( n43325 , n43324 );
xor ( n43326 , n31426 , n41287 );
xor ( n43327 , n43326 , n39935 );
and ( n43328 , n43325 , n43327 );
xor ( n43329 , n38038 , n43328 );
not ( n13601 , n29614 );
and ( n13602 , n13601 , RI173bddf0_1830);
and ( n13603 , n43329 , n29614 );
or ( n43330 , n13602 , n13603 );
not ( n13604 , RI1754c610_2);
and ( n13605 , n13604 , n43330 );
and ( n13606 , C0 , RI1754c610_2);
or ( n43331 , n13605 , n13606 );
buf ( n43332 , n43331 );
not ( n13607 , n27683 );
and ( n13608 , n13607 , RI19ab8958_2391);
and ( n13609 , RI19ac12b0_2321 , n27683 );
or ( n43333 , n13608 , n13609 );
not ( n13610 , RI1754c610_2);
and ( n13611 , n13610 , n43333 );
and ( n13612 , C0 , RI1754c610_2);
or ( n43334 , n13611 , n13612 );
buf ( n43335 , n43334 );
xor ( n43336 , n37037 , n40662 );
xor ( n43337 , n43336 , n39208 );
xor ( n43338 , n34250 , n37526 );
xor ( n43339 , n43338 , n41049 );
not ( n43340 , n43339 );
xor ( n43341 , n36112 , n39131 );
xor ( n43342 , n43341 , n39151 );
and ( n43343 , n43340 , n43342 );
xor ( n43344 , n43337 , n43343 );
not ( n13613 , n29614 );
and ( n13614 , n13613 , RI173abd30_1918);
and ( n13615 , n43344 , n29614 );
or ( n43345 , n13614 , n13615 );
not ( n13616 , RI1754c610_2);
and ( n13617 , n13616 , n43345 );
and ( n13618 , C0 , RI1754c610_2);
or ( n43346 , n13617 , n13618 );
buf ( n43347 , n43346 );
and ( n43348 , RI1754be18_19 , n34844 );
and ( n43349 , RI1754be18_19 , n34847 );
and ( n43350 , RI1754be18_19 , n34850 );
and ( n43351 , RI1754be18_19 , n34852 );
and ( n43352 , RI1754be18_19 , n34854 );
or ( n43353 , n43348 , n43349 , n43350 , n43351 , n43352 , C0 , C0 , C0 );
not ( n13619 , n34859 );
and ( n13620 , n13619 , n43353 );
and ( n13621 , RI1754be18_19 , n34859 );
or ( n43354 , n13620 , n13621 );
not ( n13622 , RI19a22f70_2797);
and ( n13623 , n13622 , n43354 );
and ( n13624 , C0 , RI19a22f70_2797);
or ( n43355 , n13623 , n13624 );
not ( n13625 , n27683 );
and ( n13626 , n13625 , RI19a981f8_2625);
and ( n13627 , n43355 , n27683 );
or ( n43356 , n13626 , n13627 );
not ( n13628 , RI1754c610_2);
and ( n13629 , n13628 , n43356 );
and ( n13630 , C0 , RI1754c610_2);
or ( n43357 , n13629 , n13630 );
buf ( n43358 , n43357 );
not ( n13631 , n27683 );
and ( n13632 , n13631 , RI19a8e478_2695);
and ( n13633 , RI19a98630_2623 , n27683 );
or ( n43359 , n13632 , n13633 );
not ( n13634 , RI1754c610_2);
and ( n13635 , n13634 , n43359 );
and ( n13636 , C0 , RI1754c610_2);
or ( n43360 , n13635 , n13636 );
buf ( n43361 , n43360 );
xor ( n43362 , n39554 , n38401 );
xor ( n43363 , n43362 , n41068 );
not ( n43364 , n42932 );
and ( n43365 , n43364 , n42947 );
xor ( n43366 , n43363 , n43365 );
not ( n13637 , n29614 );
and ( n13638 , n13637 , RI173e3338_1648);
and ( n13639 , n43366 , n29614 );
or ( n43367 , n13638 , n13639 );
not ( n13640 , RI1754c610_2);
and ( n13641 , n13640 , n43367 );
and ( n13642 , C0 , RI1754c610_2);
or ( n43368 , n13641 , n13642 );
buf ( n43369 , n43368 );
xor ( n43370 , n42503 , n30461 );
xor ( n43371 , n43370 , n39262 );
xor ( n43372 , n40270 , n37623 );
xor ( n43373 , n43372 , n37651 );
not ( n43374 , n43373 );
and ( n43375 , n43374 , n41372 );
xor ( n43376 , n43371 , n43375 );
not ( n13643 , n29614 );
and ( n13644 , n13643 , RI1749d878_968);
and ( n13645 , n43376 , n29614 );
or ( n43377 , n13644 , n13645 );
not ( n13646 , RI1754c610_2);
and ( n13647 , n13646 , n43377 );
and ( n13648 , C0 , RI1754c610_2);
or ( n43378 , n13647 , n13648 );
buf ( n43379 , n43378 );
xor ( n43380 , n40331 , n37987 );
xor ( n43381 , n43380 , n38037 );
xor ( n43382 , n39026 , n36947 );
xor ( n43383 , n43382 , n39702 );
not ( n43384 , n43383 );
and ( n43385 , n43384 , n41905 );
xor ( n43386 , n43381 , n43385 );
not ( n13649 , n29614 );
and ( n13650 , n13649 , RI173d3d20_1723);
and ( n13651 , n43386 , n29614 );
or ( n43387 , n13650 , n13651 );
not ( n13652 , RI1754c610_2);
and ( n13653 , n13652 , n43387 );
and ( n13654 , C0 , RI1754c610_2);
or ( n43388 , n13653 , n13654 );
buf ( n43389 , n43388 );
not ( n43390 , n41910 );
and ( n43391 , n43390 , n43381 );
xor ( n43392 , n41907 , n43391 );
not ( n13655 , n29614 );
and ( n13656 , n13655 , RI173ff808_1510);
and ( n13657 , n43392 , n29614 );
or ( n43393 , n13656 , n13657 );
not ( n13658 , RI1754c610_2);
and ( n13659 , n13658 , n43393 );
and ( n13660 , C0 , RI1754c610_2);
or ( n43394 , n13659 , n13660 );
buf ( n43395 , n43394 );
xor ( n43396 , n33556 , n40915 );
xor ( n43397 , n43396 , n41740 );
xor ( n43398 , n34621 , n35544 );
xor ( n43399 , n43398 , n35594 );
not ( n43400 , n43399 );
xor ( n43401 , n33347 , n39005 );
xor ( n43402 , n43401 , n39543 );
and ( n43403 , n43400 , n43402 );
xor ( n43404 , n43397 , n43403 );
not ( n13661 , n29614 );
and ( n13662 , n13661 , RI17528e68_639);
and ( n13663 , n43404 , n29614 );
or ( n43405 , n13662 , n13663 );
not ( n13664 , RI1754c610_2);
and ( n13665 , n13664 , n43405 );
and ( n13666 , C0 , RI1754c610_2);
or ( n43406 , n13665 , n13666 );
buf ( n43407 , n43406 );
xor ( n43408 , n40547 , n40966 );
xor ( n43409 , n43408 , n37460 );
xor ( n43410 , n37358 , n33505 );
xor ( n43411 , n43410 , n39635 );
not ( n43412 , n43411 );
xor ( n43413 , n39765 , n33125 );
xor ( n43414 , n43413 , n33175 );
and ( n43415 , n43412 , n43414 );
xor ( n43416 , n43409 , n43415 );
not ( n13667 , n29614 );
and ( n13668 , n13667 , RI173c8f20_1776);
and ( n13669 , n43416 , n29614 );
or ( n43417 , n13668 , n13669 );
not ( n13670 , RI1754c610_2);
and ( n13671 , n13670 , n43417 );
and ( n13672 , C0 , RI1754c610_2);
or ( n43418 , n13671 , n13672 );
buf ( n43419 , n43418 );
xor ( n43420 , n29108 , n34517 );
xor ( n43421 , n43420 , n35911 );
xor ( n43422 , n37239 , n41391 );
xor ( n43423 , n43422 , n39686 );
not ( n43424 , n43423 );
xor ( n43425 , n42609 , n39856 );
xor ( n43426 , n43425 , n39886 );
and ( n43427 , n43424 , n43426 );
xor ( n43428 , n43421 , n43427 );
not ( n13673 , n29614 );
and ( n13674 , n13673 , RI1752eb38_621);
and ( n13675 , n43428 , n29614 );
or ( n43429 , n13674 , n13675 );
not ( n13676 , RI1754c610_2);
and ( n13677 , n13676 , n43429 );
and ( n13678 , C0 , RI1754c610_2);
or ( n43430 , n13677 , n13678 );
buf ( n43431 , n43430 );
not ( n43432 , n39622 );
and ( n43433 , n43432 , n39656 );
xor ( n43434 , n34042 , n43433 );
not ( n13679 , n29614 );
and ( n13680 , n13679 , RI173b71a8_1863);
and ( n13681 , n43434 , n29614 );
or ( n43435 , n13680 , n13681 );
not ( n13682 , RI1754c610_2);
and ( n13683 , n13682 , n43435 );
and ( n13684 , C0 , RI1754c610_2);
or ( n43436 , n13683 , n13684 );
buf ( n43437 , n43436 );
xor ( n43438 , n40485 , n38933 );
xor ( n43439 , n43438 , n41430 );
not ( n43440 , n40267 );
and ( n43441 , n43440 , n40285 );
xor ( n43442 , n43439 , n43441 );
not ( n13685 , n29614 );
and ( n13686 , n13685 , RI174a20a8_946);
and ( n13687 , n43442 , n29614 );
or ( n43443 , n13686 , n13687 );
not ( n13688 , RI1754c610_2);
and ( n13689 , n13688 , n43443 );
and ( n13690 , C0 , RI1754c610_2);
or ( n43444 , n13689 , n13690 );
buf ( n43445 , n43444 );
xor ( n43446 , n39701 , n33337 );
xor ( n43447 , n43446 , n33397 );
xor ( n43448 , n38903 , n42309 );
not ( n43449 , n40933 );
and ( n43450 , n43449 , n40494 );
xor ( n43451 , n38760 , n43450 );
xor ( n43452 , n41163 , n43451 );
not ( n43453 , n40939 );
and ( n43454 , n43453 , n40500 );
xor ( n43455 , n38770 , n43454 );
xor ( n43456 , n43452 , n43455 );
not ( n43457 , n40945 );
and ( n43458 , n43457 , n40506 );
xor ( n43459 , n38780 , n43458 );
xor ( n43460 , n43456 , n43459 );
not ( n43461 , n40696 );
and ( n43462 , n43461 , n40512 );
xor ( n43463 , n38790 , n43462 );
xor ( n43464 , n43460 , n43463 );
xor ( n43465 , n43448 , n43464 );
not ( n43466 , n43465 );
xor ( n43467 , n37507 , n37942 );
xor ( n43468 , n43467 , n34395 );
and ( n43469 , n43466 , n43468 );
xor ( n43470 , n43447 , n43469 );
not ( n13691 , n29614 );
and ( n13692 , n13691 , RI17533890_606);
and ( n13693 , n43470 , n29614 );
or ( n43471 , n13692 , n13693 );
not ( n13694 , RI1754c610_2);
and ( n13695 , n13694 , n43471 );
and ( n13696 , C0 , RI1754c610_2);
or ( n43472 , n13695 , n13696 );
buf ( n43473 , n43472 );
not ( n43474 , n32056 );
and ( n43475 , n43474 , n35179 );
xor ( n43476 , n32053 , n43475 );
not ( n43477 , n32065 );
and ( n43478 , n43477 , n35186 );
xor ( n43479 , n32062 , n43478 );
xor ( n43480 , n43476 , n43479 );
not ( n43481 , n32075 );
and ( n43482 , n43481 , n35194 );
xor ( n43483 , n32072 , n43482 );
xor ( n43484 , n43480 , n43483 );
not ( n43485 , n32095 );
and ( n43486 , n43485 , n35202 );
xor ( n43487 , n32092 , n43486 );
xor ( n43488 , n43484 , n43487 );
not ( n43489 , n32105 );
and ( n43490 , n43489 , n35210 );
xor ( n43491 , n32102 , n43490 );
xor ( n43492 , n43488 , n43491 );
xor ( n43493 , n35184 , n43492 );
xor ( n43494 , n43493 , n38634 );
xor ( n43495 , n37173 , n32481 );
xor ( n43496 , n43495 , n33030 );
not ( n43497 , n43496 );
xor ( n43498 , n37282 , n34127 );
xor ( n43499 , n43498 , n40190 );
and ( n43500 , n43497 , n43499 );
xor ( n43501 , n43494 , n43500 );
not ( n13697 , n29614 );
and ( n13698 , n13697 , RI17449db8_1376);
and ( n13699 , n43501 , n29614 );
or ( n43502 , n13698 , n13699 );
not ( n13700 , RI1754c610_2);
and ( n13701 , n13700 , n43502 );
and ( n13702 , C0 , RI1754c610_2);
or ( n43503 , n13701 , n13702 );
buf ( n43504 , n43503 );
not ( n43505 , n42271 );
xor ( n43506 , n33174 , n37235 );
xor ( n43507 , n43506 , n37255 );
and ( n43508 , n43505 , n43507 );
xor ( n43509 , n42268 , n43508 );
not ( n13703 , n29614 );
and ( n13704 , n13703 , RI1750be58_729);
and ( n13705 , n43509 , n29614 );
or ( n43510 , n13704 , n13705 );
not ( n13706 , RI1754c610_2);
and ( n13707 , n13706 , n43510 );
and ( n13708 , C0 , RI1754c610_2);
or ( n43511 , n13707 , n13708 );
buf ( n43512 , n43511 );
and ( n43513 , RI1754b350_42 , n34844 );
and ( n43514 , RI1754b350_42 , n34847 );
and ( n43515 , RI1754b350_42 , n34850 );
buf ( n43516 , n34852 );
or ( n43517 , n43513 , n43514 , n43515 , n43516 , C0 , C0 , C0 , C0 );
not ( n13709 , n34859 );
and ( n13710 , n13709 , n43517 );
and ( n13711 , RI1754b350_42 , n34859 );
or ( n43518 , n13710 , n13711 );
not ( n13712 , RI19a22f70_2797);
and ( n13713 , n13712 , n43518 );
and ( n13714 , C0 , RI19a22f70_2797);
or ( n43519 , n13713 , n13714 );
not ( n13715 , n27683 );
and ( n13716 , n13715 , RI19abba90_2370);
and ( n13717 , n43519 , n27683 );
or ( n43520 , n13716 , n13717 );
not ( n13718 , RI1754c610_2);
and ( n13719 , n13718 , n43520 );
and ( n13720 , C0 , RI1754c610_2);
or ( n43521 , n13719 , n13720 );
buf ( n43522 , n43521 );
xor ( n43523 , n38494 , n39771 );
xor ( n43524 , n43523 , n39791 );
xor ( n43525 , n39919 , n40890 );
xor ( n43526 , n43525 , n38724 );
not ( n43527 , n43526 );
and ( n43528 , n43527 , n43175 );
xor ( n43529 , n43524 , n43528 );
not ( n13721 , n29614 );
and ( n13722 , n13721 , RI173341e0_2187);
and ( n13723 , n43529 , n29614 );
or ( n43530 , n13722 , n13723 );
not ( n13724 , RI1754c610_2);
and ( n13725 , n13724 , n43530 );
and ( n13726 , C0 , RI1754c610_2);
or ( n43531 , n13725 , n13726 );
buf ( n43532 , n43531 );
xor ( n43533 , n31052 , n41622 );
xor ( n43534 , n43533 , n38512 );
xor ( n43535 , n32570 , n39182 );
xor ( n43536 , n43535 , n38991 );
not ( n43537 , n43536 );
xor ( n43538 , n37396 , n38267 );
xor ( n43539 , n43538 , n38284 );
and ( n43540 , n43537 , n43539 );
xor ( n43541 , n43534 , n43540 );
not ( n13727 , n29614 );
and ( n13728 , n13727 , RI1740a2a8_1458);
and ( n13729 , n43541 , n29614 );
or ( n43542 , n13728 , n13729 );
not ( n13730 , RI1754c610_2);
and ( n13731 , n13730 , n43542 );
and ( n13732 , C0 , RI1754c610_2);
or ( n43543 , n13731 , n13732 );
buf ( n43544 , n43543 );
buf ( n43545 , RI174872d0_1077);
buf ( n43546 , RI174720d8_1180);
buf ( n43547 , RI17507628_743);
not ( n43548 , n41100 );
and ( n43549 , n43548 , n41827 );
xor ( n43550 , n41078 , n43549 );
not ( n13733 , n29614 );
and ( n13734 , n13733 , RI17401f68_1498);
and ( n13735 , n43550 , n29614 );
or ( n43551 , n13734 , n13735 );
not ( n13736 , RI1754c610_2);
and ( n13737 , n13736 , n43551 );
and ( n13738 , C0 , RI1754c610_2);
or ( n43552 , n13737 , n13738 );
buf ( n43553 , n43552 );
not ( n43554 , n43414 );
xor ( n43555 , n42375 , n36431 );
xor ( n43556 , n43555 , n34221 );
and ( n43557 , n43554 , n43556 );
xor ( n43558 , n43411 , n43557 );
not ( n13739 , n29614 );
and ( n13740 , n13739 , RI173d7b78_1704);
and ( n13741 , n43558 , n29614 );
or ( n43559 , n13740 , n13741 );
not ( n13742 , RI1754c610_2);
and ( n13743 , n13742 , n43559 );
and ( n13744 , C0 , RI1754c610_2);
or ( n43560 , n13743 , n13744 );
buf ( n43561 , n43560 );
not ( n13745 , n27683 );
and ( n13746 , n13745 , RI19ab73c8_2400);
and ( n13747 , RI19ac0338_2330 , n27683 );
or ( n43562 , n13746 , n13747 );
not ( n13748 , RI1754c610_2);
and ( n13749 , n13748 , n43562 );
and ( n13750 , C0 , RI1754c610_2);
or ( n43563 , n13749 , n13750 );
buf ( n43564 , n43563 );
xor ( n43565 , n39331 , n35416 );
xor ( n43566 , n43565 , n29843 );
xor ( n43567 , n39207 , n37676 );
xor ( n43568 , n43567 , n37696 );
not ( n43569 , n43568 );
xor ( n43570 , n35088 , n40283 );
xor ( n43571 , n43570 , n32560 );
and ( n43572 , n43569 , n43571 );
xor ( n43573 , n43566 , n43572 );
not ( n13751 , n29614 );
and ( n13752 , n13751 , RI173a9c60_1928);
and ( n13753 , n43573 , n29614 );
or ( n43574 , n13752 , n13753 );
not ( n13754 , RI1754c610_2);
and ( n13755 , n13754 , n43574 );
and ( n13756 , C0 , RI1754c610_2);
or ( n43575 , n13755 , n13756 );
buf ( n43576 , n43575 );
buf ( n43577 , RI174b0658_876);
not ( n13757 , n27683 );
and ( n13758 , n13757 , RI19ac3290_2305);
and ( n13759 , RI19acc200_2238 , n27683 );
or ( n43578 , n13758 , n13759 );
not ( n13760 , RI1754c610_2);
and ( n13761 , n13760 , n43578 );
and ( n13762 , C0 , RI1754c610_2);
or ( n43579 , n13761 , n13762 );
buf ( n43580 , n43579 );
buf ( n43581 , RI174a2738_944);
buf ( n43582 , RI17495880_1007);
xor ( n43583 , n36055 , n34475 );
xor ( n43584 , n43583 , n37371 );
xor ( n43585 , n31379 , n37074 );
xor ( n43586 , n43585 , n37104 );
not ( n43587 , n43586 );
xor ( n43588 , n35520 , n37460 );
xor ( n43589 , n43588 , n37490 );
and ( n43590 , n43587 , n43589 );
xor ( n43591 , n43584 , n43590 );
not ( n13763 , n29614 );
and ( n13764 , n13763 , RI173b1fa0_1888);
and ( n13765 , n43591 , n29614 );
or ( n43592 , n13764 , n13765 );
not ( n13766 , RI1754c610_2);
and ( n13767 , n13766 , n43592 );
and ( n13768 , C0 , RI1754c610_2);
or ( n43593 , n13767 , n13768 );
buf ( n43594 , n43593 );
buf ( n43595 , RI174c67c8_793);
xor ( n43596 , n37638 , n40149 );
xor ( n43597 , n43596 , n40166 );
not ( n43598 , n41227 );
and ( n43599 , n43598 , n41242 );
xor ( n43600 , n43597 , n43599 );
not ( n13769 , n29614 );
and ( n13770 , n13769 , RI173e1f88_1654);
and ( n13771 , n43600 , n29614 );
or ( n43601 , n13770 , n13771 );
not ( n13772 , RI1754c610_2);
and ( n13773 , n13772 , n43601 );
and ( n13774 , C0 , RI1754c610_2);
or ( n43602 , n13773 , n13774 );
buf ( n43603 , n43602 );
not ( n13775 , n27683 );
and ( n13776 , n13775 , RI19a8b700_2715);
and ( n13777 , RI19a95930_2643 , n27683 );
or ( n43604 , n13776 , n13777 );
not ( n13778 , RI1754c610_2);
and ( n13779 , n13778 , n43604 );
and ( n13780 , C0 , RI1754c610_2);
or ( n43605 , n13779 , n13780 );
buf ( n43606 , n43605 );
not ( n13781 , n27683 );
and ( n13782 , n13781 , RI19a9bfd8_2598);
and ( n13783 , RI19aa5560_2527 , n27683 );
or ( n43607 , n13782 , n13783 );
not ( n13784 , RI1754c610_2);
and ( n13785 , n13784 , n43607 );
and ( n13786 , C0 , RI1754c610_2);
or ( n43608 , n13785 , n13786 );
buf ( n43609 , n43608 );
xor ( n43610 , n33216 , n31317 );
xor ( n43611 , n43610 , n40302 );
xor ( n43612 , n34086 , n39525 );
xor ( n43613 , n43612 , n42377 );
not ( n43614 , n43613 );
and ( n43615 , n43614 , n42589 );
xor ( n43616 , n43611 , n43615 );
not ( n13787 , n29614 );
and ( n13788 , n13787 , RI173390a0_2163);
and ( n13789 , n43616 , n29614 );
or ( n43617 , n13788 , n13789 );
not ( n13790 , RI1754c610_2);
and ( n13791 , n13790 , n43617 );
and ( n13792 , C0 , RI1754c610_2);
or ( n43618 , n13791 , n13792 );
buf ( n43619 , n43618 );
xor ( n43620 , n37667 , n37549 );
xor ( n43621 , n43620 , n37579 );
xor ( n43622 , n33114 , n38244 );
xor ( n43623 , n43622 , n37235 );
not ( n43624 , n43623 );
xor ( n43625 , n36251 , n41370 );
xor ( n43626 , n43625 , n37898 );
and ( n43627 , n43624 , n43626 );
xor ( n43628 , n43621 , n43627 );
not ( n13793 , n29614 );
and ( n13794 , n13793 , RI1748e8f0_1041);
and ( n13795 , n43628 , n29614 );
or ( n43629 , n13794 , n13795 );
not ( n13796 , RI1754c610_2);
and ( n13797 , n13796 , n43629 );
and ( n13798 , C0 , RI1754c610_2);
or ( n43630 , n13797 , n13798 );
buf ( n43631 , n43630 );
xor ( n43632 , n41609 , n43278 );
xor ( n43633 , n43632 , n31664 );
xor ( n43634 , n39926 , n40890 );
xor ( n43635 , n43634 , n38724 );
not ( n43636 , n43635 );
xor ( n43637 , n30727 , n33728 );
xor ( n43638 , n43637 , n33778 );
and ( n43639 , n43636 , n43638 );
xor ( n43640 , n43633 , n43639 );
not ( n13799 , n29614 );
and ( n13800 , n13799 , RI17392650_2042);
and ( n13801 , n43640 , n29614 );
or ( n43641 , n13800 , n13801 );
not ( n13802 , RI1754c610_2);
and ( n13803 , n13802 , n43641 );
and ( n13804 , C0 , RI1754c610_2);
or ( n43642 , n13803 , n13804 );
buf ( n43643 , n43642 );
buf ( n43644 , RI174b16c0_871);
buf ( n43645 , RI174a1a18_948);
not ( n13805 , n27683 );
and ( n13806 , n13805 , RI19ac04a0_2329);
and ( n13807 , RI19ac96e0_2259 , n27683 );
or ( n43646 , n13806 , n13807 );
not ( n13808 , RI1754c610_2);
and ( n13809 , n13808 , n43646 );
and ( n13810 , C0 , RI1754c610_2);
or ( n43647 , n13809 , n13810 );
buf ( n43648 , n43647 );
xor ( n43649 , n36551 , n37438 );
xor ( n43650 , n43649 , n30247 );
xor ( n43651 , n34512 , n31380 );
xor ( n43652 , n43651 , n36463 );
not ( n43653 , n43652 );
xor ( n43654 , n35759 , n39563 );
xor ( n43655 , n43654 , n35416 );
and ( n43656 , n43653 , n43655 );
xor ( n43657 , n43650 , n43656 );
not ( n13811 , n29614 );
and ( n13812 , n13811 , RI17506bd8_745);
and ( n13813 , n43657 , n29614 );
or ( n43658 , n13812 , n13813 );
not ( n13814 , RI1754c610_2);
and ( n13815 , n13814 , n43658 );
and ( n13816 , C0 , RI1754c610_2);
or ( n43659 , n13815 , n13816 );
buf ( n43660 , n43659 );
xor ( n43661 , n37727 , n41772 );
xor ( n43662 , n43661 , n32663 );
xor ( n43663 , n36509 , n40381 );
xor ( n43664 , n43663 , n37438 );
not ( n43665 , n43664 );
xor ( n43666 , n36207 , n32923 );
xor ( n43667 , n43666 , n32973 );
and ( n43668 , n43665 , n43667 );
xor ( n43669 , n43662 , n43668 );
not ( n13817 , n29614 );
and ( n13818 , n13817 , RI17398230_2014);
and ( n13819 , n43669 , n29614 );
or ( n43670 , n13818 , n13819 );
not ( n13820 , RI1754c610_2);
and ( n13821 , n13820 , n43670 );
and ( n13822 , C0 , RI1754c610_2);
or ( n43671 , n13821 , n13822 );
buf ( n43672 , n43671 );
not ( n13823 , n27683 );
and ( n13824 , n13823 , RI19ac6620_2282);
and ( n13825 , RI19acf1d0_2217 , n27683 );
or ( n43673 , n13824 , n13825 );
not ( n13826 , RI1754c610_2);
and ( n13827 , n13826 , n43673 );
and ( n13828 , C0 , RI1754c610_2);
or ( n43674 , n13827 , n13828 );
buf ( n43675 , n43674 );
not ( n13829 , n27683 );
and ( n13830 , n13829 , RI19aa2068_2552);
and ( n13831 , RI19aac6d0_2480 , n27683 );
or ( n43676 , n13830 , n13831 );
not ( n13832 , RI1754c610_2);
and ( n13833 , n13832 , n43676 );
and ( n13834 , C0 , RI1754c610_2);
or ( n43677 , n13833 , n13834 );
buf ( n43678 , n43677 );
xor ( n43679 , n43455 , n40949 );
xor ( n43680 , n43679 , n34572 );
not ( n43681 , n43680 );
xor ( n43682 , n37455 , n36874 );
xor ( n43683 , n43682 , n42188 );
and ( n43684 , n43681 , n43683 );
xor ( n43685 , n42740 , n43684 );
not ( n13835 , n29614 );
and ( n13836 , n13835 , RI1744c860_1363);
and ( n13837 , n43685 , n29614 );
or ( n43686 , n13836 , n13837 );
not ( n13838 , RI1754c610_2);
and ( n13839 , n13838 , n43686 );
and ( n13840 , C0 , RI1754c610_2);
or ( n43687 , n13839 , n13840 );
buf ( n43688 , n43687 );
xor ( n43689 , n36973 , n41818 );
xor ( n43690 , n43689 , n40662 );
xor ( n43691 , n38918 , n42309 );
xor ( n43692 , n43691 , n43464 );
not ( n43693 , n43692 );
xor ( n43694 , n37671 , n37549 );
xor ( n43695 , n43694 , n37579 );
and ( n43696 , n43693 , n43695 );
xor ( n43697 , n43690 , n43696 );
not ( n13841 , n29614 );
and ( n13842 , n13841 , RI1738ee88_2059);
and ( n13843 , n43697 , n29614 );
or ( n43698 , n13842 , n13843 );
not ( n13844 , RI1754c610_2);
and ( n13845 , n13844 , n43698 );
and ( n13846 , C0 , RI1754c610_2);
or ( n43699 , n13845 , n13846 );
buf ( n43700 , n43699 );
not ( n13847 , n27683 );
and ( n13848 , n13847 , RI19aa10f0_2560);
and ( n13849 , RI19aab0c8_2488 , n27683 );
or ( n43701 , n13848 , n13849 );
not ( n13850 , RI1754c610_2);
and ( n13851 , n13850 , n43701 );
and ( n13852 , C0 , RI1754c610_2);
or ( n43702 , n13851 , n13852 );
buf ( n43703 , n43702 );
buf ( n43704 , RI1748fca0_1035);
buf ( n43705 , RI17494818_1012);
buf ( n43706 , RI17486c40_1079);
buf ( n43707 , RI1748b7b8_1056);
xor ( n43708 , n31652 , n30604 );
xor ( n43709 , n43708 , n30741 );
xor ( n43710 , n37027 , n40662 );
xor ( n43711 , n43710 , n39208 );
not ( n43712 , n43711 );
xor ( n43713 , n37572 , n34968 );
xor ( n43714 , n43713 , n39771 );
and ( n43715 , n43712 , n43714 );
xor ( n43716 , n43709 , n43715 );
not ( n13853 , n29614 );
and ( n13854 , n13853 , RI17456928_1314);
and ( n13855 , n43716 , n29614 );
or ( n43717 , n13854 , n13855 );
not ( n13856 , RI1754c610_2);
and ( n13857 , n13856 , n43717 );
and ( n13858 , C0 , RI1754c610_2);
or ( n43718 , n13857 , n13858 );
buf ( n43719 , n43718 );
buf ( n43720 , RI174d0278_763);
xor ( n43721 , n32761 , n37186 );
xor ( n43722 , n43721 , n37203 );
xor ( n43723 , n36225 , n31831 );
xor ( n43724 , n43723 , n31925 );
not ( n43725 , n43724 );
xor ( n43726 , n33336 , n38991 );
xor ( n43727 , n43726 , n39005 );
and ( n43728 , n43725 , n43727 );
xor ( n43729 , n43722 , n43728 );
not ( n13859 , n29614 );
and ( n13860 , n13859 , RI1745c1c0_1287);
and ( n13861 , n43729 , n29614 );
or ( n43730 , n13860 , n13861 );
not ( n13862 , RI1754c610_2);
and ( n13863 , n13862 , n43730 );
and ( n13864 , C0 , RI1754c610_2);
or ( n43731 , n13863 , n13864 );
buf ( n43732 , n43731 );
buf ( n43733 , RI1750dd48_723);
xor ( n43734 , n35442 , n32715 );
xor ( n43735 , n43734 , n36654 );
xor ( n43736 , n33251 , n40302 );
xor ( n43737 , n43736 , n40319 );
not ( n43738 , n43737 );
and ( n43739 , n43738 , n38245 );
xor ( n43740 , n43735 , n43739 );
not ( n13865 , n29614 );
and ( n13866 , n13865 , RI1733c1d8_2148);
and ( n13867 , n43740 , n29614 );
or ( n43741 , n13866 , n13867 );
not ( n13868 , RI1754c610_2);
and ( n13869 , n13868 , n43741 );
and ( n13870 , C0 , RI1754c610_2);
or ( n43742 , n13869 , n13870 );
buf ( n43743 , n43742 );
xor ( n43744 , n34040 , n34251 );
xor ( n43745 , n43744 , n42033 );
xor ( n43746 , n41727 , n34837 );
xor ( n43747 , n43746 , n33880 );
not ( n43748 , n43747 );
xor ( n43749 , n40992 , n36998 );
xor ( n43750 , n43749 , n37048 );
and ( n43751 , n43748 , n43750 );
xor ( n43752 , n43745 , n43751 );
not ( n13871 , n29614 );
and ( n13872 , n13871 , RI174122a0_1419);
and ( n13873 , n43752 , n29614 );
or ( n43753 , n13872 , n13873 );
not ( n13874 , RI1754c610_2);
and ( n13875 , n13874 , n43753 );
and ( n13876 , C0 , RI1754c610_2);
or ( n43754 , n13875 , n13876 );
buf ( n43755 , n43754 );
buf ( n43756 , RI174c24c0_806);
not ( n43757 , n42723 );
and ( n43758 , n43757 , n42725 );
xor ( n43759 , n43050 , n43758 );
not ( n13877 , n29614 );
and ( n13878 , n13877 , RI173fb668_1530);
and ( n13879 , n43759 , n29614 );
or ( n43760 , n13878 , n13879 );
not ( n13880 , RI1754c610_2);
and ( n13881 , n13880 , n43760 );
and ( n13882 , C0 , RI1754c610_2);
or ( n43761 , n13881 , n13882 );
buf ( n43762 , n43761 );
buf ( n43763 , RI174c9b58_783);
and ( n43764 , RI1754c250_10 , n34844 );
and ( n43765 , RI1754c250_10 , n34847 );
and ( n43766 , RI1754c250_10 , n34850 );
and ( n43767 , RI1754c250_10 , n34852 );
and ( n43768 , RI1754c250_10 , n34854 );
and ( n43769 , RI1754c250_10 , n34856 );
and ( n43770 , RI1754c250_10 , n39233 );
nor ( n43771 , RI1754a5b8_71 , RI1754a630_70 , RI1754a6a8_69);
buf ( n43772 , n43771 );
or ( n43773 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43772 );
not ( n13883 , n34859 );
and ( n13884 , n13883 , n43773 );
and ( n13885 , RI1754c250_10 , n34859 );
or ( n43774 , n13884 , n13885 );
not ( n13886 , RI19a22f70_2797);
and ( n13887 , n13886 , n43774 );
and ( n13888 , C0 , RI19a22f70_2797);
or ( n43775 , n13887 , n13888 );
not ( n13889 , n27683 );
and ( n13890 , n13889 , RI19a89e28_2725);
and ( n13891 , n43775 , n27683 );
or ( n43776 , n13890 , n13891 );
not ( n13892 , RI1754c610_2);
and ( n13893 , n13892 , n43776 );
and ( n13894 , C0 , RI1754c610_2);
or ( n43777 , n13893 , n13894 );
buf ( n43778 , n43777 );
not ( n43779 , n42888 );
and ( n43780 , n43779 , n42574 );
xor ( n43781 , n42885 , n43780 );
not ( n13895 , n29614 );
and ( n13896 , n13895 , RI173f7ea0_1547);
and ( n13897 , n43781 , n29614 );
or ( n43782 , n13896 , n13897 );
not ( n13898 , RI1754c610_2);
and ( n13899 , n13898 , n43782 );
and ( n13900 , C0 , RI1754c610_2);
or ( n43783 , n13899 , n13900 );
buf ( n43784 , n43783 );
not ( n13901 , n27683 );
and ( n13902 , n13901 , RI19a964e8_2638);
and ( n13903 , RI19aa0358_2567 , n27683 );
or ( n43785 , n13902 , n13903 );
not ( n13904 , RI1754c610_2);
and ( n13905 , n13904 , n43785 );
and ( n13906 , C0 , RI1754c610_2);
or ( n43786 , n13905 , n13906 );
buf ( n43787 , n43786 );
not ( n43788 , n42461 );
xor ( n43789 , n39885 , n42504 );
xor ( n43790 , n43789 , n41818 );
and ( n43791 , n43788 , n43790 );
xor ( n43792 , n42458 , n43791 );
not ( n13907 , n29614 );
and ( n13908 , n13907 , RI1739a648_2003);
and ( n13909 , n43792 , n29614 );
or ( n43793 , n13908 , n13909 );
not ( n13910 , RI1754c610_2);
and ( n13911 , n13910 , n43793 );
and ( n13912 , C0 , RI1754c610_2);
or ( n43794 , n13911 , n13912 );
buf ( n43795 , n43794 );
xor ( n43796 , n41381 , n33567 );
xor ( n43797 , n43796 , n33617 );
xor ( n43798 , n37177 , n32481 );
xor ( n43799 , n43798 , n33030 );
not ( n43800 , n43799 );
xor ( n43801 , n38366 , n33880 );
xor ( n43802 , n43801 , n33935 );
and ( n43803 , n43800 , n43802 );
xor ( n43804 , n43797 , n43803 );
not ( n13913 , n29614 );
and ( n13914 , n13913 , RI17390238_2053);
and ( n13915 , n43804 , n29614 );
or ( n43805 , n13914 , n13915 );
not ( n13916 , RI1754c610_2);
and ( n13917 , n13916 , n43805 );
and ( n13918 , C0 , RI1754c610_2);
or ( n43806 , n13917 , n13918 );
buf ( n43807 , n43806 );
xor ( n43808 , n35429 , n32663 );
xor ( n43809 , n43808 , n32715 );
xor ( n43810 , n32962 , n41659 );
xor ( n43811 , n43810 , n37800 );
not ( n43812 , n43811 );
xor ( n43813 , n37234 , n39467 );
xor ( n43814 , n43813 , n41391 );
and ( n43815 , n43812 , n43814 );
xor ( n43816 , n43809 , n43815 );
not ( n13919 , n29614 );
and ( n13920 , n13919 , RI17460018_1268);
and ( n13921 , n43816 , n29614 );
or ( n43817 , n13920 , n13921 );
not ( n13922 , RI1754c610_2);
and ( n13923 , n13922 , n43817 );
and ( n13924 , C0 , RI1754c610_2);
or ( n43818 , n13923 , n13924 );
buf ( n43819 , n43818 );
xor ( n43820 , n39847 , n36742 );
xor ( n43821 , n43820 , n42504 );
xor ( n43822 , n40803 , n40437 );
xor ( n43823 , n43822 , n42635 );
not ( n43824 , n43823 );
xor ( n43825 , n38400 , n37169 );
xor ( n43826 , n43825 , n36339 );
and ( n43827 , n43824 , n43826 );
xor ( n43828 , n43821 , n43827 );
not ( n13925 , n29614 );
and ( n13926 , n13925 , RI173a7500_1940);
and ( n13927 , n43828 , n29614 );
or ( n43829 , n13926 , n13927 );
not ( n13928 , RI1754c610_2);
and ( n13929 , n13928 , n43829 );
and ( n13930 , C0 , RI1754c610_2);
or ( n43830 , n13929 , n13930 );
buf ( n43831 , n43830 );
not ( n43832 , n43735 );
and ( n43833 , n43832 , n43737 );
xor ( n43834 , n38285 , n43833 );
not ( n13931 , n29614 );
and ( n13932 , n13931 , RI173b6b18_1865);
and ( n13933 , n43834 , n29614 );
or ( n43835 , n13932 , n13933 );
not ( n13934 , RI1754c610_2);
and ( n13935 , n13934 , n43835 );
and ( n13936 , C0 , RI1754c610_2);
or ( n43836 , n13935 , n13936 );
buf ( n43837 , n43836 );
xor ( n43838 , n37113 , n40237 );
xor ( n43839 , n43838 , n40254 );
not ( n43840 , n41267 );
and ( n43841 , n43840 , n41269 );
xor ( n43842 , n43839 , n43841 );
not ( n13937 , n29614 );
and ( n13938 , n13937 , RI17411580_1423);
and ( n13939 , n43842 , n29614 );
or ( n43843 , n13938 , n13939 );
not ( n13940 , RI1754c610_2);
and ( n13941 , n13940 , n43843 );
and ( n13942 , C0 , RI1754c610_2);
or ( n43844 , n13941 , n13942 );
buf ( n43845 , n43844 );
xor ( n43846 , n33680 , n41854 );
xor ( n43847 , n43846 , n40283 );
not ( n43848 , n43847 );
xor ( n43849 , n40144 , n38948 );
xor ( n43850 , n43849 , n39039 );
and ( n43851 , n43848 , n43850 );
xor ( n43852 , n43750 , n43851 );
not ( n13943 , n29614 );
and ( n13944 , n13943 , RI17452ad0_1333);
and ( n13945 , n43852 , n29614 );
or ( n43853 , n13944 , n13945 );
not ( n13946 , RI1754c610_2);
and ( n13947 , n13946 , n43853 );
and ( n13948 , C0 , RI1754c610_2);
or ( n43854 , n13947 , n13948 );
buf ( n43855 , n43854 );
xor ( n43856 , n42255 , n40743 );
xor ( n43857 , n43856 , n36062 );
not ( n43858 , n43857 );
xor ( n43859 , n37519 , n37942 );
xor ( n43860 , n43859 , n34395 );
and ( n43861 , n43858 , n43860 );
xor ( n43862 , n41451 , n43861 );
not ( n13949 , n29614 );
and ( n13950 , n13949 , RI17390f58_2049);
and ( n13951 , n43862 , n29614 );
or ( n43863 , n13950 , n13951 );
not ( n13952 , RI1754c610_2);
and ( n13953 , n13952 , n43863 );
and ( n13954 , C0 , RI1754c610_2);
or ( n43864 , n13953 , n13954 );
buf ( n43865 , n43864 );
buf ( n43866 , RI17491398_1028);
not ( n13955 , n27683 );
and ( n13956 , n13955 , RI19aacbf8_2477);
and ( n13957 , RI19ab65b8_2406 , n27683 );
or ( n43867 , n13956 , n13957 );
not ( n13958 , RI1754c610_2);
and ( n13959 , n13958 , n43867 );
and ( n13960 , C0 , RI1754c610_2);
or ( n43868 , n13959 , n13960 );
buf ( n43869 , n43868 );
buf ( n43870 , RI174c7740_790);
xor ( n43871 , n40209 , n34041 );
xor ( n43872 , n43871 , n41934 );
xor ( n43873 , n32635 , n36195 );
xor ( n43874 , n43873 , n36209 );
not ( n43875 , n43874 );
xor ( n43876 , n34279 , n38886 );
xor ( n43877 , n43876 , n39604 );
and ( n43878 , n43875 , n43877 );
xor ( n43879 , n43872 , n43878 );
not ( n13961 , n29614 );
and ( n13962 , n13961 , RI17335c20_2179);
and ( n13963 , n43879 , n29614 );
or ( n43880 , n13962 , n13963 );
not ( n13964 , RI1754c610_2);
and ( n13965 , n13964 , n43880 );
and ( n13966 , C0 , RI1754c610_2);
or ( n43881 , n13965 , n13966 );
buf ( n43882 , n43881 );
not ( n13967 , n27683 );
and ( n13968 , n13967 , RI19aaf088_2461);
and ( n13969 , RI19ab8d90_2389 , n27683 );
or ( n43883 , n13968 , n13969 );
not ( n13970 , RI1754c610_2);
and ( n13971 , n13970 , n43883 );
and ( n13972 , C0 , RI1754c610_2);
or ( n43884 , n13971 , n13972 );
buf ( n43885 , n43884 );
not ( n43886 , n37375 );
xor ( n43887 , n41046 , n34395 );
xor ( n43888 , n43887 , n34445 );
and ( n43889 , n43886 , n43888 );
xor ( n43890 , n37372 , n43889 );
not ( n13973 , n29614 );
and ( n13974 , n13973 , RI173caca8_1767);
and ( n13975 , n43890 , n29614 );
or ( n43891 , n13974 , n13975 );
not ( n13976 , RI1754c610_2);
and ( n13977 , n13976 , n43891 );
and ( n13978 , C0 , RI1754c610_2);
or ( n43892 , n13977 , n13978 );
buf ( n43893 , n43892 );
not ( n43894 , n39894 );
and ( n43895 , n43894 , n39915 );
xor ( n43896 , n40831 , n43895 );
not ( n13979 , n29614 );
and ( n13980 , n13979 , RI17347308_2094);
and ( n13981 , n43896 , n29614 );
or ( n43897 , n13980 , n13981 );
not ( n13982 , RI1754c610_2);
and ( n13983 , n13982 , n43897 );
and ( n13984 , C0 , RI1754c610_2);
or ( n43898 , n13983 , n13984 );
buf ( n43899 , n43898 );
xor ( n43900 , n31724 , n30741 );
xor ( n43901 , n43900 , n40769 );
xor ( n43902 , n38413 , n40585 );
xor ( n43903 , n43902 , n34918 );
not ( n43904 , n43903 );
and ( n43905 , n43904 , n43797 );
xor ( n43906 , n43901 , n43905 );
not ( n13985 , n29614 );
and ( n13986 , n13985 , RI173bc068_1839);
and ( n13987 , n43906 , n29614 );
or ( n43907 , n13986 , n13987 );
not ( n13988 , RI1754c610_2);
and ( n13989 , n13988 , n43907 );
and ( n13990 , C0 , RI1754c610_2);
or ( n43908 , n13989 , n13990 );
buf ( n43909 , n43908 );
xor ( n43910 , n32107 , n36702 );
xor ( n43911 , n43910 , n38872 );
xor ( n43912 , n30802 , n38115 );
xor ( n43913 , n43912 , n41622 );
not ( n43914 , n43913 );
xor ( n43915 , n38762 , n40516 );
xor ( n43916 , n43915 , n40966 );
and ( n43917 , n43914 , n43916 );
xor ( n43918 , n43911 , n43917 );
not ( n13991 , n29614 );
and ( n13992 , n13991 , RI173bf1a0_1824);
and ( n13993 , n43918 , n29614 );
or ( n43919 , n13992 , n13993 );
not ( n13994 , RI1754c610_2);
and ( n13995 , n13994 , n43919 );
and ( n13996 , C0 , RI1754c610_2);
or ( n43920 , n13995 , n13996 );
buf ( n43921 , n43920 );
xor ( n43922 , n38392 , n37169 );
xor ( n43923 , n43922 , n36339 );
xor ( n43924 , n38867 , n41125 );
xor ( n43925 , n43924 , n31506 );
not ( n43926 , n43925 );
xor ( n43927 , n37868 , n35128 );
xor ( n43928 , n43927 , n36917 );
and ( n43929 , n43926 , n43928 );
xor ( n43930 , n43923 , n43929 );
not ( n13997 , n29614 );
and ( n13998 , n13997 , RI17502e70_751);
and ( n13999 , n43930 , n29614 );
or ( n43931 , n13998 , n13999 );
not ( n14000 , RI1754c610_2);
and ( n14001 , n14000 , n43931 );
and ( n14002 , C0 , RI1754c610_2);
or ( n43932 , n14001 , n14002 );
buf ( n43933 , n43932 );
xor ( n43934 , n40470 , n38933 );
xor ( n43935 , n43934 , n41430 );
xor ( n43936 , n36391 , n34190 );
xor ( n43937 , n43936 , n36252 );
not ( n43938 , n43937 );
and ( n43939 , n43938 , n39210 );
xor ( n43940 , n43935 , n43939 );
not ( n14003 , n29614 );
and ( n14004 , n14003 , RI173c8890_1778);
and ( n14005 , n43940 , n29614 );
or ( n43941 , n14004 , n14005 );
not ( n14006 , RI1754c610_2);
and ( n14007 , n14006 , n43941 );
and ( n14008 , C0 , RI1754c610_2);
or ( n43942 , n14007 , n14008 );
buf ( n43943 , n43942 );
xor ( n43944 , n32559 , n37651 );
xor ( n43945 , n43944 , n39182 );
xor ( n43946 , n31647 , n30604 );
xor ( n43947 , n43946 , n30741 );
not ( n43948 , n43947 );
xor ( n43949 , n37278 , n34127 );
xor ( n43950 , n43949 , n40190 );
and ( n43951 , n43948 , n43950 );
xor ( n43952 , n43945 , n43951 );
not ( n14009 , n29614 );
and ( n14010 , n14009 , RI17532e40_608);
and ( n14011 , n43952 , n29614 );
or ( n43953 , n14010 , n14011 );
not ( n14012 , RI1754c610_2);
and ( n14013 , n14012 , n43953 );
and ( n14014 , C0 , RI1754c610_2);
or ( n43954 , n14013 , n14014 );
buf ( n43955 , n43954 );
xor ( n43956 , n40025 , n40855 );
xor ( n43957 , n43956 , n38574 );
xor ( n43958 , n30907 , n38115 );
xor ( n43959 , n43958 , n41622 );
not ( n43960 , n43959 );
xor ( n43961 , n36681 , n39635 );
xor ( n43962 , n43961 , n39655 );
and ( n43963 , n43960 , n43962 );
xor ( n43964 , n43957 , n43963 );
not ( n14015 , n29614 );
and ( n14016 , n14015 , RI175153e0_700);
and ( n14017 , n43964 , n29614 );
or ( n43965 , n14016 , n14017 );
not ( n14018 , RI1754c610_2);
and ( n14019 , n14018 , n43965 );
and ( n14020 , C0 , RI1754c610_2);
or ( n43966 , n14019 , n14020 );
buf ( n43967 , n43966 );
xor ( n43968 , n38876 , n31506 );
xor ( n43969 , n43968 , n31621 );
xor ( n43970 , n33007 , n35639 );
xor ( n43971 , n43970 , n36227 );
not ( n43972 , n43971 );
xor ( n43973 , n33914 , n37291 );
xor ( n43974 , n43973 , n37311 );
and ( n43975 , n43972 , n43974 );
xor ( n43976 , n43969 , n43975 );
not ( n14021 , n29614 );
and ( n14022 , n14021 , RI174b1030_873);
and ( n14023 , n43976 , n29614 );
or ( n43977 , n14022 , n14023 );
not ( n14024 , RI1754c610_2);
and ( n14025 , n14024 , n43977 );
and ( n14026 , C0 , RI1754c610_2);
or ( n43978 , n14025 , n14026 );
buf ( n43979 , n43978 );
xor ( n43980 , n41465 , n39686 );
xor ( n43981 , n43980 , n34087 );
not ( n43982 , n37757 );
and ( n43983 , n43982 , n37759 );
xor ( n43984 , n40416 , n43983 );
not ( n43985 , n37766 );
and ( n43986 , n43985 , n37768 );
xor ( n43987 , n40421 , n43986 );
xor ( n43988 , n43984 , n43987 );
not ( n43989 , n37776 );
and ( n43990 , n43989 , n37778 );
xor ( n43991 , n40427 , n43990 );
xor ( n43992 , n43988 , n43991 );
xor ( n43993 , n43992 , n41343 );
xor ( n43994 , n43993 , n40789 );
xor ( n43995 , n37783 , n43994 );
xor ( n43996 , n43995 , n31213 );
not ( n43997 , n43996 );
and ( n43998 , n43997 , n39831 );
xor ( n43999 , n43981 , n43998 );
not ( n14027 , n29614 );
and ( n14028 , n14027 , RI173e0f20_1659);
and ( n14029 , n43999 , n29614 );
or ( n44000 , n14028 , n14029 );
not ( n14030 , RI1754c610_2);
and ( n14031 , n14030 , n44000 );
and ( n14032 , C0 , RI1754c610_2);
or ( n44001 , n14031 , n14032 );
buf ( n44002 , n44001 );
xor ( n44003 , n32354 , n41316 );
xor ( n44004 , n44003 , n35622 );
not ( n44005 , n44004 );
and ( n44006 , n44005 , n42421 );
xor ( n44007 , n38952 , n44006 );
not ( n14033 , n29614 );
and ( n14034 , n14033 , RI174c9108_785);
and ( n14035 , n44007 , n29614 );
or ( n44008 , n14034 , n14035 );
not ( n14036 , RI1754c610_2);
and ( n14037 , n14036 , n44008 );
and ( n14038 , C0 , RI1754c610_2);
or ( n44009 , n14037 , n14038 );
buf ( n44010 , n44009 );
not ( n44011 , n34341 );
and ( n44012 , n44011 , n34446 );
xor ( n44013 , n39184 , n44012 );
not ( n14039 , n29614 );
and ( n14040 , n14039 , RI174cc9c0_774);
and ( n14041 , n44013 , n29614 );
or ( n44014 , n14040 , n14041 );
not ( n14042 , RI1754c610_2);
and ( n14043 , n14042 , n44014 );
and ( n14044 , C0 , RI1754c610_2);
or ( n44015 , n14043 , n14044 );
buf ( n44016 , n44015 );
not ( n14045 , n27683 );
and ( n14046 , n14045 , RI19ab3840_2427);
and ( n14047 , RI19abd6b0_2355 , n27683 );
or ( n44017 , n14046 , n14047 );
not ( n14048 , RI1754c610_2);
and ( n14049 , n14048 , n44017 );
and ( n14050 , C0 , RI1754c610_2);
or ( n44018 , n14049 , n14050 );
buf ( n44019 , n44018 );
and ( n44020 , RI1754b1e8_45 , n34844 );
and ( n44021 , RI1754b1e8_45 , n34847 );
or ( n44022 , n44020 , n44021 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n14051 , n34859 );
and ( n14052 , n14051 , n44022 );
and ( n14053 , RI1754b1e8_45 , n34859 );
or ( n44023 , n14052 , n14053 );
not ( n14054 , RI19a22f70_2797);
and ( n14055 , n14054 , n44023 );
and ( n14056 , C0 , RI19a22f70_2797);
or ( n44024 , n14055 , n14056 );
not ( n14057 , n27683 );
and ( n14058 , n14057 , RI19abf690_2337);
and ( n14059 , n44024 , n27683 );
or ( n44025 , n14058 , n14059 );
not ( n14060 , RI1754c610_2);
and ( n14061 , n14060 , n44025 );
and ( n14062 , C0 , RI1754c610_2);
or ( n44026 , n14061 , n14062 );
buf ( n44027 , n44026 );
not ( n44028 , n43790 );
xor ( n44029 , n40812 , n42635 );
xor ( n44030 , n44029 , n33648 );
and ( n44031 , n44028 , n44030 );
xor ( n44032 , n42461 , n44031 );
not ( n14063 , n29614 );
and ( n14064 , n14063 , RI173a8f40_1932);
and ( n14065 , n44032 , n29614 );
or ( n44033 , n14064 , n14065 );
not ( n14066 , RI1754c610_2);
and ( n14067 , n14066 , n44033 );
and ( n14068 , C0 , RI1754c610_2);
or ( n44034 , n14067 , n14068 );
buf ( n44035 , n44034 );
xor ( n44036 , n42259 , n40743 );
xor ( n44037 , n44036 , n36062 );
not ( n44038 , n44037 );
xor ( n44039 , n40562 , n40966 );
xor ( n44040 , n44039 , n37460 );
and ( n44041 , n44038 , n44040 );
xor ( n44042 , n39706 , n44041 );
not ( n14069 , n29614 );
and ( n14070 , n14069 , RI17485890_1085);
and ( n14071 , n44042 , n29614 );
or ( n44043 , n14070 , n14071 );
not ( n14072 , RI1754c610_2);
and ( n14073 , n14072 , n44043 );
and ( n14074 , C0 , RI1754c610_2);
or ( n44044 , n14073 , n14074 );
buf ( n44045 , n44044 );
not ( n14075 , n27683 );
and ( n14076 , n14075 , RI19a8ed60_2691);
and ( n14077 , RI19a98d38_2620 , n27683 );
or ( n44046 , n14076 , n14077 );
not ( n14078 , RI1754c610_2);
and ( n14079 , n14078 , n44046 );
and ( n14080 , C0 , RI1754c610_2);
or ( n44047 , n14079 , n14080 );
buf ( n44048 , n44047 );
not ( n44049 , n43877 );
xor ( n44050 , n35483 , n38512 );
xor ( n44051 , n44050 , n38532 );
and ( n44052 , n44049 , n44051 );
xor ( n44053 , n43874 , n44052 );
not ( n14081 , n29614 );
and ( n14082 , n14081 , RI174b2a70_865);
and ( n14083 , n44053 , n29614 );
or ( n44054 , n14082 , n14083 );
not ( n14084 , RI1754c610_2);
and ( n14085 , n14084 , n44054 );
and ( n14086 , C0 , RI1754c610_2);
or ( n44055 , n14085 , n14086 );
buf ( n44056 , n44055 );
xor ( n44057 , n34917 , n36772 );
xor ( n44058 , n44057 , n36802 );
not ( n44059 , n38349 );
and ( n44060 , n44059 , n38351 );
xor ( n44061 , n44058 , n44060 );
not ( n14087 , n29614 );
and ( n14088 , n14087 , RI17333b50_2189);
and ( n14089 , n44061 , n29614 );
or ( n44062 , n14088 , n14089 );
not ( n14090 , RI1754c610_2);
and ( n14091 , n14090 , n44062 );
and ( n14092 , C0 , RI1754c610_2);
or ( n44063 , n14091 , n14092 );
buf ( n44064 , n44063 );
not ( n14093 , n27683 );
and ( n14094 , n14093 , RI19aaf628_2458);
and ( n14095 , RI19ab92b8_2387 , n27683 );
or ( n44065 , n14094 , n14095 );
not ( n14096 , RI1754c610_2);
and ( n14097 , n14096 , n44065 );
and ( n14098 , C0 , RI1754c610_2);
or ( n44066 , n14097 , n14098 );
buf ( n44067 , n44066 );
xor ( n44068 , n37447 , n36874 );
xor ( n44069 , n44068 , n42188 );
not ( n44070 , n44069 );
xor ( n44071 , n42545 , n37421 );
xor ( n44072 , n44071 , n42605 );
and ( n44073 , n44070 , n44072 );
xor ( n44074 , n42163 , n44073 );
not ( n14099 , n29614 );
and ( n14100 , n14099 , RI173c74e0_1784);
and ( n14101 , n44074 , n29614 );
or ( n44075 , n14100 , n14101 );
not ( n14102 , RI1754c610_2);
and ( n14103 , n14102 , n44075 );
and ( n14104 , C0 , RI1754c610_2);
or ( n44076 , n14103 , n14104 );
buf ( n44077 , n44076 );
not ( n44078 , n40052 );
and ( n44079 , n44078 , n41327 );
xor ( n44080 , n40010 , n44079 );
not ( n14105 , n29614 );
and ( n14106 , n14105 , RI173bb9d8_1841);
and ( n14107 , n44080 , n29614 );
or ( n44081 , n14106 , n14107 );
not ( n14108 , RI1754c610_2);
and ( n14109 , n14108 , n44081 );
and ( n14110 , C0 , RI1754c610_2);
or ( n44082 , n14109 , n14110 );
buf ( n44083 , n44082 );
xor ( n44084 , n34244 , n37526 );
xor ( n44085 , n44084 , n41049 );
xor ( n44086 , n35271 , n39952 );
xor ( n44087 , n44086 , n42945 );
not ( n44088 , n44087 );
and ( n44089 , n44088 , n43494 );
xor ( n44090 , n44085 , n44089 );
not ( n14111 , n29614 );
and ( n14112 , n14111 , RI173b95c0_1852);
and ( n14113 , n44090 , n29614 );
or ( n44091 , n14112 , n14113 );
not ( n14114 , RI1754c610_2);
and ( n14115 , n14114 , n44091 );
and ( n14116 , C0 , RI1754c610_2);
or ( n44092 , n14115 , n14116 );
buf ( n44093 , n44092 );
xor ( n44094 , n37302 , n40190 );
xor ( n44095 , n44094 , n40210 );
xor ( n44096 , n39504 , n30923 );
xor ( n44097 , n44096 , n31053 );
not ( n44098 , n44097 );
xor ( n44099 , n35415 , n41068 );
xor ( n44100 , n44099 , n39091 );
and ( n44101 , n44098 , n44100 );
xor ( n44102 , n44095 , n44101 );
not ( n14117 , n29614 );
and ( n14118 , n14117 , RI173e7b68_1626);
and ( n14119 , n44102 , n29614 );
or ( n44103 , n14118 , n14119 );
not ( n14120 , RI1754c610_2);
and ( n14121 , n14120 , n44103 );
and ( n14122 , C0 , RI1754c610_2);
or ( n44104 , n14121 , n14122 );
buf ( n44105 , n44104 );
not ( n44106 , n43974 );
xor ( n44107 , n39032 , n36947 );
xor ( n44108 , n44107 , n39702 );
and ( n44109 , n44106 , n44108 );
xor ( n44110 , n43971 , n44109 );
not ( n14123 , n29614 );
and ( n14124 , n14123 , RI174c3960_802);
and ( n14125 , n44110 , n29614 );
or ( n44111 , n14124 , n14125 );
not ( n14126 , RI1754c610_2);
and ( n14127 , n14126 , n44111 );
and ( n14128 , C0 , RI1754c610_2);
or ( n44112 , n14127 , n14128 );
buf ( n44113 , n44112 );
xor ( n44114 , n39761 , n33125 );
xor ( n44115 , n44114 , n33175 );
not ( n44116 , n42235 );
and ( n44117 , n44116 , n42237 );
xor ( n44118 , n44115 , n44117 );
not ( n14129 , n29614 );
and ( n14130 , n14129 , RI1747adf0_1137);
and ( n14131 , n44118 , n29614 );
or ( n44119 , n14130 , n14131 );
not ( n14132 , RI1754c610_2);
and ( n14133 , n14132 , n44119 );
and ( n14134 , C0 , RI1754c610_2);
or ( n44120 , n14133 , n14134 );
buf ( n44121 , n44120 );
not ( n14135 , n27683 );
and ( n14136 , n14135 , RI19aab0c8_2488);
and ( n14137 , RI19ab4dd0_2417 , n27683 );
or ( n44122 , n14136 , n14137 );
not ( n14138 , RI1754c610_2);
and ( n14139 , n14138 , n44122 );
and ( n14140 , C0 , RI1754c610_2);
or ( n44123 , n14139 , n14140 );
buf ( n44124 , n44123 );
xor ( n44125 , n34001 , n34251 );
xor ( n44126 , n44125 , n42033 );
not ( n44127 , n43633 );
and ( n44128 , n44127 , n43635 );
xor ( n44129 , n44126 , n44128 );
not ( n14141 , n29614 );
and ( n14142 , n14141 , RI173434b0_2113);
and ( n14143 , n44129 , n29614 );
or ( n44130 , n14142 , n14143 );
not ( n14144 , RI1754c610_2);
and ( n14145 , n14144 , n44130 );
and ( n14146 , C0 , RI1754c610_2);
or ( n44131 , n14145 , n14146 );
buf ( n44132 , n44131 );
xor ( n44133 , n41414 , n43464 );
not ( n44134 , n34539 );
and ( n44135 , n44134 , n36818 );
xor ( n44136 , n34536 , n44135 );
xor ( n44137 , n34527 , n44136 );
not ( n44138 , n34549 );
and ( n44139 , n44138 , n36806 );
xor ( n44140 , n34546 , n44139 );
xor ( n44141 , n44137 , n44140 );
xor ( n44142 , n44141 , n43025 );
not ( n44143 , n34569 );
and ( n44144 , n44143 , n36838 );
xor ( n44145 , n34566 , n44144 );
xor ( n44146 , n44142 , n44145 );
xor ( n44147 , n44133 , n44146 );
xor ( n44148 , n41805 , n39262 );
xor ( n44149 , n44148 , n39282 );
not ( n44150 , n44149 );
xor ( n44151 , n35298 , n41990 );
xor ( n44152 , n44151 , n41005 );
and ( n44153 , n44150 , n44152 );
xor ( n44154 , n44147 , n44153 );
not ( n14147 , n29614 );
and ( n14148 , n14147 , RI1746b490_1213);
and ( n14149 , n44154 , n29614 );
or ( n44155 , n14148 , n14149 );
not ( n14150 , RI1754c610_2);
and ( n14151 , n14150 , n44155 );
and ( n14152 , C0 , RI1754c610_2);
or ( n44156 , n14151 , n14152 );
buf ( n44157 , n44156 );
xor ( n44158 , n40194 , n34041 );
xor ( n44159 , n44158 , n41934 );
xor ( n44160 , n39437 , n38495 );
xor ( n44161 , n44160 , n36611 );
not ( n44162 , n44161 );
xor ( n44163 , n41581 , n39065 );
xor ( n44164 , n44163 , n37331 );
and ( n44165 , n44162 , n44164 );
xor ( n44166 , n44159 , n44165 );
not ( n14153 , n29614 );
and ( n14154 , n14153 , RI17445240_1399);
and ( n14155 , n44166 , n29614 );
or ( n44167 , n14154 , n14155 );
not ( n14156 , RI1754c610_2);
and ( n14157 , n14156 , n44167 );
and ( n14158 , C0 , RI1754c610_2);
or ( n44168 , n14157 , n14158 );
buf ( n44169 , n44168 );
xor ( n44170 , n41210 , n39397 );
xor ( n44171 , n44170 , n39414 );
xor ( n44172 , n40301 , n37849 );
xor ( n44173 , n44172 , n37869 );
not ( n44174 , n44173 );
xor ( n44175 , n36622 , n40412 );
xor ( n44176 , n44175 , n40437 );
and ( n44177 , n44174 , n44176 );
xor ( n44178 , n44171 , n44177 );
not ( n14159 , n29614 );
and ( n14160 , n14159 , RI174ba3d8_831);
and ( n14161 , n44178 , n29614 );
or ( n44179 , n14160 , n14161 );
not ( n14162 , RI1754c610_2);
and ( n14163 , n14162 , n44179 );
and ( n14164 , C0 , RI1754c610_2);
or ( n44180 , n14163 , n14164 );
buf ( n44181 , n44180 );
xor ( n44182 , n38326 , n38872 );
xor ( n44183 , n44182 , n38886 );
xor ( n44184 , n37937 , n40210 );
xor ( n44185 , n44184 , n39989 );
not ( n44186 , n44185 );
and ( n44187 , n44186 , n40867 );
xor ( n44188 , n44183 , n44187 );
not ( n14165 , n29614 );
and ( n14166 , n14165 , RI17481a38_1104);
and ( n14167 , n44188 , n29614 );
or ( n44189 , n14166 , n14167 );
not ( n14168 , RI1754c610_2);
and ( n14169 , n14168 , n44189 );
and ( n14170 , C0 , RI1754c610_2);
or ( n44190 , n14169 , n14170 );
buf ( n44191 , n44190 );
xor ( n44192 , n38279 , n36568 );
xor ( n44193 , n44192 , n36742 );
not ( n44194 , n42201 );
and ( n44195 , n44194 , n42203 );
xor ( n44196 , n44193 , n44195 );
not ( n14171 , n29614 );
and ( n14172 , n14171 , RI17525ad8_649);
and ( n14173 , n44196 , n29614 );
or ( n44197 , n14172 , n14173 );
not ( n14174 , RI1754c610_2);
and ( n14175 , n14174 , n44197 );
and ( n14176 , C0 , RI1754c610_2);
or ( n44198 , n14175 , n14176 );
buf ( n44199 , n44198 );
xor ( n44200 , n38629 , n38347 );
xor ( n44201 , n44200 , n34300 );
xor ( n44202 , n33029 , n35639 );
xor ( n44203 , n44202 , n36227 );
not ( n44204 , n44203 );
xor ( n44205 , n34359 , n39989 );
xor ( n44206 , n44205 , n40009 );
and ( n44207 , n44204 , n44206 );
xor ( n44208 , n44201 , n44207 );
not ( n14177 , n29614 );
and ( n14178 , n14177 , RI174951f0_1009);
and ( n14179 , n44208 , n29614 );
or ( n44209 , n14178 , n14179 );
not ( n14180 , RI1754c610_2);
and ( n14181 , n14180 , n44209 );
and ( n14182 , C0 , RI1754c610_2);
or ( n44210 , n14181 , n14182 );
buf ( n44211 , n44210 );
not ( n44212 , n43242 );
xor ( n44213 , n36214 , n31831 );
xor ( n44214 , n44213 , n31925 );
and ( n44215 , n44212 , n44214 );
xor ( n44216 , n43239 , n44215 );
not ( n14183 , n29614 );
and ( n14184 , n14183 , RI174989b8_992);
and ( n14185 , n44216 , n29614 );
or ( n44217 , n14184 , n14185 );
not ( n14186 , RI1754c610_2);
and ( n14187 , n14186 , n44217 );
and ( n14188 , C0 , RI1754c610_2);
or ( n44218 , n14187 , n14188 );
buf ( n44219 , n44218 );
not ( n14189 , n27683 );
and ( n14190 , n14189 , RI19a97028_2633);
and ( n14191 , RI19aa0b50_2563 , n27683 );
or ( n44220 , n14190 , n14191 );
not ( n14192 , RI1754c610_2);
and ( n14193 , n14192 , n44220 );
and ( n14194 , C0 , RI1754c610_2);
or ( n44221 , n14193 , n14194 );
buf ( n44222 , n44221 );
xor ( n44223 , n36388 , n34190 );
xor ( n44224 , n44223 , n36252 );
xor ( n44225 , n34064 , n39525 );
xor ( n44226 , n44225 , n42377 );
not ( n44227 , n44226 );
xor ( n44228 , n41734 , n34837 );
xor ( n44229 , n44228 , n33880 );
and ( n44230 , n44227 , n44229 );
xor ( n44231 , n44224 , n44230 );
not ( n14195 , n29614 );
and ( n14196 , n14195 , RI1746d218_1204);
and ( n14197 , n44231 , n29614 );
or ( n44232 , n14196 , n14197 );
not ( n14198 , RI1754c610_2);
and ( n14199 , n14198 , n44232 );
and ( n14200 , C0 , RI1754c610_2);
or ( n44233 , n14199 , n14200 );
buf ( n44234 , n44233 );
not ( n44235 , n37491 );
xor ( n44236 , n35498 , n38532 );
xor ( n44237 , n44236 , n38933 );
and ( n44238 , n44235 , n44237 );
xor ( n44239 , n37440 , n44238 );
not ( n14201 , n29614 );
and ( n14202 , n14201 , RI173995e0_2008);
and ( n14203 , n44239 , n29614 );
or ( n44240 , n14202 , n14203 );
not ( n14204 , RI1754c610_2);
and ( n14205 , n14204 , n44240 );
and ( n14206 , C0 , RI1754c610_2);
or ( n44241 , n14205 , n14206 );
buf ( n44242 , n44241 );
xor ( n44243 , n37193 , n33030 );
xor ( n44244 , n44243 , n33069 );
not ( n44245 , n44244 );
xor ( n44246 , n41809 , n39262 );
xor ( n44247 , n44246 , n39282 );
and ( n44248 , n44245 , n44247 );
xor ( n44249 , n37267 , n44248 );
not ( n14207 , n29614 );
and ( n14208 , n14207 , RI173c8200_1780);
and ( n14209 , n44249 , n29614 );
or ( n44250 , n14208 , n14209 );
not ( n14210 , RI1754c610_2);
and ( n14211 , n14210 , n44250 );
and ( n14212 , C0 , RI1754c610_2);
or ( n44251 , n14211 , n14212 );
buf ( n44252 , n44251 );
not ( n14213 , n27683 );
and ( n14214 , n14213 , RI19abef88_2341);
and ( n14215 , RI19ac7f70_2270 , n27683 );
or ( n44253 , n14214 , n14215 );
not ( n14216 , RI1754c610_2);
and ( n14217 , n14216 , n44253 );
and ( n14218 , C0 , RI1754c610_2);
or ( n44254 , n14217 , n14218 );
buf ( n44255 , n44254 );
not ( n14219 , n27683 );
and ( n14220 , n14219 , RI19a82790_2777);
and ( n14221 , RI19aac388_2481 , n27683 );
or ( n44256 , n14220 , n14221 );
not ( n14222 , RI1754c610_2);
and ( n14223 , n14222 , n44256 );
and ( n14224 , C0 , RI1754c610_2);
or ( n44257 , n14223 , n14224 );
buf ( n44258 , n44257 );
not ( n44259 , n41827 );
and ( n44260 , n44259 , n41829 );
xor ( n44261 , n41100 , n44260 );
not ( n14225 , n29614 );
and ( n14226 , n14225 , RI173c7b70_1782);
and ( n14227 , n44261 , n29614 );
or ( n44262 , n14226 , n14227 );
not ( n14228 , RI1754c610_2);
and ( n14229 , n14228 , n44262 );
and ( n14230 , C0 , RI1754c610_2);
or ( n44263 , n14229 , n14230 );
buf ( n44264 , n44263 );
not ( n14231 , n27683 );
and ( n14232 , n14231 , RI19aa7c48_2511);
and ( n14233 , RI19ab1ba8_2441 , n27683 );
or ( n44265 , n14232 , n14233 );
not ( n14234 , RI1754c610_2);
and ( n14235 , n14234 , n44265 );
and ( n14236 , C0 , RI1754c610_2);
or ( n44266 , n14235 , n14236 );
buf ( n44267 , n44266 );
not ( n44268 , n36103 );
and ( n44269 , n44268 , n36288 );
xor ( n44270 , n36029 , n44269 );
not ( n14237 , n29614 );
and ( n14238 , n14237 , RI174a7c88_918);
and ( n14239 , n44270 , n29614 );
or ( n44271 , n14238 , n14239 );
not ( n14240 , RI1754c610_2);
and ( n14241 , n14240 , n44271 );
and ( n14242 , C0 , RI1754c610_2);
or ( n44272 , n14241 , n14242 );
buf ( n44273 , n44272 );
xor ( n44274 , n35930 , n36148 );
xor ( n44275 , n44274 , n37421 );
xor ( n44276 , n35994 , n35438 );
xor ( n44277 , n44276 , n35458 );
not ( n44278 , n44277 );
xor ( n44279 , n40509 , n41430 );
xor ( n44280 , n44279 , n36844 );
and ( n44281 , n44278 , n44280 );
xor ( n44282 , n44275 , n44281 );
not ( n14243 , n29614 );
and ( n14244 , n14243 , RI174b8650_837);
and ( n14245 , n44282 , n29614 );
or ( n44283 , n14244 , n14245 );
not ( n14246 , RI1754c610_2);
and ( n14247 , n14246 , n44283 );
and ( n14248 , C0 , RI1754c610_2);
or ( n44284 , n14247 , n14248 );
buf ( n44285 , n44284 );
xor ( n44286 , n35127 , n40283 );
xor ( n44287 , n44286 , n32560 );
not ( n44288 , n44287 );
xor ( n44289 , n39804 , n37800 );
xor ( n44290 , n44289 , n37814 );
and ( n44291 , n44288 , n44290 );
xor ( n44292 , n42973 , n44291 );
not ( n14249 , n29614 );
and ( n14250 , n14249 , RI174be1b8_819);
and ( n14251 , n44292 , n29614 );
or ( n44293 , n14250 , n14251 );
not ( n14252 , RI1754c610_2);
and ( n14253 , n14252 , n44293 );
and ( n14254 , C0 , RI1754c610_2);
or ( n44294 , n14253 , n14254 );
buf ( n44295 , n44294 );
not ( n14255 , n27683 );
and ( n14256 , n14255 , RI19a98f90_2619);
and ( n14257 , RI19aa27e8_2549 , n27683 );
or ( n44296 , n14256 , n14257 );
not ( n14258 , RI1754c610_2);
and ( n14259 , n14258 , n44296 );
and ( n14260 , C0 , RI1754c610_2);
or ( n44297 , n14259 , n14260 );
buf ( n44298 , n44297 );
not ( n14261 , n27683 );
and ( n14262 , n14261 , RI19ab5820_2412);
and ( n14263 , RI19abeda8_2342 , n27683 );
or ( n44299 , n14262 , n14263 );
not ( n14264 , RI1754c610_2);
and ( n14265 , n14264 , n44299 );
and ( n14266 , C0 , RI1754c610_2);
or ( n44300 , n14265 , n14266 );
buf ( n44301 , n44300 );
xor ( n44302 , n36190 , n32309 );
xor ( n44303 , n44302 , n32923 );
xor ( n44304 , n38932 , n42309 );
xor ( n44305 , n44304 , n43464 );
not ( n44306 , n44305 );
xor ( n44307 , n39530 , n35842 );
xor ( n44308 , n44307 , n38401 );
and ( n44309 , n44306 , n44308 );
xor ( n44310 , n44303 , n44309 );
not ( n14267 , n29614 );
and ( n14268 , n14267 , RI173fc6d0_1525);
and ( n14269 , n44310 , n29614 );
or ( n44311 , n14268 , n14269 );
not ( n14270 , RI1754c610_2);
and ( n14271 , n14270 , n44311 );
and ( n14272 , C0 , RI1754c610_2);
or ( n44312 , n14271 , n14272 );
buf ( n44313 , n44312 );
not ( n44314 , n36004 );
xor ( n44315 , n36946 , n32620 );
xor ( n44316 , n44315 , n33337 );
and ( n44317 , n44314 , n44316 );
xor ( n44318 , n35956 , n44317 );
not ( n14273 , n29614 );
and ( n14274 , n14273 , RI173a6498_1945);
and ( n14275 , n44318 , n29614 );
or ( n44319 , n14274 , n14275 );
not ( n14276 , RI1754c610_2);
and ( n14277 , n14276 , n44319 );
and ( n14278 , C0 , RI1754c610_2);
or ( n44320 , n14277 , n14278 );
buf ( n44321 , n44320 );
xor ( n44322 , n37330 , n39914 );
xor ( n44323 , n44322 , n40237 );
not ( n44324 , n44323 );
xor ( n44325 , n35236 , n39952 );
xor ( n44326 , n44325 , n42945 );
and ( n44327 , n44324 , n44326 );
xor ( n44328 , n43667 , n44327 );
not ( n14279 , n29614 );
and ( n14280 , n14279 , RI173b5420_1872);
and ( n14281 , n44328 , n29614 );
or ( n44329 , n14280 , n14281 );
not ( n14282 , RI1754c610_2);
and ( n14283 , n14282 , n44329 );
and ( n14284 , C0 , RI1754c610_2);
or ( n44330 , n14283 , n14284 );
buf ( n44331 , n44330 );
xor ( n44332 , n37715 , n40463 );
xor ( n44333 , n44332 , n41772 );
xor ( n44334 , n42172 , n41215 );
xor ( n44335 , n44334 , n33824 );
not ( n44336 , n44335 );
xor ( n44337 , n40733 , n31925 );
xor ( n44338 , n44337 , n34475 );
and ( n44339 , n44336 , n44338 );
xor ( n44340 , n44333 , n44339 );
not ( n14285 , n29614 );
and ( n14286 , n14285 , RI173c0f28_1815);
and ( n14287 , n44340 , n29614 );
or ( n44341 , n14286 , n14287 );
not ( n14288 , RI1754c610_2);
and ( n14289 , n14288 , n44341 );
and ( n14290 , C0 , RI1754c610_2);
or ( n44342 , n14289 , n14290 );
buf ( n44343 , n44342 );
buf ( n44344 , RI17467638_1232);
buf ( n44345 , RI1746f630_1193);
xor ( n44346 , n43476 , n32108 );
xor ( n44347 , n44346 , n38347 );
xor ( n44348 , n42938 , n29425 );
xor ( n44349 , n44348 , n29610 );
not ( n44350 , n44349 );
xor ( n44351 , n35399 , n41068 );
xor ( n44352 , n44351 , n39091 );
and ( n44353 , n44350 , n44352 );
xor ( n44354 , n44347 , n44353 );
not ( n14291 , n29614 );
and ( n14292 , n14291 , RI17359350_2090);
and ( n14293 , n44354 , n29614 );
or ( n44355 , n14292 , n14293 );
not ( n14294 , RI1754c610_2);
and ( n14295 , n14294 , n44355 );
and ( n14296 , C0 , RI1754c610_2);
or ( n44356 , n14295 , n14296 );
buf ( n44357 , n44356 );
not ( n44358 , n43111 );
and ( n44359 , n44358 , n43113 );
xor ( n44360 , n42556 , n44359 );
not ( n14297 , n29614 );
and ( n14298 , n14297 , RI173327a0_2195);
and ( n14299 , n44360 , n29614 );
or ( n44361 , n14298 , n14299 );
not ( n14300 , RI1754c610_2);
and ( n14301 , n14300 , n44361 );
and ( n14302 , C0 , RI1754c610_2);
or ( n44362 , n14301 , n14302 );
buf ( n44363 , n44362 );
not ( n14303 , n27683 );
and ( n14304 , n14303 , RI19aa48b8_2533);
and ( n14305 , RI19aaeb60_2463 , n27683 );
or ( n44364 , n14304 , n14305 );
not ( n14306 , RI1754c610_2);
and ( n14307 , n14306 , n44364 );
and ( n14308 , C0 , RI1754c610_2);
or ( n44365 , n14307 , n14308 );
buf ( n44366 , n44365 );
xor ( n44367 , n36085 , n37371 );
xor ( n44368 , n44367 , n36682 );
not ( n44369 , n42017 );
and ( n44370 , n44369 , n42035 );
xor ( n44371 , n44368 , n44370 );
not ( n14309 , n29614 );
and ( n14310 , n14309 , RI173ec398_1604);
and ( n14311 , n44371 , n29614 );
or ( n44372 , n14310 , n14311 );
not ( n14312 , RI1754c610_2);
and ( n14313 , n14312 , n44372 );
and ( n14314 , C0 , RI1754c610_2);
or ( n44373 , n14313 , n14314 );
buf ( n44374 , n44373 );
not ( n14315 , n27683 );
and ( n14316 , n14315 , RI19ac46b8_2296);
and ( n14317 , RI19acd358_2230 , n27683 );
or ( n44375 , n14316 , n14317 );
not ( n14318 , RI1754c610_2);
and ( n14319 , n14318 , n44375 );
and ( n14320 , C0 , RI1754c610_2);
or ( n44376 , n14319 , n14320 );
buf ( n44377 , n44376 );
xor ( n44378 , n38585 , n29109 );
xor ( n44379 , n44378 , n40463 );
not ( n44380 , n44379 );
xor ( n44381 , n36867 , n41198 );
xor ( n44382 , n44381 , n41215 );
and ( n44383 , n44380 , n44382 );
xor ( n44384 , n43916 , n44383 );
not ( n14321 , n29614 );
and ( n14322 , n14321 , RI173936b8_2037);
and ( n14323 , n44384 , n29614 );
or ( n44385 , n14322 , n14323 );
not ( n14324 , RI1754c610_2);
and ( n14325 , n14324 , n44385 );
and ( n14326 , C0 , RI1754c610_2);
or ( n44386 , n14325 , n14326 );
buf ( n44387 , n44386 );
xor ( n44388 , n36997 , n41818 );
xor ( n44389 , n44388 , n40662 );
xor ( n44390 , n31959 , n36682 );
xor ( n44391 , n44390 , n36702 );
not ( n44392 , n44391 );
xor ( n44393 , n39378 , n35594 );
xor ( n44394 , n44393 , n32403 );
and ( n44395 , n44392 , n44394 );
xor ( n44396 , n44389 , n44395 );
not ( n14327 , n29614 );
and ( n14328 , n14327 , RI173334c0_2191);
and ( n14329 , n44396 , n29614 );
or ( n44397 , n14328 , n14329 );
not ( n14330 , RI1754c610_2);
and ( n14331 , n14330 , n44397 );
and ( n14332 , C0 , RI1754c610_2);
or ( n44398 , n14331 , n14332 );
buf ( n44399 , n44398 );
not ( n14333 , n27683 );
and ( n14334 , n14333 , RI19aa8bc0_2505);
and ( n14335 , RI19ab2b98_2434 , n27683 );
or ( n44400 , n14334 , n14335 );
not ( n14336 , RI1754c610_2);
and ( n14337 , n14336 , n44400 );
and ( n14338 , C0 , RI1754c610_2);
or ( n44401 , n14337 , n14338 );
buf ( n44402 , n44401 );
buf ( n44403 , RI17492a90_1021);
buf ( n44404 , RI17481d80_1103);
buf ( n44405 , RI17510160_716);
buf ( n44406 , RI174c4e00_798);
xor ( n44407 , n37687 , n37579 );
xor ( n44408 , n44407 , n38495 );
xor ( n44409 , n41141 , n34087 );
xor ( n44410 , n44409 , n34127 );
not ( n44411 , n44410 );
and ( n44412 , n44411 , n41160 );
xor ( n44413 , n44408 , n44412 );
not ( n14339 , n29614 );
and ( n14340 , n14339 , RI173e6128_1634);
and ( n14341 , n44413 , n29614 );
or ( n44414 , n14340 , n14341 );
not ( n14342 , RI1754c610_2);
and ( n14343 , n14342 , n44414 );
and ( n14344 , C0 , RI1754c610_2);
or ( n44415 , n14343 , n14344 );
buf ( n44416 , n44415 );
not ( n44417 , n42683 );
xor ( n44418 , n35024 , n37814 );
xor ( n44419 , n44418 , n33223 );
and ( n44420 , n44417 , n44419 );
xor ( n44421 , n42680 , n44420 );
not ( n14345 , n29614 );
and ( n14346 , n14345 , RI173fa600_1535);
and ( n14347 , n44421 , n29614 );
or ( n44422 , n14346 , n14347 );
not ( n14348 , RI1754c610_2);
and ( n14349 , n14348 , n44422 );
and ( n14350 , C0 , RI1754c610_2);
or ( n44423 , n14349 , n14350 );
buf ( n44424 , n44423 );
not ( n44425 , n42556 );
and ( n44426 , n44425 , n43111 );
xor ( n44427 , n42534 , n44426 );
not ( n14351 , n29614 );
and ( n14352 , n14351 , RI1751f8e0_668);
and ( n14353 , n44427 , n29614 );
or ( n44428 , n14352 , n14353 );
not ( n14354 , RI1754c610_2);
and ( n14355 , n14354 , n44428 );
and ( n14356 , C0 , RI1754c610_2);
or ( n44429 , n14355 , n14356 );
buf ( n44430 , n44429 );
xor ( n44431 , n35000 , n42945 );
xor ( n44432 , n44431 , n34497 );
xor ( n44433 , n33504 , n40360 );
xor ( n44434 , n44433 , n35176 );
not ( n44435 , n44434 );
xor ( n44436 , n41085 , n38150 );
xor ( n44437 , n44436 , n38167 );
and ( n44438 , n44435 , n44437 );
xor ( n44439 , n44432 , n44438 );
not ( n14357 , n29614 );
and ( n14358 , n14357 , RI17496258_1004);
and ( n14359 , n44439 , n29614 );
or ( n44440 , n14358 , n14359 );
not ( n14360 , RI1754c610_2);
and ( n14361 , n14360 , n44440 );
and ( n14362 , C0 , RI1754c610_2);
or ( n44441 , n14361 , n14362 );
buf ( n44442 , n44441 );
not ( n14363 , n27683 );
and ( n14364 , n14363 , RI19a96038_2640);
and ( n14365 , RI19a9ff20_2569 , n27683 );
or ( n44443 , n14364 , n14365 );
not ( n14366 , RI1754c610_2);
and ( n14367 , n14366 , n44443 );
and ( n14368 , C0 , RI1754c610_2);
or ( n44444 , n14367 , n14368 );
buf ( n44445 , n44444 );
xor ( n44446 , n36741 , n30247 );
xor ( n44447 , n44446 , n30461 );
xor ( n44448 , n34456 , n33453 );
xor ( n44449 , n44448 , n33505 );
not ( n44450 , n44449 );
xor ( n44451 , n40550 , n40966 );
xor ( n44452 , n44451 , n37460 );
and ( n44453 , n44450 , n44452 );
xor ( n44454 , n44447 , n44453 );
not ( n14369 , n29614 );
and ( n14370 , n14369 , RI17332e30_2193);
and ( n14371 , n44454 , n29614 );
or ( n44455 , n14370 , n14371 );
not ( n14372 , RI1754c610_2);
and ( n14373 , n14372 , n44455 );
and ( n14374 , C0 , RI1754c610_2);
or ( n44456 , n14373 , n14374 );
buf ( n44457 , n44456 );
xor ( n44458 , n38258 , n36530 );
xor ( n44459 , n44458 , n36568 );
xor ( n44460 , n34748 , n42619 );
xor ( n44461 , n44460 , n41990 );
not ( n44462 , n44461 );
xor ( n44463 , n42187 , n41215 );
xor ( n44464 , n44463 , n33824 );
and ( n44465 , n44462 , n44464 );
xor ( n44466 , n44459 , n44465 );
not ( n14375 , n29614 );
and ( n14376 , n14375 , RI17480d18_1108);
and ( n14377 , n44466 , n29614 );
or ( n44467 , n14376 , n14377 );
not ( n14378 , RI1754c610_2);
and ( n14379 , n14378 , n44467 );
and ( n14380 , C0 , RI1754c610_2);
or ( n44468 , n14379 , n14380 );
buf ( n44469 , n44468 );
xor ( n44470 , n39045 , n39702 );
xor ( n44471 , n44470 , n39914 );
xor ( n44472 , n41646 , n40692 );
xor ( n44473 , n44472 , n43994 );
not ( n44474 , n44473 );
xor ( n44475 , n36221 , n31831 );
xor ( n44476 , n44475 , n31925 );
and ( n44477 , n44474 , n44476 );
xor ( n44478 , n44471 , n44477 );
not ( n14381 , n29614 );
and ( n14382 , n14381 , RI174b4e88_854);
and ( n14383 , n44478 , n29614 );
or ( n44479 , n14382 , n14383 );
not ( n14384 , RI1754c610_2);
and ( n14385 , n14384 , n44479 );
and ( n14386 , C0 , RI1754c610_2);
or ( n44480 , n14385 , n14386 );
buf ( n44481 , n44480 );
xor ( n44482 , n37864 , n35128 );
xor ( n44483 , n44482 , n36917 );
not ( n44484 , n34671 );
and ( n44485 , n44484 , n34756 );
xor ( n44486 , n44483 , n44485 );
not ( n14387 , n29614 );
and ( n14388 , n14387 , RI173fe110_1517);
and ( n14389 , n44486 , n29614 );
or ( n44487 , n14388 , n14389 );
not ( n14390 , RI1754c610_2);
and ( n14391 , n14390 , n44487 );
and ( n14392 , C0 , RI1754c610_2);
or ( n44488 , n14391 , n14392 );
buf ( n44489 , n44488 );
not ( n14393 , n27683 );
and ( n14394 , n14393 , RI19aa9d90_2497);
and ( n14395 , RI19ab3840_2427 , n27683 );
or ( n44490 , n14394 , n14395 );
not ( n14396 , RI1754c610_2);
and ( n14397 , n14396 , n44490 );
and ( n14398 , C0 , RI1754c610_2);
or ( n44491 , n14397 , n14398 );
buf ( n44492 , n44491 );
buf ( n44493 , RI174a9a10_909);
buf ( n44494 , RI17497c98_996);
buf ( n44495 , RI1747fff8_1112);
buf ( n44496 , RI17471a48_1182);
buf ( n44497 , RI1746e280_1199);
buf ( n44498 , RI175134f0_706);
not ( n44499 , n42825 );
xor ( n44500 , n39786 , n33175 );
xor ( n44501 , n44500 , n34797 );
and ( n44502 , n44499 , n44501 );
xor ( n44503 , n42822 , n44502 );
not ( n14399 , n29614 );
and ( n14400 , n14399 , RI17471a48_1182);
and ( n14401 , n44503 , n29614 );
or ( n44504 , n14400 , n14401 );
not ( n14402 , RI1754c610_2);
and ( n14403 , n14402 , n44504 );
and ( n14404 , C0 , RI1754c610_2);
or ( n44505 , n14403 , n14404 );
buf ( n44506 , n44505 );
buf ( n44507 , RI174bcd18_823);
not ( n14405 , n27683 );
and ( n14406 , n14405 , RI19a91e98_2669);
and ( n14407 , RI19a9bfd8_2598 , n27683 );
or ( n44508 , n14406 , n14407 );
not ( n14408 , RI1754c610_2);
and ( n14409 , n14408 , n44508 );
and ( n14410 , C0 , RI1754c610_2);
or ( n44509 , n14409 , n14410 );
buf ( n44510 , n44509 );
buf ( n44511 , RI174ad1d8_892);
buf ( n44512 , RI17465568_1242);
xor ( n44513 , n39445 , n38495 );
xor ( n44514 , n44513 , n36611 );
xor ( n44515 , n37437 , n34725 );
xor ( n44516 , n44515 , n34755 );
not ( n44517 , n44516 );
and ( n44518 , n44517 , n40726 );
xor ( n44519 , n44514 , n44518 );
not ( n14411 , n29614 );
and ( n14412 , n14411 , RI1748ec38_1040);
and ( n14413 , n44519 , n29614 );
or ( n44520 , n14412 , n14413 );
not ( n14414 , RI1754c610_2);
and ( n14415 , n14414 , n44520 );
and ( n14416 , C0 , RI1754c610_2);
or ( n44521 , n14415 , n14416 );
buf ( n44522 , n44521 );
xor ( n44523 , n33767 , n40486 );
xor ( n44524 , n44523 , n40516 );
xor ( n44525 , n40411 , n32973 );
xor ( n44526 , n44525 , n39816 );
not ( n44527 , n44526 );
xor ( n44528 , n36439 , n37104 );
xor ( n44529 , n44528 , n35986 );
and ( n44530 , n44527 , n44529 );
xor ( n44531 , n44524 , n44530 );
not ( n14417 , n29614 );
and ( n14418 , n14417 , RI174b09a0_875);
and ( n14419 , n44531 , n29614 );
or ( n44532 , n14418 , n14419 );
not ( n14420 , RI1754c610_2);
and ( n14421 , n14420 , n44532 );
and ( n14422 , C0 , RI1754c610_2);
or ( n44533 , n14421 , n14422 );
buf ( n44534 , n44533 );
xor ( n44535 , n33596 , n41740 );
xor ( n44536 , n44535 , n38371 );
not ( n44537 , n38402 );
and ( n44538 , n44537 , n38446 );
xor ( n44539 , n44536 , n44538 );
not ( n14423 , n29614 );
and ( n14424 , n14423 , RI1739a990_2002);
and ( n14425 , n44539 , n29614 );
or ( n44540 , n14424 , n14425 );
not ( n14426 , RI1754c610_2);
and ( n14427 , n14426 , n44540 );
and ( n14428 , C0 , RI1754c610_2);
or ( n44541 , n14427 , n14428 );
buf ( n44542 , n44541 );
not ( n14429 , n27683 );
and ( n14430 , n14429 , RI19aced20_2219);
and ( n14431 , RI19a9cc08_2592 , n27683 );
or ( n44543 , n14430 , n14431 );
not ( n14432 , RI1754c610_2);
and ( n14433 , n14432 , n44543 );
and ( n14434 , C0 , RI1754c610_2);
or ( n44544 , n14433 , n14434 );
buf ( n44545 , n44544 );
xor ( n44546 , n37764 , n43994 );
xor ( n44547 , n44546 , n31213 );
not ( n44548 , n44547 );
xor ( n44549 , n32528 , n37651 );
xor ( n44550 , n44549 , n39182 );
and ( n44551 , n44548 , n44550 );
xor ( n44552 , n42915 , n44551 );
not ( n14435 , n29614 );
and ( n14436 , n14435 , RI173b7838_1861);
and ( n14437 , n44552 , n29614 );
or ( n44553 , n14436 , n14437 );
not ( n14438 , RI1754c610_2);
and ( n14439 , n14438 , n44553 );
and ( n14440 , C0 , RI1754c610_2);
or ( n44554 , n14439 , n14440 );
buf ( n44555 , n44554 );
xor ( n44556 , n39735 , n39506 );
xor ( n44557 , n44556 , n38150 );
xor ( n44558 , n38370 , n33880 );
xor ( n44559 , n44558 , n33935 );
not ( n44560 , n44559 );
and ( n44561 , n44560 , n28469 );
xor ( n44562 , n44557 , n44561 );
not ( n14441 , n29614 );
and ( n14442 , n14441 , RI17491398_1028);
and ( n14443 , n44562 , n29614 );
or ( n44563 , n14442 , n14443 );
not ( n14444 , RI1754c610_2);
and ( n14445 , n14444 , n44563 );
and ( n14446 , C0 , RI1754c610_2);
or ( n44564 , n14445 , n14446 );
buf ( n44565 , n44564 );
not ( n14447 , n27683 );
and ( n14448 , n14447 , RI19a8f8a0_2686);
and ( n14449 , RI19a998f0_2615 , n27683 );
or ( n44566 , n14448 , n14449 );
not ( n14450 , RI1754c610_2);
and ( n14451 , n14450 , n44566 );
and ( n14452 , C0 , RI1754c610_2);
or ( n44567 , n14451 , n14452 );
buf ( n44568 , n44567 );
xor ( n44569 , n34668 , n32863 );
xor ( n44570 , n44569 , n34644 );
xor ( n44571 , n36345 , n38676 );
xor ( n44572 , n44571 , n28111 );
not ( n44573 , n44572 );
xor ( n44574 , n37600 , n40319 );
xor ( n44575 , n44574 , n40149 );
and ( n44576 , n44573 , n44575 );
xor ( n44577 , n44570 , n44576 );
not ( n14453 , n29614 );
and ( n14454 , n14453 , RI173393e8_2162);
and ( n14455 , n44577 , n29614 );
or ( n44578 , n14454 , n14455 );
not ( n14456 , RI1754c610_2);
and ( n14457 , n14456 , n44578 );
and ( n14458 , C0 , RI1754c610_2);
or ( n44579 , n14457 , n14458 );
buf ( n44580 , n44579 );
xor ( n44581 , n34232 , n37526 );
xor ( n44582 , n44581 , n41049 );
not ( n44583 , n44582 );
xor ( n44584 , n35107 , n40283 );
xor ( n44585 , n44584 , n32560 );
and ( n44586 , n44583 , n44585 );
xor ( n44587 , n40260 , n44586 );
not ( n14459 , n29614 );
and ( n14460 , n14459 , RI173c4d80_1796);
and ( n14461 , n44587 , n29614 );
or ( n44588 , n14460 , n14461 );
not ( n14462 , RI1754c610_2);
and ( n14463 , n14462 , n44588 );
and ( n14464 , C0 , RI1754c610_2);
or ( n44589 , n14463 , n14464 );
buf ( n44590 , n44589 );
xor ( n44591 , n40716 , n39333 );
xor ( n44592 , n44591 , n39347 );
not ( n44593 , n44592 );
and ( n44594 , n44593 , n43004 );
xor ( n44595 , n42362 , n44594 );
not ( n14465 , n29614 );
and ( n14466 , n14465 , RI17473140_1175);
and ( n14467 , n44595 , n29614 );
or ( n44596 , n14466 , n14467 );
not ( n14468 , RI1754c610_2);
and ( n14469 , n14468 , n44596 );
and ( n14470 , C0 , RI1754c610_2);
or ( n44597 , n14469 , n14470 );
buf ( n44598 , n44597 );
xor ( n44599 , n33062 , n36227 );
xor ( n44600 , n44599 , n40743 );
not ( n44601 , n44600 );
xor ( n44602 , n38552 , n35458 );
xor ( n44603 , n44602 , n40692 );
and ( n44604 , n44601 , n44603 );
xor ( n44605 , n37652 , n44604 );
not ( n14471 , n29614 );
and ( n14472 , n14471 , RI17500a58_758);
and ( n14473 , n44605 , n29614 );
or ( n44606 , n14472 , n14473 );
not ( n14474 , RI1754c610_2);
and ( n14475 , n14474 , n44606 );
and ( n14476 , C0 , RI1754c610_2);
or ( n44607 , n14475 , n14476 );
buf ( n44608 , n44607 );
not ( n14477 , n27683 );
and ( n14478 , n14477 , RI19ab36d8_2428);
and ( n14479 , RI19abd4d0_2356 , n27683 );
or ( n44609 , n14478 , n14479 );
not ( n14480 , RI1754c610_2);
and ( n14481 , n14480 , n44609 );
and ( n14482 , C0 , RI1754c610_2);
or ( n44610 , n14481 , n14482 );
buf ( n44611 , n44610 );
xor ( n44612 , n38149 , n31053 );
xor ( n44613 , n44612 , n35494 );
xor ( n44614 , n39195 , n37676 );
xor ( n44615 , n44614 , n37696 );
not ( n44616 , n44615 );
xor ( n44617 , n40815 , n42635 );
xor ( n44618 , n44617 , n33648 );
and ( n44619 , n44616 , n44618 );
xor ( n44620 , n44613 , n44619 );
not ( n14483 , n29614 );
and ( n14484 , n14483 , RI174a16d0_949);
and ( n14485 , n44620 , n29614 );
or ( n44621 , n14484 , n14485 );
not ( n14486 , RI1754c610_2);
and ( n14487 , n14486 , n44621 );
and ( n14488 , C0 , RI1754c610_2);
or ( n44622 , n14487 , n14488 );
buf ( n44623 , n44622 );
xor ( n44624 , n36217 , n31831 );
xor ( n44625 , n44624 , n31925 );
xor ( n44626 , n38428 , n40585 );
xor ( n44627 , n44626 , n34918 );
not ( n44628 , n44627 );
and ( n44629 , n44628 , n33618 );
xor ( n44630 , n44625 , n44629 );
not ( n14489 , n29614 );
and ( n14490 , n14489 , RI173d71a0_1707);
and ( n14491 , n44630 , n29614 );
or ( n44631 , n14490 , n14491 );
not ( n14492 , RI1754c610_2);
and ( n14493 , n14492 , n44631 );
and ( n14494 , C0 , RI1754c610_2);
or ( n44632 , n14493 , n14494 );
buf ( n44633 , n44632 );
and ( n44634 , RI19a24578_2786 , n43086 );
not ( n14495 , n43088 );
and ( n14496 , n14495 , RI19a24320_2787);
and ( n14497 , n44634 , n43088 );
or ( n44635 , n14496 , n14497 );
not ( n14498 , RI1754c610_2);
and ( n14499 , n14498 , n44635 );
and ( n14500 , C0 , RI1754c610_2);
or ( n44636 , n14499 , n14500 );
buf ( n44637 , n44636 );
not ( n44638 , n42728 );
and ( n44639 , n44638 , n43047 );
xor ( n44640 , n42725 , n44639 );
not ( n14501 , n29614 );
and ( n14502 , n14501 , RI174506b8_1344);
and ( n14503 , n44640 , n29614 );
or ( n44641 , n14502 , n14503 );
not ( n14504 , RI1754c610_2);
and ( n14505 , n14504 , n44641 );
and ( n14506 , C0 , RI1754c610_2);
or ( n44642 , n14505 , n14506 );
buf ( n44643 , n44642 );
xor ( n44644 , n41613 , n43278 );
xor ( n44645 , n44644 , n31664 );
xor ( n44646 , n42342 , n29981 );
xor ( n44647 , n44646 , n35955 );
not ( n44648 , n44647 );
and ( n44649 , n44648 , n40839 );
xor ( n44650 , n44645 , n44649 );
not ( n14507 , n29614 );
and ( n14508 , n14507 , RI1748c4d8_1052);
and ( n14509 , n44650 , n29614 );
or ( n44651 , n14508 , n14509 );
not ( n14510 , RI1754c610_2);
and ( n14511 , n14510 , n44651 );
and ( n14512 , C0 , RI1754c610_2);
or ( n44652 , n14511 , n14512 );
buf ( n44653 , n44652 );
buf ( n44654 , RI17478348_1150);
not ( n44655 , n43494 );
and ( n44656 , n44655 , n43496 );
xor ( n44657 , n44087 , n44656 );
not ( n14513 , n29614 );
and ( n14514 , n14513 , RI173e46e8_1642);
and ( n14515 , n44657 , n29614 );
or ( n44658 , n14514 , n14515 );
not ( n14516 , RI1754c610_2);
and ( n14517 , n14516 , n44658 );
and ( n14518 , C0 , RI1754c610_2);
or ( n44659 , n14517 , n14518 );
buf ( n44660 , n44659 );
xor ( n44661 , n41390 , n33567 );
xor ( n44662 , n44661 , n33617 );
not ( n44663 , n44662 );
xor ( n44664 , n34979 , n42945 );
xor ( n44665 , n44664 , n34497 );
and ( n44666 , n44663 , n44665 );
xor ( n44667 , n40070 , n44666 );
not ( n14519 , n29614 );
and ( n14520 , n14519 , RI17523198_657);
and ( n14521 , n44667 , n29614 );
or ( n44668 , n14520 , n14521 );
not ( n14522 , RI1754c610_2);
and ( n14523 , n14522 , n44668 );
and ( n14524 , C0 , RI1754c610_2);
or ( n44669 , n14523 , n14524 );
buf ( n44670 , n44669 );
buf ( n44671 , RI174972c0_999);
buf ( n44672 , RI1748be48_1054);
buf ( n44673 , RI174cf300_766);
not ( n14525 , n27683 );
and ( n14526 , n14525 , RI19a852b0_2758);
and ( n14527 , RI19ac6878_2281 , n27683 );
or ( n44674 , n14526 , n14527 );
not ( n14528 , RI1754c610_2);
and ( n14529 , n14528 , n44674 );
and ( n14530 , C0 , RI1754c610_2);
or ( n44675 , n14529 , n14530 );
buf ( n44676 , n44675 );
buf ( n44677 , RI174c3960_802);
not ( n14531 , n27683 );
and ( n14532 , n14531 , RI19abfd98_2333);
and ( n14533 , RI19ac8e70_2263 , n27683 );
or ( n44678 , n14532 , n14533 );
not ( n14534 , RI1754c610_2);
and ( n14535 , n14534 , n44678 );
and ( n14536 , C0 , RI1754c610_2);
or ( n44679 , n14535 , n14536 );
buf ( n44680 , n44679 );
not ( n14537 , n27683 );
and ( n14538 , n14537 , RI19a95b88_2642);
and ( n14539 , RI19a9f908_2572 , n27683 );
or ( n44681 , n14538 , n14539 );
not ( n14540 , RI1754c610_2);
and ( n14541 , n14540 , n44681 );
and ( n14542 , C0 , RI1754c610_2);
or ( n44682 , n14541 , n14542 );
buf ( n44683 , n44682 );
xor ( n44684 , n33301 , n38991 );
xor ( n44685 , n44684 , n39005 );
xor ( n44686 , n38663 , n39347 );
xor ( n44687 , n44686 , n42344 );
not ( n44688 , n44687 );
xor ( n44689 , n41925 , n42033 );
xor ( n44690 , n44689 , n37987 );
and ( n44691 , n44688 , n44690 );
xor ( n44692 , n44685 , n44691 );
not ( n14543 , n29614 );
and ( n14544 , n14543 , RI1733e2a8_2138);
and ( n14545 , n44692 , n29614 );
or ( n44693 , n14544 , n14545 );
not ( n14546 , RI1754c610_2);
and ( n14547 , n14546 , n44693 );
and ( n14548 , C0 , RI1754c610_2);
or ( n44694 , n14547 , n14548 );
buf ( n44695 , n44694 );
not ( n44696 , n37341 );
xor ( n44697 , n40358 , n37898 );
xor ( n44698 , n44697 , n37915 );
and ( n44699 , n44696 , n44698 );
xor ( n44700 , n37333 , n44699 );
not ( n14549 , n29614 );
and ( n14550 , n14549 , RI174772e0_1155);
and ( n14551 , n44700 , n29614 );
or ( n44701 , n14550 , n14551 );
not ( n14552 , RI1754c610_2);
and ( n14553 , n14552 , n44701 );
and ( n14554 , C0 , RI1754c610_2);
or ( n44702 , n14553 , n14554 );
buf ( n44703 , n44702 );
not ( n44704 , n42510 );
xor ( n44705 , n43269 , n41099 );
xor ( n44706 , n44705 , n30604 );
and ( n44707 , n44704 , n44706 );
xor ( n44708 , n42507 , n44707 );
not ( n14555 , n29614 );
and ( n14556 , n14555 , RI173cbd10_1762);
and ( n14557 , n44708 , n29614 );
or ( n44709 , n14556 , n14557 );
not ( n14558 , RI1754c610_2);
and ( n14559 , n14558 , n44709 );
and ( n14560 , C0 , RI1754c610_2);
or ( n44710 , n14559 , n14560 );
buf ( n44711 , n44710 );
not ( n44712 , n43426 );
xor ( n44713 , n43991 , n40808 );
xor ( n44714 , n44713 , n40828 );
and ( n44715 , n44712 , n44714 );
xor ( n44716 , n43423 , n44715 );
not ( n14561 , n29614 );
and ( n14562 , n14561 , RI174aaa78_904);
and ( n14563 , n44716 , n29614 );
or ( n44717 , n14562 , n14563 );
not ( n14564 , RI1754c610_2);
and ( n14565 , n14564 , n44717 );
and ( n14566 , C0 , RI1754c610_2);
or ( n44718 , n14565 , n14566 );
buf ( n44719 , n44718 );
not ( n44720 , n38373 );
xor ( n44721 , n37644 , n40149 );
xor ( n44722 , n44721 , n40166 );
and ( n44723 , n44720 , n44722 );
xor ( n44724 , n38351 , n44723 );
not ( n14567 , n29614 );
and ( n14568 , n14567 , RI174c3438_803);
and ( n14569 , n44724 , n29614 );
or ( n44725 , n14568 , n14569 );
not ( n14570 , RI1754c610_2);
and ( n14571 , n14570 , n44725 );
and ( n14572 , C0 , RI1754c610_2);
or ( n44726 , n14571 , n14572 );
buf ( n44727 , n44726 );
xor ( n44728 , n41090 , n38150 );
xor ( n44729 , n44728 , n38167 );
xor ( n44730 , n40231 , n35710 );
xor ( n44731 , n44730 , n35760 );
not ( n44732 , n44731 );
and ( n44733 , n44732 , n42788 );
xor ( n44734 , n44729 , n44733 );
not ( n14573 , n29614 );
and ( n14574 , n14573 , RI173d46f8_1720);
and ( n14575 , n44734 , n29614 );
or ( n44735 , n14574 , n14575 );
not ( n14576 , RI1754c610_2);
and ( n14577 , n14576 , n44735 );
and ( n14578 , C0 , RI1754c610_2);
or ( n44736 , n14577 , n14578 );
buf ( n44737 , n44736 );
xor ( n44738 , n34492 , n29610 );
xor ( n44739 , n44738 , n31380 );
not ( n44740 , n35129 );
and ( n44741 , n44740 , n35217 );
xor ( n44742 , n44739 , n44741 );
not ( n14579 , n29614 );
and ( n14580 , n14579 , RI173b4070_1878);
and ( n14581 , n44742 , n29614 );
or ( n44743 , n14580 , n14581 );
not ( n14582 , RI1754c610_2);
and ( n14583 , n14582 , n44743 );
and ( n14584 , C0 , RI1754c610_2);
or ( n44744 , n14583 , n14584 );
buf ( n44745 , n44744 );
xor ( n44746 , n35583 , n37490 );
xor ( n44747 , n44746 , n41316 );
not ( n44748 , n44613 );
and ( n44749 , n44748 , n44615 );
xor ( n44750 , n44747 , n44749 );
not ( n14585 , n29614 );
and ( n14586 , n14585 , RI17492dd8_1020);
and ( n14587 , n44750 , n29614 );
or ( n44751 , n14586 , n14587 );
not ( n14588 , RI1754c610_2);
and ( n14589 , n14588 , n44751 );
and ( n14590 , C0 , RI1754c610_2);
or ( n44752 , n14589 , n14590 );
buf ( n44753 , n44752 );
xor ( n44754 , n39118 , n28111 );
xor ( n44755 , n44754 , n28468 );
xor ( n44756 , n43483 , n32108 );
xor ( n44757 , n44756 , n38347 );
not ( n44758 , n44757 );
xor ( n44759 , n42943 , n29425 );
xor ( n44760 , n44759 , n29610 );
and ( n44761 , n44758 , n44760 );
xor ( n44762 , n44755 , n44761 );
not ( n14591 , n29614 );
and ( n14592 , n14591 , RI173de130_1673);
and ( n14593 , n44762 , n29614 );
or ( n44763 , n14592 , n14593 );
not ( n14594 , RI1754c610_2);
and ( n14595 , n14594 , n44763 );
and ( n14596 , C0 , RI1754c610_2);
or ( n44764 , n14595 , n14596 );
buf ( n44765 , n44764 );
and ( n44766 , RI1754b5a8_37 , n34844 );
and ( n44767 , RI1754b5a8_37 , n34847 );
and ( n44768 , RI1754b5a8_37 , n34850 );
or ( n44769 , n44766 , n44767 , n44768 , C0 , C0 , C0 , C0 , C0 );
not ( n14597 , n34859 );
and ( n14598 , n14597 , n44769 );
and ( n14599 , RI1754b5a8_37 , n34859 );
or ( n44770 , n14598 , n14599 );
not ( n14600 , RI19a22f70_2797);
and ( n14601 , n14600 , n44770 );
and ( n14602 , C0 , RI19a22f70_2797);
or ( n44771 , n14601 , n14602 );
not ( n14603 , n27683 );
and ( n14604 , n14603 , RI19ab3c00_2425);
and ( n14605 , n44771 , n27683 );
or ( n44772 , n14604 , n14605 );
not ( n14606 , RI1754c610_2);
and ( n14607 , n14606 , n44772 );
and ( n14608 , C0 , RI1754c610_2);
or ( n44773 , n14607 , n14608 );
buf ( n44774 , n44773 );
not ( n14609 , n27683 );
and ( n14610 , n14609 , RI19a85e68_2753);
and ( n14611 , RI19a23858_2792 , n27683 );
or ( n44775 , n14610 , n14611 );
not ( n14612 , RI1754c610_2);
and ( n14613 , n14612 , n44775 );
and ( n14614 , C0 , RI1754c610_2);
or ( n44776 , n14613 , n14614 );
buf ( n44777 , n44776 );
xor ( n44778 , n36093 , n37371 );
xor ( n44779 , n44778 , n36682 );
xor ( n44780 , n31212 , n40828 );
xor ( n44781 , n44780 , n42049 );
not ( n44782 , n44781 );
xor ( n44783 , n41488 , n34445 );
xor ( n44784 , n44783 , n41885 );
and ( n44785 , n44782 , n44784 );
xor ( n44786 , n44779 , n44785 );
not ( n14615 , n29614 );
and ( n14616 , n14615 , RI1751ab88_683);
and ( n14617 , n44786 , n29614 );
or ( n44787 , n14616 , n14617 );
not ( n14618 , RI1754c610_2);
and ( n14619 , n14618 , n44787 );
and ( n14620 , C0 , RI1754c610_2);
or ( n44788 , n14619 , n14620 );
buf ( n44789 , n44788 );
xor ( n44790 , n35261 , n39952 );
xor ( n44791 , n44790 , n42945 );
not ( n44792 , n43447 );
and ( n44793 , n44792 , n43465 );
xor ( n44794 , n44791 , n44793 );
not ( n14621 , n29614 );
and ( n14622 , n14621 , RI1751ca78_677);
and ( n14623 , n44794 , n29614 );
or ( n44795 , n14622 , n14623 );
not ( n14624 , RI1754c610_2);
and ( n14625 , n14624 , n44795 );
and ( n14626 , C0 , RI1754c610_2);
or ( n44796 , n14625 , n14626 );
buf ( n44797 , n44796 );
xor ( n44798 , n36418 , n33935 );
xor ( n44799 , n44798 , n36287 );
not ( n44800 , n44799 );
xor ( n44801 , n40081 , n38037 );
xor ( n44802 , n44801 , n39740 );
and ( n44803 , n44800 , n44802 );
xor ( n44804 , n39307 , n44803 );
not ( n14627 , n29614 );
and ( n14628 , n14627 , RI173bdaa8_1831);
and ( n14629 , n44804 , n29614 );
or ( n44805 , n14628 , n14629 );
not ( n14630 , RI1754c610_2);
and ( n14631 , n14630 , n44805 );
and ( n14632 , C0 , RI1754c610_2);
or ( n44806 , n14631 , n14632 );
buf ( n44807 , n44806 );
xor ( n44808 , n33738 , n40486 );
xor ( n44809 , n44808 , n40516 );
xor ( n44810 , n41977 , n39886 );
xor ( n44811 , n44810 , n36998 );
not ( n44812 , n44811 );
and ( n44813 , n44812 , n38602 );
xor ( n44814 , n44809 , n44813 );
not ( n14633 , n29614 );
and ( n14634 , n14633 , RI1746b148_1214);
and ( n14635 , n44814 , n29614 );
or ( n44815 , n14634 , n14635 );
not ( n14636 , RI1754c610_2);
and ( n14637 , n14636 , n44815 );
and ( n14638 , C0 , RI1754c610_2);
or ( n44816 , n14637 , n14638 );
buf ( n44817 , n44816 );
not ( n14639 , n27683 );
and ( n14640 , n14639 , RI19a91100_2675);
and ( n14641 , RI19a9b1c8_2604 , n27683 );
or ( n44818 , n14640 , n14641 );
not ( n14642 , RI1754c610_2);
and ( n14643 , n14642 , n44818 );
and ( n14644 , C0 , RI1754c610_2);
or ( n44819 , n14643 , n14644 );
buf ( n44820 , n44819 );
not ( n14645 , n27683 );
and ( n14646 , n14645 , RI19ac40a0_2299);
and ( n14647 , RI19accc50_2233 , n27683 );
or ( n44821 , n14646 , n14647 );
not ( n14648 , RI1754c610_2);
and ( n14649 , n14648 , n44821 );
and ( n14650 , C0 , RI1754c610_2);
or ( n44822 , n14649 , n14650 );
buf ( n44823 , n44822 );
not ( n14651 , n27683 );
and ( n14652 , n14651 , RI19a9d400_2589);
and ( n14653 , RI19aa6b68_2518 , n27683 );
or ( n44824 , n14652 , n14653 );
not ( n14654 , RI1754c610_2);
and ( n14655 , n14654 , n44824 );
and ( n14656 , C0 , RI1754c610_2);
or ( n44825 , n14655 , n14656 );
buf ( n44826 , n44825 );
not ( n14657 , n27683 );
and ( n14658 , n14657 , RI19a952a0_2646);
and ( n14659 , RI19a9f188_2576 , n27683 );
or ( n44827 , n14658 , n14659 );
not ( n14660 , RI1754c610_2);
and ( n14661 , n14660 , n44827 );
and ( n14662 , C0 , RI1754c610_2);
or ( n44828 , n14661 , n14662 );
buf ( n44829 , n44828 );
xor ( n44830 , n32012 , n36682 );
xor ( n44831 , n44830 , n36702 );
not ( n44832 , n42832 );
and ( n44833 , n44832 , n42834 );
xor ( n44834 , n44831 , n44833 );
not ( n14663 , n29614 );
and ( n14664 , n14663 , RI1739fee0_1976);
and ( n14665 , n44834 , n29614 );
or ( n44835 , n14664 , n14665 );
not ( n14666 , RI1754c610_2);
and ( n14667 , n14666 , n44835 );
and ( n14668 , C0 , RI1754c610_2);
or ( n44836 , n14667 , n14668 );
buf ( n44837 , n44836 );
not ( n14669 , n27683 );
and ( n14670 , n14669 , RI19aaf790_2457);
and ( n14671 , RI19ab9498_2386 , n27683 );
or ( n44838 , n14670 , n14671 );
not ( n14672 , RI1754c610_2);
and ( n14673 , n14672 , n44838 );
and ( n14674 , C0 , RI1754c610_2);
or ( n44839 , n14673 , n14674 );
buf ( n44840 , n44839 );
not ( n14675 , n27683 );
and ( n14676 , n14675 , RI19aaf268_2460);
and ( n14677 , RI19ab8f70_2388 , n27683 );
or ( n44841 , n14676 , n14677 );
not ( n14678 , RI1754c610_2);
and ( n14679 , n14678 , n44841 );
and ( n14680 , C0 , RI1754c610_2);
or ( n44842 , n14679 , n14680 );
buf ( n44843 , n44842 );
xor ( n44844 , n34126 , n42377 );
xor ( n44845 , n44844 , n33991 );
xor ( n44846 , n41643 , n40692 );
xor ( n44847 , n44846 , n43994 );
not ( n44848 , n44847 );
xor ( n44849 , n37318 , n39914 );
xor ( n44850 , n44849 , n40237 );
and ( n44851 , n44848 , n44850 );
xor ( n44852 , n44845 , n44851 );
not ( n14681 , n29614 );
and ( n14682 , n14681 , RI17408868_1466);
and ( n14683 , n44852 , n29614 );
or ( n44853 , n14682 , n14683 );
not ( n14684 , RI1754c610_2);
and ( n14685 , n14684 , n44853 );
and ( n14686 , C0 , RI1754c610_2);
or ( n44854 , n14685 , n14686 );
buf ( n44855 , n44854 );
xor ( n44856 , n31657 , n30604 );
xor ( n44857 , n44856 , n30741 );
not ( n44858 , n42992 );
and ( n44859 , n44858 , n42994 );
xor ( n44860 , n44857 , n44859 );
not ( n14687 , n29614 );
and ( n14688 , n14687 , RI17491a28_1026);
and ( n14689 , n44860 , n29614 );
or ( n44861 , n14688 , n14689 );
not ( n14690 , RI1754c610_2);
and ( n14691 , n14690 , n44861 );
and ( n14692 , C0 , RI1754c610_2);
or ( n44862 , n14691 , n14692 );
buf ( n44863 , n44862 );
not ( n14693 , n27683 );
and ( n14694 , n14693 , RI19abc4e0_2365);
and ( n14695 , RI19ac4b68_2294 , n27683 );
or ( n44864 , n14694 , n14695 );
not ( n14696 , RI1754c610_2);
and ( n14697 , n14696 , n44864 );
and ( n14698 , C0 , RI1754c610_2);
or ( n44865 , n14697 , n14698 );
buf ( n44866 , n44865 );
not ( n14699 , n27683 );
and ( n14700 , n14699 , RI19a95750_2644);
and ( n14701 , RI19a9f548_2574 , n27683 );
or ( n44867 , n14700 , n14701 );
not ( n14702 , RI1754c610_2);
and ( n14703 , n14702 , n44867 );
and ( n14704 , C0 , RI1754c610_2);
or ( n44868 , n14703 , n14704 );
buf ( n44869 , n44868 );
not ( n14705 , n27683 );
and ( n14706 , n14705 , RI19aca9a0_2251);
and ( n14707 , RI19a85e68_2753 , n27683 );
or ( n44870 , n14706 , n14707 );
not ( n14708 , RI1754c610_2);
and ( n14709 , n14708 , n44870 );
and ( n14710 , C0 , RI1754c610_2);
or ( n44871 , n14709 , n14710 );
buf ( n44872 , n44871 );
xor ( n44873 , n40880 , n34340 );
xor ( n44874 , n44873 , n38817 );
xor ( n44875 , n35825 , n37129 );
xor ( n44876 , n44875 , n37169 );
not ( n44877 , n44876 );
xor ( n44878 , n40850 , n35009 );
xor ( n44879 , n44878 , n28816 );
and ( n44880 , n44877 , n44879 );
xor ( n44881 , n44874 , n44880 );
not ( n14711 , n29614 );
and ( n14712 , n14711 , RI17396b38_2021);
and ( n14713 , n44881 , n29614 );
or ( n44882 , n14712 , n14713 );
not ( n14714 , RI1754c610_2);
and ( n14715 , n14714 , n44882 );
and ( n14716 , C0 , RI1754c610_2);
or ( n44883 , n14715 , n14716 );
buf ( n44884 , n44883 );
xor ( n44885 , n39346 , n29843 );
xor ( n44886 , n44885 , n29981 );
xor ( n44887 , n38995 , n35804 );
xor ( n44888 , n44887 , n35842 );
not ( n44889 , n44888 );
xor ( n44890 , n37804 , n31213 );
xor ( n44891 , n44890 , n31317 );
and ( n44892 , n44889 , n44891 );
xor ( n44893 , n44886 , n44892 );
not ( n14717 , n29614 );
and ( n14718 , n14717 , RI173e9260_1619);
and ( n14719 , n44893 , n29614 );
or ( n44894 , n14718 , n14719 );
not ( n14720 , RI1754c610_2);
and ( n14721 , n14720 , n44894 );
and ( n14722 , C0 , RI1754c610_2);
or ( n44895 , n14721 , n14722 );
buf ( n44896 , n44895 );
xor ( n44897 , n36182 , n32309 );
xor ( n44898 , n44897 , n32923 );
xor ( n44899 , n34704 , n42605 );
xor ( n44900 , n44899 , n42619 );
not ( n44901 , n44900 );
xor ( n44902 , n41654 , n40692 );
xor ( n44903 , n44902 , n43994 );
and ( n44904 , n44901 , n44903 );
xor ( n44905 , n44898 , n44904 );
not ( n14723 , n29614 );
and ( n14724 , n14723 , RI17398578_2013);
and ( n14725 , n44905 , n29614 );
or ( n44906 , n14724 , n14725 );
not ( n14726 , RI1754c610_2);
and ( n14727 , n14726 , n44906 );
and ( n14728 , C0 , RI1754c610_2);
or ( n44907 , n14727 , n14728 );
buf ( n44908 , n44907 );
xor ( n44909 , n38396 , n37169 );
xor ( n44910 , n44909 , n36339 );
xor ( n44911 , n43277 , n41099 );
xor ( n44912 , n44911 , n30604 );
not ( n44913 , n44912 );
xor ( n44914 , n42020 , n41049 );
xor ( n44915 , n44914 , n41504 );
and ( n44916 , n44913 , n44915 );
xor ( n44917 , n44910 , n44916 );
not ( n14729 , n29614 );
and ( n14730 , n14729 , RI1738bd50_2074);
and ( n14731 , n44917 , n29614 );
or ( n44918 , n14730 , n14731 );
not ( n14732 , RI1754c610_2);
and ( n14733 , n14732 , n44918 );
and ( n14734 , C0 , RI1754c610_2);
or ( n44919 , n14733 , n14734 );
buf ( n44920 , n44919 );
xor ( n44921 , n40763 , n33778 );
xor ( n44922 , n44921 , n38793 );
not ( n44923 , n42112 );
and ( n44924 , n44923 , n42114 );
xor ( n44925 , n44922 , n44924 );
not ( n14735 , n29614 );
and ( n14736 , n14735 , RI173e9c38_1616);
and ( n14737 , n44925 , n29614 );
or ( n44926 , n14736 , n14737 );
not ( n14738 , RI1754c610_2);
and ( n14739 , n14738 , n44926 );
and ( n14740 , C0 , RI1754c610_2);
or ( n44927 , n14739 , n14740 );
buf ( n44928 , n44927 );
xor ( n44929 , n36352 , n38676 );
xor ( n44930 , n44929 , n28111 );
xor ( n44931 , n32185 , n35986 );
xor ( n44932 , n44931 , n36003 );
not ( n44933 , n44932 );
xor ( n44934 , n32704 , n36209 );
xor ( n44935 , n44934 , n40412 );
and ( n44936 , n44933 , n44935 );
xor ( n44937 , n44930 , n44936 );
not ( n14741 , n29614 );
and ( n14742 , n14741 , RI174513d8_1340);
and ( n14743 , n44937 , n29614 );
or ( n44938 , n14742 , n14743 );
not ( n14744 , RI1754c610_2);
and ( n14745 , n14744 , n44938 );
and ( n14746 , C0 , RI1754c610_2);
or ( n44939 , n14745 , n14746 );
buf ( n44940 , n44939 );
xor ( n44941 , n37230 , n39467 );
xor ( n44942 , n44941 , n41391 );
not ( n44943 , n44942 );
xor ( n44944 , n36843 , n44146 );
xor ( n44945 , n44944 , n41198 );
and ( n44946 , n44943 , n44945 );
xor ( n44947 , n44476 , n44946 );
not ( n14747 , n29614 );
and ( n14748 , n14747 , RI17511600_712);
and ( n14749 , n44947 , n29614 );
or ( n44948 , n14748 , n14749 );
not ( n14750 , RI1754c610_2);
and ( n14751 , n14750 , n44948 );
and ( n14752 , C0 , RI1754c610_2);
or ( n44949 , n14751 , n14752 );
buf ( n44950 , n44949 );
not ( n44951 , n42283 );
xor ( n44952 , n39384 , n35594 );
xor ( n44953 , n44952 , n32403 );
and ( n44954 , n44951 , n44953 );
xor ( n44955 , n42280 , n44954 );
not ( n14753 , n29614 );
and ( n14754 , n14753 , RI1740f7f8_1432);
and ( n14755 , n44955 , n29614 );
or ( n44956 , n14754 , n14755 );
not ( n14756 , RI1754c610_2);
and ( n14757 , n14756 , n44956 );
and ( n14758 , C0 , RI1754c610_2);
or ( n44957 , n14757 , n14758 );
buf ( n44958 , n44957 );
not ( n14759 , n27683 );
and ( n14760 , n14759 , RI19ac3920_2302);
and ( n14761 , RI19acc5c0_2236 , n27683 );
or ( n44959 , n14760 , n14761 );
not ( n14762 , RI1754c610_2);
and ( n14763 , n14762 , n44959 );
and ( n14764 , C0 , RI1754c610_2);
or ( n44960 , n14763 , n14764 );
buf ( n44961 , n44960 );
xor ( n44962 , n36795 , n38214 );
xor ( n44963 , n44962 , n38244 );
not ( n44964 , n38830 );
and ( n44965 , n44964 , n38835 );
xor ( n44966 , n44963 , n44965 );
not ( n14765 , n29614 );
and ( n14766 , n14765 , RI1748e260_1043);
and ( n14767 , n44966 , n29614 );
or ( n44967 , n14766 , n14767 );
not ( n14768 , RI1754c610_2);
and ( n14769 , n14768 , n44967 );
and ( n14770 , C0 , RI1754c610_2);
or ( n44968 , n14769 , n14770 );
buf ( n44969 , n44968 );
xor ( n44970 , n40961 , n36844 );
xor ( n44971 , n44970 , n36874 );
xor ( n44972 , n41884 , n38085 );
xor ( n44973 , n44972 , n38115 );
not ( n44974 , n44973 );
xor ( n44975 , n39249 , n35361 );
xor ( n44976 , n44975 , n38445 );
and ( n44977 , n44974 , n44976 );
xor ( n44978 , n44971 , n44977 );
not ( n14771 , n29614 );
and ( n14772 , n14771 , RI17492748_1022);
and ( n14773 , n44978 , n29614 );
or ( n44979 , n14772 , n14773 );
not ( n14774 , RI1754c610_2);
and ( n14775 , n14774 , n44979 );
and ( n14776 , C0 , RI1754c610_2);
or ( n44980 , n14775 , n14776 );
buf ( n44981 , n44980 );
xor ( n44982 , n39913 , n33397 );
xor ( n44983 , n44982 , n35710 );
xor ( n44984 , n31335 , n37074 );
xor ( n44985 , n44984 , n37104 );
not ( n44986 , n44985 );
xor ( n44987 , n40759 , n33778 );
xor ( n44988 , n44987 , n38793 );
and ( n44989 , n44986 , n44988 );
xor ( n44990 , n44983 , n44989 );
not ( n14777 , n29614 );
and ( n14778 , n14777 , RI1749b460_979);
and ( n14779 , n44990 , n29614 );
or ( n44991 , n14778 , n14779 );
not ( n14780 , RI1754c610_2);
and ( n14781 , n14780 , n44991 );
and ( n14782 , C0 , RI1754c610_2);
or ( n44992 , n14781 , n14782 );
buf ( n44993 , n44992 );
buf ( n44994 , RI174a16d0_949);
not ( n44995 , n43928 );
xor ( n44996 , n30962 , n41622 );
xor ( n44997 , n44996 , n38512 );
and ( n44998 , n44995 , n44997 );
xor ( n44999 , n43925 , n44998 );
not ( n14783 , n29614 );
and ( n14784 , n14783 , RI1751bb00_680);
and ( n14785 , n44999 , n29614 );
or ( n45000 , n14784 , n14785 );
not ( n14786 , RI1754c610_2);
and ( n14787 , n14786 , n45000 );
and ( n14788 , C0 , RI1754c610_2);
or ( n45001 , n14787 , n14788 );
buf ( n45002 , n45001 );
xor ( n45003 , n38924 , n42309 );
xor ( n45004 , n45003 , n43464 );
xor ( n45005 , n39988 , n41934 );
xor ( n45006 , n45005 , n40341 );
not ( n45007 , n45006 );
xor ( n45008 , n34731 , n42619 );
xor ( n45009 , n45008 , n41990 );
and ( n45010 , n45007 , n45009 );
xor ( n45011 , n45004 , n45010 );
not ( n14789 , n29614 );
and ( n14790 , n14789 , RI174920b8_1024);
and ( n14791 , n45011 , n29614 );
or ( n45012 , n14790 , n14791 );
not ( n14792 , RI1754c610_2);
and ( n14793 , n14792 , n45012 );
and ( n14794 , C0 , RI1754c610_2);
or ( n45013 , n14793 , n14794 );
buf ( n45014 , n45013 );
buf ( n45015 , RI174b1a08_870);
xor ( n45016 , n39492 , n30923 );
xor ( n45017 , n45016 , n31053 );
not ( n45018 , n41148 );
and ( n45019 , n45018 , n41150 );
xor ( n45020 , n45017 , n45019 );
not ( n14795 , n29614 );
and ( n14796 , n14795 , RI174462a8_1394);
and ( n14797 , n45020 , n29614 );
or ( n45021 , n14796 , n14797 );
not ( n14798 , RI1754c610_2);
and ( n14799 , n14798 , n45021 );
and ( n14800 , C0 , RI1754c610_2);
or ( n45022 , n14799 , n14800 );
buf ( n45023 , n45022 );
xor ( n45024 , n37929 , n40210 );
xor ( n45025 , n45024 , n39989 );
not ( n45026 , n37422 );
and ( n45027 , n45026 , n37440 );
xor ( n45028 , n45025 , n45027 );
not ( n14801 , n29614 );
and ( n14802 , n14801 , RI17455230_1321);
and ( n14803 , n45028 , n29614 );
or ( n45029 , n14802 , n14803 );
not ( n14804 , RI1754c610_2);
and ( n14805 , n14804 , n45029 );
and ( n14806 , C0 , RI1754c610_2);
or ( n45030 , n14805 , n14806 );
buf ( n45031 , n45030 );
not ( n14807 , n27683 );
and ( n14808 , n14807 , RI19ab34f8_2429);
and ( n14809 , RI19abd2f0_2357 , n27683 );
or ( n45032 , n14808 , n14809 );
not ( n14810 , RI1754c610_2);
and ( n14811 , n14810 , n45032 );
and ( n14812 , C0 , RI1754c610_2);
or ( n45033 , n14811 , n14812 );
buf ( n45034 , n45033 );
not ( n14813 , n27683 );
and ( n14814 , n14813 , RI19a83690_2770);
and ( n14815 , RI19ab6cc0_2403 , n27683 );
or ( n45035 , n14814 , n14815 );
not ( n14816 , RI1754c610_2);
and ( n14817 , n14816 , n45035 );
and ( n14818 , C0 , RI1754c610_2);
or ( n45036 , n14817 , n14818 );
buf ( n45037 , n45036 );
xor ( n45038 , n36061 , n34475 );
xor ( n45039 , n45038 , n37371 );
xor ( n45040 , n38091 , n40111 );
xor ( n45041 , n45040 , n43278 );
not ( n45042 , n45041 );
xor ( n45043 , n28265 , n41799 );
xor ( n45044 , n45043 , n40381 );
and ( n45045 , n45042 , n45044 );
xor ( n45046 , n45039 , n45045 );
not ( n14819 , n29614 );
and ( n14820 , n14819 , RI174a44c0_935);
and ( n14821 , n45046 , n29614 );
or ( n45047 , n14820 , n14821 );
not ( n14822 , RI1754c610_2);
and ( n14823 , n14822 , n45047 );
and ( n14824 , C0 , RI1754c610_2);
or ( n45048 , n14823 , n14824 );
buf ( n45049 , n45048 );
not ( n45050 , n43022 );
and ( n45051 , n45050 , n43027 );
xor ( n45052 , n42325 , n45051 );
not ( n14825 , n29614 );
and ( n14826 , n14825 , RI174b8a10_836);
and ( n14827 , n45052 , n29614 );
or ( n45053 , n14826 , n14827 );
not ( n14828 , RI1754c610_2);
and ( n14829 , n14828 , n45053 );
and ( n14830 , C0 , RI1754c610_2);
or ( n45054 , n14829 , n14830 );
buf ( n45055 , n45054 );
not ( n14831 , n27683 );
and ( n14832 , n14831 , RI19abdf98_2350);
and ( n14833 , RI19ac6e18_2278 , n27683 );
or ( n45056 , n14832 , n14833 );
not ( n14834 , RI1754c610_2);
and ( n14835 , n14834 , n45056 );
and ( n14836 , C0 , RI1754c610_2);
or ( n45057 , n14835 , n14836 );
buf ( n45058 , n45057 );
not ( n14837 , RI1754c610_2);
and ( n14838 , n14837 , RI17539218_590);
and ( n14839 , C0 , RI1754c610_2);
or ( n45059 , n14838 , n14839 );
buf ( n45060 , n45059 );
not ( n45061 , n35598 );
xor ( n45062 , n34272 , n38886 );
xor ( n45063 , n45062 , n39604 );
and ( n45064 , n45061 , n45063 );
xor ( n45065 , n35595 , n45064 );
not ( n14840 , n29614 );
and ( n14841 , n14840 , RI173f7b58_1548);
and ( n14842 , n45065 , n29614 );
or ( n45066 , n14841 , n14842 );
not ( n14843 , RI1754c610_2);
and ( n14844 , n14843 , n45066 );
and ( n14845 , C0 , RI1754c610_2);
or ( n45067 , n14844 , n14845 );
buf ( n45068 , n45067 );
xor ( n45069 , n40515 , n41430 );
xor ( n45070 , n45069 , n36844 );
xor ( n45071 , n41606 , n43278 );
xor ( n45072 , n45071 , n31664 );
not ( n45073 , n45072 );
xor ( n45074 , n34102 , n42377 );
xor ( n45075 , n45074 , n33991 );
and ( n45076 , n45073 , n45075 );
xor ( n45077 , n45070 , n45076 );
not ( n14846 , n29614 );
and ( n14847 , n14846 , RI17455578_1320);
and ( n14848 , n45077 , n29614 );
or ( n45078 , n14847 , n14848 );
not ( n14849 , RI1754c610_2);
and ( n14850 , n14849 , n45078 );
and ( n14851 , C0 , RI1754c610_2);
or ( n45079 , n14850 , n14851 );
buf ( n45080 , n45079 );
xor ( n45081 , n41206 , n39397 );
xor ( n45082 , n45081 , n39414 );
xor ( n45083 , n38436 , n40585 );
xor ( n45084 , n45083 , n34918 );
not ( n45085 , n45084 );
xor ( n45086 , n30603 , n38167 );
xor ( n45087 , n45086 , n33728 );
and ( n45088 , n45085 , n45087 );
xor ( n45089 , n45082 , n45088 );
not ( n14852 , n29614 );
and ( n14853 , n14852 , RI17510160_716);
and ( n14854 , n45089 , n29614 );
or ( n45090 , n14853 , n14854 );
not ( n14855 , RI1754c610_2);
and ( n14856 , n14855 , n45090 );
and ( n14857 , C0 , RI1754c610_2);
or ( n45091 , n14856 , n14857 );
buf ( n45092 , n45091 );
not ( n45093 , n36465 );
xor ( n45094 , n36689 , n39655 );
xor ( n45095 , n45094 , n41125 );
and ( n45096 , n45093 , n45095 );
xor ( n45097 , n36433 , n45096 );
not ( n14858 , n29614 );
and ( n14859 , n14858 , RI17335590_2181);
and ( n14860 , n45097 , n29614 );
or ( n45098 , n14859 , n14860 );
not ( n14861 , RI1754c610_2);
and ( n14862 , n14861 , n45098 );
and ( n14863 , C0 , RI1754c610_2);
or ( n45099 , n14862 , n14863 );
buf ( n45100 , n45099 );
not ( n45101 , n42320 );
and ( n45102 , n45101 , n42322 );
xor ( n45103 , n43027 , n45102 );
not ( n14864 , n29614 );
and ( n14865 , n14864 , RI175177f8_693);
and ( n14866 , n45103 , n29614 );
or ( n45104 , n14865 , n14866 );
not ( n14867 , RI1754c610_2);
and ( n14868 , n14867 , n45104 );
and ( n14869 , C0 , RI1754c610_2);
or ( n45105 , n14868 , n14869 );
buf ( n45106 , n45105 );
xor ( n45107 , n33068 , n36227 );
xor ( n45108 , n45107 , n40743 );
xor ( n45109 , n37466 , n42188 );
xor ( n45110 , n45109 , n41526 );
not ( n45111 , n45110 );
xor ( n45112 , n30989 , n41622 );
xor ( n45113 , n45112 , n38512 );
and ( n45114 , n45111 , n45113 );
xor ( n45115 , n45108 , n45114 );
not ( n14870 , n29614 );
and ( n14871 , n14870 , RI1748e5a8_1042);
and ( n14872 , n45115 , n29614 );
or ( n45116 , n14871 , n14872 );
not ( n14873 , RI1754c610_2);
and ( n14874 , n14873 , n45116 );
and ( n14875 , C0 , RI1754c610_2);
or ( n45117 , n14874 , n14875 );
buf ( n45118 , n45117 );
not ( n45119 , n43015 );
and ( n45120 , n45119 , n40770 );
xor ( n45121 , n43012 , n45120 );
not ( n14876 , n29614 );
and ( n14877 , n14876 , RI17400bb8_1504);
and ( n14878 , n45121 , n29614 );
or ( n45122 , n14877 , n14878 );
not ( n14879 , RI1754c610_2);
and ( n14880 , n14879 , n45122 );
and ( n14881 , C0 , RI1754c610_2);
or ( n45123 , n14880 , n14881 );
buf ( n45124 , n45123 );
not ( n14882 , n27683 );
and ( n14883 , n14882 , RI19aba8c0_2377);
and ( n14884 , RI19ac30b0_2306 , n27683 );
or ( n45125 , n14883 , n14884 );
not ( n14885 , RI1754c610_2);
and ( n14886 , n14885 , n45125 );
and ( n14887 , C0 , RI1754c610_2);
or ( n45126 , n14886 , n14887 );
buf ( n45127 , n45126 );
xor ( n45128 , n37675 , n37549 );
xor ( n45129 , n45128 , n37579 );
xor ( n45130 , n38967 , n41590 );
xor ( n45131 , n45130 , n35804 );
not ( n45132 , n45131 );
xor ( n45133 , n43479 , n32108 );
xor ( n45134 , n45133 , n38347 );
and ( n45135 , n45132 , n45134 );
xor ( n45136 , n45129 , n45135 );
not ( n14888 , n29614 );
and ( n14889 , n14888 , RI1749e250_965);
and ( n14890 , n45136 , n29614 );
or ( n45137 , n14889 , n14890 );
not ( n14891 , RI1754c610_2);
and ( n14892 , n14891 , n45137 );
and ( n14893 , C0 , RI1754c610_2);
or ( n45138 , n14892 , n14893 );
buf ( n45139 , n45138 );
xor ( n45140 , n37926 , n40210 );
xor ( n45141 , n45140 , n39989 );
xor ( n45142 , n34937 , n36802 );
xor ( n45143 , n45142 , n33125 );
not ( n45144 , n45143 );
and ( n45145 , n45144 , n40390 );
xor ( n45146 , n45141 , n45145 );
not ( n14894 , n29614 );
and ( n14895 , n14894 , RI174abae0_899);
and ( n14896 , n45146 , n29614 );
or ( n45147 , n14895 , n14896 );
not ( n14897 , RI1754c610_2);
and ( n14898 , n14897 , n45147 );
and ( n14899 , C0 , RI1754c610_2);
or ( n45148 , n14898 , n14899 );
buf ( n45149 , n45148 );
not ( n14900 , n27683 );
and ( n14901 , n14900 , RI19a96bf0_2635);
and ( n14902 , RI19aa0790_2565 , n27683 );
or ( n45150 , n14901 , n14902 );
not ( n14903 , RI1754c610_2);
and ( n14904 , n14903 , n45150 );
and ( n14905 , C0 , RI1754c610_2);
or ( n45151 , n14904 , n14905 );
buf ( n45152 , n45151 );
xor ( n45153 , n37160 , n40254 );
xor ( n45154 , n45153 , n40718 );
not ( n45155 , n45154 );
xor ( n45156 , n40584 , n37048 );
xor ( n45157 , n45156 , n36772 );
and ( n45158 , n45155 , n45157 );
xor ( n45159 , n41705 , n45158 );
not ( n14906 , n29614 );
and ( n14907 , n14906 , RI1739acd8_2001);
and ( n14908 , n45159 , n29614 );
or ( n45160 , n14907 , n14908 );
not ( n14909 , RI1754c610_2);
and ( n14910 , n14909 , n45160 );
and ( n14911 , C0 , RI1754c610_2);
or ( n45161 , n14910 , n14911 );
buf ( n45162 , n45161 );
xor ( n45163 , n32443 , n35622 );
xor ( n45164 , n45163 , n35639 );
not ( n45165 , n44963 );
and ( n45166 , n45165 , n38830 );
xor ( n45167 , n45164 , n45166 );
not ( n14912 , n29614 );
and ( n14913 , n14912 , RI1747fcb0_1113);
and ( n14914 , n45167 , n29614 );
or ( n45168 , n14913 , n14914 );
not ( n14915 , RI1754c610_2);
and ( n14916 , n14915 , n45168 );
and ( n14917 , C0 , RI1754c610_2);
or ( n45169 , n14916 , n14917 );
buf ( n45170 , n45169 );
xor ( n45171 , n33696 , n41854 );
xor ( n45172 , n45171 , n40283 );
not ( n45173 , n45172 );
xor ( n45174 , n38638 , n34300 );
xor ( n45175 , n45174 , n34340 );
and ( n45176 , n45173 , n45175 );
xor ( n45177 , n42985 , n45176 );
not ( n14918 , n29614 );
and ( n14919 , n14918 , RI1749a3f8_984);
and ( n14920 , n45177 , n29614 );
or ( n45178 , n14919 , n14920 );
not ( n14921 , RI1754c610_2);
and ( n14922 , n14921 , n45178 );
and ( n14923 , C0 , RI1754c610_2);
or ( n45179 , n14922 , n14923 );
buf ( n45180 , n45179 );
xor ( n45181 , n31771 , n34644 );
xor ( n45182 , n45181 , n36401 );
xor ( n45183 , n39939 , n38724 );
xor ( n45184 , n45183 , n29425 );
not ( n45185 , n45184 );
and ( n45186 , n45185 , n44095 );
xor ( n45187 , n45182 , n45186 );
not ( n14924 , n29614 );
and ( n14925 , n14924 , RI173ca618_1769);
and ( n14926 , n45187 , n29614 );
or ( n45188 , n14925 , n14926 );
not ( n14927 , RI1754c610_2);
and ( n14928 , n14927 , n45188 );
and ( n14929 , C0 , RI1754c610_2);
or ( n45189 , n14928 , n14929 );
buf ( n45190 , n45189 );
xor ( n45191 , n37986 , n41504 );
xor ( n45192 , n45191 , n41690 );
xor ( n45193 , n39862 , n42504 );
xor ( n45194 , n45193 , n41818 );
not ( n45195 , n45194 );
xor ( n45196 , n35445 , n32715 );
xor ( n45197 , n45196 , n36654 );
and ( n45198 , n45195 , n45197 );
xor ( n45199 , n45192 , n45198 );
not ( n14930 , n29614 );
and ( n14931 , n14930 , RI174a0cf8_952);
and ( n14932 , n45199 , n29614 );
or ( n45200 , n14931 , n14932 );
not ( n14933 , RI1754c610_2);
and ( n14934 , n14933 , n45200 );
and ( n14935 , C0 , RI1754c610_2);
or ( n45201 , n14934 , n14935 );
buf ( n45202 , n45201 );
xor ( n45203 , n38361 , n33880 );
xor ( n45204 , n45203 , n33935 );
not ( n45205 , n45204 );
and ( n45206 , n45205 , n43923 );
xor ( n45207 , n44997 , n45206 );
not ( n14936 , n29614 );
and ( n14937 , n14936 , RI174ace90_893);
and ( n14938 , n45207 , n29614 );
or ( n45208 , n14937 , n14938 );
not ( n14939 , RI1754c610_2);
and ( n14940 , n14939 , n45208 );
and ( n14941 , C0 , RI1754c610_2);
or ( n45209 , n14940 , n14941 );
buf ( n45210 , n45209 );
buf ( n45211 , RI17475f30_1161);
buf ( n45212 , RI1747adf0_1137);
xor ( n45213 , n40996 , n36998 );
xor ( n45214 , n45213 , n37048 );
not ( n45215 , n45214 );
xor ( n45216 , n31294 , n42049 );
xor ( n45217 , n45216 , n37849 );
and ( n45218 , n45215 , n45217 );
xor ( n45219 , n39103 , n45218 );
not ( n14942 , n29614 );
and ( n14943 , n14942 , RI1738a9a0_2080);
and ( n14944 , n45219 , n29614 );
or ( n45220 , n14943 , n14944 );
not ( n14945 , RI1754c610_2);
and ( n14946 , n14945 , n45220 );
and ( n14947 , C0 , RI1754c610_2);
or ( n45221 , n14946 , n14947 );
buf ( n45222 , n45221 );
xor ( n45223 , n41989 , n39886 );
xor ( n45224 , n45223 , n36998 );
xor ( n45225 , n39135 , n28468 );
xor ( n45226 , n45225 , n36530 );
not ( n45227 , n45226 );
xor ( n45228 , n39050 , n39702 );
xor ( n45229 , n45228 , n39914 );
and ( n45230 , n45227 , n45229 );
xor ( n45231 , n45224 , n45230 );
not ( n14948 , n29614 );
and ( n14949 , n14948 , RI173f6af0_1553);
and ( n14950 , n45231 , n29614 );
or ( n45232 , n14949 , n14950 );
not ( n14951 , RI1754c610_2);
and ( n14952 , n14951 , n45232 );
and ( n14953 , C0 , RI1754c610_2);
or ( n45233 , n14952 , n14953 );
buf ( n45234 , n45233 );
not ( n14954 , n27683 );
and ( n14955 , n14954 , RI19a83f78_2766);
and ( n14956 , RI19abba90_2370 , n27683 );
or ( n45235 , n14955 , n14956 );
not ( n14957 , RI1754c610_2);
and ( n14958 , n14957 , n45235 );
and ( n14959 , C0 , RI1754c610_2);
or ( n45236 , n14958 , n14959 );
buf ( n45237 , n45236 );
xor ( n45238 , n34308 , n39604 );
xor ( n45239 , n45238 , n39621 );
not ( n45240 , n45239 );
and ( n45241 , n45240 , n42125 );
xor ( n45242 , n41592 , n45241 );
not ( n14960 , n29614 );
and ( n14961 , n14960 , RI173c39d0_1802);
and ( n14962 , n45242 , n29614 );
or ( n45243 , n14961 , n14962 );
not ( n14963 , RI1754c610_2);
and ( n14964 , n14963 , n45243 );
and ( n14965 , C0 , RI1754c610_2);
or ( n45244 , n14964 , n14965 );
buf ( n45245 , n45244 );
buf ( n45246 , RI1746ced0_1205);
xor ( n45247 , n41197 , n34622 );
xor ( n45248 , n45247 , n39397 );
xor ( n45249 , n39075 , n36377 );
xor ( n45250 , n45249 , n39131 );
not ( n45251 , n45250 );
and ( n45252 , n45251 , n37697 );
xor ( n45253 , n45248 , n45252 );
not ( n14966 , n29614 );
and ( n14967 , n14966 , RI1740b9a0_1451);
and ( n14968 , n45253 , n29614 );
or ( n45254 , n14967 , n14968 );
not ( n14969 , RI1754c610_2);
and ( n14970 , n14969 , n45254 );
and ( n14971 , C0 , RI1754c610_2);
or ( n45255 , n14970 , n14971 );
buf ( n45256 , n45255 );
not ( n14972 , n27683 );
and ( n14973 , n14972 , RI19aa2c20_2547);
and ( n14974 , RI19aacdd8_2476 , n27683 );
or ( n45257 , n14973 , n14974 );
not ( n14975 , RI1754c610_2);
and ( n14976 , n14975 , n45257 );
and ( n14977 , C0 , RI1754c610_2);
or ( n45258 , n14976 , n14977 );
buf ( n45259 , n45258 );
not ( n45260 , n39479 );
xor ( n45261 , n34134 , n33069 );
xor ( n45262 , n45261 , n42264 );
and ( n45263 , n45260 , n45262 );
xor ( n45264 , n39473 , n45263 );
not ( n14978 , n29614 );
and ( n14979 , n14978 , RI173ade00_1908);
and ( n14980 , n45264 , n29614 );
or ( n45265 , n14979 , n14980 );
not ( n14981 , RI1754c610_2);
and ( n14982 , n14981 , n45265 );
and ( n14983 , C0 , RI1754c610_2);
or ( n45266 , n14982 , n14983 );
buf ( n45267 , n45266 );
xor ( n45268 , n34812 , n41478 );
xor ( n45269 , n45268 , n41146 );
not ( n45270 , n45269 );
and ( n45271 , n45270 , n43237 );
xor ( n45272 , n44214 , n45271 );
not ( n14984 , n29614 );
and ( n14985 , n14984 , RI1746ced0_1205);
and ( n14986 , n45272 , n29614 );
or ( n45273 , n14985 , n14986 );
not ( n14987 , RI1754c610_2);
and ( n14988 , n14987 , n45273 );
and ( n14989 , C0 , RI1754c610_2);
or ( n45274 , n14988 , n14989 );
buf ( n45275 , n45274 );
buf ( n45276 , RI17485bd8_1084);
buf ( n45277 , RI17509f68_735);
xor ( n45278 , n34561 , n40563 );
xor ( n45279 , n45278 , n35544 );
xor ( n45280 , n40827 , n42635 );
xor ( n45281 , n45280 , n33648 );
not ( n45282 , n45281 );
xor ( n45283 , n36179 , n32309 );
xor ( n45284 , n45283 , n32923 );
and ( n45285 , n45282 , n45284 );
xor ( n45286 , n45279 , n45285 );
not ( n14990 , n29614 );
and ( n14991 , n14990 , RI174b51d0_853);
and ( n14992 , n45286 , n29614 );
or ( n45287 , n14991 , n14992 );
not ( n14993 , RI1754c610_2);
and ( n14994 , n14993 , n45287 );
and ( n14995 , C0 , RI1754c610_2);
or ( n45288 , n14994 , n14995 );
buf ( n45289 , n45288 );
xor ( n45290 , n41303 , n41526 );
xor ( n45291 , n45290 , n41543 );
not ( n45292 , n43071 );
and ( n45293 , n45292 , n42844 );
xor ( n45294 , n45291 , n45293 );
not ( n14996 , n29614 );
and ( n14997 , n14996 , RI174c2f10_804);
and ( n14998 , n45294 , n29614 );
or ( n45295 , n14997 , n14998 );
not ( n14999 , RI1754c610_2);
and ( n15000 , n14999 , n45295 );
and ( n15001 , C0 , RI1754c610_2);
or ( n45296 , n15000 , n15001 );
buf ( n45297 , n45296 );
xor ( n45298 , n40935 , n38793 );
xor ( n45299 , n45298 , n40563 );
not ( n45300 , n39468 );
and ( n45301 , n45300 , n39473 );
xor ( n45302 , n45299 , n45301 );
not ( n15002 , n29614 );
and ( n15003 , n15002 , RI17457300_1311);
and ( n15004 , n45302 , n29614 );
or ( n45303 , n15003 , n15004 );
not ( n15005 , RI1754c610_2);
and ( n15006 , n15005 , n45303 );
and ( n15007 , C0 , RI1754c610_2);
or ( n45304 , n15006 , n15007 );
buf ( n45305 , n45304 );
xor ( n45306 , n37489 , n42188 );
xor ( n45307 , n45306 , n41526 );
xor ( n45308 , n35812 , n37129 );
xor ( n45309 , n45308 , n37169 );
not ( n45310 , n45309 );
xor ( n45311 , n35027 , n37814 );
xor ( n45312 , n45311 , n33223 );
and ( n45313 , n45310 , n45312 );
xor ( n45314 , n45307 , n45313 );
not ( n15008 , n29614 );
and ( n15009 , n15008 , RI173386c8_2166);
and ( n15010 , n45314 , n29614 );
or ( n45315 , n15009 , n15010 );
not ( n15011 , RI1754c610_2);
and ( n15012 , n15011 , n45315 );
and ( n15013 , C0 , RI1754c610_2);
or ( n45316 , n15012 , n15013 );
buf ( n45317 , n45316 );
xor ( n45318 , n40354 , n37898 );
xor ( n45319 , n45318 , n37915 );
xor ( n45320 , n37978 , n41504 );
xor ( n45321 , n45320 , n41690 );
not ( n45322 , n45321 );
xor ( n45323 , n41214 , n39397 );
xor ( n45324 , n45323 , n39414 );
and ( n45325 , n45322 , n45324 );
xor ( n45326 , n45319 , n45325 );
not ( n15014 , n29614 );
and ( n15015 , n15014 , RI1739fb98_1977);
and ( n15016 , n45326 , n29614 );
or ( n45327 , n15015 , n15016 );
not ( n15017 , RI1754c610_2);
and ( n15018 , n15017 , n45327 );
and ( n15019 , C0 , RI1754c610_2);
or ( n45328 , n15018 , n15019 );
buf ( n45329 , n45328 );
xor ( n45330 , n33396 , n39005 );
xor ( n45331 , n45330 , n39543 );
xor ( n45332 , n41300 , n41526 );
xor ( n45333 , n45332 , n41543 );
not ( n45334 , n45333 );
and ( n45335 , n45334 , n41462 );
xor ( n45336 , n45331 , n45335 );
not ( n15020 , n29614 );
and ( n15021 , n15020 , RI17404038_1488);
and ( n15022 , n45336 , n29614 );
or ( n45337 , n15021 , n15022 );
not ( n15023 , RI1754c610_2);
and ( n15024 , n15023 , n45337 );
and ( n15025 , C0 , RI1754c610_2);
or ( n45338 , n15024 , n15025 );
buf ( n45339 , n45338 );
not ( n45340 , n42564 );
and ( n45341 , n45340 , n35656 );
xor ( n45342 , n36703 , n45341 );
not ( n15026 , n29614 );
and ( n15027 , n15026 , RI17494b60_1011);
and ( n15028 , n45342 , n29614 );
or ( n45343 , n15027 , n15028 );
not ( n15029 , RI1754c610_2);
and ( n15030 , n15029 , n45343 );
and ( n15031 , C0 , RI1754c610_2);
or ( n45344 , n15030 , n15031 );
buf ( n45345 , n45344 );
not ( n15032 , n27683 );
and ( n15033 , n15032 , RI19ab71e8_2401);
and ( n15034 , RI19ac0158_2331 , n27683 );
or ( n45346 , n15033 , n15034 );
not ( n15035 , RI1754c610_2);
and ( n15036 , n15035 , n45346 );
and ( n15037 , C0 , RI1754c610_2);
or ( n45347 , n15036 , n15037 );
buf ( n45348 , n45347 );
not ( n15038 , n27683 );
and ( n15039 , n15038 , RI19ab5640_2413);
and ( n15040 , RI19abebc8_2343 , n27683 );
or ( n45349 , n15039 , n15040 );
not ( n15041 , RI1754c610_2);
and ( n15042 , n15041 , n45349 );
and ( n15043 , C0 , RI1754c610_2);
or ( n45350 , n15042 , n15043 );
buf ( n45351 , n45350 );
not ( n45352 , n42973 );
and ( n45353 , n45352 , n44287 );
xor ( n45354 , n42970 , n45353 );
not ( n15044 , n29614 );
and ( n15045 , n15044 , RI1745b7e8_1290);
and ( n15046 , n45354 , n29614 );
or ( n45355 , n15045 , n15046 );
not ( n15047 , RI1754c610_2);
and ( n15048 , n15047 , n45355 );
and ( n15049 , C0 , RI1754c610_2);
or ( n45356 , n15048 , n15049 );
buf ( n45357 , n45356 );
not ( n45358 , n44338 );
xor ( n45359 , n42043 , n33648 );
xor ( n45360 , n45359 , n33697 );
and ( n45361 , n45358 , n45360 );
xor ( n45362 , n44335 , n45361 );
not ( n15050 , n29614 );
and ( n15051 , n15050 , RI17345f58_2100);
and ( n15052 , n45362 , n29614 );
or ( n45363 , n15051 , n15052 );
not ( n15053 , RI1754c610_2);
and ( n15054 , n15053 , n45363 );
and ( n15055 , C0 , RI1754c610_2);
or ( n45364 , n15054 , n15055 );
buf ( n45365 , n45364 );
xor ( n45366 , n42614 , n39856 );
xor ( n45367 , n45366 , n39886 );
xor ( n45368 , n39524 , n38371 );
xor ( n45369 , n45368 , n36431 );
not ( n45370 , n45369 );
xor ( n45371 , n39547 , n38401 );
xor ( n45372 , n45371 , n41068 );
and ( n45373 , n45370 , n45372 );
xor ( n45374 , n45367 , n45373 );
not ( n15056 , n29614 );
and ( n15057 , n15056 , RI173ab010_1922);
and ( n15058 , n45374 , n29614 );
or ( n45375 , n15057 , n15058 );
not ( n15059 , RI1754c610_2);
and ( n15060 , n15059 , n45375 );
and ( n15061 , C0 , RI1754c610_2);
or ( n45376 , n15060 , n15061 );
buf ( n45377 , n45376 );
not ( n15062 , n27683 );
and ( n15063 , n15062 , RI19ac8510_2267);
and ( n15064 , RI19a83438_2771 , n27683 );
or ( n45378 , n15063 , n15064 );
not ( n15065 , RI1754c610_2);
and ( n15066 , n15065 , n45378 );
and ( n15067 , C0 , RI1754c610_2);
or ( n45379 , n15066 , n15067 );
buf ( n45380 , n45379 );
buf ( n45381 , RI174a8318_916);
buf ( n45382 , RI17474b80_1167);
buf ( n45383 , RI174ab108_902);
xor ( n45384 , n34059 , n39525 );
xor ( n45385 , n45384 , n42377 );
xor ( n45386 , n34414 , n40009 );
xor ( n45387 , n45386 , n38085 );
not ( n45388 , n45387 );
and ( n45389 , n45388 , n41712 );
xor ( n45390 , n45385 , n45389 );
not ( n15068 , n29614 );
and ( n15069 , n15068 , RI17342ad8_2116);
and ( n15070 , n45390 , n29614 );
or ( n45391 , n15069 , n15070 );
not ( n15071 , RI1754c610_2);
and ( n15072 , n15071 , n45391 );
and ( n15073 , C0 , RI1754c610_2);
or ( n45392 , n15072 , n15073 );
buf ( n45393 , n45392 );
not ( n15074 , n27683 );
and ( n15075 , n15074 , RI19ac1148_2322);
and ( n15076 , RI19aca4f0_2253 , n27683 );
or ( n45394 , n15075 , n15076 );
not ( n15077 , RI1754c610_2);
and ( n15078 , n15077 , n45394 );
and ( n15079 , C0 , RI1754c610_2);
or ( n45395 , n15078 , n15079 );
buf ( n45396 , n45395 );
not ( n45397 , n44280 );
xor ( n45398 , n39620 , n35272 );
xor ( n45399 , n45398 , n35009 );
and ( n45400 , n45397 , n45399 );
xor ( n45401 , n44277 , n45400 );
not ( n15080 , n29614 );
and ( n15081 , n15080 , RI174cf300_766);
and ( n15082 , n45401 , n29614 );
or ( n45402 , n15081 , n15082 );
not ( n15083 , RI1754c610_2);
and ( n15084 , n15083 , n45402 );
and ( n15085 , C0 , RI1754c610_2);
or ( n45403 , n15084 , n15085 );
buf ( n45404 , n45403 );
not ( n15086 , n27683 );
and ( n15087 , n15086 , RI19ab3318_2430);
and ( n15088 , RI19abd188_2358 , n27683 );
or ( n45405 , n15087 , n15088 );
not ( n15089 , RI1754c610_2);
and ( n15090 , n15089 , n45405 );
and ( n15091 , C0 , RI1754c610_2);
or ( n45406 , n15090 , n15091 );
buf ( n45407 , n45406 );
not ( n45408 , n41131 );
and ( n45409 , n45408 , n43228 );
xor ( n45410 , n41128 , n45409 );
not ( n15092 , n29614 );
and ( n15093 , n15092 , RI1746ae00_1215);
and ( n15094 , n45410 , n29614 );
or ( n45411 , n15093 , n15094 );
not ( n15095 , RI1754c610_2);
and ( n15096 , n15095 , n45411 );
and ( n15097 , C0 , RI1754c610_2);
or ( n45412 , n15096 , n15097 );
buf ( n45413 , n45412 );
xor ( n45414 , n35059 , n33223 );
xor ( n45415 , n45414 , n33282 );
xor ( n45416 , n31170 , n40828 );
xor ( n45417 , n45416 , n42049 );
not ( n45418 , n45417 );
xor ( n45419 , n41521 , n33824 );
xor ( n45420 , n45419 , n32786 );
and ( n45421 , n45418 , n45420 );
xor ( n45422 , n45415 , n45421 );
not ( n15098 , n29614 );
and ( n15099 , n15098 , RI17475f30_1161);
and ( n15100 , n45422 , n29614 );
or ( n45423 , n15099 , n15100 );
not ( n15101 , RI1754c610_2);
and ( n15102 , n15101 , n45423 );
and ( n15103 , C0 , RI1754c610_2);
or ( n45424 , n15102 , n15103 );
buf ( n45425 , n45424 );
not ( n45426 , n42985 );
and ( n45427 , n45426 , n45172 );
xor ( n45428 , n42982 , n45427 );
not ( n15104 , n29614 );
and ( n15105 , n15104 , RI1748b7b8_1056);
and ( n15106 , n45428 , n29614 );
or ( n45429 , n15105 , n15106 );
not ( n15107 , RI1754c610_2);
and ( n15108 , n15107 , n45429 );
and ( n15109 , C0 , RI1754c610_2);
or ( n45430 , n15108 , n15109 );
buf ( n45431 , n45430 );
not ( n15110 , n27683 );
and ( n15111 , n15110 , RI19aa3c88_2539);
and ( n15112 , RI19aae110_2467 , n27683 );
or ( n45432 , n15111 , n15112 );
not ( n15113 , RI1754c610_2);
and ( n15114 , n15113 , n45432 );
and ( n15115 , C0 , RI1754c610_2);
or ( n45433 , n15114 , n15115 );
buf ( n45434 , n45433 );
buf ( n45435 , RI174a6248_926);
buf ( n45436 , RI1748d1f8_1048);
xor ( n45437 , n39401 , n32403 );
xor ( n45438 , n45437 , n32481 );
xor ( n45439 , n37477 , n42188 );
xor ( n45440 , n45439 , n41526 );
not ( n45441 , n45440 );
and ( n45442 , n45441 , n43057 );
xor ( n45443 , n45438 , n45442 );
not ( n15116 , n29614 );
and ( n15117 , n15116 , RI174709e0_1187);
and ( n15118 , n45443 , n29614 );
or ( n45444 , n15117 , n15118 );
not ( n15119 , RI1754c610_2);
and ( n15120 , n15119 , n45444 );
and ( n15121 , C0 , RI1754c610_2);
or ( n45445 , n15120 , n15121 );
buf ( n45446 , n45445 );
buf ( n45447 , RI174cd938_771);
not ( n15122 , n27683 );
and ( n15123 , n15122 , RI19ac9500_2260);
and ( n15124 , RI19a846f8_2763 , n27683 );
or ( n45448 , n15123 , n15124 );
not ( n15125 , RI1754c610_2);
and ( n15126 , n15125 , n45448 );
and ( n15127 , C0 , RI1754c610_2);
or ( n45449 , n15126 , n15127 );
buf ( n45450 , n45449 );
buf ( n45451 , RI174b0ce8_874);
xor ( n45452 , n39616 , n35272 );
xor ( n45453 , n45452 , n35009 );
not ( n45454 , n45453 );
xor ( n45455 , n41503 , n34445 );
xor ( n45456 , n45455 , n41885 );
and ( n45457 , n45454 , n45456 );
xor ( n45458 , n42076 , n45457 );
not ( n15128 , n29614 );
and ( n15129 , n15128 , RI173ec6e0_1603);
and ( n15130 , n45458 , n29614 );
or ( n45459 , n15129 , n15130 );
not ( n15131 , RI1754c610_2);
and ( n15132 , n15131 , n45459 );
and ( n15133 , C0 , RI1754c610_2);
or ( n45460 , n15132 , n15133 );
buf ( n45461 , n45460 );
xor ( n45462 , n34639 , n34150 );
xor ( n45463 , n45462 , n34190 );
not ( n45464 , n45463 );
xor ( n45465 , n43463 , n40949 );
xor ( n45466 , n45465 , n34572 );
and ( n45467 , n45464 , n45466 );
xor ( n45468 , n40170 , n45467 );
not ( n15134 , n29614 );
and ( n15135 , n15134 , RI17485200_1087);
and ( n15136 , n45468 , n29614 );
or ( n45469 , n15135 , n15136 );
not ( n15137 , RI1754c610_2);
and ( n15138 , n15137 , n45469 );
and ( n15139 , C0 , RI1754c610_2);
or ( n45470 , n15138 , n15139 );
buf ( n45471 , n45470 );
xor ( n45472 , n39612 , n35272 );
xor ( n45473 , n45472 , n35009 );
xor ( n45474 , n38076 , n40091 );
xor ( n45475 , n45474 , n40111 );
not ( n45476 , n45475 );
and ( n45477 , n45476 , n42444 );
xor ( n45478 , n45473 , n45477 );
not ( n15140 , n29614 );
and ( n15141 , n15140 , RI17482410_1101);
and ( n15142 , n45478 , n29614 );
or ( n45479 , n15141 , n15142 );
not ( n15143 , RI1754c610_2);
and ( n15144 , n15143 , n45479 );
and ( n15145 , C0 , RI1754c610_2);
or ( n45480 , n15144 , n15145 );
buf ( n45481 , n45480 );
xor ( n45482 , n34291 , n38886 );
xor ( n45483 , n45482 , n39604 );
xor ( n45484 , n32972 , n41659 );
xor ( n45485 , n45484 , n37800 );
not ( n45486 , n45485 );
xor ( n45487 , n33038 , n36227 );
xor ( n45488 , n45487 , n40743 );
and ( n45489 , n45486 , n45488 );
xor ( n45490 , n45483 , n45489 );
not ( n15146 , n29614 );
and ( n15147 , n15146 , RI173b3350_1882);
and ( n15148 , n45490 , n29614 );
or ( n45491 , n15147 , n15148 );
not ( n15149 , RI1754c610_2);
and ( n15150 , n15149 , n45491 );
and ( n15151 , C0 , RI1754c610_2);
or ( n45492 , n15150 , n15151 );
buf ( n45493 , n45492 );
not ( n15152 , n27683 );
and ( n15153 , n15152 , RI19aacdd8_2476);
and ( n15154 , RI19ab6900_2405 , n27683 );
or ( n45494 , n15153 , n15154 );
not ( n15155 , RI1754c610_2);
and ( n15156 , n15155 , n45494 );
and ( n15157 , C0 , RI1754c610_2);
or ( n45495 , n15156 , n15157 );
buf ( n45496 , n45495 );
xor ( n45497 , n42935 , n29425 );
xor ( n45498 , n45497 , n29610 );
xor ( n45499 , n40350 , n37898 );
xor ( n45500 , n45499 , n37915 );
not ( n45501 , n45500 );
and ( n45502 , n45501 , n38116 );
xor ( n45503 , n45498 , n45502 );
not ( n15158 , n29614 );
and ( n15159 , n15158 , RI1740da70_1441);
and ( n15160 , n45503 , n29614 );
or ( n45504 , n15159 , n15160 );
not ( n15161 , RI1754c610_2);
and ( n15162 , n15161 , n45504 );
and ( n15163 , C0 , RI1754c610_2);
or ( n45505 , n15162 , n15163 );
buf ( n45506 , n45505 );
not ( n45507 , n42740 );
and ( n45508 , n45507 , n43680 );
xor ( n45509 , n42737 , n45508 );
not ( n15164 , n29614 );
and ( n15165 , n15164 , RI1740ee20_1435);
and ( n15166 , n45509 , n29614 );
or ( n45510 , n15165 , n15166 );
not ( n15167 , RI1754c610_2);
and ( n15168 , n15167 , n45510 );
and ( n15169 , C0 , RI1754c610_2);
or ( n45511 , n15168 , n15169 );
buf ( n45512 , n45511 );
xor ( n45513 , n36376 , n38676 );
xor ( n45514 , n45513 , n28111 );
xor ( n45515 , n34158 , n42264 );
xor ( n45516 , n45515 , n41370 );
not ( n45517 , n45516 );
xor ( n45518 , n40021 , n40855 );
xor ( n45519 , n45518 , n38574 );
and ( n45520 , n45517 , n45519 );
xor ( n45521 , n45514 , n45520 );
not ( n15170 , n29614 );
and ( n15171 , n15170 , RI174050a0_1483);
and ( n15172 , n45521 , n29614 );
or ( n45522 , n15171 , n15172 );
not ( n15173 , RI1754c610_2);
and ( n15174 , n15173 , n45522 );
and ( n15175 , C0 , RI1754c610_2);
or ( n45523 , n15174 , n15175 );
buf ( n45524 , n45523 );
not ( n15176 , n27683 );
and ( n15177 , n15176 , RI19aafad8_2456);
and ( n15178 , RI19ab96f0_2385 , n27683 );
or ( n45525 , n15177 , n15178 );
not ( n15179 , RI1754c610_2);
and ( n15180 , n15179 , n45525 );
and ( n15181 , C0 , RI1754c610_2);
or ( n45526 , n15180 , n15181 );
buf ( n45527 , n45526 );
xor ( n45528 , n39790 , n33175 );
xor ( n45529 , n45528 , n34797 );
xor ( n45530 , n40447 , n35911 );
xor ( n45531 , n45530 , n38188 );
not ( n45532 , n45531 );
xor ( n45533 , n40273 , n37623 );
xor ( n45534 , n45533 , n37651 );
and ( n45535 , n45532 , n45534 );
xor ( n45536 , n45529 , n45535 );
not ( n15182 , n29614 );
and ( n15183 , n15182 , RI17407b48_1470);
and ( n15184 , n45536 , n29614 );
or ( n45537 , n15183 , n15184 );
not ( n15185 , RI1754c610_2);
and ( n15186 , n15185 , n45537 );
and ( n15187 , C0 , RI1754c610_2);
or ( n45538 , n15186 , n15187 );
buf ( n45539 , n45538 );
xor ( n45540 , n27795 , n42344 );
xor ( n45541 , n45540 , n41799 );
xor ( n45542 , n37560 , n34968 );
xor ( n45543 , n45542 , n39771 );
not ( n45544 , n45543 );
xor ( n45545 , n41766 , n38188 );
xor ( n45546 , n45545 , n36195 );
and ( n45547 , n45544 , n45546 );
xor ( n45548 , n45541 , n45547 );
not ( n15188 , n29614 );
and ( n15189 , n15188 , RI173d1908_1734);
and ( n15190 , n45548 , n29614 );
or ( n45549 , n15189 , n15190 );
not ( n15191 , RI1754c610_2);
and ( n15192 , n15191 , n45549 );
and ( n15193 , C0 , RI1754c610_2);
or ( n45550 , n15192 , n15193 );
buf ( n45551 , n45550 );
not ( n15194 , n27683 );
and ( n15195 , n15194 , RI19a9a160_2611);
and ( n15196 , RI19aa38c8_2541 , n27683 );
or ( n45552 , n15195 , n15196 );
not ( n15197 , RI1754c610_2);
and ( n15198 , n15197 , n45552 );
and ( n15199 , C0 , RI1754c610_2);
or ( n45553 , n15198 , n15199 );
buf ( n45554 , n45553 );
not ( n45555 , n44229 );
xor ( n45556 , n40314 , n37869 );
xor ( n45557 , n45556 , n38948 );
and ( n45558 , n45555 , n45557 );
xor ( n45559 , n44226 , n45558 );
not ( n15200 , n29614 );
and ( n15201 , n15200 , RI1747bb10_1133);
and ( n15202 , n45559 , n29614 );
or ( n45560 , n15201 , n15202 );
not ( n15203 , RI1754c610_2);
and ( n15204 , n15203 , n45560 );
and ( n15205 , C0 , RI1754c610_2);
or ( n45561 , n15204 , n15205 );
buf ( n45562 , n45561 );
not ( n45563 , n42117 );
xor ( n45564 , n43987 , n40808 );
xor ( n45565 , n45564 , n40828 );
and ( n45566 , n45563 , n45565 );
xor ( n45567 , n42114 , n45566 );
not ( n15206 , n29614 );
and ( n15207 , n15206 , RI17406e28_1474);
and ( n15208 , n45567 , n29614 );
or ( n45568 , n15207 , n15208 );
not ( n15209 , RI1754c610_2);
and ( n15210 , n15209 , n45568 );
and ( n15211 , C0 , RI1754c610_2);
or ( n45569 , n15210 , n15211 );
buf ( n45570 , n45569 );
xor ( n45571 , n38388 , n37169 );
xor ( n45572 , n45571 , n36339 );
not ( n45573 , n45572 );
and ( n45574 , n45573 , n42678 );
xor ( n45575 , n44419 , n45574 );
not ( n15212 , n29614 );
and ( n15213 , n15212 , RI173cee48_1747);
and ( n15214 , n45575 , n29614 );
or ( n45576 , n15213 , n15214 );
not ( n15215 , RI1754c610_2);
and ( n15216 , n15215 , n45576 );
and ( n15217 , C0 , RI1754c610_2);
or ( n45577 , n15216 , n15217 );
buf ( n45578 , n45577 );
buf ( n45579 , RI1749cea0_971);
buf ( n45580 , RI1749cb58_972);
buf ( n45581 , RI17493af8_1016);
buf ( n45582 , RI17487ca8_1074);
buf ( n45583 , RI17461da0_1259);
buf ( n45584 , RI174613c8_1262);
buf ( n45585 , RI17506bd8_745);
buf ( n45586 , RI174c9630_784);
xor ( n45587 , n40679 , n36654 );
xor ( n45588 , n45587 , n40808 );
not ( n45589 , n45588 );
xor ( n45590 , n34173 , n42264 );
xor ( n45591 , n45590 , n41370 );
and ( n45592 , n45589 , n45591 );
xor ( n45593 , n43165 , n45592 );
not ( n15218 , n29614 );
and ( n15219 , n15218 , RI17410ba8_1426);
and ( n15220 , n45593 , n29614 );
or ( n45594 , n15219 , n15220 );
not ( n15221 , RI1754c610_2);
and ( n15222 , n15221 , n45594 );
and ( n15223 , C0 , RI1754c610_2);
or ( n45595 , n15222 , n15223 );
buf ( n45596 , n45595 );
buf ( n45597 , RI174b68c8_846);
buf ( n45598 , RI1749c810_973);
buf ( n45599 , RI174a7c88_918);
buf ( n45600 , RI1748c820_1051);
buf ( n45601 , RI17503398_750);
xor ( n45602 , n34110 , n42377 );
xor ( n45603 , n45602 , n33991 );
not ( n45604 , n43566 );
and ( n45605 , n45604 , n43568 );
xor ( n45606 , n45603 , n45605 );
not ( n15224 , n29614 );
and ( n15225 , n15224 , RI1739b020_2000);
and ( n15226 , n45606 , n29614 );
or ( n45607 , n15225 , n15226 );
not ( n15227 , RI1754c610_2);
and ( n15228 , n15227 , n45607 );
and ( n15229 , C0 , RI1754c610_2);
or ( n45608 , n15228 , n15229 );
buf ( n45609 , n45608 );
buf ( n45610 , RI174af2a8_882);
xor ( n45611 , n36450 , n37104 );
xor ( n45612 , n45611 , n35986 );
xor ( n45613 , n33721 , n35514 );
xor ( n45614 , n45613 , n40486 );
not ( n45615 , n45614 );
xor ( n45616 , n37525 , n37942 );
xor ( n45617 , n45616 , n34395 );
and ( n45618 , n45615 , n45617 );
xor ( n45619 , n45612 , n45618 );
not ( n15230 , n29614 );
and ( n15231 , n15230 , RI17483478_1096);
and ( n15232 , n45619 , n29614 );
or ( n45620 , n15231 , n15232 );
not ( n15233 , RI1754c610_2);
and ( n15234 , n15233 , n45620 );
and ( n15235 , C0 , RI1754c610_2);
or ( n45621 , n15234 , n15235 );
buf ( n45622 , n45621 );
xor ( n45623 , n41770 , n38188 );
xor ( n45624 , n45623 , n36195 );
xor ( n45625 , n38675 , n39347 );
xor ( n45626 , n45625 , n42344 );
not ( n45627 , n45626 );
xor ( n45628 , n41516 , n33824 );
xor ( n45629 , n45628 , n32786 );
and ( n45630 , n45627 , n45629 );
xor ( n45631 , n45624 , n45630 );
not ( n15236 , n29614 );
and ( n15237 , n15236 , RI1751e968_671);
and ( n15238 , n45631 , n29614 );
or ( n45632 , n15237 , n15238 );
not ( n15239 , RI1754c610_2);
and ( n15240 , n15239 , n45632 );
and ( n15241 , C0 , RI1754c610_2);
or ( n45633 , n15240 , n15241 );
buf ( n45634 , n45633 );
not ( n15242 , n27683 );
and ( n15243 , n15242 , RI19a8cd80_2705);
and ( n15244 , RI19a97028_2633 , n27683 );
or ( n45635 , n15243 , n15244 );
not ( n15245 , RI1754c610_2);
and ( n15246 , n15245 , n45635 );
and ( n15247 , C0 , RI1754c610_2);
or ( n45636 , n15246 , n15247 );
buf ( n45637 , n45636 );
not ( n15248 , n27683 );
and ( n15249 , n15248 , RI19aa3418_2543);
and ( n15250 , RI19aad648_2472 , n27683 );
or ( n45638 , n15249 , n15250 );
not ( n15251 , RI1754c610_2);
and ( n15252 , n15251 , n45638 );
and ( n15253 , C0 , RI1754c610_2);
or ( n45639 , n15252 , n15253 );
buf ( n45640 , n45639 );
not ( n45641 , n42051 );
xor ( n45642 , n40708 , n39333 );
xor ( n45643 , n45642 , n39347 );
and ( n45644 , n45641 , n45643 );
xor ( n45645 , n42035 , n45644 );
not ( n15254 , n29614 );
and ( n15255 , n15254 , RI17409588_1462);
and ( n15256 , n45645 , n29614 );
or ( n45646 , n15255 , n15256 );
not ( n15257 , RI1754c610_2);
and ( n15258 , n15257 , n45646 );
and ( n15259 , C0 , RI1754c610_2);
or ( n45647 , n15258 , n15259 );
buf ( n45648 , n45647 );
not ( n45649 , n41964 );
xor ( n45650 , n32058 , n36702 );
xor ( n45651 , n45650 , n38872 );
and ( n45652 , n45649 , n45651 );
xor ( n45653 , n41961 , n45652 );
not ( n15260 , n29614 );
and ( n15261 , n15260 , RI17499a20_987);
and ( n15262 , n45653 , n29614 );
or ( n45654 , n15261 , n15262 );
not ( n15263 , RI1754c610_2);
and ( n15264 , n15263 , n45654 );
and ( n15265 , C0 , RI1754c610_2);
or ( n45655 , n15264 , n15265 );
buf ( n45656 , n45655 );
not ( n45657 , n43381 );
and ( n45658 , n45657 , n43383 );
xor ( n45659 , n41910 , n45658 );
not ( n15266 , n29614 );
and ( n15267 , n15266 , RI173c5410_1794);
and ( n15268 , n45659 , n29614 );
or ( n45660 , n15267 , n15268 );
not ( n15269 , RI1754c610_2);
and ( n15270 , n15269 , n45660 );
and ( n15271 , C0 , RI1754c610_2);
or ( n45661 , n15270 , n15271 );
buf ( n45662 , n45661 );
not ( n15272 , n27683 );
and ( n15273 , n15272 , RI19ab98d0_2384);
and ( n15274 , RI19ac2390_2312 , n27683 );
or ( n45663 , n15273 , n15274 );
not ( n15275 , RI1754c610_2);
and ( n15276 , n15275 , n45663 );
and ( n15277 , C0 , RI1754c610_2);
or ( n45664 , n15276 , n15277 );
buf ( n45665 , n45664 );
xor ( n45666 , n34467 , n33453 );
xor ( n45667 , n45666 , n33505 );
xor ( n45668 , n39982 , n41934 );
xor ( n45669 , n45668 , n40341 );
not ( n45670 , n45669 );
xor ( n45671 , n37459 , n36874 );
xor ( n45672 , n45671 , n42188 );
and ( n45673 , n45670 , n45672 );
xor ( n45674 , n45667 , n45673 );
not ( n15278 , n29614 );
and ( n15279 , n15278 , RI1739f850_1978);
and ( n15280 , n45674 , n29614 );
or ( n45675 , n15279 , n15280 );
not ( n15281 , RI1754c610_2);
and ( n15282 , n15281 , n45675 );
and ( n15283 , C0 , RI1754c610_2);
or ( n45676 , n15282 , n15283 );
buf ( n45677 , n45676 );
xor ( n45678 , n32654 , n36195 );
xor ( n45679 , n45678 , n36209 );
not ( n45680 , n45679 );
and ( n45681 , n45680 , n40544 );
xor ( n45682 , n43188 , n45681 );
not ( n15284 , n29614 );
and ( n15285 , n15284 , RI174889c8_1070);
and ( n15286 , n45682 , n29614 );
or ( n45683 , n15285 , n15286 );
not ( n15287 , RI1754c610_2);
and ( n15288 , n15287 , n45683 );
and ( n15289 , C0 , RI1754c610_2);
or ( n45684 , n15288 , n15289 );
buf ( n45685 , n45684 );
xor ( n45686 , n38617 , n38347 );
xor ( n45687 , n45686 , n34300 );
not ( n45688 , n45687 );
xor ( n45689 , n38506 , n31664 );
xor ( n45690 , n45689 , n31725 );
and ( n45691 , n45688 , n45690 );
xor ( n45692 , n44529 , n45691 );
not ( n15290 , n29614 );
and ( n15291 , n15290 , RI1740e448_1438);
and ( n15292 , n45692 , n29614 );
or ( n45693 , n15291 , n15292 );
not ( n15293 , RI1754c610_2);
and ( n15294 , n15293 , n45693 );
and ( n15295 , C0 , RI1754c610_2);
or ( n45694 , n15294 , n15295 );
buf ( n45695 , n45694 );
buf ( n45696 , RI174b6c10_845);
buf ( n45697 , RI1749c4c8_974);
xor ( n45698 , n38102 , n40111 );
xor ( n45699 , n45698 , n43278 );
not ( n45700 , n36412 );
and ( n45701 , n45700 , n36433 );
xor ( n45702 , n45699 , n45701 );
not ( n15296 , n29614 );
and ( n15297 , n15296 , RI1750d2f8_725);
and ( n15298 , n45702 , n29614 );
or ( n45703 , n15297 , n15298 );
not ( n15299 , RI1754c610_2);
and ( n15300 , n15299 , n45703 );
and ( n15301 , C0 , RI1754c610_2);
or ( n45704 , n15300 , n15301 );
buf ( n45705 , n45704 );
not ( n15302 , n27683 );
and ( n15303 , n15302 , RI19aa0b50_2563);
and ( n15304 , RI19aaaa38_2491 , n27683 );
or ( n45706 , n15303 , n15304 );
not ( n15305 , RI1754c610_2);
and ( n15306 , n15305 , n45706 );
and ( n15307 , C0 , RI1754c610_2);
or ( n45707 , n15306 , n15307 );
buf ( n45708 , n45707 );
not ( n45709 , n41700 );
and ( n45710 , n45709 , n41702 );
xor ( n45711 , n45157 , n45710 );
not ( n15308 , n29614 );
and ( n15309 , n15308 , RI173b8210_1858);
and ( n15310 , n45711 , n29614 );
or ( n45712 , n15309 , n15310 );
not ( n15311 , RI1754c610_2);
and ( n15312 , n15311 , n45712 );
and ( n15313 , C0 , RI1754c610_2);
or ( n45713 , n15312 , n15313 );
buf ( n45714 , n45713 );
xor ( n45715 , n37425 , n34725 );
xor ( n45716 , n45715 , n34755 );
xor ( n45717 , n32952 , n41659 );
xor ( n45718 , n45717 , n37800 );
not ( n45719 , n45718 );
xor ( n45720 , n35537 , n37460 );
xor ( n45721 , n45720 , n37490 );
and ( n45722 , n45719 , n45721 );
xor ( n45723 , n45716 , n45722 );
not ( n15314 , n29614 );
and ( n15315 , n15314 , RI174b8f38_835);
and ( n15316 , n45723 , n29614 );
or ( n45724 , n15315 , n15316 );
not ( n15317 , RI1754c610_2);
and ( n15318 , n15317 , n45724 );
and ( n15319 , C0 , RI1754c610_2);
or ( n45725 , n15318 , n15319 );
buf ( n45726 , n45725 );
xor ( n45727 , n43262 , n41099 );
xor ( n45728 , n45727 , n30604 );
xor ( n45729 , n36823 , n44146 );
xor ( n45730 , n45729 , n41198 );
not ( n45731 , n45730 );
xor ( n45732 , n35890 , n36463 );
xor ( n45733 , n45732 , n32220 );
and ( n45734 , n45731 , n45733 );
xor ( n45735 , n45728 , n45734 );
not ( n15320 , n29614 );
and ( n15321 , n15320 , RI17344860_2107);
and ( n15322 , n45735 , n29614 );
or ( n45736 , n15321 , n15322 );
not ( n15323 , RI1754c610_2);
and ( n15324 , n15323 , n45736 );
and ( n15325 , C0 , RI1754c610_2);
or ( n45737 , n15324 , n15325 );
buf ( n45738 , n45737 );
not ( n45739 , n43935 );
and ( n45740 , n45739 , n43937 );
xor ( n45741 , n39221 , n45740 );
not ( n15326 , n29614 );
and ( n15327 , n15326 , RI17402fd0_1493);
and ( n15328 , n45741 , n29614 );
or ( n45742 , n15327 , n15328 );
not ( n15329 , RI1754c610_2);
and ( n15330 , n15329 , n45742 );
and ( n15331 , C0 , RI1754c610_2);
or ( n45743 , n15330 , n15331 );
buf ( n45744 , n45743 );
not ( n15332 , n27683 );
and ( n15333 , n15332 , RI19a8dd70_2698);
and ( n15334 , RI19a97dc0_2627 , n27683 );
or ( n45745 , n15333 , n15334 );
not ( n15335 , RI1754c610_2);
and ( n15336 , n15335 , n45745 );
and ( n15337 , C0 , RI1754c610_2);
or ( n45746 , n15336 , n15337 );
buf ( n45747 , n45746 );
not ( n15338 , n27683 );
and ( n15339 , n15338 , RI19ab3138_2431);
and ( n15340 , RI19abcdc8_2360 , n27683 );
or ( n45748 , n15339 , n15340 );
not ( n15341 , RI1754c610_2);
and ( n15342 , n15341 , n45748 );
and ( n15343 , C0 , RI1754c610_2);
or ( n45749 , n15342 , n15343 );
buf ( n45750 , n45749 );
xor ( n45751 , n40795 , n40437 );
xor ( n45752 , n45751 , n42635 );
not ( n45753 , n45752 );
xor ( n45754 , n36395 , n34190 );
xor ( n45755 , n45754 , n36252 );
and ( n45756 , n45753 , n45755 );
xor ( n45757 , n43402 , n45756 );
not ( n15344 , n29614 );
and ( n15345 , n15344 , RI174b5518_852);
and ( n15346 , n45757 , n29614 );
or ( n45758 , n15345 , n15346 );
not ( n15347 , RI1754c610_2);
and ( n15348 , n15347 , n45758 );
and ( n15349 , C0 , RI1754c610_2);
or ( n45759 , n15348 , n15349 );
buf ( n45760 , n45759 );
xor ( n45761 , n40909 , n34797 );
xor ( n45762 , n45761 , n34837 );
not ( n45763 , n45762 );
xor ( n45764 , n40297 , n37849 );
xor ( n45765 , n45764 , n37869 );
and ( n45766 , n45763 , n45765 );
xor ( n45767 , n44394 , n45766 );
not ( n15350 , n29614 );
and ( n15351 , n15350 , RI174c29e8_805);
and ( n15352 , n45767 , n29614 );
or ( n45768 , n15351 , n15352 );
not ( n15353 , RI1754c610_2);
and ( n15354 , n15353 , n45768 );
and ( n15355 , C0 , RI1754c610_2);
or ( n45769 , n15354 , n15355 );
buf ( n45770 , n45769 );
not ( n45771 , n43371 );
and ( n45772 , n45771 , n43373 );
xor ( n45773 , n41393 , n45772 );
not ( n15356 , n29614 );
and ( n15357 , n15356 , RI1748f2c8_1038);
and ( n15358 , n45773 , n29614 );
or ( n45774 , n15357 , n15358 );
not ( n15359 , RI1754c610_2);
and ( n15360 , n15359 , n45774 );
and ( n15361 , C0 , RI1754c610_2);
or ( n45775 , n15360 , n15361 );
buf ( n45776 , n45775 );
buf ( n45777 , RI174689e8_1226);
xor ( n45778 , n33242 , n40302 );
xor ( n45779 , n45778 , n40319 );
not ( n45780 , n45779 );
xor ( n45781 , n35967 , n37744 );
xor ( n45782 , n45781 , n35438 );
and ( n45783 , n45780 , n45782 );
xor ( n45784 , n43727 , n45783 );
not ( n15362 , n29614 );
and ( n15363 , n15362 , RI173ddaa0_1675);
and ( n15364 , n45784 , n29614 );
or ( n45785 , n15363 , n15364 );
not ( n15365 , RI1754c610_2);
and ( n15366 , n15365 , n45785 );
and ( n15367 , C0 , RI1754c610_2);
or ( n45786 , n15366 , n15367 );
buf ( n45787 , n45786 );
xor ( n45788 , n34788 , n37255 );
xor ( n45789 , n45788 , n41478 );
xor ( n45790 , n41098 , n38150 );
xor ( n45791 , n45790 , n38167 );
not ( n45792 , n45791 );
xor ( n45793 , n41974 , n39886 );
xor ( n45794 , n45793 , n36998 );
and ( n45795 , n45792 , n45794 );
xor ( n45796 , n45789 , n45795 );
not ( n15368 , n29614 );
and ( n15369 , n15368 , RI173acd98_1913);
and ( n15370 , n45796 , n29614 );
or ( n45797 , n15369 , n15370 );
not ( n15371 , RI1754c610_2);
and ( n15372 , n15371 , n45797 );
and ( n15373 , C0 , RI1754c610_2);
or ( n45798 , n15372 , n15373 );
buf ( n45799 , n45798 );
not ( n15374 , n27683 );
and ( n15375 , n15374 , RI19ace870_2221);
and ( n15376 , RI19a99ad0_2614 , n27683 );
or ( n45800 , n15375 , n15376 );
not ( n15377 , RI1754c610_2);
and ( n15378 , n15377 , n45800 );
and ( n15379 , C0 , RI1754c610_2);
or ( n45801 , n15378 , n15379 );
buf ( n45802 , n45801 );
xor ( n45803 , n29860 , n36128 );
xor ( n45804 , n45803 , n36148 );
xor ( n45805 , n39169 , n40166 );
xor ( n45806 , n45805 , n41590 );
not ( n45807 , n45806 );
xor ( n45808 , n31567 , n39935 );
xor ( n45809 , n45808 , n39952 );
and ( n45810 , n45807 , n45809 );
xor ( n45811 , n45804 , n45810 );
not ( n15380 , n29614 );
and ( n15381 , n15380 , RI17412930_1417);
and ( n15382 , n45811 , n29614 );
or ( n45812 , n15381 , n15382 );
not ( n15383 , RI1754c610_2);
and ( n15384 , n15383 , n45812 );
and ( n15385 , C0 , RI1754c610_2);
or ( n45813 , n15384 , n15385 );
buf ( n45814 , n45813 );
buf ( n45815 , RI174b6f58_844);
buf ( n45816 , RI1749be38_976);
not ( n45817 , n42138 );
xor ( n45818 , n42304 , n40769 );
xor ( n45819 , n45818 , n40949 );
and ( n45820 , n45817 , n45819 );
xor ( n45821 , n42135 , n45820 );
not ( n15386 , n29614 );
and ( n15387 , n15386 , RI173d9f90_1693);
and ( n15388 , n45821 , n29614 );
or ( n45822 , n15387 , n15388 );
not ( n15389 , RI1754c610_2);
and ( n15390 , n15389 , n45822 );
and ( n15391 , C0 , RI1754c610_2);
or ( n45823 , n15390 , n15391 );
buf ( n45824 , n45823 );
xor ( n45825 , n39930 , n40890 );
xor ( n45826 , n45825 , n38724 );
xor ( n45827 , n34189 , n42264 );
xor ( n45828 , n45827 , n41370 );
not ( n45829 , n45828 );
xor ( n45830 , n41674 , n41885 );
xor ( n45831 , n45830 , n30923 );
and ( n45832 , n45829 , n45831 );
xor ( n45833 , n45826 , n45832 );
not ( n15392 , n29614 );
and ( n15393 , n15392 , RI17495bc8_1006);
and ( n15394 , n45833 , n29614 );
or ( n45834 , n15393 , n15394 );
not ( n15395 , RI1754c610_2);
and ( n15396 , n15395 , n45834 );
and ( n15397 , C0 , RI1754c610_2);
or ( n45835 , n15396 , n15397 );
buf ( n45836 , n45835 );
not ( n45837 , n42381 );
xor ( n45838 , n40241 , n35760 );
xor ( n45839 , n45838 , n39333 );
and ( n45840 , n45837 , n45839 );
xor ( n45841 , n42378 , n45840 );
not ( n15398 , n29614 );
and ( n15399 , n15398 , RI175298b8_637);
and ( n15400 , n45841 , n29614 );
or ( n45842 , n15399 , n15400 );
not ( n15401 , RI1754c610_2);
and ( n15402 , n15401 , n45842 );
and ( n15403 , C0 , RI1754c610_2);
or ( n45843 , n15402 , n15403 );
buf ( n45844 , n45843 );
xor ( n45845 , n33484 , n40360 );
xor ( n45846 , n45845 , n35176 );
xor ( n45847 , n32097 , n36702 );
xor ( n45848 , n45847 , n38872 );
not ( n45849 , n45848 );
and ( n45850 , n45849 , n44886 );
xor ( n45851 , n45846 , n45850 );
not ( n15404 , n29614 );
and ( n15405 , n15404 , RI1745d570_1281);
and ( n15406 , n45851 , n29614 );
or ( n45852 , n15405 , n15406 );
not ( n15407 , RI1754c610_2);
and ( n15408 , n15407 , n45852 );
and ( n15409 , C0 , RI1754c610_2);
or ( n45853 , n15408 , n15409 );
buf ( n45854 , n45853 );
xor ( n45855 , n37606 , n40319 );
xor ( n45856 , n45855 , n40149 );
not ( n45857 , n43304 );
and ( n45858 , n45857 , n40621 );
xor ( n45859 , n45856 , n45858 );
not ( n15410 , n29614 );
and ( n15411 , n15410 , RI17467cc8_1230);
and ( n15412 , n45859 , n29614 );
or ( n45860 , n15411 , n15412 );
not ( n15413 , RI1754c610_2);
and ( n15414 , n15413 , n45860 );
and ( n15415 , C0 , RI1754c610_2);
or ( n45861 , n15414 , n15415 );
buf ( n45862 , n45861 );
not ( n45863 , n29611 );
and ( n45864 , n45863 , n44557 );
xor ( n45865 , n29110 , n45864 );
not ( n15416 , n29614 );
and ( n15417 , n15416 , RI17473e60_1171);
and ( n15418 , n45865 , n29614 );
or ( n45866 , n15417 , n15418 );
not ( n15419 , RI1754c610_2);
and ( n15420 , n15419 , n45866 );
and ( n15421 , C0 , RI1754c610_2);
or ( n45867 , n15420 , n15421 );
buf ( n45868 , n45867 );
not ( n15422 , n27683 );
and ( n15423 , n15422 , RI19abb748_2371);
and ( n15424 , RI19ac40a0_2299 , n27683 );
or ( n45869 , n15423 , n15424 );
not ( n15425 , RI1754c610_2);
and ( n15426 , n15425 , n45869 );
and ( n15427 , C0 , RI1754c610_2);
or ( n45870 , n15426 , n15427 );
buf ( n45871 , n45870 );
xor ( n45872 , n41739 , n34837 );
xor ( n45873 , n45872 , n33880 );
xor ( n45874 , n29478 , n40051 );
xor ( n45875 , n45874 , n37074 );
not ( n45876 , n45875 );
xor ( n45877 , n33474 , n40360 );
xor ( n45878 , n45877 , n35176 );
and ( n45879 , n45876 , n45878 );
xor ( n45880 , n45873 , n45879 );
not ( n15428 , n29614 );
and ( n15429 , n15428 , RI17334f00_2183);
and ( n15430 , n45880 , n29614 );
or ( n45881 , n15429 , n15430 );
not ( n15431 , RI1754c610_2);
and ( n15432 , n15431 , n45881 );
and ( n15433 , C0 , RI1754c610_2);
or ( n45882 , n15432 , n15433 );
buf ( n45883 , n45882 );
not ( n45884 , n45420 );
xor ( n45885 , n38511 , n31664 );
xor ( n45886 , n45885 , n31725 );
and ( n45887 , n45884 , n45886 );
xor ( n45888 , n45417 , n45887 );
not ( n15434 , n29614 );
and ( n15435 , n15434 , RI17484828_1090);
and ( n15436 , n45888 , n29614 );
or ( n45889 , n15435 , n15436 );
not ( n15437 , RI1754c610_2);
and ( n15438 , n15437 , n45889 );
and ( n15439 , C0 , RI1754c610_2);
or ( n45890 , n15438 , n15439 );
buf ( n45891 , n45890 );
not ( n15440 , n27683 );
and ( n15441 , n15440 , RI19abd6b0_2355);
and ( n15442 , RI19ac6080_2284 , n27683 );
or ( n45892 , n15441 , n15442 );
not ( n15443 , RI1754c610_2);
and ( n15444 , n15443 , n45892 );
and ( n15445 , C0 , RI1754c610_2);
or ( n45893 , n15444 , n15445 );
buf ( n45894 , n45893 );
xor ( n45895 , n38540 , n35458 );
xor ( n45896 , n45895 , n40692 );
not ( n45897 , n43821 );
and ( n45898 , n45897 , n43823 );
xor ( n45899 , n45896 , n45898 );
not ( n15446 , n29614 );
and ( n15447 , n15446 , RI173988c0_2012);
and ( n15448 , n45899 , n29614 );
or ( n45900 , n15447 , n15448 );
not ( n15449 , RI1754c610_2);
and ( n15450 , n15449 , n45900 );
and ( n15451 , C0 , RI1754c610_2);
or ( n45901 , n15450 , n15451 );
buf ( n45902 , n45901 );
not ( n45903 , n44308 );
xor ( n45904 , n39867 , n42504 );
xor ( n45905 , n45904 , n41818 );
and ( n45906 , n45903 , n45905 );
xor ( n45907 , n44305 , n45906 );
not ( n15452 , n29614 );
and ( n15453 , n15452 , RI1740ac80_1455);
and ( n15454 , n45907 , n29614 );
or ( n45908 , n15453 , n15454 );
not ( n15455 , RI1754c610_2);
and ( n15456 , n15455 , n45908 );
and ( n15457 , C0 , RI1754c610_2);
or ( n45909 , n15456 , n15457 );
buf ( n45910 , n45909 );
xor ( n45911 , n36360 , n38676 );
xor ( n45912 , n45911 , n28111 );
xor ( n45913 , n40458 , n35911 );
xor ( n45914 , n45913 , n38188 );
not ( n45915 , n45914 );
and ( n45916 , n45915 , n43094 );
xor ( n45917 , n45912 , n45916 );
not ( n15458 , n29614 );
and ( n15459 , n15458 , RI173a6150_1946);
and ( n15460 , n45917 , n29614 );
or ( n45918 , n15459 , n15460 );
not ( n15461 , RI1754c610_2);
and ( n15462 , n15461 , n45918 );
and ( n15463 , C0 , RI1754c610_2);
or ( n45919 , n15462 , n15463 );
buf ( n45920 , n45919 );
xor ( n45921 , n42248 , n40743 );
xor ( n45922 , n45921 , n36062 );
xor ( n45923 , n43451 , n40949 );
xor ( n45924 , n45923 , n34572 );
not ( n45925 , n45924 );
xor ( n45926 , n37566 , n34968 );
xor ( n45927 , n45926 , n39771 );
and ( n45928 , n45925 , n45927 );
xor ( n45929 , n45922 , n45928 );
not ( n15464 , n29614 );
and ( n15465 , n15464 , RI174af938_880);
and ( n15466 , n45929 , n29614 );
or ( n45930 , n15465 , n15466 );
not ( n15467 , RI1754c610_2);
and ( n15468 , n15467 , n45930 );
and ( n15469 , C0 , RI1754c610_2);
or ( n45931 , n15468 , n15469 );
buf ( n45932 , n45931 );
xor ( n45933 , n38275 , n36568 );
xor ( n45934 , n45933 , n36742 );
not ( n45935 , n41639 );
and ( n45936 , n45935 , n41660 );
xor ( n45937 , n45934 , n45936 );
not ( n15470 , n29614 );
and ( n15471 , n15470 , RI173e4d78_1640);
and ( n15472 , n45937 , n29614 );
or ( n45938 , n15471 , n15472 );
not ( n15473 , RI1754c610_2);
and ( n15474 , n15473 , n45938 );
and ( n15475 , C0 , RI1754c610_2);
or ( n45939 , n15474 , n15475 );
buf ( n45940 , n45939 );
xor ( n45941 , n35474 , n38512 );
xor ( n45942 , n45941 , n38532 );
xor ( n45943 , n38271 , n36568 );
xor ( n45944 , n45943 , n36742 );
not ( n45945 , n45944 );
xor ( n45946 , n40372 , n42554 );
xor ( n45947 , n45946 , n34725 );
and ( n45948 , n45945 , n45947 );
xor ( n45949 , n45942 , n45948 );
not ( n15476 , n29614 );
and ( n15477 , n15476 , RI1746aab8_1216);
and ( n15478 , n45949 , n29614 );
or ( n45950 , n15477 , n15478 );
not ( n15479 , RI1754c610_2);
and ( n15480 , n15479 , n45950 );
and ( n15481 , C0 , RI1754c610_2);
or ( n45951 , n15480 , n15481 );
buf ( n45952 , n45951 );
xor ( n45953 , n38544 , n35458 );
xor ( n45954 , n45953 , n40692 );
not ( n45955 , n44971 );
and ( n45956 , n45955 , n44973 );
xor ( n45957 , n45954 , n45956 );
not ( n15482 , n29614 );
and ( n15483 , n15482 , RI17483e50_1093);
and ( n15484 , n45957 , n29614 );
or ( n45958 , n15483 , n15484 );
not ( n15485 , RI1754c610_2);
and ( n15486 , n15485 , n45958 );
and ( n15487 , C0 , RI1754c610_2);
or ( n45959 , n15486 , n15487 );
buf ( n45960 , n45959 );
xor ( n45961 , n41689 , n41885 );
xor ( n45962 , n45961 , n30923 );
not ( n45963 , n36743 );
and ( n45964 , n45963 , n36803 );
xor ( n45965 , n45962 , n45964 );
not ( n15488 , n29614 );
and ( n15489 , n15488 , RI173bb000_1844);
and ( n15490 , n45965 , n29614 );
or ( n45966 , n15489 , n15490 );
not ( n15491 , RI1754c610_2);
and ( n15492 , n15491 , n45966 );
and ( n15493 , C0 , RI1754c610_2);
or ( n45967 , n15492 , n15493 );
buf ( n45968 , n45967 );
not ( n15494 , n27683 );
and ( n15495 , n15494 , RI19abcdc8_2360);
and ( n15496 , RI19ac5720_2288 , n27683 );
or ( n45969 , n15495 , n15496 );
not ( n15497 , RI1754c610_2);
and ( n15498 , n15497 , n45969 );
and ( n15499 , C0 , RI1754c610_2);
or ( n45970 , n15498 , n15499 );
buf ( n45971 , n45970 );
not ( n45972 , n42362 );
and ( n45973 , n45972 , n44592 );
xor ( n45974 , n42359 , n45973 );
not ( n15500 , n29614 );
and ( n15501 , n15500 , RI174541c8_1326);
and ( n15502 , n45974 , n29614 );
or ( n45975 , n15501 , n15502 );
not ( n15503 , RI1754c610_2);
and ( n15504 , n15503 , n45975 );
and ( n15505 , C0 , RI1754c610_2);
or ( n45976 , n15504 , n15505 );
buf ( n45977 , n45976 );
buf ( n45978 , RI17462778_1256);
buf ( n45979 , RI174641b8_1248);
not ( n45980 , n38890 );
xor ( n45981 , n40792 , n40437 );
xor ( n45982 , n45981 , n42635 );
and ( n45983 , n45980 , n45982 );
xor ( n45984 , n38887 , n45983 );
not ( n15506 , n29614 );
and ( n15507 , n15506 , RI173fa2b8_1536);
and ( n15508 , n45984 , n29614 );
or ( n45985 , n15507 , n15508 );
not ( n15509 , RI1754c610_2);
and ( n15510 , n15509 , n45985 );
and ( n15511 , C0 , RI1754c610_2);
or ( n45986 , n15510 , n15511 );
buf ( n45987 , n45986 );
not ( n45988 , n43727 );
and ( n45989 , n45988 , n45779 );
xor ( n45990 , n43724 , n45989 );
not ( n15512 , n29614 );
and ( n15513 , n15512 , RI174c8be0_786);
and ( n15514 , n45990 , n29614 );
or ( n45991 , n15513 , n15514 );
not ( n15515 , RI1754c610_2);
and ( n15516 , n15515 , n45991 );
and ( n15517 , C0 , RI1754c610_2);
or ( n45992 , n15516 , n15517 );
buf ( n45993 , n45992 );
xor ( n45994 , n41378 , n33567 );
xor ( n45995 , n45994 , n33617 );
xor ( n45996 , n30335 , n35311 );
xor ( n45997 , n45996 , n35361 );
not ( n45998 , n45997 );
xor ( n45999 , n31264 , n42049 );
xor ( n46000 , n45999 , n37849 );
and ( n46001 , n45998 , n46000 );
xor ( n46002 , n45995 , n46001 );
not ( n15518 , n29614 );
and ( n15519 , n15518 , RI174153d8_1404);
and ( n15520 , n46002 , n29614 );
or ( n46003 , n15519 , n15520 );
not ( n15521 , RI1754c610_2);
and ( n15522 , n15521 , n46003 );
and ( n15523 , C0 , RI1754c610_2);
or ( n46004 , n15522 , n15523 );
buf ( n46005 , n46004 );
buf ( n46006 , RI174b72a0_843);
xor ( n46007 , n41589 , n39065 );
xor ( n46008 , n46007 , n37331 );
xor ( n46009 , n28606 , n34497 );
xor ( n46010 , n46009 , n34517 );
not ( n46011 , n46010 );
and ( n46012 , n46011 , n42409 );
xor ( n46013 , n46008 , n46012 );
not ( n15524 , n29614 );
and ( n15525 , n15524 , RI174a9a10_909);
and ( n15526 , n46013 , n29614 );
or ( n46014 , n15525 , n15526 );
not ( n15527 , RI1754c610_2);
and ( n15528 , n15527 , n46014 );
and ( n15529 , C0 , RI1754c610_2);
or ( n46015 , n15528 , n15529 );
buf ( n46016 , n46015 );
buf ( n46017 , RI1749baf0_977);
not ( n46018 , n37210 );
xor ( n46019 , n34070 , n39525 );
xor ( n46020 , n46019 , n42377 );
and ( n46021 , n46018 , n46020 );
xor ( n46022 , n37204 , n46021 );
not ( n15530 , n29614 );
and ( n15531 , n15530 , RI173c9f88_1771);
and ( n15532 , n46022 , n29614 );
or ( n46023 , n15531 , n15532 );
not ( n15533 , RI1754c610_2);
and ( n15534 , n15533 , n46023 );
and ( n15535 , C0 , RI1754c610_2);
or ( n46024 , n15534 , n15535 );
buf ( n46025 , n46024 );
not ( n46026 , n44085 );
and ( n46027 , n46026 , n44087 );
xor ( n46028 , n43499 , n46027 );
not ( n15536 , n29614 );
and ( n15537 , n15536 , RI1749e598_964);
and ( n15538 , n46028 , n29614 );
or ( n46029 , n15537 , n15538 );
not ( n15539 , RI1754c610_2);
and ( n15540 , n15539 , n46029 );
and ( n15541 , C0 , RI1754c610_2);
or ( n46030 , n15540 , n15541 );
buf ( n46031 , n46030 );
not ( n15542 , RI1754c610_2);
and ( n15543 , n15542 , RI175379b8_594);
and ( n15544 , C0 , RI1754c610_2);
or ( n46032 , n15543 , n15544 );
buf ( n46033 , n46032 );
xor ( n46034 , n41116 , n41241 );
xor ( n46035 , n46034 , n41287 );
xor ( n46036 , n34030 , n34251 );
xor ( n46037 , n46036 , n42033 );
not ( n46038 , n46037 );
xor ( n46039 , n34149 , n33069 );
xor ( n46040 , n46039 , n42264 );
and ( n46041 , n46038 , n46040 );
xor ( n46042 , n46035 , n46041 );
not ( n15545 , n29614 );
and ( n15546 , n15545 , RI17513f40_704);
and ( n15547 , n46042 , n29614 );
or ( n46043 , n15546 , n15547 );
not ( n15548 , RI1754c610_2);
and ( n15549 , n15548 , n46043 );
and ( n15550 , C0 , RI1754c610_2);
or ( n46044 , n15549 , n15550 );
buf ( n46045 , n46044 );
not ( n46046 , n43062 );
and ( n46047 , n46046 , n45438 );
xor ( n46048 , n43059 , n46047 );
not ( n15551 , n29614 );
and ( n15552 , n15551 , RI1749c810_973);
and ( n15553 , n46048 , n29614 );
or ( n46049 , n15552 , n15553 );
not ( n15554 , RI1754c610_2);
and ( n15555 , n15554 , n46049 );
and ( n15556 , C0 , RI1754c610_2);
or ( n46050 , n15555 , n15556 );
buf ( n46051 , n46050 );
not ( n46052 , n43860 );
and ( n46053 , n46052 , n41443 );
xor ( n46054 , n43857 , n46053 );
not ( n15557 , n29614 );
and ( n15558 , n15557 , RI1739f508_1979);
and ( n15559 , n46054 , n29614 );
or ( n46055 , n15558 , n15559 );
not ( n15560 , RI1754c610_2);
and ( n15561 , n15560 , n46055 );
and ( n15562 , C0 , RI1754c610_2);
or ( n46056 , n15561 , n15562 );
buf ( n46057 , n46056 );
xor ( n46058 , n29896 , n36128 );
xor ( n46059 , n46058 , n36148 );
xor ( n46060 , n38812 , n39621 );
xor ( n46061 , n46060 , n40855 );
not ( n46062 , n46061 );
and ( n46063 , n46062 , n45039 );
xor ( n46064 , n46059 , n46063 );
not ( n15563 , n29614 );
and ( n15564 , n15563 , RI174872d0_1077);
and ( n15565 , n46064 , n29614 );
or ( n46065 , n15564 , n15565 );
not ( n15566 , RI1754c610_2);
and ( n15567 , n15566 , n46065 );
and ( n15568 , C0 , RI1754c610_2);
or ( n46066 , n15567 , n15568 );
buf ( n46067 , n46066 );
xor ( n46068 , n41182 , n34622 );
xor ( n46069 , n46068 , n39397 );
xor ( n46070 , n41875 , n38085 );
xor ( n46071 , n46070 , n38115 );
not ( n46072 , n46071 );
and ( n46073 , n46072 , n43650 );
xor ( n46074 , n46069 , n46073 );
not ( n15569 , n29614 );
and ( n15570 , n15569 , RI174ae240_887);
and ( n15571 , n46074 , n29614 );
or ( n46075 , n15570 , n15571 );
not ( n15572 , RI1754c610_2);
and ( n15573 , n15572 , n46075 );
and ( n15574 , C0 , RI1754c610_2);
or ( n46076 , n15573 , n15574 );
buf ( n46077 , n46076 );
not ( n15575 , n27683 );
and ( n15576 , n15575 , RI19ab2f58_2432);
and ( n15577 , RI19abcbe8_2361 , n27683 );
or ( n46078 , n15576 , n15577 );
not ( n15578 , RI1754c610_2);
and ( n15579 , n15578 , n46078 );
and ( n15580 , C0 , RI1754c610_2);
or ( n46079 , n15579 , n15580 );
buf ( n46080 , n46079 );
xor ( n46081 , n36400 , n34190 );
xor ( n46082 , n46081 , n36252 );
not ( n46083 , n46082 );
and ( n46084 , n46083 , n44126 );
xor ( n46085 , n43638 , n46084 );
not ( n15581 , n29614 );
and ( n15582 , n15581 , RI173af840_1900);
and ( n15583 , n46085 , n29614 );
or ( n46086 , n15582 , n15583 );
not ( n15584 , RI1754c610_2);
and ( n15585 , n15584 , n46086 );
and ( n15586 , C0 , RI1754c610_2);
or ( n46087 , n15585 , n15586 );
buf ( n46088 , n46087 );
not ( n15587 , n27683 );
and ( n15588 , n15587 , RI19ac5e28_2285);
and ( n15589 , RI19aceac8_2220 , n27683 );
or ( n46089 , n15588 , n15589 );
not ( n15590 , RI1754c610_2);
and ( n15591 , n15590 , n46089 );
and ( n15592 , C0 , RI1754c610_2);
or ( n46090 , n15591 , n15592 );
buf ( n46091 , n46090 );
xor ( n46092 , n36835 , n44146 );
xor ( n46093 , n46092 , n41198 );
not ( n46094 , n42505 );
and ( n46095 , n46094 , n42507 );
xor ( n46096 , n46093 , n46095 );
not ( n15593 , n29614 );
and ( n15594 , n15593 , RI173f7810_1549);
and ( n15595 , n46096 , n29614 );
or ( n46097 , n15594 , n15595 );
not ( n15596 , RI1754c610_2);
and ( n15597 , n15596 , n46097 );
and ( n15598 , C0 , RI1754c610_2);
or ( n46098 , n15597 , n15598 );
buf ( n46099 , n46098 );
xor ( n46100 , n39840 , n36742 );
xor ( n46101 , n46100 , n42504 );
not ( n46102 , n46101 );
xor ( n46103 , n39533 , n35842 );
xor ( n46104 , n46103 , n38401 );
and ( n46105 , n46102 , n46104 );
xor ( n46106 , n43962 , n46105 );
not ( n15599 , n29614 );
and ( n15600 , n15599 , RI1733a450_2157);
and ( n15601 , n46106 , n29614 );
or ( n46107 , n15600 , n15601 );
not ( n15602 , RI1754c610_2);
and ( n15603 , n15602 , n46107 );
and ( n15604 , C0 , RI1754c610_2);
or ( n46108 , n15603 , n15604 );
buf ( n46109 , n46108 );
xor ( n46110 , n34208 , n36287 );
xor ( n46111 , n46110 , n37526 );
xor ( n46112 , n39086 , n36377 );
xor ( n46113 , n46112 , n39131 );
not ( n46114 , n46113 );
xor ( n46115 , n37578 , n34968 );
xor ( n46116 , n46115 , n39771 );
and ( n46117 , n46114 , n46116 );
xor ( n46118 , n46111 , n46117 );
not ( n15605 , n29614 );
and ( n15606 , n15605 , RI1739b368_1999);
and ( n15607 , n46118 , n29614 );
or ( n46119 , n15606 , n15607 );
not ( n15608 , RI1754c610_2);
and ( n15609 , n15608 , n46119 );
and ( n15610 , C0 , RI1754c610_2);
or ( n46120 , n15609 , n15610 );
buf ( n46121 , n46120 );
not ( n46122 , n45157 );
and ( n46123 , n46122 , n41700 );
xor ( n46124 , n45154 , n46123 );
not ( n15611 , n29614 );
and ( n15612 , n15611 , RI173a9918_1929);
and ( n15613 , n46124 , n29614 );
or ( n46125 , n15612 , n15613 );
not ( n15614 , RI1754c610_2);
and ( n15615 , n15614 , n46125 );
and ( n15616 , C0 , RI1754c610_2);
or ( n46126 , n15615 , n15616 );
buf ( n46127 , n46126 );
not ( n15617 , n27683 );
and ( n15618 , n15617 , RI19aab410_2487);
and ( n15619 , RI19ab5118_2416 , n27683 );
or ( n46128 , n15618 , n15619 );
not ( n15620 , RI1754c610_2);
and ( n15621 , n15620 , n46128 );
and ( n15622 , C0 , RI1754c610_2);
or ( n46129 , n15621 , n15622 );
buf ( n46130 , n46129 );
not ( n15623 , n27683 );
and ( n15624 , n15623 , RI19acadd8_2249);
and ( n15625 , RI19a86318_2751 , n27683 );
or ( n46131 , n15624 , n15625 );
not ( n15626 , RI1754c610_2);
and ( n15627 , n15626 , n46131 );
and ( n15628 , C0 , RI1754c610_2);
or ( n46132 , n15627 , n15628 );
buf ( n46133 , n46132 );
xor ( n46134 , n32885 , n38553 );
xor ( n46135 , n46134 , n41659 );
xor ( n46136 , n31548 , n39935 );
xor ( n46137 , n46136 , n39952 );
not ( n46138 , n46137 );
xor ( n46139 , n31700 , n30741 );
xor ( n46140 , n46139 , n40769 );
and ( n46141 , n46138 , n46140 );
xor ( n46142 , n46135 , n46141 );
not ( n15629 , n29614 );
and ( n15630 , n15629 , RI174b3100_863);
and ( n15631 , n46142 , n29614 );
or ( n46143 , n15630 , n15631 );
not ( n15632 , RI1754c610_2);
and ( n15633 , n15632 , n46143 );
and ( n15634 , C0 , RI1754c610_2);
or ( n46144 , n15633 , n15634 );
buf ( n46145 , n46144 );
buf ( n46146 , RI174965a0_1003);
buf ( n46147 , RI1746b490_1213);
buf ( n46148 , RI174bf658_815);
not ( n15635 , n27683 );
and ( n15636 , n15635 , RI19aa53f8_2528);
and ( n15637 , RI19aaf790_2457 , n27683 );
or ( n46149 , n15636 , n15637 );
not ( n15638 , RI1754c610_2);
and ( n15639 , n15638 , n46149 );
and ( n15640 , C0 , RI1754c610_2);
or ( n46150 , n15639 , n15640 );
buf ( n46151 , n46150 );
xor ( n46152 , n34020 , n34251 );
xor ( n46153 , n46152 , n42033 );
xor ( n46154 , n41617 , n43278 );
xor ( n46155 , n46154 , n31664 );
not ( n46156 , n46155 );
and ( n46157 , n46156 , n45514 );
xor ( n46158 , n46153 , n46157 );
not ( n15641 , n29614 );
and ( n15642 , n15641 , RI173e7eb0_1625);
and ( n15643 , n46158 , n29614 );
or ( n46159 , n15642 , n15643 );
not ( n15644 , RI1754c610_2);
and ( n15645 , n15644 , n46159 );
and ( n15646 , C0 , RI1754c610_2);
or ( n46160 , n15645 , n15646 );
buf ( n46161 , n46160 );
not ( n15647 , n27683 );
and ( n15648 , n15647 , RI19a9dbf8_2586);
and ( n15649 , RI19aa71f8_2515 , n27683 );
or ( n46162 , n15648 , n15649 );
not ( n15650 , RI1754c610_2);
and ( n15651 , n15650 , n46162 );
and ( n15652 , C0 , RI1754c610_2);
or ( n46163 , n15651 , n15652 );
buf ( n46164 , n46163 );
buf ( n46165 , RI17498670_993);
buf ( n46166 , RI17482de8_1098);
buf ( n46167 , RI1747a418_1140);
buf ( n46168 , RI17469708_1222);
buf ( n46169 , RI1750e270_722);
xor ( n46170 , n40368 , n42554 );
xor ( n46171 , n46170 , n34725 );
not ( n46172 , n46171 );
xor ( n46173 , n39731 , n39506 );
xor ( n46174 , n46173 , n38150 );
and ( n46175 , n46172 , n46174 );
xor ( n46176 , n45372 , n46175 );
not ( n15653 , n29614 );
and ( n15654 , n15653 , RI1733ec80_2135);
and ( n15655 , n46176 , n29614 );
or ( n46177 , n15654 , n15655 );
not ( n15656 , RI1754c610_2);
and ( n15657 , n15656 , n46177 );
and ( n15658 , C0 , RI1754c610_2);
or ( n46178 , n15657 , n15658 );
buf ( n46179 , n46178 );
xor ( n46180 , n37190 , n33030 );
xor ( n46181 , n46180 , n33069 );
xor ( n46182 , n33538 , n40915 );
xor ( n46183 , n46182 , n41740 );
not ( n46184 , n46183 );
xor ( n46185 , n33154 , n37235 );
xor ( n46186 , n46185 , n37255 );
and ( n46187 , n46184 , n46186 );
xor ( n46188 , n46181 , n46187 );
not ( n15659 , n29614 );
and ( n15660 , n15659 , RI1746cb88_1206);
and ( n15661 , n46188 , n29614 );
or ( n46189 , n15660 , n15661 );
not ( n15662 , RI1754c610_2);
and ( n15663 , n15662 , n46189 );
and ( n15664 , C0 , RI1754c610_2);
or ( n46190 , n15663 , n15664 );
buf ( n46191 , n46190 );
buf ( n46192 , RI174bbda0_826);
buf ( n46193 , RI174b1d50_869);
buf ( n46194 , RI174a1388_950);
buf ( n46195 , RI17479068_1146);
xor ( n46196 , n40576 , n37048 );
xor ( n46197 , n46196 , n36772 );
xor ( n46198 , n35453 , n32715 );
xor ( n46199 , n46198 , n36654 );
not ( n46200 , n46199 );
xor ( n46201 , n39150 , n28468 );
xor ( n46202 , n46201 , n36530 );
and ( n46203 , n46200 , n46202 );
xor ( n46204 , n46197 , n46203 );
not ( n15665 , n29614 );
and ( n15666 , n15665 , RI175085a0_740);
and ( n15667 , n46204 , n29614 );
or ( n46205 , n15666 , n15667 );
not ( n15668 , RI1754c610_2);
and ( n15669 , n15668 , n46205 );
and ( n15670 , C0 , RI1754c610_2);
or ( n46206 , n15669 , n15670 );
buf ( n46207 , n46206 );
not ( n15671 , n27683 );
and ( n15672 , n15671 , RI19aafcb8_2455);
and ( n15673 , RI19ab98d0_2384 , n27683 );
or ( n46208 , n15672 , n15673 );
not ( n15674 , RI1754c610_2);
and ( n15675 , n15674 , n46208 );
and ( n15676 , C0 , RI1754c610_2);
or ( n46209 , n15675 , n15676 );
buf ( n46210 , n46209 );
xor ( n46211 , n34473 , n33453 );
xor ( n46212 , n46211 , n33505 );
not ( n46213 , n41216 );
and ( n46214 , n46213 , n38962 );
xor ( n46215 , n46212 , n46214 );
not ( n15677 , n29614 );
and ( n15678 , n15677 , RI174944d0_1013);
and ( n15679 , n46215 , n29614 );
or ( n46216 , n15678 , n15679 );
not ( n15680 , RI1754c610_2);
and ( n15681 , n15680 , n46216 );
and ( n15682 , C0 , RI1754c610_2);
or ( n46217 , n15681 , n15682 );
buf ( n46218 , n46217 );
xor ( n46219 , n39898 , n33397 );
xor ( n46220 , n46219 , n35710 );
not ( n46221 , n43312 );
and ( n46222 , n46221 , n43314 );
xor ( n46223 , n46220 , n46222 );
not ( n15683 , n29614 );
and ( n15684 , n15683 , RI173d0888_1739);
and ( n15685 , n46223 , n29614 );
or ( n46224 , n15684 , n15685 );
not ( n15686 , RI1754c610_2);
and ( n15687 , n15686 , n46224 );
and ( n15688 , C0 , RI1754c610_2);
or ( n46225 , n15687 , n15688 );
buf ( n46226 , n46225 );
buf ( n46227 , RI174b7930_841);
buf ( n46228 , RI1749b7a8_978);
and ( n46229 , RI19a22f70_2797 , RI19a23e70_2789);
not ( n15689 , n46229 );
and ( n15690 , n15689 , RI19ad04a8_2209);
and ( n15691 , C1 , n46229 );
or ( n46230 , n15690 , n15691 );
not ( n46231 , RI1754c610_2);
and ( n46232 , n46230 , n46231 );
buf ( n46233 , n46232 );
xor ( n46234 , n40248 , n35760 );
xor ( n46235 , n46234 , n39333 );
not ( n46236 , n46235 );
and ( n46237 , n46236 , n44739 );
xor ( n46238 , n35274 , n46237 );
not ( n15692 , n29614 );
and ( n15693 , n15692 , RI17396e80_2020);
and ( n15694 , n46238 , n29614 );
or ( n46239 , n15693 , n15694 );
not ( n15695 , RI1754c610_2);
and ( n15696 , n15695 , n46239 );
and ( n15697 , C0 , RI1754c610_2);
or ( n46240 , n15696 , n15697 );
buf ( n46241 , n46240 );
not ( n15698 , n27683 );
and ( n15699 , n15698 , RI19a9c5f0_2595);
and ( n15700 , RI19aa5fb0_2523 , n27683 );
or ( n46242 , n15699 , n15700 );
not ( n15701 , RI1754c610_2);
and ( n15702 , n15701 , n46242 );
and ( n15703 , C0 , RI1754c610_2);
or ( n46243 , n15702 , n15703 );
buf ( n46244 , n46243 );
xor ( n46245 , n41921 , n42033 );
xor ( n46246 , n46245 , n37987 );
not ( n46247 , n44459 );
and ( n46248 , n46247 , n44461 );
xor ( n46249 , n46246 , n46248 );
not ( n15704 , n29614 );
and ( n15705 , n15704 , RI174558c0_1319);
and ( n15706 , n46249 , n29614 );
or ( n46250 , n15705 , n15706 );
not ( n15707 , RI1754c610_2);
and ( n15708 , n15707 , n46250 );
and ( n15709 , C0 , RI1754c610_2);
or ( n46251 , n15708 , n15709 );
buf ( n46252 , n46251 );
xor ( n46253 , n42047 , n33648 );
xor ( n46254 , n46253 , n33697 );
not ( n46255 , n46254 );
xor ( n46256 , n40462 , n35911 );
xor ( n46257 , n46256 , n38188 );
and ( n46258 , n46255 , n46257 );
xor ( n46259 , n46186 , n46258 );
not ( n15710 , n29614 );
and ( n15711 , n15710 , RI17489a30_1065);
and ( n15712 , n46259 , n29614 );
or ( n46260 , n15711 , n15712 );
not ( n15713 , RI1754c610_2);
and ( n15714 , n15713 , n46260 );
and ( n15715 , C0 , RI1754c610_2);
or ( n46261 , n15714 , n15715 );
buf ( n46262 , n46261 );
not ( n15716 , n27683 );
and ( n15717 , n15716 , RI19aa6d48_2517);
and ( n15718 , RI19ab0ff0_2446 , n27683 );
or ( n46263 , n15717 , n15718 );
not ( n15719 , RI1754c610_2);
and ( n15720 , n15719 , n46263 );
and ( n15721 , C0 , RI1754c610_2);
or ( n46264 , n15720 , n15721 );
buf ( n46265 , n46264 );
xor ( n46266 , n36855 , n41198 );
xor ( n46267 , n46266 , n41215 );
xor ( n46268 , n39458 , n36611 );
xor ( n46269 , n46268 , n33567 );
not ( n46270 , n46269 );
and ( n46271 , n46270 , n41971 );
xor ( n46272 , n46267 , n46271 );
not ( n15722 , n29614 );
and ( n15723 , n15722 , RI174c24c0_806);
and ( n15724 , n46272 , n29614 );
or ( n46273 , n15723 , n15724 );
not ( n15725 , RI1754c610_2);
and ( n15726 , n15725 , n46273 );
and ( n15727 , C0 , RI1754c610_2);
or ( n46274 , n15726 , n15727 );
buf ( n46275 , n46274 );
xor ( n46276 , n33727 , n35514 );
xor ( n46277 , n46276 , n40486 );
not ( n46278 , n46277 );
and ( n46279 , n46278 , n46220 );
xor ( n46280 , n43317 , n46279 );
not ( n15728 , n29614 );
and ( n15729 , n15728 , RI173fc388_1526);
and ( n15730 , n46280 , n29614 );
or ( n46281 , n15729 , n15730 );
not ( n15731 , RI1754c610_2);
and ( n15732 , n15731 , n46281 );
and ( n15733 , C0 , RI1754c610_2);
or ( n46282 , n15732 , n15733 );
buf ( n46283 , n46282 );
not ( n15734 , n27683 );
and ( n15735 , n15734 , RI19a98ae0_2621);
and ( n15736 , RI19aa2248_2551 , n27683 );
or ( n46284 , n15735 , n15736 );
not ( n15737 , RI1754c610_2);
and ( n15738 , n15737 , n46284 );
and ( n15739 , C0 , RI1754c610_2);
or ( n46285 , n15738 , n15739 );
buf ( n46286 , n46285 );
not ( n46287 , n41245 );
xor ( n46288 , n34368 , n39989 );
xor ( n46289 , n46288 , n40009 );
and ( n46290 , n46287 , n46289 );
xor ( n46291 , n41242 , n46290 );
not ( n15740 , n29614 );
and ( n15741 , n15740 , RI173ff4c0_1511);
and ( n15742 , n46291 , n29614 );
or ( n46292 , n15741 , n15742 );
not ( n15743 , RI1754c610_2);
and ( n15744 , n15743 , n46292 );
and ( n15745 , C0 , RI1754c610_2);
or ( n46293 , n15744 , n15745 );
buf ( n46294 , n46293 );
not ( n46295 , n42915 );
and ( n46296 , n46295 , n44547 );
xor ( n46297 , n42912 , n46296 );
not ( n15746 , n29614 );
and ( n15747 , n15746 , RI173a8bf8_1933);
and ( n15748 , n46297 , n29614 );
or ( n46298 , n15747 , n15748 );
not ( n15749 , RI1754c610_2);
and ( n15750 , n15749 , n46298 );
and ( n15751 , C0 , RI1754c610_2);
or ( n46299 , n15750 , n15751 );
buf ( n46300 , n46299 );
not ( n15752 , n27683 );
and ( n15753 , n15752 , RI19a922d0_2667);
and ( n15754 , RI19a9c398_2596 , n27683 );
or ( n46301 , n15753 , n15754 );
not ( n15755 , RI1754c610_2);
and ( n15756 , n15755 , n46301 );
and ( n15757 , C0 , RI1754c610_2);
or ( n46302 , n15756 , n15757 );
buf ( n46303 , n46302 );
not ( n46304 , n43175 );
and ( n46305 , n46304 , n43177 );
xor ( n46306 , n43526 , n46305 );
not ( n15758 , n29614 );
and ( n15759 , n15758 , RI174b1378_872);
and ( n15760 , n46306 , n29614 );
or ( n46307 , n15759 , n15760 );
not ( n15761 , RI1754c610_2);
and ( n15762 , n15761 , n46307 );
and ( n15763 , C0 , RI1754c610_2);
or ( n46308 , n15762 , n15763 );
buf ( n46309 , n46308 );
xor ( n46310 , n41794 , n35955 );
xor ( n46311 , n46310 , n42554 );
not ( n46312 , n45070 );
and ( n46313 , n46312 , n45072 );
xor ( n46314 , n46311 , n46313 );
not ( n15764 , n29614 );
and ( n15765 , n15764 , RI17394db0_2030);
and ( n15766 , n46314 , n29614 );
or ( n46315 , n15765 , n15766 );
not ( n15767 , RI1754c610_2);
and ( n15768 , n15767 , n46315 );
and ( n15769 , C0 , RI1754c610_2);
or ( n46316 , n15768 , n15769 );
buf ( n46317 , n46316 );
not ( n46318 , n45733 );
xor ( n46319 , n39390 , n35594 );
xor ( n46320 , n46319 , n32403 );
and ( n46321 , n46318 , n46320 );
xor ( n46322 , n45730 , n46321 );
not ( n15770 , n29614 );
and ( n15771 , n15770 , RI17393a00_2036);
and ( n15772 , n46322 , n29614 );
or ( n46323 , n15771 , n15772 );
not ( n15773 , RI1754c610_2);
and ( n15774 , n15773 , n46323 );
and ( n15775 , C0 , RI1754c610_2);
or ( n46324 , n15774 , n15775 );
buf ( n46325 , n46324 );
not ( n46326 , n40747 );
and ( n46327 , n46326 , n44514 );
xor ( n46328 , n40744 , n46327 );
not ( n15776 , n29614 );
and ( n15777 , n15776 , RI17471700_1183);
and ( n15778 , n46328 , n29614 );
or ( n46329 , n15777 , n15778 );
not ( n15779 , RI1754c610_2);
and ( n15780 , n15779 , n46329 );
and ( n15781 , C0 , RI1754c610_2);
or ( n46330 , n15780 , n15781 );
buf ( n46331 , n46330 );
not ( n15782 , n27683 );
and ( n15783 , n15782 , RI19ab2d78_2433);
and ( n15784 , RI19abca80_2362 , n27683 );
or ( n46332 , n15783 , n15784 );
not ( n15785 , RI1754c610_2);
and ( n15786 , n15785 , n46332 );
and ( n15787 , C0 , RI1754c610_2);
or ( n46333 , n15786 , n15787 );
buf ( n46334 , n46333 );
not ( n46335 , n43662 );
and ( n46336 , n46335 , n43664 );
xor ( n46337 , n44326 , n46336 );
not ( n15788 , n29614 );
and ( n15789 , n15788 , RI17389c80_2084);
and ( n15790 , n46337 , n29614 );
or ( n46338 , n15789 , n15790 );
not ( n15791 , RI1754c610_2);
and ( n15792 , n15791 , n46338 );
and ( n15793 , C0 , RI1754c610_2);
or ( n46339 , n15792 , n15793 );
buf ( n46340 , n46339 );
not ( n46341 , n34252 );
xor ( n46342 , n41429 , n43464 );
xor ( n46343 , n46342 , n44146 );
and ( n46344 , n46341 , n46343 );
xor ( n46345 , n34191 , n46344 );
not ( n15794 , n29614 );
and ( n15795 , n15794 , RI1739f1c0_1980);
and ( n15796 , n46345 , n29614 );
or ( n46346 , n15795 , n15796 );
not ( n15797 , RI1754c610_2);
and ( n15798 , n15797 , n46346 );
and ( n15799 , C0 , RI1754c610_2);
or ( n46347 , n15798 , n15799 );
buf ( n46348 , n46347 );
xor ( n46349 , n28998 , n34517 );
xor ( n46350 , n46349 , n35911 );
not ( n46351 , n44857 );
and ( n46352 , n46351 , n42992 );
xor ( n46353 , n46350 , n46352 );
not ( n15800 , n29614 );
and ( n15801 , n15800 , RI17482de8_1098);
and ( n15802 , n46353 , n29614 );
or ( n46354 , n15801 , n15802 );
not ( n15803 , RI1754c610_2);
and ( n15804 , n15803 , n46354 );
and ( n15805 , C0 , RI1754c610_2);
or ( n46355 , n15804 , n15805 );
buf ( n46356 , n46355 );
not ( n15806 , n27683 );
and ( n15807 , n15806 , RI19ac6ff8_2277);
and ( n15808 , RI19acfb30_2213 , n27683 );
or ( n46357 , n15807 , n15808 );
not ( n15809 , RI1754c610_2);
and ( n15810 , n15809 , n46357 );
and ( n15811 , C0 , RI1754c610_2);
or ( n46358 , n15810 , n15811 );
buf ( n46359 , n46358 );
not ( n15812 , n27683 );
and ( n15813 , n15812 , RI19ac7b38_2272);
and ( n15814 , RI19a82970_2776 , n27683 );
or ( n46360 , n15813 , n15814 );
not ( n15815 , RI1754c610_2);
and ( n15816 , n15815 , n46360 );
and ( n15817 , C0 , RI1754c610_2);
or ( n46361 , n15816 , n15817 );
buf ( n46362 , n46361 );
not ( n46363 , n44714 );
xor ( n46364 , n42183 , n41215 );
xor ( n46365 , n46364 , n33824 );
and ( n46366 , n46363 , n46365 );
xor ( n46367 , n43426 , n46366 );
not ( n15818 , n29614 );
and ( n15819 , n15818 , RI174b9460_834);
and ( n15820 , n46367 , n29614 );
or ( n46368 , n15819 , n15820 );
not ( n15821 , RI1754c610_2);
and ( n15822 , n15821 , n46368 );
and ( n15823 , C0 , RI1754c610_2);
or ( n46369 , n15822 , n15823 );
buf ( n46370 , n46369 );
xor ( n46371 , n40477 , n38933 );
xor ( n46372 , n46371 , n41430 );
not ( n46373 , n45279 );
and ( n46374 , n46373 , n45281 );
xor ( n46375 , n46372 , n46374 );
not ( n15824 , n29614 );
and ( n15825 , n15824 , RI1745ae10_1293);
and ( n15826 , n46375 , n29614 );
or ( n46376 , n15825 , n15826 );
not ( n15827 , RI1754c610_2);
and ( n15828 , n15827 , n46376 );
and ( n15829 , C0 , RI1754c610_2);
or ( n46377 , n15828 , n15829 );
buf ( n46378 , n46377 );
not ( n15830 , n27683 );
and ( n15831 , n15830 , RI19a860c0_2752);
and ( n15832 , RI19a23a38_2791 , n27683 );
or ( n46379 , n15831 , n15832 );
not ( n15833 , RI1754c610_2);
and ( n15834 , n15833 , n46379 );
and ( n15835 , C0 , RI1754c610_2);
or ( n46380 , n15834 , n15835 );
buf ( n46381 , n46380 );
xor ( n46382 , n36270 , n37311 );
xor ( n46383 , n46382 , n37942 );
not ( n46384 , n45667 );
and ( n46385 , n46384 , n45669 );
xor ( n46386 , n46383 , n46385 );
not ( n15836 , n29614 );
and ( n15837 , n15836 , RI173912a0_2048);
and ( n15838 , n46386 , n29614 );
or ( n46387 , n15837 , n15838 );
not ( n15839 , RI1754c610_2);
and ( n15840 , n15839 , n46387 );
and ( n15841 , C0 , RI1754c610_2);
or ( n46388 , n15840 , n15841 );
buf ( n46389 , n46388 );
xor ( n46390 , n39409 , n32403 );
xor ( n46391 , n46390 , n32481 );
xor ( n46392 , n36462 , n37104 );
xor ( n46393 , n46392 , n35986 );
not ( n46394 , n46393 );
xor ( n46395 , n33577 , n41740 );
xor ( n46396 , n46395 , n38371 );
and ( n46397 , n46394 , n46396 );
xor ( n46398 , n46391 , n46397 );
not ( n15842 , n29614 );
and ( n15843 , n15842 , RI17518770_690);
and ( n15844 , n46398 , n29614 );
or ( n46399 , n15843 , n15844 );
not ( n15845 , RI1754c610_2);
and ( n15846 , n15845 , n46399 );
and ( n15847 , C0 , RI1754c610_2);
or ( n46400 , n15846 , n15847 );
buf ( n46401 , n46400 );
xor ( n46402 , n40278 , n37623 );
xor ( n46403 , n46402 , n37651 );
not ( n46404 , n46403 );
xor ( n46405 , n37310 , n40190 );
xor ( n46406 , n46405 , n40210 );
and ( n46407 , n46404 , n46406 );
xor ( n46408 , n46000 , n46407 );
not ( n15848 , n29614 );
and ( n15849 , n15848 , RI17463498_1252);
and ( n15850 , n46408 , n29614 );
or ( n46409 , n15849 , n15850 );
not ( n15851 , RI1754c610_2);
and ( n15852 , n15851 , n46409 );
and ( n15853 , C0 , RI1754c610_2);
or ( n46410 , n15852 , n15853 );
buf ( n46411 , n46410 );
buf ( n46412 , RI174744f0_1169);
xor ( n46413 , n39695 , n33337 );
xor ( n46414 , n46413 , n33397 );
not ( n46415 , n44536 );
and ( n46416 , n46415 , n38402 );
xor ( n46417 , n46414 , n46416 );
not ( n15854 , n29614 );
and ( n15855 , n15854 , RI1738c3e0_2072);
and ( n15856 , n46417 , n29614 );
or ( n46418 , n15855 , n15856 );
not ( n15857 , RI1754c610_2);
and ( n15858 , n15857 , n46418 );
and ( n15859 , C0 , RI1754c610_2);
or ( n46419 , n15858 , n15859 );
buf ( n46420 , n46419 );
not ( n15860 , n27683 );
and ( n15861 , n15860 , RI19a93950_2657);
and ( n15862 , RI19a9dbf8_2586 , n27683 );
or ( n46421 , n15861 , n15862 );
not ( n15863 , RI1754c610_2);
and ( n15864 , n15863 , n46421 );
and ( n15865 , C0 , RI1754c610_2);
or ( n46422 , n15864 , n15865 );
buf ( n46423 , n46422 );
buf ( n46424 , RI174b7c78_840);
buf ( n46425 , RI1749b460_979);
xor ( n46426 , n41185 , n34622 );
xor ( n46427 , n46426 , n39397 );
xor ( n46428 , n34782 , n37255 );
xor ( n46429 , n46428 , n41478 );
not ( n46430 , n46429 );
xor ( n46431 , n39520 , n38371 );
xor ( n46432 , n46431 , n36431 );
and ( n46433 , n46430 , n46432 );
xor ( n46434 , n46427 , n46433 );
not ( n15866 , n29614 );
and ( n15867 , n15866 , RI17458020_1307);
and ( n15868 , n46434 , n29614 );
or ( n46435 , n15867 , n15868 );
not ( n15869 , RI1754c610_2);
and ( n15870 , n15869 , n46435 );
and ( n15871 , C0 , RI1754c610_2);
or ( n46436 , n15870 , n15871 );
buf ( n46437 , n46436 );
xor ( n46438 , n42541 , n37421 );
xor ( n46439 , n46438 , n42605 );
not ( n46440 , n46439 );
xor ( n46441 , n39142 , n28468 );
xor ( n46442 , n46441 , n36530 );
and ( n46443 , n46440 , n46442 );
xor ( n46444 , n44437 , n46443 );
not ( n15872 , n29614 );
and ( n15873 , n15872 , RI1746a770_1217);
and ( n15874 , n46444 , n29614 );
or ( n46445 , n15873 , n15874 );
not ( n15875 , RI1754c610_2);
and ( n15876 , n15875 , n46445 );
and ( n15877 , C0 , RI1754c610_2);
or ( n46446 , n15876 , n15877 );
buf ( n46447 , n46446 );
not ( n46448 , n43342 );
xor ( n46449 , n35292 , n41990 );
xor ( n46450 , n46449 , n41005 );
and ( n46451 , n46448 , n46450 );
xor ( n46452 , n43339 , n46451 );
not ( n15878 , n29614 );
and ( n15879 , n15878 , RI173ba628_1847);
and ( n15880 , n46452 , n29614 );
or ( n46453 , n15879 , n15880 );
not ( n15881 , RI1754c610_2);
and ( n15882 , n15881 , n46453 );
and ( n15883 , C0 , RI1754c610_2);
or ( n46454 , n15882 , n15883 );
buf ( n46455 , n46454 );
not ( n15884 , n27683 );
and ( n15885 , n15884 , RI19a9ad18_2606);
and ( n15886 , RI19aa46d8_2534 , n27683 );
or ( n46456 , n15885 , n15886 );
not ( n15887 , RI1754c610_2);
and ( n15888 , n15887 , n46456 );
and ( n15889 , C0 , RI1754c610_2);
or ( n46457 , n15888 , n15889 );
buf ( n46458 , n46457 );
not ( n46459 , n44690 );
xor ( n46460 , n35946 , n36148 );
xor ( n46461 , n46460 , n37421 );
and ( n46462 , n46459 , n46461 );
xor ( n46463 , n44687 , n46462 );
not ( n15890 , n29614 );
and ( n15891 , n15890 , RI1738d448_2067);
and ( n15892 , n46463 , n29614 );
or ( n46464 , n15891 , n15892 );
not ( n15893 , RI1754c610_2);
and ( n15894 , n15893 , n46464 );
and ( n15895 , C0 , RI1754c610_2);
or ( n46465 , n15894 , n15895 );
buf ( n46466 , n46465 );
not ( n46467 , n43539 );
xor ( n46468 , n41278 , n38648 );
xor ( n46469 , n46468 , n40890 );
and ( n46470 , n46467 , n46469 );
xor ( n46471 , n43536 , n46470 );
not ( n15896 , n29614 );
and ( n15897 , n15896 , RI173cfeb0_1742);
and ( n15898 , n46471 , n29614 );
or ( n46472 , n15897 , n15898 );
not ( n15899 , RI1754c610_2);
and ( n15900 , n15899 , n46472 );
and ( n15901 , C0 , RI1754c610_2);
or ( n46473 , n15900 , n15901 );
buf ( n46474 , n46473 );
not ( n15902 , n27683 );
and ( n15903 , n15902 , RI19a89270_2730);
and ( n15904 , RI19a932c0_2660 , n27683 );
or ( n46475 , n15903 , n15904 );
not ( n15905 , RI1754c610_2);
and ( n15906 , n15905 , n46475 );
and ( n15907 , C0 , RI1754c610_2);
or ( n46476 , n15906 , n15907 );
buf ( n46477 , n46476 );
buf ( n46478 , RI17464b90_1245);
xor ( n46479 , n38569 , n28816 );
xor ( n46480 , n46479 , n29109 );
not ( n46481 , n42749 );
and ( n46482 , n46481 , n42751 );
xor ( n46483 , n46480 , n46482 );
not ( n15908 , n29614 );
and ( n15909 , n15908 , RI1751d9f0_674);
and ( n15910 , n46483 , n29614 );
or ( n46484 , n15909 , n15910 );
not ( n15911 , RI1754c610_2);
and ( n15912 , n15911 , n46484 );
and ( n15913 , C0 , RI1754c610_2);
or ( n46485 , n15912 , n15913 );
buf ( n46486 , n46485 );
not ( n15914 , n27683 );
and ( n15915 , n15914 , RI19a8c6f0_2708);
and ( n15916 , RI19a96740_2637 , n27683 );
or ( n46487 , n15915 , n15916 );
not ( n15917 , RI1754c610_2);
and ( n15918 , n15917 , n46487 );
and ( n15919 , C0 , RI1754c610_2);
or ( n46488 , n15918 , n15919 );
buf ( n46489 , n46488 );
not ( n46490 , n40778 );
and ( n46491 , n46490 , n43012 );
xor ( n46492 , n40772 , n46491 );
not ( n15920 , n29614 );
and ( n15921 , n15920 , RI173e3680_1647);
and ( n15922 , n46492 , n29614 );
or ( n46493 , n15921 , n15922 );
not ( n15923 , RI1754c610_2);
and ( n15924 , n15923 , n46493 );
and ( n15925 , C0 , RI1754c610_2);
or ( n46494 , n15924 , n15925 );
buf ( n46495 , n46494 );
xor ( n46496 , n38707 , n38817 );
xor ( n46497 , n46496 , n40034 );
not ( n46498 , n46497 );
xor ( n46499 , n28745 , n34497 );
xor ( n46500 , n46499 , n34517 );
and ( n46501 , n46498 , n46500 );
xor ( n46502 , n45229 , n46501 );
not ( n15926 , n29614 );
and ( n15927 , n15926 , RI17450028_1346);
and ( n15928 , n46502 , n29614 );
or ( n46503 , n15927 , n15928 );
not ( n15929 , RI1754c610_2);
and ( n15930 , n15929 , n46503 );
and ( n15931 , C0 , RI1754c610_2);
or ( n46504 , n15930 , n15931 );
buf ( n46505 , n46504 );
xor ( n46506 , n40503 , n41430 );
xor ( n46507 , n46506 , n36844 );
not ( n46508 , n35640 );
and ( n46509 , n46508 , n34969 );
xor ( n46510 , n46507 , n46509 );
not ( n15932 , n29614 );
and ( n15933 , n15932 , RI173e9f80_1615);
and ( n15934 , n46510 , n29614 );
or ( n46511 , n15933 , n15934 );
not ( n15935 , RI1754c610_2);
and ( n15936 , n15935 , n46511 );
and ( n15937 , C0 , RI1754c610_2);
or ( n46512 , n15936 , n15937 );
buf ( n46513 , n46512 );
not ( n46514 , n44760 );
xor ( n46515 , n38084 , n40091 );
xor ( n46516 , n46515 , n40111 );
and ( n46517 , n46514 , n46516 );
xor ( n46518 , n44757 , n46517 );
not ( n15938 , n29614 );
and ( n15939 , n15938 , RI173eca28_1602);
and ( n15940 , n46518 , n29614 );
or ( n46519 , n15939 , n15940 );
not ( n15941 , RI1754c610_2);
and ( n15942 , n15941 , n46519 );
and ( n15943 , C0 , RI1754c610_2);
or ( n46520 , n15942 , n15943 );
buf ( n46521 , n46520 );
xor ( n46522 , n29796 , n39091 );
xor ( n46523 , n46522 , n36128 );
xor ( n46524 , n38531 , n31725 );
xor ( n46525 , n46524 , n42309 );
not ( n46526 , n46525 );
xor ( n46527 , n40078 , n38037 );
xor ( n46528 , n46527 , n39740 );
and ( n46529 , n46526 , n46528 );
xor ( n46530 , n46523 , n46529 );
not ( n15944 , n29614 );
and ( n15945 , n15944 , RI17390580_2052);
and ( n15946 , n46530 , n29614 );
or ( n46531 , n15945 , n15946 );
not ( n15947 , RI1754c610_2);
and ( n15948 , n15947 , n46531 );
and ( n15949 , C0 , RI1754c610_2);
or ( n46532 , n15948 , n15949 );
buf ( n46533 , n46532 );
not ( n46534 , n42456 );
and ( n46535 , n46534 , n42458 );
xor ( n46536 , n44030 , n46535 );
not ( n15950 , n29614 );
and ( n15951 , n15950 , RI1733cbb0_2145);
and ( n15952 , n46536 , n29614 );
or ( n46537 , n15951 , n15952 );
not ( n15953 , RI1754c610_2);
and ( n15954 , n15953 , n46537 );
and ( n15955 , C0 , RI1754c610_2);
or ( n46538 , n15954 , n15955 );
buf ( n46539 , n46538 );
not ( n46540 , n42903 );
xor ( n46541 , n33124 , n38244 );
xor ( n46542 , n46541 , n37235 );
and ( n46543 , n46540 , n46542 );
xor ( n46544 , n42900 , n46543 );
not ( n15956 , n29614 );
and ( n15957 , n15956 , RI1739b6b0_1998);
and ( n15958 , n46544 , n29614 );
or ( n46545 , n15957 , n15958 );
not ( n15959 , RI1754c610_2);
and ( n15960 , n15959 , n46545 );
and ( n15961 , C0 , RI1754c610_2);
or ( n46546 , n15960 , n15961 );
buf ( n46547 , n46546 );
not ( n46548 , n45324 );
xor ( n46549 , n33529 , n40915 );
xor ( n46550 , n46549 , n41740 );
and ( n46551 , n46548 , n46550 );
xor ( n46552 , n45321 , n46551 );
not ( n15962 , n29614 );
and ( n15963 , n15962 , RI173ae7d8_1905);
and ( n15964 , n46552 , n29614 );
or ( n46553 , n15963 , n15964 );
not ( n15965 , RI1754c610_2);
and ( n15966 , n15965 , n46553 );
and ( n15967 , C0 , RI1754c610_2);
or ( n46554 , n15966 , n15967 );
buf ( n46555 , n46554 );
xor ( n46556 , n39017 , n36947 );
xor ( n46557 , n46556 , n39702 );
not ( n46558 , n46557 );
and ( n46559 , n46558 , n42898 );
xor ( n46560 , n46542 , n46559 );
not ( n15968 , n29614 );
and ( n15969 , n15968 , RI173b8be8_1855);
and ( n15970 , n46560 , n29614 );
or ( n46561 , n15969 , n15970 );
not ( n15971 , RI1754c610_2);
and ( n15972 , n15971 , n46561 );
and ( n15973 , C0 , RI1754c610_2);
or ( n46562 , n15972 , n15973 );
buf ( n46563 , n46562 );
not ( n46564 , n45534 );
xor ( n46565 , n42179 , n41215 );
xor ( n46566 , n46565 , n33824 );
and ( n46567 , n46564 , n46566 );
xor ( n46568 , n45531 , n46567 );
not ( n15974 , n29614 );
and ( n15975 , n15974 , RI173cd408_1755);
and ( n15976 , n46568 , n29614 );
or ( n46569 , n15975 , n15976 );
not ( n15977 , RI1754c610_2);
and ( n15978 , n15977 , n46569 );
and ( n15979 , C0 , RI1754c610_2);
or ( n46570 , n15978 , n15979 );
buf ( n46571 , n46570 );
xor ( n46572 , n42494 , n30461 );
xor ( n46573 , n46572 , n39262 );
xor ( n46574 , n39515 , n38371 );
xor ( n46575 , n46574 , n36431 );
not ( n46576 , n46575 );
xor ( n46577 , n40819 , n42635 );
xor ( n46578 , n46577 , n33648 );
and ( n46579 , n46576 , n46578 );
xor ( n46580 , n46573 , n46579 );
not ( n15980 , n29614 );
and ( n15981 , n15980 , RI173d2cb8_1728);
and ( n15982 , n46580 , n29614 );
or ( n46581 , n15981 , n15982 );
not ( n15983 , RI1754c610_2);
and ( n15984 , n15983 , n46581 );
and ( n15985 , C0 , RI1754c610_2);
or ( n46582 , n15984 , n15985 );
buf ( n46583 , n46582 );
xor ( n46584 , n38723 , n38817 );
xor ( n46585 , n46584 , n40034 );
not ( n46586 , n42189 );
and ( n46587 , n46586 , n42191 );
xor ( n46588 , n46585 , n46587 );
not ( n15986 , n29614 );
and ( n15987 , n15986 , RI174a6248_926);
and ( n15988 , n46588 , n29614 );
or ( n46589 , n15987 , n15988 );
not ( n15989 , RI1754c610_2);
and ( n15990 , n15989 , n46589 );
and ( n15991 , C0 , RI1754c610_2);
or ( n46590 , n15990 , n15991 );
buf ( n46591 , n46590 );
xor ( n46592 , n37429 , n34725 );
xor ( n46593 , n46592 , n34755 );
xor ( n46594 , n39879 , n42504 );
xor ( n46595 , n46594 , n41818 );
not ( n46596 , n46595 );
and ( n46597 , n46596 , n41868 );
xor ( n46598 , n46593 , n46597 );
not ( n15992 , n29614 );
and ( n15993 , n15992 , RI17483130_1097);
and ( n15994 , n46598 , n29614 );
or ( n46599 , n15993 , n15994 );
not ( n15995 , RI1754c610_2);
and ( n15996 , n15995 , n46599 );
and ( n15997 , C0 , RI1754c610_2);
or ( n46600 , n15996 , n15997 );
buf ( n46601 , n46600 );
not ( n15998 , n27683 );
and ( n15999 , n15998 , RI19ab2b98_2434);
and ( n16000 , RI19abc8a0_2363 , n27683 );
or ( n46602 , n15999 , n16000 );
not ( n16001 , RI1754c610_2);
and ( n16002 , n16001 , n46602 );
and ( n16003 , C0 , RI1754c610_2);
or ( n46603 , n16002 , n16003 );
buf ( n46604 , n46603 );
not ( n46605 , n45372 );
and ( n46606 , n46605 , n46171 );
xor ( n46607 , n45369 , n46606 );
not ( n16004 , n29614 );
and ( n16005 , n16004 , RI173b9c50_1850);
and ( n16006 , n46607 , n29614 );
or ( n46608 , n16005 , n16006 );
not ( n16007 , RI1754c610_2);
and ( n16008 , n16007 , n46608 );
and ( n16009 , C0 , RI1754c610_2);
or ( n46609 , n16008 , n16009 );
buf ( n46610 , n46609 );
not ( n16010 , n27683 );
and ( n16011 , n16010 , RI19a905c0_2680);
and ( n16012 , RI19a9a610_2609 , n27683 );
or ( n46611 , n16011 , n16012 );
not ( n16013 , RI1754c610_2);
and ( n16014 , n16013 , n46611 );
and ( n16015 , C0 , RI1754c610_2);
or ( n46612 , n16014 , n16015 );
buf ( n46613 , n46612 );
xor ( n46614 , n37185 , n32481 );
xor ( n46615 , n46614 , n33030 );
not ( n46616 , n36569 );
and ( n46617 , n46616 , n36613 );
xor ( n46618 , n46615 , n46617 );
not ( n16016 , n29614 );
and ( n16017 , n16016 , RI1740c378_1448);
and ( n16018 , n46618 , n29614 );
or ( n46619 , n16017 , n16018 );
not ( n16019 , RI1754c610_2);
and ( n16020 , n16019 , n46619 );
and ( n16021 , C0 , RI1754c610_2);
or ( n46620 , n16020 , n16021 );
buf ( n46621 , n46620 );
not ( n16022 , RI19ad21b8_2198);
and ( n16023 , n16022 , RI19ad0700_2208);
and ( n16024 , C1 , RI19ad21b8_2198);
or ( n46622 , n16023 , n16024 );
not ( n46623 , RI1754c610_2);
and ( n46624 , n46622 , n46623 );
buf ( n46625 , n46624 );
xor ( n46626 , n44145 , n34572 );
xor ( n46627 , n46626 , n34622 );
xor ( n46628 , n30525 , n38167 );
xor ( n46629 , n46628 , n33728 );
not ( n46630 , n46629 );
xor ( n46631 , n34202 , n36287 );
xor ( n46632 , n46631 , n37526 );
and ( n46633 , n46630 , n46632 );
xor ( n46634 , n46627 , n46633 );
not ( n16025 , n29614 );
and ( n16026 , n16025 , RI17457cd8_1308);
and ( n16027 , n46634 , n29614 );
or ( n46635 , n16026 , n16027 );
not ( n16028 , RI1754c610_2);
and ( n16029 , n16028 , n46635 );
and ( n16030 , C0 , RI1754c610_2);
or ( n46636 , n16029 , n16030 );
buf ( n46637 , n46636 );
not ( n46638 , n43165 );
and ( n46639 , n46638 , n45588 );
xor ( n46640 , n43162 , n46639 );
not ( n16031 , n29614 );
and ( n16032 , n16031 , RI173e4a30_1641);
and ( n16033 , n46640 , n29614 );
or ( n46641 , n16032 , n16033 );
not ( n16034 , RI1754c610_2);
and ( n16035 , n16034 , n46641 );
and ( n16036 , C0 , RI1754c610_2);
or ( n46642 , n16035 , n16036 );
buf ( n46643 , n46642 );
xor ( n46644 , n38096 , n40111 );
xor ( n46645 , n46644 , n43278 );
not ( n46646 , n46645 );
xor ( n46647 , n35787 , n37331 );
xor ( n46648 , n46647 , n37129 );
and ( n46649 , n46646 , n46648 );
xor ( n46650 , n42525 , n46649 );
not ( n16037 , n29614 );
and ( n16038 , n16037 , RI173c5aa0_1792);
and ( n16039 , n46650 , n29614 );
or ( n46651 , n16038 , n16039 );
not ( n16040 , RI1754c610_2);
and ( n16041 , n16040 , n46651 );
and ( n16042 , C0 , RI1754c610_2);
or ( n46652 , n16041 , n16042 );
buf ( n46653 , n46652 );
not ( n16043 , n27683 );
and ( n16044 , n16043 , RI19aa6190_2522);
and ( n16045 , RI19ab03c0_2452 , n27683 );
or ( n46654 , n16044 , n16045 );
not ( n16046 , RI1754c610_2);
and ( n16047 , n16046 , n46654 );
and ( n16048 , C0 , RI1754c610_2);
or ( n46655 , n16047 , n16048 );
buf ( n46656 , n46655 );
xor ( n46657 , n35633 , n34669 );
xor ( n46658 , n46657 , n31831 );
xor ( n46659 , n37286 , n34127 );
xor ( n46660 , n46659 , n40190 );
not ( n46661 , n46660 );
xor ( n46662 , n33777 , n40486 );
xor ( n46663 , n46662 , n40516 );
and ( n46664 , n46661 , n46663 );
xor ( n46665 , n46658 , n46664 );
not ( n16049 , n29614 );
and ( n16050 , n16049 , RI1739ee78_1981);
and ( n16051 , n46665 , n29614 );
or ( n46666 , n16050 , n16051 );
not ( n16052 , RI1754c610_2);
and ( n16053 , n16052 , n46666 );
and ( n16054 , C0 , RI1754c610_2);
or ( n46667 , n16053 , n16054 );
buf ( n46668 , n46667 );
xor ( n46669 , n37812 , n31213 );
xor ( n46670 , n46669 , n31317 );
not ( n46671 , n42429 );
and ( n46672 , n46671 , n42431 );
xor ( n46673 , n46670 , n46672 );
not ( n16055 , n29614 );
and ( n16056 , n16055 , RI17498328_994);
and ( n16057 , n46673 , n29614 );
or ( n46674 , n16056 , n16057 );
not ( n16058 , RI1754c610_2);
and ( n16059 , n16058 , n46674 );
and ( n16060 , C0 , RI1754c610_2);
or ( n46675 , n16059 , n16060 );
buf ( n46676 , n46675 );
xor ( n46677 , n40450 , n35911 );
xor ( n46678 , n46677 , n38188 );
not ( n46679 , n45082 );
and ( n46680 , n46679 , n45084 );
xor ( n46681 , n46678 , n46680 );
not ( n16061 , n29614 );
and ( n16062 , n16061 , RI174c86b8_787);
and ( n16063 , n46681 , n29614 );
or ( n46682 , n16062 , n16063 );
not ( n16064 , RI1754c610_2);
and ( n16065 , n16064 , n46682 );
and ( n16066 , C0 , RI1754c610_2);
or ( n46683 , n16065 , n16066 );
buf ( n46684 , n46683 );
not ( n46685 , n36024 );
and ( n46686 , n46685 , n36029 );
xor ( n46687 , n36293 , n46686 );
not ( n16067 , n29614 );
and ( n16068 , n16067 , RI1748a750_1061);
and ( n16069 , n46687 , n29614 );
or ( n46688 , n16068 , n16069 );
not ( n16070 , RI1754c610_2);
and ( n16071 , n16070 , n46688 );
and ( n16072 , C0 , RI1754c610_2);
or ( n46689 , n16071 , n16072 );
buf ( n46690 , n46689 );
not ( n16073 , n27683 );
and ( n16074 , n16073 , RI19aa19d8_2555);
and ( n16075 , RI19aabb90_2484 , n27683 );
or ( n46691 , n16074 , n16075 );
not ( n16076 , RI1754c610_2);
and ( n16077 , n16076 , n46691 );
and ( n16078 , C0 , RI1754c610_2);
or ( n46692 , n16077 , n16078 );
buf ( n46693 , n46692 );
xor ( n46694 , n33108 , n38244 );
xor ( n46695 , n46694 , n37235 );
not ( n46696 , n46695 );
xor ( n46697 , n40823 , n42635 );
xor ( n46698 , n46697 , n33648 );
and ( n46699 , n46696 , n46698 );
xor ( n46700 , n44452 , n46699 );
not ( n16079 , n29614 );
and ( n16080 , n16079 , RI174c1f98_807);
and ( n16081 , n46700 , n29614 );
or ( n46701 , n16080 , n16081 );
not ( n16082 , RI1754c610_2);
and ( n16083 , n16082 , n46701 );
and ( n16084 , C0 , RI1754c610_2);
or ( n46702 , n16083 , n16084 );
buf ( n46703 , n46702 );
xor ( n46704 , n43487 , n32108 );
xor ( n46705 , n46704 , n38347 );
not ( n46706 , n46705 );
xor ( n46707 , n33281 , n40302 );
xor ( n46708 , n46707 , n40319 );
and ( n46709 , n46706 , n46708 );
xor ( n46710 , n39564 , n46709 );
not ( n16085 , n29614 );
and ( n16086 , n16085 , RI17502948_752);
and ( n16087 , n46710 , n29614 );
or ( n46711 , n16086 , n16087 );
not ( n16088 , RI1754c610_2);
and ( n16089 , n16088 , n46711 );
and ( n16090 , C0 , RI1754c610_2);
or ( n46712 , n16089 , n16090 );
buf ( n46713 , n46712 );
not ( n46714 , n45765 );
and ( n46715 , n46714 , n44389 );
xor ( n46716 , n45762 , n46715 );
not ( n16091 , n29614 );
and ( n16092 , n16091 , RI17509f68_735);
and ( n16093 , n46716 , n29614 );
or ( n46717 , n16092 , n16093 );
not ( n16094 , RI1754c610_2);
and ( n16095 , n16094 , n46717 );
and ( n16096 , C0 , RI1754c610_2);
or ( n46718 , n16095 , n16096 );
buf ( n46719 , n46718 );
xor ( n46720 , n41311 , n41526 );
xor ( n46721 , n46720 , n41543 );
xor ( n46722 , n38647 , n34300 );
xor ( n46723 , n46722 , n34340 );
not ( n46724 , n46723 );
xor ( n46725 , n38154 , n35494 );
xor ( n46726 , n46725 , n35514 );
and ( n46727 , n46724 , n46726 );
xor ( n46728 , n46721 , n46727 );
not ( n16097 , n29614 );
and ( n16098 , n16097 , RI173b0f38_1893);
and ( n16099 , n46728 , n29614 );
or ( n46729 , n16098 , n16099 );
not ( n16100 , RI1754c610_2);
and ( n16101 , n16100 , n46729 );
and ( n16102 , C0 , RI1754c610_2);
or ( n46730 , n16101 , n16102 );
buf ( n46731 , n46730 );
xor ( n46732 , n35287 , n41990 );
xor ( n46733 , n46732 , n41005 );
xor ( n46734 , n35389 , n41068 );
xor ( n46735 , n46734 , n39091 );
not ( n46736 , n46735 );
xor ( n46737 , n40454 , n35911 );
xor ( n46738 , n46737 , n38188 );
and ( n46739 , n46736 , n46738 );
xor ( n46740 , n46733 , n46739 );
not ( n16103 , n29614 );
and ( n16104 , n16103 , RI17413998_1412);
and ( n16105 , n46740 , n29614 );
or ( n46741 , n16104 , n16105 );
not ( n16106 , RI1754c610_2);
and ( n16107 , n16106 , n46741 );
and ( n16108 , C0 , RI1754c610_2);
or ( n46742 , n16107 , n16108 );
buf ( n46743 , n46742 );
not ( n46744 , n43556 );
xor ( n46745 , n36916 , n32560 );
xor ( n46746 , n46745 , n32620 );
and ( n46747 , n46744 , n46746 );
xor ( n46748 , n43414 , n46747 );
not ( n16109 , n29614 );
and ( n16110 , n16109 , RI173e6470_1633);
and ( n16111 , n46748 , n29614 );
or ( n46749 , n16110 , n16111 );
not ( n16112 , RI1754c610_2);
and ( n16113 , n16112 , n46749 );
and ( n16114 , C0 , RI1754c610_2);
or ( n46750 , n16113 , n16114 );
buf ( n46751 , n46750 );
buf ( n46752 , RI174920b8_1024);
buf ( n46753 , RI174893a0_1067);
buf ( n46754 , RI17502948_752);
buf ( n46755 , RI1747cb78_1128);
not ( n46756 , n46480 );
and ( n46757 , n46756 , n42749 );
xor ( n46758 , n42866 , n46757 );
not ( n16115 , n29614 );
and ( n16116 , n16115 , RI175066b0_746);
and ( n16117 , n46758 , n29614 );
or ( n46759 , n16116 , n16117 );
not ( n16118 , RI1754c610_2);
and ( n16119 , n16118 , n46759 );
and ( n16120 , C0 , RI1754c610_2);
or ( n46760 , n16119 , n16120 );
buf ( n46761 , n46760 );
buf ( n46762 , RI174637e0_1251);
xor ( n46763 , n33271 , n40302 );
xor ( n46764 , n46763 , n40319 );
not ( n46765 , n46615 );
and ( n46766 , n46765 , n36569 );
xor ( n46767 , n46764 , n46766 );
not ( n16121 , n29614 );
and ( n16122 , n16121 , RI173fddc8_1518);
and ( n16123 , n46767 , n29614 );
or ( n46768 , n16122 , n16123 );
not ( n16124 , RI1754c610_2);
and ( n16125 , n16124 , n46768 );
and ( n16126 , C0 , RI1754c610_2);
or ( n46769 , n16125 , n16126 );
buf ( n46770 , n46769 );
not ( n46771 , n42910 );
and ( n46772 , n46771 , n42912 );
xor ( n46773 , n44550 , n46772 );
not ( n16127 , n29614 );
and ( n16128 , n16127 , RI1738ba08_2075);
and ( n16129 , n46773 , n29614 );
or ( n46774 , n16128 , n16129 );
not ( n16130 , RI1754c610_2);
and ( n16131 , n16130 , n46774 );
and ( n16132 , C0 , RI1754c610_2);
or ( n46775 , n16131 , n16132 );
buf ( n46776 , n46775 );
xor ( n46777 , n39269 , n38445 );
xor ( n46778 , n46777 , n37549 );
xor ( n46779 , n40941 , n38793 );
xor ( n46780 , n46779 , n40563 );
not ( n46781 , n46780 );
xor ( n46782 , n34957 , n36802 );
xor ( n46783 , n46782 , n33125 );
and ( n46784 , n46781 , n46783 );
xor ( n46785 , n46778 , n46784 );
not ( n16133 , n29614 );
and ( n16134 , n16133 , RI1738f1d0_2058);
and ( n16135 , n46785 , n29614 );
or ( n46786 , n16134 , n16135 );
not ( n16136 , RI1754c610_2);
and ( n16137 , n16136 , n46786 );
and ( n16138 , C0 , RI1754c610_2);
or ( n46787 , n16137 , n16138 );
buf ( n46788 , n46787 );
not ( n46789 , n39348 );
xor ( n46790 , n34501 , n31380 );
xor ( n46791 , n46790 , n36463 );
and ( n46792 , n46789 , n46791 );
xor ( n46793 , n39316 , n46792 );
not ( n16139 , n29614 );
and ( n16140 , n16139 , RI173b5df8_1869);
and ( n16141 , n46793 , n29614 );
or ( n46794 , n16140 , n16141 );
not ( n16142 , RI1754c610_2);
and ( n16143 , n16142 , n46794 );
and ( n16144 , C0 , RI1754c610_2);
or ( n46795 , n16143 , n16144 );
buf ( n46796 , n46795 );
buf ( n46797 , RI174cba48_777);
not ( n16145 , n27683 );
and ( n16146 , n16145 , RI19aa9f70_2496);
and ( n16147 , RI19ab3de0_2424 , n27683 );
or ( n46798 , n16146 , n16147 );
not ( n16148 , RI1754c610_2);
and ( n16149 , n16148 , n46798 );
and ( n16150 , C0 , RI1754c610_2);
or ( n46799 , n16149 , n16150 );
buf ( n46800 , n46799 );
xor ( n46801 , n35709 , n39543 );
xor ( n46802 , n46801 , n39563 );
xor ( n46803 , n29238 , n40034 );
xor ( n46804 , n46803 , n40051 );
not ( n46805 , n46804 );
and ( n46806 , n46805 , n44898 );
xor ( n46807 , n46802 , n46806 );
not ( n16151 , n29614 );
and ( n16152 , n16151 , RI173c4060_1800);
and ( n16153 , n46807 , n29614 );
or ( n46808 , n16152 , n16153 );
not ( n16154 , RI1754c610_2);
and ( n16155 , n16154 , n46808 );
and ( n16156 , C0 , RI1754c610_2);
or ( n46809 , n16155 , n16156 );
buf ( n46810 , n46809 );
xor ( n46811 , n39373 , n35594 );
xor ( n46812 , n46811 , n32403 );
xor ( n46813 , n32067 , n36702 );
xor ( n46814 , n46813 , n38872 );
not ( n46815 , n46814 );
xor ( n46816 , n33550 , n40915 );
xor ( n46817 , n46816 , n41740 );
and ( n46818 , n46815 , n46817 );
xor ( n46819 , n46812 , n46818 );
not ( n16157 , n29614 );
and ( n16158 , n16157 , RI173c98f8_1773);
and ( n16159 , n46819 , n29614 );
or ( n46820 , n16158 , n16159 );
not ( n16160 , RI1754c610_2);
and ( n16161 , n16160 , n46820 );
and ( n16162 , C0 , RI1754c610_2);
or ( n46821 , n16161 , n16162 );
buf ( n46822 , n46821 );
buf ( n46823 , RI174b7fc0_839);
buf ( n46824 , RI1749ec28_962);
xor ( n46825 , n33206 , n31317 );
xor ( n46826 , n46825 , n40302 );
xor ( n46827 , n44140 , n34572 );
xor ( n46828 , n46827 , n34622 );
not ( n46829 , n46828 );
xor ( n46830 , n34664 , n32863 );
xor ( n46831 , n46830 , n34644 );
and ( n46832 , n46829 , n46831 );
xor ( n46833 , n46826 , n46832 );
not ( n16163 , n29614 );
and ( n16164 , n16163 , RI173db9d0_1685);
and ( n16165 , n46833 , n29614 );
or ( n46834 , n16164 , n16165 );
not ( n16166 , RI1754c610_2);
and ( n16167 , n16166 , n46834 );
and ( n16168 , C0 , RI1754c610_2);
or ( n46835 , n16167 , n16168 );
buf ( n46836 , n46835 );
xor ( n46837 , n36318 , n40718 );
xor ( n46838 , n46837 , n38676 );
xor ( n46839 , n35739 , n39563 );
xor ( n46840 , n46839 , n35416 );
not ( n46841 , n46840 );
and ( n46842 , n46841 , n44201 );
xor ( n46843 , n46838 , n46842 );
not ( n16169 , n29614 );
and ( n16170 , n16169 , RI17478348_1150);
and ( n16171 , n46843 , n29614 );
or ( n46844 , n16170 , n16171 );
not ( n16172 , RI1754c610_2);
and ( n16173 , n16172 , n46844 );
and ( n16174 , C0 , RI1754c610_2);
or ( n46845 , n16173 , n16174 );
buf ( n46846 , n46845 );
not ( n16175 , n27683 );
and ( n16176 , n16175 , RI19ab29b8_2435);
and ( n16177 , RI19abc6c0_2364 , n27683 );
or ( n46847 , n16176 , n16177 );
not ( n16178 , RI1754c610_2);
and ( n16179 , n16178 , n46847 );
and ( n16180 , C0 , RI1754c610_2);
or ( n46848 , n16179 , n16180 );
buf ( n46849 , n46848 );
xor ( n46850 , n39843 , n36742 );
xor ( n46851 , n46850 , n42504 );
xor ( n46852 , n35035 , n37814 );
xor ( n46853 , n46852 , n33223 );
not ( n46854 , n46853 );
xor ( n46855 , n37847 , n33697 );
xor ( n46856 , n46855 , n35128 );
and ( n46857 , n46854 , n46856 );
xor ( n46858 , n46851 , n46857 );
not ( n16181 , n29614 );
and ( n16182 , n16181 , RI17452440_1335);
and ( n16183 , n46858 , n29614 );
or ( n46859 , n16182 , n16183 );
not ( n16184 , RI1754c610_2);
and ( n16185 , n16184 , n46859 );
and ( n16186 , C0 , RI1754c610_2);
or ( n46860 , n16185 , n16186 );
buf ( n46861 , n46860 );
not ( n16187 , n27683 );
and ( n16188 , n16187 , RI19ab7008_2402);
and ( n16189 , RI19abff78_2332 , n27683 );
or ( n46862 , n16188 , n16189 );
not ( n16190 , RI1754c610_2);
and ( n16191 , n16190 , n46862 );
and ( n16192 , C0 , RI1754c610_2);
or ( n46863 , n16191 , n16192 );
buf ( n46864 , n46863 );
not ( n16193 , n27683 );
and ( n16194 , n16193 , RI19ab0000_2454);
and ( n16195 , RI19ab9a38_2383 , n27683 );
or ( n46865 , n16194 , n16195 );
not ( n16196 , RI1754c610_2);
and ( n16197 , n16196 , n46865 );
and ( n16198 , C0 , RI1754c610_2);
or ( n46866 , n16197 , n16198 );
buf ( n46867 , n46866 );
not ( n46868 , n41666 );
xor ( n46869 , n41202 , n39397 );
xor ( n46870 , n46869 , n39414 );
and ( n46871 , n46868 , n46870 );
xor ( n46872 , n41660 , n46871 );
not ( n16199 , n29614 );
and ( n16200 , n16199 , RI17401c20_1499);
and ( n16201 , n46872 , n29614 );
or ( n46873 , n16200 , n16201 );
not ( n16202 , RI1754c610_2);
and ( n16203 , n16202 , n46873 );
and ( n16204 , C0 , RI1754c610_2);
or ( n46874 , n16203 , n16204 );
buf ( n46875 , n46874 );
xor ( n46876 , n36519 , n40381 );
xor ( n46877 , n46876 , n37438 );
not ( n46878 , n44983 );
and ( n46879 , n46878 , n44985 );
xor ( n46880 , n46877 , n46879 );
not ( n16205 , n29614 );
and ( n16206 , n16205 , RI1748cb68_1050);
and ( n16207 , n46880 , n29614 );
or ( n46881 , n16206 , n16207 );
not ( n16208 , RI1754c610_2);
and ( n16209 , n16208 , n46881 );
and ( n16210 , C0 , RI1754c610_2);
or ( n46882 , n16209 , n16210 );
buf ( n46883 , n46882 );
buf ( n46884 , RI174ad520_891);
buf ( n46885 , RI174a96c8_910);
xor ( n46886 , n42630 , n35052 );
xor ( n46887 , n46886 , n35069 );
xor ( n46888 , n34836 , n41478 );
xor ( n46889 , n46888 , n41146 );
not ( n46890 , n46889 );
xor ( n46891 , n38198 , n37696 );
xor ( n46892 , n46891 , n39450 );
and ( n46893 , n46890 , n46892 );
xor ( n46894 , n46887 , n46893 );
not ( n16211 , n29614 );
and ( n16212 , n16211 , RI17336c88_2174);
and ( n16213 , n46894 , n29614 );
or ( n46895 , n16212 , n16213 );
not ( n16214 , RI1754c610_2);
and ( n16215 , n16214 , n46895 );
and ( n16216 , C0 , RI1754c610_2);
or ( n46896 , n16215 , n16216 );
buf ( n46897 , n46896 );
not ( n16217 , n27683 );
and ( n16218 , n16217 , RI19a82970_2776);
and ( n16219 , RI19aadb70_2470 , n27683 );
or ( n46898 , n16218 , n16219 );
not ( n16220 , RI1754c610_2);
and ( n16221 , n16220 , n46898 );
and ( n16222 , C0 , RI1754c610_2);
or ( n46899 , n16221 , n16222 );
buf ( n46900 , n46899 );
not ( n46901 , n45546 );
xor ( n46902 , n31200 , n40828 );
xor ( n46903 , n46902 , n42049 );
and ( n46904 , n46901 , n46903 );
xor ( n46905 , n45543 , n46904 );
not ( n16223 , n29614 );
and ( n16224 , n16223 , RI173e0200_1663);
and ( n16225 , n46905 , n29614 );
or ( n46906 , n16224 , n16225 );
not ( n16226 , RI1754c610_2);
and ( n16227 , n16226 , n46906 );
and ( n16228 , C0 , RI1754c610_2);
or ( n46907 , n16227 , n16228 );
buf ( n46908 , n46907 );
not ( n46909 , n43802 );
and ( n46910 , n46909 , n43901 );
xor ( n46911 , n43799 , n46910 );
not ( n16229 , n29614 );
and ( n16230 , n16229 , RI1739eb30_1982);
and ( n16231 , n46911 , n29614 );
or ( n46912 , n16230 , n16231 );
not ( n16232 , RI1754c610_2);
and ( n16233 , n16232 , n46912 );
and ( n16234 , C0 , RI1754c610_2);
or ( n46913 , n16233 , n16234 );
buf ( n46914 , n46913 );
xor ( n46915 , n36771 , n39208 );
xor ( n46916 , n46915 , n38214 );
xor ( n46917 , n36723 , n30247 );
xor ( n46918 , n46917 , n30461 );
not ( n46919 , n46918 );
xor ( n46920 , n40244 , n35760 );
xor ( n46921 , n46920 , n39333 );
and ( n46922 , n46919 , n46921 );
xor ( n46923 , n46916 , n46922 );
not ( n16235 , n29614 );
and ( n16236 , n16235 , RI173fda80_1519);
and ( n16237 , n46923 , n29614 );
or ( n46924 , n16236 , n16237 );
not ( n16238 , RI1754c610_2);
and ( n16239 , n16238 , n46924 );
and ( n16240 , C0 , RI1754c610_2);
or ( n46925 , n16239 , n16240 );
buf ( n46926 , n46925 );
not ( n46927 , n45782 );
and ( n46928 , n46927 , n43722 );
xor ( n46929 , n45779 , n46928 );
not ( n16241 , n29614 );
and ( n16242 , n16241 , RI174101d0_1429);
and ( n16243 , n46929 , n29614 );
or ( n46930 , n16242 , n16243 );
not ( n16244 , RI1754c610_2);
and ( n16245 , n16244 , n46930 );
and ( n16246 , C0 , RI1754c610_2);
or ( n46931 , n16245 , n16246 );
buf ( n46932 , n46931 );
xor ( n46933 , n36629 , n40412 );
xor ( n46934 , n46933 , n40437 );
not ( n46935 , n39314 );
and ( n46936 , n46935 , n39316 );
xor ( n46937 , n46934 , n46936 );
not ( n16247 , n29614 );
and ( n16248 , n16247 , RI17398c08_2011);
and ( n16249 , n46937 , n29614 );
or ( n46938 , n16248 , n16249 );
not ( n16250 , RI1754c610_2);
and ( n16251 , n16250 , n46938 );
and ( n16252 , C0 , RI1754c610_2);
or ( n46939 , n16251 , n16252 );
buf ( n46940 , n46939 );
xor ( n46941 , n36827 , n44146 );
xor ( n46942 , n46941 , n41198 );
not ( n46943 , n35362 );
and ( n46944 , n46943 , n35418 );
xor ( n46945 , n46942 , n46944 );
not ( n16253 , n29614 );
and ( n16254 , n16253 , RI1747ef90_1117);
and ( n16255 , n46945 , n29614 );
or ( n46946 , n16254 , n16255 );
not ( n16256 , RI1754c610_2);
and ( n16257 , n16256 , n46946 );
and ( n16258 , C0 , RI1754c610_2);
or ( n46947 , n16257 , n16258 );
buf ( n46948 , n46947 );
not ( n46949 , n46550 );
xor ( n46950 , n40197 , n34041 );
xor ( n46951 , n46950 , n41934 );
and ( n46952 , n46949 , n46951 );
xor ( n46953 , n45324 , n46952 );
not ( n16259 , n29614 );
and ( n16260 , n16259 , RI173bd0d0_1834);
and ( n16261 , n46953 , n29614 );
or ( n46954 , n16260 , n16261 );
not ( n16262 , RI1754c610_2);
and ( n16263 , n16262 , n46954 );
and ( n16264 , C0 , RI1754c610_2);
or ( n46955 , n16263 , n16264 );
buf ( n46956 , n46955 );
not ( n46957 , n41405 );
xor ( n46958 , n36923 , n32620 );
xor ( n46959 , n46958 , n33337 );
and ( n46960 , n46957 , n46959 );
xor ( n46961 , n41402 , n46960 );
not ( n16265 , n29614 );
and ( n16266 , n16265 , RI1748f958_1036);
and ( n16267 , n46961 , n29614 );
or ( n46962 , n16266 , n16267 );
not ( n16268 , RI1754c610_2);
and ( n16269 , n16268 , n46962 );
and ( n16270 , C0 , RI1754c610_2);
or ( n46963 , n16269 , n16270 );
buf ( n46964 , n46963 );
xor ( n46965 , n36002 , n35438 );
xor ( n46966 , n46965 , n35458 );
xor ( n46967 , n35606 , n41543 );
xor ( n46968 , n46967 , n34669 );
not ( n46969 , n46968 );
xor ( n46970 , n37885 , n36102 );
xor ( n46971 , n46970 , n32048 );
and ( n46972 , n46969 , n46971 );
xor ( n46973 , n46966 , n46972 );
not ( n16271 , n29614 );
and ( n16272 , n16271 , RI173c15b8_1813);
and ( n16273 , n46973 , n29614 );
or ( n46974 , n16272 , n16273 );
not ( n16274 , RI1754c610_2);
and ( n16275 , n16274 , n46974 );
and ( n16276 , C0 , RI1754c610_2);
or ( n46975 , n16275 , n16276 );
buf ( n46976 , n46975 );
xor ( n46977 , n37843 , n33697 );
xor ( n46978 , n46977 , n35128 );
xor ( n46979 , n32852 , n37203 );
xor ( n46980 , n46979 , n34150 );
not ( n46981 , n46980 );
xor ( n46982 , n36194 , n32309 );
xor ( n46983 , n46982 , n32923 );
and ( n46984 , n46981 , n46983 );
xor ( n46985 , n46978 , n46984 );
not ( n16277 , n29614 );
and ( n16278 , n16277 , RI17500530_759);
and ( n16279 , n46985 , n29614 );
or ( n46986 , n16278 , n16279 );
not ( n16280 , RI1754c610_2);
and ( n16281 , n16280 , n46986 );
and ( n16282 , C0 , RI1754c610_2);
or ( n46987 , n16281 , n16282 );
buf ( n46988 , n46987 );
and ( n46989 , RI1754c160_12 , n34844 );
and ( n46990 , RI1754c160_12 , n34847 );
and ( n46991 , RI1754c160_12 , n34850 );
and ( n46992 , RI1754c160_12 , n34852 );
and ( n46993 , RI1754c160_12 , n34854 );
and ( n46994 , RI1754c160_12 , n34856 );
or ( n46995 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , C0 , C0 );
not ( n16283 , n34859 );
and ( n16284 , n16283 , n46995 );
and ( n16285 , RI1754c160_12 , n34859 );
or ( n46996 , n16284 , n16285 );
not ( n16286 , RI19a22f70_2797);
and ( n16287 , n16286 , n46996 );
and ( n16288 , C0 , RI19a22f70_2797);
or ( n46997 , n16287 , n16288 );
not ( n16289 , n27683 );
and ( n16290 , n16289 , RI19a8d230_2703);
and ( n16291 , n46997 , n27683 );
or ( n46998 , n16290 , n16291 );
not ( n16292 , RI1754c610_2);
and ( n16293 , n16292 , n46998 );
and ( n16294 , C0 , RI1754c610_2);
or ( n46999 , n16293 , n16294 );
buf ( n47000 , n46999 );
not ( n16295 , n27683 );
and ( n16296 , n16295 , RI19ab2670_2436);
and ( n16297 , RI19abc4e0_2365 , n27683 );
or ( n47001 , n16296 , n16297 );
not ( n16298 , RI1754c610_2);
and ( n16299 , n16298 , n47001 );
and ( n16300 , C0 , RI1754c610_2);
or ( n47002 , n16299 , n16300 );
buf ( n47003 , n47002 );
not ( n47004 , n45044 );
and ( n47005 , n47004 , n46059 );
xor ( n47006 , n45041 , n47005 );
not ( n16301 , n29614 );
and ( n16302 , n16301 , RI1746a428_1218);
and ( n16303 , n47006 , n29614 );
or ( n47007 , n16302 , n16303 );
not ( n16304 , RI1754c610_2);
and ( n16305 , n16304 , n47007 );
and ( n16306 , C0 , RI1754c610_2);
or ( n47008 , n16305 , n16306 );
buf ( n47009 , n47008 );
not ( n47010 , n45947 );
xor ( n47011 , n29591 , n40051 );
xor ( n47012 , n47011 , n37074 );
and ( n47013 , n47010 , n47012 );
xor ( n47014 , n45944 , n47013 );
not ( n16307 , n29614 );
and ( n16308 , n16307 , RI174793b0_1145);
and ( n16309 , n47014 , n29614 );
or ( n47015 , n16308 , n16309 );
not ( n16310 , RI1754c610_2);
and ( n16311 , n16310 , n47015 );
and ( n16312 , C0 , RI1754c610_2);
or ( n47016 , n16311 , n16312 );
buf ( n47017 , n47016 );
xor ( n47018 , n40236 , n35710 );
xor ( n47019 , n47018 , n35760 );
xor ( n47020 , n32518 , n37651 );
xor ( n47021 , n47020 , n39182 );
not ( n47022 , n47021 );
xor ( n47023 , n32898 , n38553 );
xor ( n47024 , n47023 , n41659 );
and ( n47025 , n47022 , n47024 );
xor ( n47026 , n47019 , n47025 );
not ( n16313 , n29614 );
and ( n16314 , n16313 , RI173e22d0_1653);
and ( n16315 , n47026 , n29614 );
or ( n47027 , n16314 , n16315 );
not ( n16316 , RI1754c610_2);
and ( n16317 , n16316 , n47027 );
and ( n16318 , C0 , RI1754c610_2);
or ( n47028 , n16317 , n16318 );
buf ( n47029 , n47028 );
xor ( n47030 , n34724 , n42605 );
xor ( n47031 , n47030 , n42619 );
xor ( n47032 , n36686 , n39655 );
xor ( n47033 , n47032 , n41125 );
not ( n47034 , n47033 );
xor ( n47035 , n38178 , n32220 );
xor ( n47036 , n47035 , n32309 );
and ( n47037 , n47034 , n47036 );
xor ( n47038 , n47031 , n47037 );
not ( n16319 , n29614 );
and ( n16320 , n16319 , RI17405dc0_1479);
and ( n16321 , n47038 , n29614 );
or ( n47039 , n16320 , n16321 );
not ( n16322 , RI1754c610_2);
and ( n16323 , n16322 , n47039 );
and ( n16324 , C0 , RI1754c610_2);
or ( n47040 , n16323 , n16324 );
buf ( n47041 , n47040 );
not ( n16325 , n27683 );
and ( n16326 , n16325 , RI19aad120_2475);
and ( n16327 , RI19ab6ae0_2404 , n27683 );
or ( n47042 , n16326 , n16327 );
not ( n16328 , RI1754c610_2);
and ( n16329 , n16328 , n47042 );
and ( n16330 , C0 , RI1754c610_2);
or ( n47043 , n16329 , n16330 );
buf ( n47044 , n47043 );
not ( n16331 , n27683 );
and ( n16332 , n16331 , RI19ace3c0_2223);
and ( n16333 , RI19a96998_2636 , n27683 );
or ( n47045 , n16332 , n16333 );
not ( n16334 , RI1754c610_2);
and ( n16335 , n16334 , n47045 );
and ( n16336 , C0 , RI1754c610_2);
or ( n47046 , n16335 , n16336 );
buf ( n47047 , n47046 );
not ( n47048 , n41436 );
xor ( n47049 , n30555 , n38167 );
xor ( n47050 , n47049 , n33728 );
and ( n47051 , n47048 , n47050 );
xor ( n47052 , n41433 , n47051 );
not ( n16337 , n29614 );
and ( n16338 , n16337 , RI173be7c8_1827);
and ( n16339 , n47052 , n29614 );
or ( n47053 , n16338 , n16339 );
not ( n16340 , RI1754c610_2);
and ( n16341 , n16340 , n47053 );
and ( n16342 , C0 , RI1754c610_2);
or ( n47054 , n16341 , n16342 );
buf ( n47055 , n47054 );
not ( n47056 , n45466 );
and ( n47057 , n47056 , n40130 );
xor ( n47058 , n45463 , n47057 );
not ( n16343 , n29614 );
and ( n16344 , n16343 , RI17493e40_1015);
and ( n16345 , n47058 , n29614 );
or ( n47059 , n16344 , n16345 );
not ( n16346 , RI1754c610_2);
and ( n16347 , n16346 , n47059 );
and ( n16348 , C0 , RI1754c610_2);
or ( n47060 , n16347 , n16348 );
buf ( n47061 , n47060 );
xor ( n47062 , n38026 , n41690 );
xor ( n47063 , n47062 , n39506 );
xor ( n47064 , n37897 , n36102 );
xor ( n47065 , n47064 , n32048 );
not ( n47066 , n47065 );
xor ( n47067 , n34685 , n42605 );
xor ( n47068 , n47067 , n42619 );
and ( n47069 , n47066 , n47068 );
xor ( n47070 , n47063 , n47069 );
not ( n16349 , n29614 );
and ( n16350 , n16349 , RI1752bcd0_630);
and ( n16351 , n47070 , n29614 );
or ( n47071 , n16350 , n16351 );
not ( n16352 , RI1754c610_2);
and ( n16353 , n16352 , n47071 );
and ( n16354 , C0 , RI1754c610_2);
or ( n47072 , n16353 , n16354 );
buf ( n47073 , n47072 );
not ( n47074 , n46632 );
xor ( n47075 , n27951 , n42344 );
xor ( n47076 , n47075 , n41799 );
and ( n47077 , n47074 , n47076 );
xor ( n47078 , n46629 , n47077 );
not ( n16355 , n29614 );
and ( n16356 , n16355 , RI17446938_1392);
and ( n16357 , n47078 , n29614 );
or ( n47079 , n16356 , n16357 );
not ( n16358 , RI1754c610_2);
and ( n16359 , n16358 , n47079 );
and ( n16360 , C0 , RI1754c610_2);
or ( n47080 , n16359 , n16360 );
buf ( n47081 , n47080 );
not ( n16361 , n27683 );
and ( n16362 , n16361 , RI19abe6a0_2346);
and ( n16363 , RI19ac74a8_2275 , n27683 );
or ( n47082 , n16362 , n16363 );
not ( n16364 , RI1754c610_2);
and ( n16365 , n16364 , n47082 );
and ( n16366 , C0 , RI1754c610_2);
or ( n47083 , n16365 , n16366 );
buf ( n47084 , n47083 );
buf ( n47085 , RI1747ef90_1117);
buf ( n47086 , RI17483b08_1094);
buf ( n47087 , RI1750d2f8_725);
buf ( n47088 , RI17514eb8_701);
not ( n16367 , n27683 );
and ( n16368 , n16367 , RI19acfd88_2212);
and ( n16369 , RI19aa7540_2514 , n27683 );
or ( n47089 , n16368 , n16369 );
not ( n16370 , RI1754c610_2);
and ( n16371 , n16370 , n47089 );
and ( n16372 , C0 , RI1754c610_2);
or ( n47090 , n16371 , n16372 );
buf ( n47091 , n47090 );
not ( n16373 , n27683 );
and ( n16374 , n16373 , RI19aa8da0_2504);
and ( n16375 , RI19ab2d78_2433 , n27683 );
or ( n47092 , n16374 , n16375 );
not ( n16376 , RI1754c610_2);
and ( n16377 , n16376 , n47092 );
and ( n16378 , C0 , RI1754c610_2);
or ( n47093 , n16377 , n16378 );
buf ( n47094 , n47093 );
not ( n16379 , n34859 );
and ( n16380 , n16379 , C0 );
and ( n16381 , RI1754a900_64 , n34859 );
or ( n47095 , n16380 , n16381 );
not ( n16382 , RI19a22f70_2797);
and ( n16383 , n16382 , n47095 );
and ( n16384 , C0 , RI19a22f70_2797);
or ( n47096 , n16383 , n16384 );
not ( n16385 , n27683 );
and ( n16386 , n16385 , RI19ab3a20_2426);
and ( n16387 , n47096 , n27683 );
or ( n47097 , n16386 , n16387 );
not ( n16388 , RI1754c610_2);
and ( n16389 , n16388 , n47097 );
and ( n16390 , C0 , RI1754c610_2);
or ( n47098 , n16389 , n16390 );
buf ( n47099 , n47098 );
buf ( n47100 , RI1747f968_1114);
buf ( n47101 , RI174bae28_829);
buf ( n47102 , RI174ca080_782);
and ( n47103 , RI19a24ed8_2782 , n43086 );
not ( n16391 , n43088 );
and ( n16392 , n16391 , RI19a24c80_2783);
and ( n16393 , n47103 , n43088 );
or ( n47104 , n16392 , n16393 );
not ( n16394 , RI1754c610_2);
and ( n16395 , n16394 , n47104 );
and ( n16396 , C0 , RI1754c610_2);
or ( n47105 , n16395 , n16396 );
buf ( n47106 , n47105 );
buf ( n47107 , RI1748f958_1036);
xor ( n47108 , n33757 , n40486 );
xor ( n47109 , n47108 , n40516 );
not ( n47110 , n44193 );
and ( n47111 , n47110 , n42201 );
xor ( n47112 , n47109 , n47111 );
not ( n16397 , n29614 );
and ( n16398 , n16397 , RI1750e798_721);
and ( n16399 , n47112 , n29614 );
or ( n47113 , n16398 , n16399 );
not ( n16400 , RI1754c610_2);
and ( n16401 , n16400 , n47113 );
and ( n16402 , C0 , RI1754c610_2);
or ( n47114 , n16401 , n16402 );
buf ( n47115 , n47114 );
not ( n16403 , n27683 );
and ( n16404 , n16403 , RI19a8bfe8_2711);
and ( n16405 , RI19a96038_2640 , n27683 );
or ( n47116 , n16404 , n16405 );
not ( n16406 , RI1754c610_2);
and ( n16407 , n16406 , n47116 );
and ( n16408 , C0 , RI1754c610_2);
or ( n47117 , n16407 , n16408 );
buf ( n47118 , n47117 );
not ( n47119 , n42225 );
and ( n47120 , n47119 , n42227 );
xor ( n47121 , n39291 , n47120 );
not ( n16409 , n29614 );
and ( n16410 , n16409 , RI1739e7e8_1983);
and ( n16411 , n47121 , n29614 );
or ( n47122 , n16410 , n16411 );
not ( n16412 , RI1754c610_2);
and ( n16413 , n16412 , n47122 );
and ( n16414 , C0 , RI1754c610_2);
or ( n47123 , n16413 , n16414 );
buf ( n47124 , n47123 );
xor ( n47125 , n42497 , n30461 );
xor ( n47126 , n47125 , n39262 );
xor ( n47127 , n42626 , n35052 );
xor ( n47128 , n47127 , n35069 );
not ( n47129 , n47128 );
and ( n47130 , n47129 , n46391 );
xor ( n47131 , n47126 , n47130 );
not ( n16415 , n29614 );
and ( n16416 , n16415 , RI174b9988_833);
and ( n16417 , n47131 , n29614 );
or ( n47132 , n16416 , n16417 );
not ( n16418 , RI1754c610_2);
and ( n16419 , n16418 , n47132 );
and ( n16420 , C0 , RI1754c610_2);
or ( n47133 , n16419 , n16420 );
buf ( n47134 , n47133 );
buf ( n47135 , RI17484b70_1089);
buf ( n47136 , RI1750b930_730);
not ( n47137 , n42434 );
xor ( n47138 , n38484 , n39771 );
xor ( n47139 , n47138 , n39791 );
and ( n47140 , n47137 , n47139 );
xor ( n47141 , n42431 , n47140 );
not ( n16421 , n29614 );
and ( n16422 , n16421 , RI1746c840_1207);
and ( n16423 , n47141 , n29614 );
or ( n47142 , n16422 , n16423 );
not ( n16424 , RI1754c610_2);
and ( n16425 , n16424 , n47142 );
and ( n16426 , C0 , RI1754c610_2);
or ( n47143 , n16425 , n16426 );
buf ( n47144 , n47143 );
buf ( n47145 , RI174b8308_838);
buf ( n47146 , RI1749e8e0_963);
not ( n47147 , n43499 );
and ( n47148 , n47147 , n44085 );
xor ( n47149 , n43496 , n47148 );
not ( n16427 , n29614 );
and ( n16428 , n16427 , RI174589f8_1304);
and ( n16429 , n47149 , n29614 );
or ( n47150 , n16428 , n16429 );
not ( n16430 , RI1754c610_2);
and ( n16431 , n16430 , n47150 );
and ( n16432 , C0 , RI1754c610_2);
or ( n47151 , n16431 , n16432 );
buf ( n47152 , n47151 );
not ( n16433 , n27683 );
and ( n16434 , n16433 , RI19a9e288_2583);
and ( n16435 , RI19aa7c48_2511 , n27683 );
or ( n47153 , n16434 , n16435 );
not ( n16436 , RI1754c610_2);
and ( n16437 , n16436 , n47153 );
and ( n16438 , C0 , RI1754c610_2);
or ( n47154 , n16437 , n16438 );
buf ( n47155 , n47154 );
xor ( n47156 , n41055 , n36339 );
xor ( n47157 , n47156 , n36377 );
not ( n47158 , n47157 );
xor ( n47159 , n40306 , n37869 );
xor ( n47160 , n47159 , n38948 );
and ( n47161 , n47158 , n47160 );
xor ( n47162 , n43040 , n47161 );
not ( n16439 , n29614 );
and ( n16440 , n16439 , RI173efea8_1586);
and ( n16441 , n47162 , n29614 );
or ( n47163 , n16440 , n16441 );
not ( n16442 , RI1754c610_2);
and ( n16443 , n16442 , n47163 );
and ( n16444 , C0 , RI1754c610_2);
or ( n47164 , n16443 , n16444 );
buf ( n47165 , n47164 );
buf ( n47166 , RI174758a0_1163);
xor ( n47167 , n38139 , n31053 );
xor ( n47168 , n47167 , n35494 );
xor ( n47169 , n31718 , n30741 );
xor ( n47170 , n47169 , n40769 );
not ( n47171 , n47170 );
xor ( n47172 , n35457 , n32715 );
xor ( n47173 , n47172 , n36654 );
and ( n47174 , n47171 , n47173 );
xor ( n47175 , n47168 , n47174 );
not ( n16445 , n29614 );
and ( n16446 , n16445 , RI1745a438_1296);
and ( n16447 , n47175 , n29614 );
or ( n47176 , n16446 , n16447 );
not ( n16448 , RI1754c610_2);
and ( n16449 , n16448 , n47176 );
and ( n16450 , C0 , RI1754c610_2);
or ( n47177 , n16449 , n16450 );
buf ( n47178 , n47177 );
buf ( n47179 , RI1746a770_1217);
xor ( n47180 , n42175 , n41215 );
xor ( n47181 , n47180 , n33824 );
not ( n47182 , n41017 );
and ( n47183 , n47182 , n41019 );
xor ( n47184 , n47181 , n47183 );
not ( n16451 , n29614 );
and ( n16452 , n16451 , RI17470698_1188);
and ( n16453 , n47184 , n29614 );
or ( n47185 , n16452 , n16453 );
not ( n16454 , RI1754c610_2);
and ( n16455 , n16454 , n47185 );
and ( n16456 , C0 , RI1754c610_2);
or ( n47186 , n16455 , n16456 );
buf ( n47187 , n47186 );
not ( n16457 , n27683 );
and ( n16458 , n16457 , RI19a915b0_2673);
and ( n16459 , RI19a9b8d0_2601 , n27683 );
or ( n47188 , n16458 , n16459 );
not ( n16460 , RI1754c610_2);
and ( n16461 , n16460 , n47188 );
and ( n16462 , C0 , RI1754c610_2);
or ( n47189 , n16461 , n16462 );
buf ( n47190 , n47189 );
buf ( n47191 , RI174b1030_873);
buf ( n47192 , RI174a5f00_927);
xor ( n47193 , n38782 , n40516 );
xor ( n47194 , n47193 , n40966 );
not ( n47195 , n47031 );
and ( n47196 , n47195 , n47033 );
xor ( n47197 , n47194 , n47196 );
not ( n16463 , n29614 );
and ( n16464 , n16463 , RI173f74c8_1550);
and ( n16465 , n47197 , n29614 );
or ( n47198 , n16464 , n16465 );
not ( n16466 , RI1754c610_2);
and ( n16467 , n16466 , n47198 );
and ( n16468 , C0 , RI1754c610_2);
or ( n47199 , n16467 , n16468 );
buf ( n47200 , n47199 );
xor ( n47201 , n41985 , n39886 );
xor ( n47202 , n47201 , n36998 );
not ( n47203 , n31054 );
and ( n47204 , n47203 , n31318 );
xor ( n47205 , n47202 , n47204 );
not ( n16469 , n29614 );
and ( n16470 , n16469 , RI17526528_647);
and ( n16471 , n47205 , n29614 );
or ( n47206 , n16470 , n16471 );
not ( n16472 , RI1754c610_2);
and ( n16473 , n16472 , n47206 );
and ( n16474 , C0 , RI1754c610_2);
or ( n47207 , n16473 , n16474 );
buf ( n47208 , n47207 );
not ( n16475 , n27683 );
and ( n16476 , n16475 , RI19aa7e28_2510);
and ( n16477 , RI19ab1ef0_2440 , n27683 );
or ( n47209 , n16476 , n16477 );
not ( n16478 , RI1754c610_2);
and ( n16479 , n16478 , n47209 );
and ( n16480 , C0 , RI1754c610_2);
or ( n47210 , n16479 , n16480 );
buf ( n47211 , n47210 );
and ( n47212 , RI1754bf08_17 , n34844 );
and ( n47213 , RI1754bf08_17 , n34847 );
and ( n47214 , RI1754bf08_17 , n34850 );
and ( n47215 , RI1754bf08_17 , n34852 );
and ( n47216 , RI1754bf08_17 , n34854 );
and ( n47217 , RI1754bf08_17 , n34856 );
or ( n47218 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , C0 , C0 );
not ( n16481 , n34859 );
and ( n16482 , n16481 , n47218 );
and ( n16483 , RI1754bf08_17 , n34859 );
or ( n47219 , n16482 , n16483 );
not ( n16484 , RI19a22f70_2797);
and ( n16485 , n16484 , n47219 );
and ( n16486 , C0 , RI19a22f70_2797);
or ( n47220 , n16485 , n16486 );
not ( n16487 , n27683 );
and ( n16488 , n16487 , RI19a95048_2647);
and ( n16489 , n47220 , n27683 );
or ( n47221 , n16488 , n16489 );
not ( n16490 , RI1754c610_2);
and ( n16491 , n16490 , n47221 );
and ( n16492 , C0 , RI1754c610_2);
or ( n47222 , n16491 , n16492 );
buf ( n47223 , n47222 );
not ( n47224 , n45312 );
xor ( n47225 , n41361 , n36062 );
xor ( n47226 , n47225 , n36102 );
and ( n47227 , n47224 , n47226 );
xor ( n47228 , n45309 , n47227 );
not ( n16493 , n29614 );
and ( n16494 , n16493 , RI174b5860_851);
and ( n16495 , n47228 , n29614 );
or ( n47229 , n16494 , n16495 );
not ( n16496 , RI1754c610_2);
and ( n16497 , n16496 , n47229 );
and ( n16498 , C0 , RI1754c610_2);
or ( n47230 , n16497 , n16498 );
buf ( n47231 , n47230 );
not ( n16499 , n27683 );
and ( n16500 , n16499 , RI19acb120_2247);
and ( n16501 , RI19a86750_2749 , n27683 );
or ( n47232 , n16500 , n16501 );
not ( n16502 , RI1754c610_2);
and ( n16503 , n16502 , n47232 );
and ( n16504 , C0 , RI1754c610_2);
or ( n47233 , n16503 , n16504 );
buf ( n47234 , n47233 );
not ( n47235 , n46181 );
and ( n47236 , n47235 , n46183 );
xor ( n47237 , n46257 , n47236 );
not ( n16505 , n29614 );
and ( n16506 , n16505 , RI174a6f68_922);
and ( n16507 , n47237 , n29614 );
or ( n47238 , n16506 , n16507 );
not ( n16508 , RI1754c610_2);
and ( n16509 , n16508 , n47238 );
and ( n16510 , C0 , RI1754c610_2);
or ( n47239 , n16509 , n16510 );
buf ( n47240 , n47239 );
not ( n16511 , n27683 );
and ( n16512 , n16511 , RI19aa05b0_2566);
and ( n16513 , RI19aaa150_2495 , n27683 );
or ( n47241 , n16512 , n16513 );
not ( n16514 , RI1754c610_2);
and ( n16515 , n16514 , n47241 );
and ( n16516 , C0 , RI1754c610_2);
or ( n47242 , n16515 , n16516 );
buf ( n47243 , n47242 );
buf ( n47244 , RI17477628_1154);
buf ( n47245 , RI17466c60_1235);
xor ( n47246 , n35573 , n37490 );
xor ( n47247 , n47246 , n41316 );
not ( n47248 , n45789 );
and ( n47249 , n47248 , n45791 );
xor ( n47250 , n47247 , n47249 );
not ( n16517 , n29614 );
and ( n16518 , n16517 , RI1739e4a0_1984);
and ( n16519 , n47250 , n29614 );
or ( n47251 , n16518 , n16519 );
not ( n16520 , RI1754c610_2);
and ( n16521 , n16520 , n47251 );
and ( n16522 , C0 , RI1754c610_2);
or ( n47252 , n16521 , n16522 );
buf ( n47253 , n47252 );
xor ( n47254 , n40102 , n39740 );
xor ( n47255 , n47254 , n41099 );
not ( n47256 , n38533 );
and ( n47257 , n47256 , n38554 );
xor ( n47258 , n47255 , n47257 );
not ( n16523 , n29614 );
and ( n16524 , n16523 , RI17459da8_1298);
and ( n16525 , n47258 , n29614 );
or ( n47259 , n16524 , n16525 );
not ( n16526 , RI1754c610_2);
and ( n16527 , n16526 , n47259 );
and ( n16528 , C0 , RI1754c610_2);
or ( n47260 , n16527 , n16528 );
buf ( n47261 , n47260 );
not ( n47262 , n43180 );
and ( n47263 , n47262 , n43524 );
xor ( n47264 , n43177 , n47263 );
not ( n16529 , n29614 );
and ( n16530 , n16529 , RI1750b930_730);
and ( n16531 , n47264 , n29614 );
or ( n47265 , n16530 , n16531 );
not ( n16532 , RI1754c610_2);
and ( n16533 , n16532 , n47265 );
and ( n16534 , C0 , RI1754c610_2);
or ( n47266 , n16533 , n16534 );
buf ( n47267 , n47266 );
not ( n47268 , n44645 );
and ( n47269 , n47268 , n44647 );
xor ( n47270 , n40860 , n47269 );
not ( n16535 , n29614 );
and ( n16536 , n16535 , RI1747dbe0_1123);
and ( n16537 , n47270 , n29614 );
or ( n47271 , n16536 , n16537 );
not ( n16538 , RI1754c610_2);
and ( n16539 , n16538 , n47271 );
and ( n16540 , C0 , RI1754c610_2);
or ( n47272 , n16539 , n16540 );
buf ( n47273 , n47272 );
not ( n47274 , n44206 );
and ( n47275 , n47274 , n46838 );
xor ( n47276 , n44203 , n47275 );
not ( n16541 , n29614 );
and ( n16542 , n16541 , RI174a3ae8_938);
and ( n16543 , n47276 , n29614 );
or ( n47277 , n16542 , n16543 );
not ( n16544 , RI1754c610_2);
and ( n16545 , n16544 , n47277 );
and ( n16546 , C0 , RI1754c610_2);
or ( n47278 , n16545 , n16546 );
buf ( n47279 , n47278 );
not ( n47280 , n41451 );
and ( n47281 , n47280 , n43857 );
xor ( n47282 , n41445 , n47281 );
not ( n16547 , n29614 );
and ( n16548 , n16547 , RI17341a70_2121);
and ( n16549 , n47282 , n29614 );
or ( n47283 , n16548 , n16549 );
not ( n16550 , RI1754c610_2);
and ( n16551 , n16550 , n47283 );
and ( n16552 , C0 , RI1754c610_2);
or ( n47284 , n16551 , n16552 );
buf ( n47285 , n47284 );
not ( n47286 , n46450 );
xor ( n47287 , n33715 , n35514 );
xor ( n47288 , n47287 , n40486 );
and ( n47289 , n47286 , n47288 );
xor ( n47290 , n43342 , n47289 );
not ( n16553 , n29614 );
and ( n16554 , n16553 , RI1733f658_2132);
and ( n16555 , n47290 , n29614 );
or ( n47291 , n16554 , n16555 );
not ( n16556 , RI1754c610_2);
and ( n16557 , n16556 , n47291 );
and ( n16558 , C0 , RI1754c610_2);
or ( n47292 , n16557 , n16558 );
buf ( n47293 , n47292 );
xor ( n47294 , n38213 , n37696 );
xor ( n47295 , n47294 , n39450 );
not ( n47296 , n47295 );
and ( n47297 , n47296 , n43969 );
xor ( n47298 , n44108 , n47297 );
not ( n16559 , n29614 );
and ( n16560 , n16559 , RI17522220_660);
and ( n16561 , n47298 , n29614 );
or ( n47299 , n16560 , n16561 );
not ( n16562 , RI1754c610_2);
and ( n16563 , n16562 , n47299 );
and ( n16564 , C0 , RI1754c610_2);
or ( n47300 , n16563 , n16564 );
buf ( n47301 , n47300 );
buf ( n47302 , RI1747e270_1121);
buf ( n47303 , RI1747b7c8_1134);
buf ( n47304 , RI17515e30_698);
xor ( n47305 , n35167 , n37915 );
xor ( n47306 , n47305 , n43492 );
xor ( n47307 , n36338 , n40718 );
xor ( n47308 , n47307 , n38676 );
not ( n47309 , n47308 );
xor ( n47310 , n39692 , n33337 );
xor ( n47311 , n47310 , n33397 );
and ( n47312 , n47309 , n47311 );
xor ( n47313 , n47306 , n47312 );
not ( n16565 , n29614 );
and ( n16566 , n16565 , RI17507b50_742);
and ( n16567 , n47313 , n29614 );
or ( n47314 , n16566 , n16567 );
not ( n16568 , RI1754c610_2);
and ( n16569 , n16568 , n47314 );
and ( n16570 , C0 , RI1754c610_2);
or ( n47315 , n16569 , n16570 );
buf ( n47316 , n47315 );
xor ( n47317 , n38944 , n36917 );
xor ( n47318 , n47317 , n36947 );
not ( n47319 , n46035 );
and ( n47320 , n47319 , n46037 );
xor ( n47321 , n47318 , n47320 );
not ( n16571 , n29614 );
and ( n16572 , n16571 , RI174cbf70_776);
and ( n16573 , n47321 , n29614 );
or ( n47322 , n16572 , n16573 );
not ( n16574 , RI1754c610_2);
and ( n16575 , n16574 , n47322 );
and ( n16576 , C0 , RI1754c610_2);
or ( n47323 , n16575 , n16576 );
buf ( n47324 , n47323 );
not ( n16577 , n27683 );
and ( n16578 , n16577 , RI19a841d0_2765);
and ( n16579 , RI19abcfa8_2359 , n27683 );
or ( n47325 , n16578 , n16579 );
not ( n16580 , RI1754c610_2);
and ( n16581 , n16580 , n47325 );
and ( n16582 , C0 , RI1754c610_2);
or ( n47326 , n16581 , n16582 );
buf ( n47327 , n47326 );
not ( n16583 , n27683 );
and ( n16584 , n16583 , RI19a838e8_2769);
and ( n16585 , RI19ab8778_2392 , n27683 );
or ( n47328 , n16584 , n16585 );
not ( n16586 , RI1754c610_2);
and ( n16587 , n16586 , n47328 );
and ( n16588 , C0 , RI1754c610_2);
or ( n47329 , n16587 , n16588 );
buf ( n47330 , n47329 );
xor ( n47331 , n41189 , n34622 );
xor ( n47332 , n47331 , n39397 );
xor ( n47333 , n36602 , n39791 );
xor ( n47334 , n47333 , n40915 );
not ( n47335 , n47334 );
xor ( n47336 , n38114 , n40111 );
xor ( n47337 , n47336 , n43278 );
and ( n47338 , n47335 , n47337 );
xor ( n47339 , n47332 , n47338 );
not ( n16589 , n29614 );
and ( n16590 , n16589 , RI1739e158_1985);
and ( n16591 , n47339 , n29614 );
or ( n47340 , n16590 , n16591 );
not ( n16592 , RI1754c610_2);
and ( n16593 , n16592 , n47340 );
and ( n16594 , C0 , RI1754c610_2);
or ( n47341 , n16593 , n16594 );
buf ( n47342 , n47341 );
not ( n16595 , n27683 );
and ( n16596 , n16595 , RI19a93d88_2655);
and ( n16597 , RI19a9e030_2584 , n27683 );
or ( n47343 , n16596 , n16597 );
not ( n16598 , RI1754c610_2);
and ( n16599 , n16598 , n47343 );
and ( n16600 , C0 , RI1754c610_2);
or ( n47344 , n16599 , n16600 );
buf ( n47345 , n47344 );
and ( n47346 , RI1754ac48_57 , n34844 );
buf ( n47347 , n47346 );
not ( n16601 , n34859 );
and ( n16602 , n16601 , n47347 );
and ( n16603 , RI1754ac48_57 , n34859 );
or ( n47348 , n16602 , n16603 );
not ( n16604 , RI19a22f70_2797);
and ( n16605 , n16604 , n47348 );
and ( n16606 , C0 , RI19a22f70_2797);
or ( n47349 , n16605 , n16606 );
not ( n16607 , n27683 );
and ( n16608 , n16607 , RI19a23150_2796);
and ( n16609 , n47349 , n27683 );
or ( n47350 , n16608 , n16609 );
not ( n16610 , RI1754c610_2);
and ( n16611 , n16610 , n47350 );
and ( n16612 , C0 , RI1754c610_2);
or ( n47351 , n16611 , n16612 );
buf ( n47352 , n47351 );
not ( n47353 , n44915 );
xor ( n47354 , n39778 , n33175 );
xor ( n47355 , n47354 , n34797 );
and ( n47356 , n47353 , n47355 );
xor ( n47357 , n44912 , n47356 );
not ( n16613 , n29614 );
and ( n16614 , n16613 , RI1744c518_1364);
and ( n16615 , n47357 , n29614 );
or ( n47358 , n16614 , n16615 );
not ( n16616 , RI1754c610_2);
and ( n16617 , n16616 , n47358 );
and ( n16618 , C0 , RI1754c610_2);
or ( n47359 , n16617 , n16618 );
buf ( n47360 , n47359 );
xor ( n47361 , n42251 , n40743 );
xor ( n47362 , n47361 , n36062 );
not ( n47363 , n41936 );
and ( n47364 , n47363 , n41893 );
xor ( n47365 , n47362 , n47364 );
not ( n16619 , n29614 );
and ( n16620 , n16619 , RI174593d0_1301);
and ( n16621 , n47365 , n29614 );
or ( n47366 , n16620 , n16621 );
not ( n16622 , RI1754c610_2);
and ( n16623 , n16622 , n47366 );
and ( n16624 , C0 , RI1754c610_2);
or ( n47367 , n16623 , n16624 );
buf ( n47368 , n47367 );
xor ( n47369 , n30072 , n34755 );
xor ( n47370 , n47369 , n35311 );
xor ( n47371 , n38201 , n37696 );
xor ( n47372 , n47371 , n39450 );
not ( n47373 , n47372 );
and ( n47374 , n47373 , n47332 );
xor ( n47375 , n47370 , n47374 );
not ( n16625 , n29614 );
and ( n16626 , n16625 , RI173406c0_2127);
and ( n16627 , n47375 , n29614 );
or ( n47376 , n16626 , n16627 );
not ( n16628 , RI1754c610_2);
and ( n16629 , n16628 , n47376 );
and ( n16630 , C0 , RI1754c610_2);
or ( n47377 , n16629 , n16630 );
buf ( n47378 , n47377 );
not ( n47379 , n44471 );
and ( n47380 , n47379 , n44473 );
xor ( n47381 , n44945 , n47380 );
not ( n16631 , n29614 );
and ( n16632 , n16631 , RI17338038_2168);
and ( n16633 , n47381 , n29614 );
or ( n47382 , n16632 , n16633 );
not ( n16634 , RI1754c610_2);
and ( n16635 , n16634 , n47382 );
and ( n16636 , C0 , RI1754c610_2);
or ( n47383 , n16635 , n16636 );
buf ( n47384 , n47383 );
not ( n16637 , n27683 );
and ( n16638 , n16637 , RI19ab01e0_2453);
and ( n16639 , RI19ab9c18_2382 , n27683 );
or ( n47385 , n16638 , n16639 );
not ( n16640 , RI1754c610_2);
and ( n16641 , n16640 , n47385 );
and ( n16642 , C0 , RI1754c610_2);
or ( n47386 , n16641 , n16642 );
buf ( n47387 , n47386 );
not ( n47388 , n46726 );
xor ( n47389 , n34591 , n35544 );
xor ( n47390 , n47389 , n35594 );
and ( n47391 , n47388 , n47390 );
xor ( n47392 , n46723 , n47391 );
not ( n16643 , n29614 );
and ( n16644 , n16643 , RI173bf830_1822);
and ( n16645 , n47392 , n29614 );
or ( n47393 , n16644 , n16645 );
not ( n16646 , RI1754c610_2);
and ( n16647 , n16646 , n47393 );
and ( n16648 , C0 , RI1754c610_2);
or ( n47394 , n16647 , n16648 );
buf ( n47395 , n47394 );
not ( n16649 , n27683 );
and ( n16650 , n16649 , RI19ac2390_2312);
and ( n16651 , RI19acb4e0_2245 , n27683 );
or ( n47396 , n16650 , n16651 );
not ( n16652 , RI1754c610_2);
and ( n16653 , n16652 , n47396 );
and ( n16654 , C0 , RI1754c610_2);
or ( n47397 , n16653 , n16654 );
buf ( n47398 , n47397 );
xor ( n47399 , n29295 , n40034 );
xor ( n47400 , n47399 , n40051 );
not ( n47401 , n47400 );
and ( n47402 , n47401 , n44303 );
xor ( n47403 , n45905 , n47402 );
not ( n16655 , n29614 );
and ( n16656 , n16655 , RI173df198_1668);
and ( n16657 , n47403 , n29614 );
or ( n47404 , n16656 , n16657 );
not ( n16658 , RI1754c610_2);
and ( n16659 , n16658 , n47404 );
and ( n16660 , C0 , RI1754c610_2);
or ( n47405 , n16659 , n16660 );
buf ( n47406 , n47405 );
and ( n47407 , RI1754bf80_16 , n34844 );
and ( n47408 , RI1754bf80_16 , n34847 );
and ( n47409 , RI1754bf80_16 , n34850 );
and ( n47410 , RI1754bf80_16 , n34852 );
and ( n47411 , RI1754bf80_16 , n34854 );
and ( n47412 , RI1754bf80_16 , n34856 );
or ( n47413 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , C0 , C0 );
not ( n16661 , n34859 );
and ( n16662 , n16661 , n47413 );
and ( n16663 , RI1754bf80_16 , n34859 );
or ( n47414 , n16662 , n16663 );
not ( n16664 , RI19a22f70_2797);
and ( n16665 , n16664 , n47414 );
and ( n16666 , C0 , RI19a22f70_2797);
or ( n47415 , n16665 , n16666 );
not ( n16667 , n27683 );
and ( n16668 , n16667 , RI19a93518_2659);
and ( n16669 , n47415 , n27683 );
or ( n47416 , n16668 , n16669 );
not ( n16670 , RI1754c610_2);
and ( n16671 , n16670 , n47416 );
and ( n16672 , C0 , RI1754c610_2);
or ( n47417 , n16671 , n16672 );
buf ( n47418 , n47417 );
xor ( n47419 , n35479 , n38512 );
xor ( n47420 , n47419 , n38532 );
not ( n47421 , n47420 );
and ( n47422 , n47421 , n43363 );
xor ( n47423 , n42950 , n47422 );
not ( n16673 , n29614 );
and ( n16674 , n16673 , RI173c6130_1790);
and ( n16675 , n47423 , n29614 );
or ( n47424 , n16674 , n16675 );
not ( n16676 , RI1754c610_2);
and ( n16677 , n16676 , n47424 );
and ( n16678 , C0 , RI1754c610_2);
or ( n47425 , n16677 , n16678 );
buf ( n47426 , n47425 );
buf ( n47427 , RI174b2098_868);
buf ( n47428 , RI174a1040_951);
xor ( n47429 , n41759 , n38188 );
xor ( n47430 , n47429 , n36195 );
xor ( n47431 , n31140 , n40828 );
xor ( n47432 , n47431 , n42049 );
not ( n47433 , n47432 );
xor ( n47434 , n40653 , n39282 );
xor ( n47435 , n47434 , n37676 );
and ( n47436 , n47433 , n47435 );
xor ( n47437 , n47430 , n47436 );
not ( n16679 , n29614 );
and ( n16680 , n16679 , RI1733bb48_2150);
and ( n16681 , n47437 , n29614 );
or ( n47438 , n16680 , n16681 );
not ( n16682 , RI1754c610_2);
and ( n16683 , n16682 , n47438 );
and ( n16684 , C0 , RI1754c610_2);
or ( n47439 , n16683 , n16684 );
buf ( n47440 , n47439 );
xor ( n47441 , n42027 , n41049 );
xor ( n47442 , n47441 , n41504 );
not ( n47443 , n47442 );
xor ( n47444 , n35833 , n37129 );
xor ( n47445 , n47444 , n37169 );
and ( n47446 , n47443 , n47445 );
xor ( n47447 , n43297 , n47446 );
not ( n16685 , n29614 );
and ( n16686 , n16685 , RI1747cec0_1127);
and ( n16687 , n47447 , n29614 );
or ( n47448 , n16686 , n16687 );
not ( n16688 , RI1754c610_2);
and ( n16689 , n16688 , n47448 );
and ( n16690 , C0 , RI1754c610_2);
or ( n47449 , n16689 , n16690 );
buf ( n47450 , n47449 );
not ( n47451 , n46578 );
xor ( n47452 , n40161 , n39039 );
xor ( n47453 , n47452 , n39065 );
and ( n47454 , n47451 , n47453 );
xor ( n47455 , n46575 , n47454 );
not ( n16691 , n29614 );
and ( n16692 , n16691 , RI173e1268_1658);
and ( n16693 , n47455 , n29614 );
or ( n47456 , n16692 , n16693 );
not ( n16694 , RI1754c610_2);
and ( n16695 , n16694 , n47456 );
and ( n16696 , C0 , RI1754c610_2);
or ( n47457 , n16695 , n16696 );
buf ( n47458 , n47457 );
not ( n47459 , n44603 );
and ( n47460 , n47459 , n37527 );
xor ( n47461 , n44600 , n47460 );
not ( n16697 , n29614 );
and ( n16698 , n16697 , RI175196e8_687);
and ( n16699 , n47461 , n29614 );
or ( n47462 , n16698 , n16699 );
not ( n16700 , RI1754c610_2);
and ( n16701 , n16700 , n47462 );
and ( n16702 , C0 , RI1754c610_2);
or ( n47463 , n16701 , n16702 );
buf ( n47464 , n47463 );
not ( n47465 , n41393 );
and ( n47466 , n47465 , n43371 );
xor ( n47467 , n41374 , n47466 );
not ( n16703 , n29614 );
and ( n16704 , n16703 , RI17480688_1110);
and ( n16705 , n47467 , n29614 );
or ( n47468 , n16704 , n16705 );
not ( n16706 , RI1754c610_2);
and ( n16707 , n16706 , n47468 );
and ( n16708 , C0 , RI1754c610_2);
or ( n47469 , n16707 , n16708 );
buf ( n47470 , n47469 );
not ( n16709 , n27683 );
and ( n16710 , n16709 , RI19ac9938_2258);
and ( n16711 , RI19a84ba8_2761 , n27683 );
or ( n47471 , n16710 , n16711 );
not ( n16712 , RI1754c610_2);
and ( n16713 , n16712 , n47471 );
and ( n16714 , C0 , RI1754c610_2);
or ( n47472 , n16713 , n16714 );
buf ( n47473 , n47472 );
buf ( n47474 , RI17499a20_987);
not ( n47475 , n43141 );
and ( n47476 , n47475 , n38794 );
xor ( n47477 , n43138 , n47476 );
not ( n16715 , n29614 );
and ( n16716 , n16715 , RI174cedd8_767);
and ( n16717 , n47477 , n29614 );
or ( n47478 , n16716 , n16717 );
not ( n16718 , RI1754c610_2);
and ( n16719 , n16718 , n47478 );
and ( n16720 , C0 , RI1754c610_2);
or ( n47479 , n16719 , n16720 );
buf ( n47480 , n47479 );
buf ( n47481 , RI174b9988_833);
not ( n16721 , n27683 );
and ( n16722 , n16721 , RI19a8d668_2701);
and ( n16723 , RI19a976b8_2630 , n27683 );
or ( n47482 , n16722 , n16723 );
not ( n16724 , RI1754c610_2);
and ( n16725 , n16724 , n47482 );
and ( n16726 , C0 , RI1754c610_2);
or ( n47483 , n16725 , n16726 );
buf ( n47484 , n47483 );
buf ( n47485 , RI174b4b40_855);
buf ( n47486 , RI1749e250_965);
not ( n47487 , n45175 );
and ( n47488 , n47487 , n42980 );
xor ( n47489 , n45172 , n47488 );
not ( n16727 , n29614 );
and ( n16728 , n16727 , RI174a8cf0_913);
and ( n16729 , n47489 , n29614 );
or ( n47490 , n16728 , n16729 );
not ( n16730 , RI1754c610_2);
and ( n16731 , n16730 , n47490 );
and ( n16732 , C0 , RI1754c610_2);
or ( n47491 , n16731 , n16732 );
buf ( n47492 , n47491 );
not ( n47493 , n43916 );
and ( n47494 , n47493 , n44379 );
xor ( n47495 , n43913 , n47494 );
not ( n16733 , n29614 );
and ( n16734 , n16733 , RI173441d0_2109);
and ( n16735 , n47495 , n29614 );
or ( n47496 , n16734 , n16735 );
not ( n16736 , RI1754c610_2);
and ( n16737 , n16736 , n47496 );
and ( n16738 , C0 , RI1754c610_2);
or ( n47497 , n16737 , n16738 );
buf ( n47498 , n47497 );
not ( n47499 , n43797 );
and ( n47500 , n47499 , n43799 );
xor ( n47501 , n43903 , n47500 );
not ( n16739 , n29614 );
and ( n16740 , n16739 , RI17341098_2124);
and ( n16741 , n47501 , n29614 );
or ( n47502 , n16740 , n16741 );
not ( n16742 , RI1754c610_2);
and ( n16743 , n16742 , n47502 );
and ( n16744 , C0 , RI1754c610_2);
or ( n47503 , n16743 , n16744 );
buf ( n47504 , n47503 );
not ( n47505 , n44529 );
and ( n47506 , n47505 , n45687 );
xor ( n47507 , n44526 , n47506 );
not ( n16745 , n29614 );
and ( n16746 , n16745 , RI173cb680_1764);
and ( n16747 , n47507 , n29614 );
or ( n47508 , n16746 , n16747 );
not ( n16748 , RI1754c610_2);
and ( n16749 , n16748 , n47508 );
and ( n16750 , C0 , RI1754c610_2);
or ( n47509 , n16749 , n16750 );
buf ( n47510 , n47509 );
xor ( n47511 , n30740 , n33728 );
xor ( n47512 , n47511 , n33778 );
not ( n47513 , n47512 );
xor ( n47514 , n33089 , n38244 );
xor ( n47515 , n47514 , n37235 );
and ( n47516 , n47513 , n47515 );
xor ( n47517 , n41858 , n47516 );
not ( n16751 , n29614 );
and ( n16752 , n16751 , RI174937b0_1017);
and ( n16753 , n47517 , n29614 );
or ( n47518 , n16752 , n16753 );
not ( n16754 , RI1754c610_2);
and ( n16755 , n16754 , n47518 );
and ( n16756 , C0 , RI1754c610_2);
or ( n47519 , n16755 , n16756 );
buf ( n47520 , n47519 );
not ( n16757 , RI1754c610_2);
and ( n16758 , n16757 , n27689 );
and ( n16759 , C0 , RI1754c610_2);
or ( n47521 , n16758 , n16759 );
buf ( n47522 , n47521 );
not ( n16760 , n27683 );
and ( n16761 , n16760 , RI19a9bb28_2600);
and ( n16762 , RI19aa5218_2529 , n27683 );
or ( n47523 , n16761 , n16762 );
not ( n16763 , RI1754c610_2);
and ( n16764 , n16763 , n47523 );
and ( n16765 , C0 , RI1754c610_2);
or ( n47524 , n16764 , n16765 );
buf ( n47525 , n47524 );
buf ( n47526 , RI174c7c68_789);
xor ( n47527 , n36928 , n32620 );
xor ( n47528 , n47527 , n33337 );
xor ( n47529 , n35613 , n41543 );
xor ( n47530 , n47529 , n34669 );
not ( n47531 , n47530 );
xor ( n47532 , n37893 , n36102 );
xor ( n47533 , n47532 , n32048 );
and ( n47534 , n47531 , n47533 );
xor ( n47535 , n47528 , n47534 );
not ( n16766 , n29614 );
and ( n16767 , n16766 , RI173dc6f0_1681);
and ( n16768 , n47535 , n29614 );
or ( n47536 , n16767 , n16768 );
not ( n16769 , RI1754c610_2);
and ( n16770 , n16769 , n47536 );
and ( n16771 , C0 , RI1754c610_2);
or ( n47537 , n16770 , n16771 );
buf ( n47538 , n47537 );
buf ( n47539 , RI17491050_1029);
not ( n16772 , n27683 );
and ( n16773 , n16772 , RI19aba578_2378);
and ( n16774 , RI19ac2f48_2307 , n27683 );
or ( n47540 , n16773 , n16774 );
not ( n16775 , RI1754c610_2);
and ( n16776 , n16775 , n47540 );
and ( n16777 , C0 , RI1754c610_2);
or ( n47541 , n16776 , n16777 );
buf ( n47542 , n47541 );
xor ( n47543 , n35207 , n43492 );
xor ( n47544 , n47543 , n38634 );
not ( n47545 , n44845 );
and ( n47546 , n47545 , n44847 );
xor ( n47547 , n47544 , n47546 );
not ( n16778 , n29614 );
and ( n16779 , n16778 , RI173f9f70_1537);
and ( n16780 , n47547 , n29614 );
or ( n47548 , n16779 , n16780 );
not ( n16781 , RI1754c610_2);
and ( n16782 , n16781 , n47548 );
and ( n16783 , C0 , RI1754c610_2);
or ( n47549 , n16782 , n16783 );
buf ( n47550 , n47549 );
xor ( n47551 , n41473 , n39686 );
xor ( n47552 , n47551 , n34087 );
xor ( n47553 , n43491 , n32108 );
xor ( n47554 , n47553 , n38347 );
not ( n47555 , n47554 );
and ( n47556 , n47555 , n40898 );
xor ( n47557 , n47552 , n47556 );
not ( n16784 , n29614 );
and ( n16785 , n16784 , RI173b0218_1897);
and ( n16786 , n47557 , n29614 );
or ( n47558 , n16785 , n16786 );
not ( n16787 , RI1754c610_2);
and ( n16788 , n16787 , n47558 );
and ( n16789 , C0 , RI1754c610_2);
or ( n47559 , n16788 , n16789 );
buf ( n47560 , n47559 );
and ( n47561 , RI1754bc38_23 , n34844 );
and ( n47562 , RI1754bc38_23 , n34847 );
and ( n47563 , RI1754bc38_23 , n34850 );
and ( n47564 , RI1754bc38_23 , n34852 );
and ( n47565 , RI1754bc38_23 , n34854 );
or ( n47566 , n47561 , n47562 , n47563 , n47564 , n47565 , C0 , C0 , C0 );
not ( n16790 , n34859 );
and ( n16791 , n16790 , n47566 );
and ( n16792 , RI1754bc38_23 , n34859 );
or ( n47567 , n16791 , n16792 );
not ( n16793 , RI19a22f70_2797);
and ( n16794 , n16793 , n47567 );
and ( n16795 , C0 , RI19a22f70_2797);
or ( n47568 , n16794 , n16795 );
not ( n16796 , n27683 );
and ( n16797 , n16796 , RI19a9e6c0_2581);
and ( n16798 , n47568 , n27683 );
or ( n47569 , n16797 , n16798 );
not ( n16799 , RI1754c610_2);
and ( n16800 , n16799 , n47569 );
and ( n16801 , C0 , RI1754c610_2);
or ( n47570 , n16800 , n16801 );
buf ( n47571 , n47570 );
xor ( n47572 , n37069 , n38594 );
xor ( n47573 , n47572 , n37716 );
not ( n47574 , n47573 );
xor ( n47575 , n40282 , n37623 );
xor ( n47576 , n47575 , n37651 );
and ( n47577 , n47574 , n47576 );
xor ( n47578 , n44352 , n47577 );
not ( n16802 , n29614 );
and ( n16803 , n16802 , RI173a5e08_1947);
and ( n16804 , n47578 , n29614 );
or ( n47579 , n16803 , n16804 );
not ( n16805 , RI1754c610_2);
and ( n16806 , n16805 , n47579 );
and ( n16807 , C0 , RI1754c610_2);
or ( n47580 , n16806 , n16807 );
buf ( n47581 , n47580 );
not ( n16808 , n27683 );
and ( n16809 , n16808 , RI19a8e8b0_2693);
and ( n16810 , RI19a98ae0_2621 , n27683 );
or ( n47582 , n16809 , n16810 );
not ( n16811 , RI1754c610_2);
and ( n16812 , n16811 , n47582 );
and ( n16813 , C0 , RI1754c610_2);
or ( n47583 , n16812 , n16813 );
buf ( n47584 , n47583 );
xor ( n47585 , n40399 , n32973 );
xor ( n47586 , n47585 , n39816 );
not ( n47587 , n45954 );
and ( n47588 , n47587 , n44971 );
xor ( n47589 , n47586 , n47588 );
not ( n16814 , n29614 );
and ( n16815 , n16814 , RI17475210_1165);
and ( n16816 , n47589 , n29614 );
or ( n47590 , n16815 , n16816 );
not ( n16817 , RI1754c610_2);
and ( n16818 , n16817 , n47590 );
and ( n16819 , C0 , RI1754c610_2);
or ( n47591 , n16818 , n16819 );
buf ( n47592 , n47591 );
not ( n47593 , n46020 );
xor ( n47594 , n34434 , n40009 );
xor ( n47595 , n47594 , n38085 );
and ( n47596 , n47593 , n47595 );
xor ( n47597 , n37210 , n47596 );
not ( n16820 , n29614 );
and ( n16821 , n16820 , RI173d8898_1700);
and ( n16822 , n47597 , n29614 );
or ( n47598 , n16821 , n16822 );
not ( n16823 , RI1754c610_2);
and ( n16824 , n16823 , n47598 );
and ( n16825 , C0 , RI1754c610_2);
or ( n47599 , n16824 , n16825 );
buf ( n47600 , n47599 );
xor ( n47601 , n38861 , n41125 );
xor ( n47602 , n47601 , n31506 );
xor ( n47603 , n40046 , n38574 );
xor ( n47604 , n47603 , n38594 );
not ( n47605 , n47604 );
xor ( n47606 , n39739 , n39506 );
xor ( n47607 , n47606 , n38150 );
and ( n47608 , n47605 , n47607 );
xor ( n47609 , n47602 , n47608 );
not ( n16826 , n29614 );
and ( n16827 , n16826 , RI173ecd70_1601);
and ( n16828 , n47609 , n29614 );
or ( n47610 , n16827 , n16828 );
not ( n16829 , RI1754c610_2);
and ( n16830 , n16829 , n47610 );
and ( n16831 , C0 , RI1754c610_2);
or ( n47611 , n16830 , n16831 );
buf ( n47612 , n47611 );
xor ( n47613 , n42263 , n40743 );
xor ( n47614 , n47613 , n36062 );
not ( n47615 , n46573 );
and ( n47616 , n47615 , n46575 );
xor ( n47617 , n47614 , n47616 );
not ( n16832 , n29614 );
and ( n16833 , n16832 , RI1740cd50_1445);
and ( n16834 , n47617 , n29614 );
or ( n47618 , n16833 , n16834 );
not ( n16835 , RI1754c610_2);
and ( n16836 , n16835 , n47618 );
and ( n16837 , C0 , RI1754c610_2);
or ( n47619 , n16836 , n16837 );
buf ( n47620 , n47619 );
not ( n16838 , n27683 );
and ( n16839 , n16838 , RI19ac1670_2319);
and ( n16840 , RI19acabf8_2250 , n27683 );
or ( n47621 , n16839 , n16840 );
not ( n16841 , RI1754c610_2);
and ( n16842 , n16841 , n47621 );
and ( n16843 , C0 , RI1754c610_2);
or ( n47622 , n16842 , n16843 );
buf ( n47623 , n47622 );
not ( n47624 , n42678 );
and ( n47625 , n47624 , n42680 );
xor ( n47626 , n45572 , n47625 );
not ( n16844 , n29614 );
and ( n16845 , n16844 , RI173dd410_1677);
and ( n16846 , n47626 , n29614 );
or ( n47627 , n16845 , n16846 );
not ( n16847 , RI1754c610_2);
and ( n16848 , n16847 , n47627 );
and ( n16849 , C0 , RI1754c610_2);
or ( n47628 , n16848 , n16849 );
buf ( n47629 , n47628 );
buf ( n47630 , RI17488338_1072);
buf ( n47631 , RI17506188_747);
buf ( n47632 , RI1746e5c8_1198);
xor ( n47633 , n35330 , n41005 );
xor ( n47634 , n47633 , n40585 );
xor ( n47635 , n33210 , n31317 );
xor ( n47636 , n47635 , n40302 );
not ( n47637 , n47636 );
xor ( n47638 , n35617 , n41543 );
xor ( n47639 , n47638 , n34669 );
and ( n47640 , n47637 , n47639 );
xor ( n47641 , n47634 , n47640 );
not ( n16850 , n29614 );
and ( n16851 , n16850 , RI174b9eb0_832);
and ( n16852 , n47641 , n29614 );
or ( n47642 , n16851 , n16852 );
not ( n16853 , RI1754c610_2);
and ( n16854 , n16853 , n47642 );
and ( n16855 , C0 , RI1754c610_2);
or ( n47643 , n16854 , n16855 );
buf ( n47644 , n47643 );
xor ( n47645 , n37065 , n38594 );
xor ( n47646 , n47645 , n37716 );
xor ( n47647 , n38186 , n32220 );
xor ( n47648 , n47647 , n32309 );
not ( n47649 , n47648 );
and ( n47650 , n47649 , n46916 );
xor ( n47651 , n47646 , n47650 );
not ( n16856 , n29614 );
and ( n16857 , n16856 , RI1745f640_1271);
and ( n16858 , n47651 , n29614 );
or ( n47652 , n16857 , n16858 );
not ( n16859 , RI1754c610_2);
and ( n16860 , n16859 , n47652 );
and ( n16861 , C0 , RI1754c610_2);
or ( n47653 , n16860 , n16861 );
buf ( n47654 , n47653 );
buf ( n47655 , RI17473e60_1171);
buf ( n47656 , RI1746be68_1210);
not ( n47657 , n41153 );
xor ( n47658 , n40768 , n33778 );
xor ( n47659 , n47658 , n38793 );
and ( n47660 , n47657 , n47659 );
xor ( n47661 , n41150 , n47660 );
not ( n16862 , n29614 );
and ( n16863 , n16862 , RI17477cb8_1152);
and ( n16864 , n47661 , n29614 );
or ( n47662 , n16863 , n16864 );
not ( n16865 , RI1754c610_2);
and ( n16866 , n16865 , n47662 );
and ( n16867 , C0 , RI1754c610_2);
or ( n47663 , n16866 , n16867 );
buf ( n47664 , n47663 );
not ( n47665 , n39066 );
and ( n47666 , n47665 , n46212 );
xor ( n47667 , n39006 , n47666 );
not ( n16868 , n29614 );
and ( n16869 , n16868 , RI17476f98_1156);
and ( n16870 , n47667 , n29614 );
or ( n47668 , n16869 , n16870 );
not ( n16871 , RI1754c610_2);
and ( n16872 , n16871 , n47668 );
and ( n16873 , C0 , RI1754c610_2);
or ( n47669 , n16872 , n16873 );
buf ( n47670 , n47669 );
not ( n47671 , n44201 );
and ( n47672 , n47671 , n44203 );
xor ( n47673 , n46840 , n47672 );
not ( n16874 , n29614 );
and ( n16875 , n16874 , RI174868f8_1080);
and ( n16876 , n47673 , n29614 );
or ( n47674 , n16875 , n16876 );
not ( n16877 , RI1754c610_2);
and ( n16878 , n16877 , n47674 );
and ( n16879 , C0 , RI1754c610_2);
or ( n47675 , n16878 , n16879 );
buf ( n47676 , n47675 );
not ( n16880 , n27683 );
and ( n16881 , n16880 , RI19a8f210_2689);
and ( n16882 , RI19a991e8_2618 , n27683 );
or ( n47677 , n16881 , n16882 );
not ( n16883 , RI1754c610_2);
and ( n16884 , n16883 , n47677 );
and ( n16885 , C0 , RI1754c610_2);
or ( n47678 , n16884 , n16885 );
buf ( n47679 , n47678 );
not ( n47680 , n35459 );
xor ( n47681 , n35525 , n37460 );
xor ( n47682 , n47681 , n37490 );
and ( n47683 , n47680 , n47682 );
xor ( n47684 , n35418 , n47683 );
not ( n16886 , n29614 );
and ( n16887 , n16886 , RI1749be38_976);
and ( n16888 , n47684 , n29614 );
or ( n47685 , n16887 , n16888 );
not ( n16889 , RI1754c610_2);
and ( n16890 , n16889 , n47685 );
and ( n16891 , C0 , RI1754c610_2);
or ( n47686 , n16890 , n16891 );
buf ( n47687 , n47686 );
buf ( n47688 , RI174abae0_899);
buf ( n47689 , RI174a75f8_920);
not ( n16892 , n27683 );
and ( n16893 , n16892 , RI19a8fd50_2684);
and ( n16894 , RI19a99f80_2612 , n27683 );
or ( n47690 , n16893 , n16894 );
not ( n16895 , RI1754c610_2);
and ( n16896 , n16895 , n47690 );
and ( n16897 , C0 , RI1754c610_2);
or ( n47691 , n16896 , n16897 );
buf ( n47692 , n47691 );
xor ( n47693 , n37017 , n40662 );
xor ( n47694 , n47693 , n39208 );
not ( n47695 , n46978 );
and ( n47696 , n47695 , n46980 );
xor ( n47697 , n47694 , n47696 );
not ( n16898 , n29614 );
and ( n16899 , n16898 , RI174ba900_830);
and ( n16900 , n47697 , n29614 );
or ( n47698 , n16899 , n16900 );
not ( n16901 , RI1754c610_2);
and ( n16902 , n16901 , n47698 );
and ( n16903 , C0 , RI1754c610_2);
or ( n47699 , n16902 , n16903 );
buf ( n47700 , n47699 );
xor ( n47701 , n34181 , n42264 );
xor ( n47702 , n47701 , n41370 );
not ( n47703 , n34518 );
and ( n47704 , n47703 , n34623 );
xor ( n47705 , n47702 , n47704 );
not ( n16904 , n29614 );
and ( n16905 , n16904 , RI173b1c58_1889);
and ( n16906 , n47705 , n29614 );
or ( n47706 , n16905 , n16906 );
not ( n16907 , RI1754c610_2);
and ( n16908 , n16907 , n47706 );
and ( n16909 , C0 , RI1754c610_2);
or ( n47707 , n16908 , n16909 );
buf ( n47708 , n47707 );
not ( n47709 , n39155 );
and ( n47710 , n47709 , n40595 );
xor ( n47711 , n39152 , n47710 );
not ( n16910 , n29614 );
and ( n16911 , n16910 , RI17524b60_652);
and ( n16912 , n47711 , n29614 );
or ( n47712 , n16911 , n16912 );
not ( n16913 , RI1754c610_2);
and ( n16914 , n16913 , n47712 );
and ( n16915 , C0 , RI1754c610_2);
or ( n47713 , n16914 , n16915 );
buf ( n47714 , n47713 );
xor ( n47715 , n37306 , n40190 );
xor ( n47716 , n47715 , n40210 );
not ( n47717 , n44570 );
and ( n47718 , n47717 , n44572 );
xor ( n47719 , n47716 , n47718 );
not ( n16916 , n29614 );
and ( n16917 , n16916 , RI1752a308_635);
and ( n16918 , n47719 , n29614 );
or ( n47720 , n16917 , n16918 );
not ( n16919 , RI1754c610_2);
and ( n16920 , n16919 , n47720 );
and ( n16921 , C0 , RI1754c610_2);
or ( n47721 , n16920 , n16921 );
buf ( n47722 , n47721 );
not ( n47723 , n45217 );
and ( n47724 , n47723 , n39093 );
xor ( n47725 , n45214 , n47724 );
not ( n16922 , n29614 );
and ( n16923 , n16922 , RI17398f50_2010);
and ( n16924 , n47725 , n29614 );
or ( n47726 , n16923 , n16924 );
not ( n16925 , RI1754c610_2);
and ( n16926 , n16925 , n47726 );
and ( n16927 , C0 , RI1754c610_2);
or ( n47727 , n16926 , n16927 );
buf ( n47728 , n47727 );
not ( n47729 , n39420 );
xor ( n47730 , n40687 , n36654 );
xor ( n47731 , n47730 , n40808 );
and ( n47732 , n47729 , n47731 );
xor ( n47733 , n39417 , n47732 );
not ( n16928 , n29614 );
and ( n16929 , n16928 , RI1747aaa8_1138);
and ( n16930 , n47733 , n29614 );
or ( n47734 , n16929 , n16930 );
not ( n16931 , RI1754c610_2);
and ( n16932 , n16931 , n47734 );
and ( n16933 , C0 , RI1754c610_2);
or ( n47735 , n16932 , n16933 );
buf ( n47736 , n47735 );
not ( n47737 , n46396 );
and ( n47738 , n47737 , n47126 );
xor ( n47739 , n46393 , n47738 );
not ( n16934 , n29614 );
and ( n16935 , n16934 , RI1752f588_619);
and ( n16936 , n47739 , n29614 );
or ( n47740 , n16935 , n16936 );
not ( n16937 , RI1754c610_2);
and ( n16938 , n16937 , n47740 );
and ( n16939 , C0 , RI1754c610_2);
or ( n47741 , n16938 , n16939 );
buf ( n47742 , n47741 );
xor ( n47743 , n39203 , n37676 );
xor ( n47744 , n47743 , n37696 );
not ( n47745 , n45108 );
and ( n47746 , n47745 , n45110 );
xor ( n47747 , n47744 , n47746 );
not ( n16940 , n29614 );
and ( n16941 , n16940 , RI173a4da0_1952);
and ( n16942 , n47747 , n29614 );
or ( n47748 , n16941 , n16942 );
not ( n16943 , RI1754c610_2);
and ( n16944 , n16943 , n47748 );
and ( n16945 , C0 , RI1754c610_2);
or ( n47749 , n16944 , n16945 );
buf ( n47750 , n47749 );
not ( n16946 , RI1754c610_2);
and ( n16947 , n16946 , RI17536770_597);
and ( n16948 , C0 , RI1754c610_2);
or ( n47751 , n16947 , n16948 );
buf ( n47752 , n47751 );
not ( n16949 , n27683 );
and ( n16950 , n16949 , RI19abc378_2366);
and ( n16951 , RI19ac4910_2295 , n27683 );
or ( n47753 , n16950 , n16951 );
not ( n16952 , RI1754c610_2);
and ( n16953 , n16952 , n47753 );
and ( n16954 , C0 , RI1754c610_2);
or ( n47754 , n16953 , n16954 );
buf ( n47755 , n47754 );
not ( n16955 , n27683 );
and ( n16956 , n16955 , RI19ab0e10_2447);
and ( n16957 , RI19abaa28_2376 , n27683 );
or ( n47756 , n16956 , n16957 );
not ( n16958 , RI1754c610_2);
and ( n16959 , n16958 , n47756 );
and ( n16960 , C0 , RI1754c610_2);
or ( n47757 , n16959 , n16960 );
buf ( n47758 , n47757 );
not ( n47759 , n45284 );
xor ( n47760 , n39922 , n40890 );
xor ( n47761 , n47760 , n38724 );
and ( n47762 , n47759 , n47761 );
xor ( n47763 , n45281 , n47762 );
not ( n16961 , n29614 );
and ( n16962 , n16961 , RI173d01f8_1741);
and ( n16963 , n47763 , n29614 );
or ( n47764 , n16962 , n16963 );
not ( n16964 , RI1754c610_2);
and ( n16965 , n16964 , n47764 );
and ( n16966 , C0 , RI1754c610_2);
or ( n47765 , n16965 , n16966 );
buf ( n47766 , n47765 );
xor ( n47767 , n37451 , n36874 );
xor ( n47768 , n47767 , n42188 );
not ( n47769 , n47768 );
xor ( n47770 , n41813 , n39262 );
xor ( n47771 , n47770 , n39282 );
and ( n47772 , n47769 , n47771 );
xor ( n47773 , n43285 , n47772 );
not ( n16967 , n29614 );
and ( n16968 , n16967 , RI174c8190_788);
and ( n16969 , n47773 , n29614 );
or ( n47774 , n16968 , n16969 );
not ( n16970 , RI1754c610_2);
and ( n16971 , n16970 , n47774 );
and ( n16972 , C0 , RI1754c610_2);
or ( n47775 , n16971 , n16972 );
buf ( n47776 , n47775 );
xor ( n47777 , n34214 , n36287 );
xor ( n47778 , n47777 , n37526 );
xor ( n47779 , n34967 , n36802 );
xor ( n47780 , n47779 , n33125 );
not ( n47781 , n47780 );
xor ( n47782 , n37315 , n39914 );
xor ( n47783 , n47782 , n40237 );
and ( n47784 , n47781 , n47783 );
xor ( n47785 , n47778 , n47784 );
not ( n16973 , n29614 );
and ( n16974 , n16973 , RI1748ffe8_1034);
and ( n16975 , n47785 , n29614 );
or ( n47786 , n16974 , n16975 );
not ( n16976 , RI1754c610_2);
and ( n16977 , n16976 , n47786 );
and ( n16978 , C0 , RI1754c610_2);
or ( n47787 , n16977 , n16978 );
buf ( n47788 , n47787 );
not ( n16979 , n27683 );
and ( n16980 , n16979 , RI19ab96f0_2385);
and ( n16981 , RI19ac21b0_2313 , n27683 );
or ( n47789 , n16980 , n16981 );
not ( n16982 , RI1754c610_2);
and ( n16983 , n16982 , n47789 );
and ( n16984 , C0 , RI1754c610_2);
or ( n47790 , n16983 , n16984 );
buf ( n47791 , n47790 );
buf ( n47792 , RI17486268_1082);
buf ( n47793 , RI1747d550_1125);
buf ( n47794 , RI174665d0_1237);
buf ( n47795 , RI17509518_737);
not ( n47796 , n42950 );
and ( n47797 , n47796 , n47420 );
xor ( n47798 , n42947 , n47797 );
not ( n16985 , n29614 );
and ( n16986 , n16985 , RI17400870_1505);
and ( n16987 , n47798 , n29614 );
or ( n47799 , n16986 , n16987 );
not ( n16988 , RI1754c610_2);
and ( n16989 , n16988 , n47799 );
and ( n16990 , C0 , RI1754c610_2);
or ( n47800 , n16989 , n16990 );
buf ( n47801 , n47800 );
not ( n16991 , n27683 );
and ( n16992 , n16991 , RI19acdf10_2225);
and ( n16993 , RI19a93518_2659 , n27683 );
or ( n47802 , n16992 , n16993 );
not ( n16994 , RI1754c610_2);
and ( n16995 , n16994 , n47802 );
and ( n16996 , C0 , RI1754c610_2);
or ( n47803 , n16995 , n16996 );
buf ( n47804 , n47803 );
buf ( n47805 , RI174c1020_810);
buf ( n47806 , RI174b4e88_854);
buf ( n47807 , RI1749df08_966);
not ( n47808 , n42579 );
and ( n47809 , n47808 , n42885 );
xor ( n47810 , n42576 , n47809 );
not ( n16997 , n29614 );
and ( n16998 , n16997 , RI173dacb0_1689);
and ( n16999 , n47810 , n29614 );
or ( n47811 , n16998 , n16999 );
not ( n17000 , RI1754c610_2);
and ( n17001 , n17000 , n47811 );
and ( n17002 , C0 , RI1754c610_2);
or ( n47812 , n17001 , n17002 );
buf ( n47813 , n47812 );
not ( n47814 , n45113 );
xor ( n47815 , n35340 , n41005 );
xor ( n47816 , n47815 , n40585 );
and ( n47817 , n47814 , n47816 );
xor ( n47818 , n45110 , n47817 );
not ( n17003 , n29614 );
and ( n17004 , n17003 , RI17448030_1385);
and ( n17005 , n47818 , n29614 );
or ( n47819 , n17004 , n17005 );
not ( n17006 , RI1754c610_2);
and ( n17007 , n17006 , n47819 );
and ( n17008 , C0 , RI1754c610_2);
or ( n47820 , n17007 , n17008 );
buf ( n47821 , n47820 );
buf ( n47822 , RI174951f0_1009);
xor ( n47823 , n34283 , n38886 );
xor ( n47824 , n47823 , n39604 );
xor ( n47825 , n39947 , n38724 );
xor ( n47826 , n47825 , n29425 );
not ( n47827 , n47826 );
xor ( n47828 , n38283 , n36568 );
xor ( n47829 , n47828 , n36742 );
and ( n47830 , n47827 , n47829 );
xor ( n47831 , n47824 , n47830 );
not ( n17009 , n29614 );
and ( n17010 , n17009 , RI1745e290_1277);
and ( n17011 , n47831 , n29614 );
or ( n47832 , n17010 , n17011 );
not ( n17012 , RI1754c610_2);
and ( n17013 , n17012 , n47832 );
and ( n17014 , C0 , RI1754c610_2);
or ( n47833 , n17013 , n17014 );
buf ( n47834 , n47833 );
not ( n17015 , n27683 );
and ( n17016 , n17015 , RI19ab03c0_2452);
and ( n17017 , RI19aba050_2380 , n27683 );
or ( n47835 , n17016 , n17017 );
not ( n17018 , RI1754c610_2);
and ( n17019 , n17018 , n47835 );
and ( n17020 , C0 , RI1754c610_2);
or ( n47836 , n17019 , n17020 );
buf ( n47837 , n47836 );
xor ( n47838 , n39498 , n30923 );
xor ( n47839 , n47838 , n31053 );
not ( n47840 , n38678 );
and ( n47841 , n47840 , n38683 );
xor ( n47842 , n47839 , n47841 );
not ( n17021 , n29614 );
and ( n17022 , n17021 , RI1748be48_1054);
and ( n17023 , n47842 , n29614 );
or ( n47843 , n17022 , n17023 );
not ( n17024 , RI1754c610_2);
and ( n17025 , n17024 , n47843 );
and ( n17026 , C0 , RI1754c610_2);
or ( n47844 , n17025 , n17026 );
buf ( n47845 , n47844 );
not ( n17027 , n27683 );
and ( n17028 , n17027 , RI19ac5720_2288);
and ( n17029 , RI19ace3c0_2223 , n27683 );
or ( n47846 , n17028 , n17029 );
not ( n17030 , RI1754c610_2);
and ( n17031 , n17030 , n47846 );
and ( n17032 , C0 , RI1754c610_2);
or ( n47847 , n17031 , n17032 );
buf ( n47848 , n47847 );
xor ( n47849 , n37433 , n34725 );
xor ( n47850 , n47849 , n34755 );
xor ( n47851 , n41477 , n39686 );
xor ( n47852 , n47851 , n34087 );
not ( n47853 , n47852 );
xor ( n47854 , n40227 , n35710 );
xor ( n47855 , n47854 , n35760 );
and ( n47856 , n47853 , n47855 );
xor ( n47857 , n47850 , n47856 );
not ( n17033 , n29614 );
and ( n17034 , n17033 , RI173aacc8_1923);
and ( n17035 , n47857 , n29614 );
or ( n47858 , n17034 , n17035 );
not ( n17036 , RI1754c610_2);
and ( n17037 , n17036 , n47858 );
and ( n17038 , C0 , RI1754c610_2);
or ( n47859 , n17037 , n17038 );
buf ( n47860 , n47859 );
not ( n17039 , n27683 );
and ( n17040 , n17039 , RI19ac89c0_2265);
and ( n17041 , RI19a838e8_2769 , n27683 );
or ( n47861 , n17040 , n17041 );
not ( n17042 , RI1754c610_2);
and ( n17043 , n17042 , n47861 );
and ( n17044 , C0 , RI1754c610_2);
or ( n47862 , n17043 , n17044 );
buf ( n47863 , n47862 );
not ( n47864 , n34838 );
xor ( n47865 , n40403 , n32973 );
xor ( n47866 , n47865 , n39816 );
and ( n47867 , n47864 , n47866 );
xor ( n47868 , n34756 , n47867 );
not ( n17045 , n29614 );
and ( n17046 , n17045 , RI173d22e0_1731);
and ( n17047 , n47868 , n29614 );
or ( n47869 , n17046 , n17047 );
not ( n17048 , RI1754c610_2);
and ( n17049 , n17048 , n47869 );
and ( n17050 , C0 , RI1754c610_2);
or ( n47870 , n17049 , n17050 );
buf ( n47871 , n47870 );
xor ( n47872 , n39341 , n29843 );
xor ( n47873 , n47872 , n29981 );
not ( n47874 , n47873 );
and ( n47875 , n47874 , n42655 );
xor ( n47876 , n40517 , n47875 );
not ( n17051 , n29614 );
and ( n17052 , n17051 , RI173d5418_1716);
and ( n17053 , n47876 , n29614 );
or ( n47877 , n17052 , n17053 );
not ( n17054 , RI1754c610_2);
and ( n17055 , n17054 , n47877 );
and ( n17056 , C0 , RI1754c610_2);
or ( n47878 , n17055 , n17056 );
buf ( n47879 , n47878 );
not ( n47880 , n42206 );
and ( n47881 , n47880 , n47109 );
xor ( n47882 , n42203 , n47881 );
not ( n17057 , n29614 );
and ( n17058 , n17057 , RI174b3448_862);
and ( n17059 , n47882 , n29614 );
or ( n47883 , n17058 , n17059 );
not ( n17060 , RI1754c610_2);
and ( n17061 , n17060 , n47883 );
and ( n17062 , C0 , RI1754c610_2);
or ( n47884 , n17061 , n17062 );
buf ( n47885 , n47884 );
not ( n47886 , n45927 );
xor ( n47887 , n37789 , n43994 );
xor ( n47888 , n47887 , n31213 );
and ( n47889 , n47886 , n47888 );
xor ( n47890 , n45924 , n47889 );
not ( n17063 , n29614 );
and ( n17064 , n17063 , RI174c1548_809);
and ( n17065 , n47890 , n29614 );
or ( n47891 , n17064 , n17065 );
not ( n17066 , RI1754c610_2);
and ( n17067 , n17066 , n47891 );
and ( n17068 , C0 , RI1754c610_2);
or ( n47892 , n17067 , n17068 );
buf ( n47893 , n47892 );
buf ( n47894 , RI175110d8_713);
not ( n17069 , n27683 );
and ( n17070 , n17069 , RI19a92708_2665);
and ( n17071 , RI19a9c848_2594 , n27683 );
or ( n47895 , n17070 , n17071 );
not ( n17072 , RI1754c610_2);
and ( n17073 , n17072 , n47895 );
and ( n17074 , C0 , RI1754c610_2);
or ( n47896 , n17073 , n17074 );
buf ( n47897 , n47896 );
buf ( n47898 , RI174813a8_1106);
not ( n47899 , n46153 );
and ( n47900 , n47899 , n46155 );
xor ( n47901 , n45519 , n47900 );
not ( n17075 , n29614 );
and ( n17076 , n17075 , RI173d95b8_1696);
and ( n17077 , n47901 , n29614 );
or ( n47902 , n17076 , n17077 );
not ( n17078 , RI1754c610_2);
and ( n17079 , n17078 , n47902 );
and ( n17080 , C0 , RI1754c610_2);
or ( n47903 , n17079 , n17080 );
buf ( n47904 , n47903 );
xor ( n47905 , n31804 , n34644 );
xor ( n47906 , n47905 , n36401 );
xor ( n47907 , n41365 , n36062 );
xor ( n47908 , n47907 , n36102 );
not ( n47909 , n47908 );
and ( n47910 , n47909 , n47019 );
xor ( n47911 , n47906 , n47910 );
not ( n17081 , n29614 );
and ( n17082 , n17081 , RI1745cb98_1284);
and ( n17083 , n47911 , n29614 );
or ( n47912 , n17082 , n17083 );
not ( n17084 , RI1754c610_2);
and ( n17085 , n17084 , n47912 );
and ( n17086 , C0 , RI1754c610_2);
or ( n47913 , n17085 , n17086 );
buf ( n47914 , n47913 );
not ( n17087 , n27683 );
and ( n17088 , n17087 , RI19a86318_2751);
and ( n17089 , RI19a23c18_2790 , n27683 );
or ( n47915 , n17088 , n17089 );
not ( n17090 , RI1754c610_2);
and ( n17091 , n17090 , n47915 );
and ( n17092 , C0 , RI1754c610_2);
or ( n47916 , n17091 , n17092 );
buf ( n47917 , n47916 );
not ( n17093 , n27683 );
and ( n17094 , n17093 , RI19a94238_2653);
and ( n17095 , RI19a9e468_2582 , n27683 );
or ( n47918 , n17094 , n17095 );
not ( n17096 , RI1754c610_2);
and ( n17097 , n17096 , n47918 );
and ( n17098 , C0 , RI1754c610_2);
or ( n47919 , n17097 , n17098 );
buf ( n47920 , n47919 );
not ( n17099 , n27683 );
and ( n17100 , n17099 , RI19aab5f0_2486);
and ( n17101 , RI19ab52f8_2415 , n27683 );
or ( n47921 , n17100 , n17101 );
not ( n17102 , RI1754c610_2);
and ( n17103 , n17102 , n47921 );
and ( n17104 , C0 , RI1754c610_2);
or ( n47922 , n17103 , n17104 );
buf ( n47923 , n47922 );
not ( n47924 , n40517 );
and ( n47925 , n47924 , n47873 );
xor ( n47926 , n40466 , n47925 );
not ( n17105 , n29614 );
and ( n17106 , n17105 , RI173c67c0_1788);
and ( n17107 , n47926 , n29614 );
or ( n47927 , n17106 , n17107 );
not ( n17108 , RI1754c610_2);
and ( n17109 , n17108 , n47927 );
and ( n17110 , C0 , RI1754c610_2);
or ( n47928 , n17109 , n17110 );
buf ( n47929 , n47928 );
not ( n17111 , n27683 );
and ( n17112 , n17111 , RI19a8a530_2722);
and ( n17113 , RI19a94490_2652 , n27683 );
or ( n47930 , n17112 , n17113 );
not ( n17114 , RI1754c610_2);
and ( n17115 , n17114 , n47930 );
and ( n17116 , C0 , RI1754c610_2);
or ( n47931 , n17115 , n17116 );
buf ( n47932 , n47931 );
and ( n47933 , RI19a24320_2787 , n43086 );
not ( n17117 , n43088 );
and ( n17118 , n17117 , RI19a240c8_2788);
and ( n17119 , n47933 , n43088 );
or ( n47934 , n17118 , n17119 );
not ( n17120 , RI1754c610_2);
and ( n17121 , n17120 , n47934 );
and ( n17122 , C0 , RI1754c610_2);
or ( n47935 , n17121 , n17122 );
buf ( n47936 , n47935 );
buf ( n47937 , RI17489a30_1065);
buf ( n47938 , RI175019d0_755);
buf ( n47939 , RI174ab450_901);
buf ( n47940 , RI1748e260_1043);
not ( n47941 , n40726 );
and ( n47942 , n47941 , n40744 );
xor ( n47943 , n44516 , n47942 );
not ( n17123 , n29614 );
and ( n17124 , n17123 , RI1749d1e8_970);
and ( n17125 , n47943 , n29614 );
or ( n47944 , n17124 , n17125 );
not ( n17126 , RI1754c610_2);
and ( n17127 , n17126 , n47944 );
and ( n17128 , C0 , RI1754c610_2);
or ( n47945 , n17127 , n17128 );
buf ( n47946 , n47945 );
xor ( n47947 , n39173 , n40166 );
xor ( n47948 , n47947 , n41590 );
not ( n47949 , n45483 );
and ( n47950 , n47949 , n45485 );
xor ( n47951 , n47948 , n47950 );
not ( n17129 , n29614 );
and ( n17130 , n17129 , RI173a4a58_1953);
and ( n17131 , n47951 , n29614 );
or ( n47952 , n17130 , n17131 );
not ( n17132 , RI1754c610_2);
and ( n17133 , n17132 , n47952 );
and ( n17134 , C0 , RI1754c610_2);
or ( n47953 , n17133 , n17134 );
buf ( n47954 , n47953 );
not ( n17135 , n27683 );
and ( n17136 , n17135 , RI19aa4a98_2532);
and ( n17137 , RI19aaeea8_2462 , n27683 );
or ( n47955 , n17136 , n17137 );
not ( n17138 , RI1754c610_2);
and ( n17139 , n17138 , n47955 );
and ( n17140 , C0 , RI1754c610_2);
or ( n47956 , n17139 , n17140 );
buf ( n47957 , n47956 );
xor ( n47958 , n41533 , n32786 );
xor ( n47959 , n47958 , n32863 );
xor ( n47960 , n41981 , n39886 );
xor ( n47961 , n47960 , n36998 );
not ( n47962 , n47961 );
and ( n47963 , n47962 , n39792 );
xor ( n47964 , n47959 , n47963 );
not ( n17141 , n29614 );
and ( n17142 , n17141 , RI173d67c8_1710);
and ( n17143 , n47964 , n29614 );
or ( n47965 , n17142 , n17143 );
not ( n17144 , RI1754c610_2);
and ( n17145 , n17144 , n47965 );
and ( n17146 , C0 , RI1754c610_2);
or ( n47966 , n17145 , n17146 );
buf ( n47967 , n47966 );
and ( n47968 , RI1754c070_14 , n34844 );
and ( n47969 , RI1754c070_14 , n34847 );
and ( n47970 , RI1754c070_14 , n34850 );
and ( n47971 , RI1754c070_14 , n34852 );
and ( n47972 , RI1754c070_14 , n34854 );
and ( n47973 , RI1754c070_14 , n34856 );
or ( n47974 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , C0 , C0 );
not ( n17147 , n34859 );
and ( n17148 , n17147 , n47974 );
and ( n17149 , RI1754c070_14 , n34859 );
or ( n47975 , n17148 , n17149 );
not ( n17150 , RI19a22f70_2797);
and ( n17151 , n17150 , n47975 );
and ( n17152 , C0 , RI19a22f70_2797);
or ( n47976 , n17151 , n17152 );
not ( n17153 , n27683 );
and ( n17154 , n17153 , RI19a90368_2681);
and ( n17155 , n47976 , n27683 );
or ( n47977 , n17154 , n17155 );
not ( n17156 , RI1754c610_2);
and ( n17157 , n17156 , n47977 );
and ( n17158 , C0 , RI1754c610_2);
or ( n47978 , n17157 , n17158 );
buf ( n47979 , n47978 );
not ( n17159 , n27683 );
and ( n17160 , n17159 , RI19acb4e0_2245);
and ( n17161 , RI19a86c00_2747 , n27683 );
or ( n47980 , n17160 , n17161 );
not ( n17162 , RI1754c610_2);
and ( n17163 , n17162 , n47980 );
and ( n17164 , C0 , RI1754c610_2);
or ( n47981 , n17163 , n17164 );
buf ( n47982 , n47981 );
xor ( n47983 , n36610 , n39791 );
xor ( n47984 , n47983 , n40915 );
xor ( n47985 , n38385 , n37169 );
xor ( n47986 , n47985 , n36339 );
not ( n47987 , n47986 );
xor ( n47988 , n34315 , n39604 );
xor ( n47989 , n47988 , n39621 );
and ( n47990 , n47987 , n47989 );
xor ( n47991 , n47984 , n47990 );
not ( n17165 , n29614 );
and ( n17166 , n17165 , RI1749ef70_961);
and ( n17167 , n47991 , n29614 );
or ( n47992 , n17166 , n17167 );
not ( n17168 , RI1754c610_2);
and ( n17169 , n17168 , n47992 );
and ( n17170 , C0 , RI1754c610_2);
or ( n47993 , n17169 , n17170 );
buf ( n47994 , n47993 );
not ( n17171 , n27683 );
and ( n17172 , n17171 , RI19a98630_2623);
and ( n17173 , RI19aa1f00_2553 , n27683 );
or ( n47995 , n17172 , n17173 );
not ( n17174 , RI1754c610_2);
and ( n17175 , n17174 , n47995 );
and ( n17176 , C0 , RI1754c610_2);
or ( n47996 , n17175 , n17176 );
buf ( n47997 , n47996 );
not ( n47998 , n38190 );
and ( n47999 , n47998 , n45498 );
xor ( n48000 , n38168 , n47999 );
not ( n17177 , n29614 );
and ( n17178 , n17177 , RI174a9d58_908);
and ( n17179 , n48000 , n29614 );
or ( n48001 , n17178 , n17179 );
not ( n17180 , RI1754c610_2);
and ( n17181 , n17180 , n48001 );
and ( n17182 , C0 , RI1754c610_2);
or ( n48002 , n17181 , n17182 );
buf ( n48003 , n48002 );
not ( n48004 , n41345 );
xor ( n48005 , n33566 , n40915 );
xor ( n48006 , n48005 , n41740 );
and ( n48007 , n48004 , n48006 );
xor ( n48008 , n41339 , n48007 );
not ( n17183 , n29614 );
and ( n17184 , n17183 , RI17460360_1267);
and ( n17185 , n48008 , n29614 );
or ( n48009 , n17184 , n17185 );
not ( n17186 , RI1754c610_2);
and ( n17187 , n17186 , n48009 );
and ( n17188 , C0 , RI1754c610_2);
or ( n48010 , n17187 , n17188 );
buf ( n48011 , n48010 );
xor ( n48012 , n36529 , n40381 );
xor ( n48013 , n48012 , n37438 );
not ( n48014 , n48013 );
and ( n48015 , n48014 , n42133 );
xor ( n48016 , n45819 , n48015 );
not ( n17189 , n29614 );
and ( n17190 , n17189 , RI173f7180_1551);
and ( n17191 , n48016 , n29614 );
or ( n48017 , n17190 , n17191 );
not ( n17192 , RI1754c610_2);
and ( n17193 , n17192 , n48017 );
and ( n17194 , C0 , RI1754c610_2);
or ( n48018 , n17193 , n17194 );
buf ( n48019 , n48018 );
not ( n17195 , n27683 );
and ( n17196 , n17195 , RI19a98018_2626);
and ( n17197 , RI19aa19d8_2555 , n27683 );
or ( n48020 , n17196 , n17197 );
not ( n17198 , RI1754c610_2);
and ( n17199 , n17198 , n48020 );
and ( n17200 , C0 , RI1754c610_2);
or ( n48021 , n17199 , n17200 );
buf ( n48022 , n48021 );
xor ( n48023 , n40492 , n41430 );
xor ( n48024 , n48023 , n36844 );
xor ( n48025 , n32433 , n35622 );
xor ( n48026 , n48025 , n35639 );
not ( n48027 , n48026 );
xor ( n48028 , n40683 , n36654 );
xor ( n48029 , n48028 , n40808 );
and ( n48030 , n48027 , n48029 );
xor ( n48031 , n48024 , n48030 );
not ( n17201 , n29614 );
and ( n17202 , n17201 , RI17345580_2103);
and ( n17203 , n48031 , n29614 );
or ( n48032 , n17202 , n17203 );
not ( n17204 , RI1754c610_2);
and ( n17205 , n17204 , n48032 );
and ( n17206 , C0 , RI1754c610_2);
or ( n48033 , n17205 , n17206 );
buf ( n48034 , n48033 );
not ( n17207 , n27683 );
and ( n17208 , n17207 , RI19ab0ff0_2446);
and ( n17209 , RI19abad70_2375 , n27683 );
or ( n48035 , n17208 , n17209 );
not ( n17210 , RI1754c610_2);
and ( n17211 , n17210 , n48035 );
and ( n17212 , C0 , RI1754c610_2);
or ( n48036 , n17211 , n17212 );
buf ( n48037 , n48036 );
xor ( n48038 , n39810 , n37800 );
xor ( n48039 , n48038 , n37814 );
not ( n48040 , n48039 );
and ( n48041 , n48040 , n44747 );
xor ( n48042 , n44618 , n48041 );
not ( n17213 , n29614 );
and ( n17214 , n17213 , RI17475be8_1162);
and ( n17215 , n48042 , n29614 );
or ( n48043 , n17214 , n17215 );
not ( n17216 , RI1754c610_2);
and ( n17217 , n17216 , n48043 );
and ( n17218 , C0 , RI1754c610_2);
or ( n48044 , n17217 , n17218 );
buf ( n48045 , n48044 );
not ( n48046 , n43950 );
xor ( n48047 , n40712 , n39333 );
xor ( n48048 , n48047 , n39347 );
and ( n48049 , n48046 , n48048 );
xor ( n48050 , n43947 , n48049 );
not ( n17219 , n29614 );
and ( n17220 , n17219 , RI174ad1d8_892);
and ( n17221 , n48050 , n29614 );
or ( n48051 , n17220 , n17221 );
not ( n17222 , RI1754c610_2);
and ( n17223 , n17222 , n48051 );
and ( n17224 , C0 , RI1754c610_2);
or ( n48052 , n17223 , n17224 );
buf ( n48053 , n48052 );
not ( n48054 , n46831 );
xor ( n48055 , n36801 , n38214 );
xor ( n48056 , n48055 , n38244 );
and ( n48057 , n48054 , n48056 );
xor ( n48058 , n46828 , n48057 );
not ( n17225 , n29614 );
and ( n17226 , n17225 , RI173ea2c8_1614);
and ( n17227 , n48058 , n29614 );
or ( n48059 , n17226 , n17227 );
not ( n17228 , RI1754c610_2);
and ( n17229 , n17228 , n48059 );
and ( n17230 , C0 , RI1754c610_2);
or ( n48060 , n17229 , n17230 );
buf ( n48061 , n48060 );
and ( n48062 , RI1754b3c8_41 , n34844 );
and ( n48063 , RI1754b3c8_41 , n34847 );
and ( n48064 , RI1754b3c8_41 , n34850 );
or ( n48065 , n48062 , n48063 , n48064 , C0 , C0 , C0 , C0 , C0 );
not ( n17231 , n34859 );
and ( n17232 , n17231 , n48065 );
and ( n17233 , RI1754b3c8_41 , n34859 );
or ( n48066 , n17232 , n17233 );
not ( n17234 , RI19a22f70_2797);
and ( n17235 , n17234 , n48066 );
and ( n17236 , C0 , RI19a22f70_2797);
or ( n48067 , n17235 , n17236 );
not ( n17237 , n27683 );
and ( n17238 , n17237 , RI19ab9df8_2381);
and ( n17239 , n48067 , n27683 );
or ( n48068 , n17238 , n17239 );
not ( n17240 , RI1754c610_2);
and ( n17241 , n17240 , n48068 );
and ( n17242 , C0 , RI1754c610_2);
or ( n48069 , n17241 , n17242 );
buf ( n48070 , n48069 );
not ( n48071 , n42058 );
and ( n48072 , n48071 , n41126 );
xor ( n48073 , n43228 , n48072 );
not ( n17243 , n29614 );
and ( n17244 , n17243 , RI17487ff0_1073);
and ( n17245 , n48073 , n29614 );
or ( n48074 , n17244 , n17245 );
not ( n17246 , RI1754c610_2);
and ( n17247 , n17246 , n48074 );
and ( n17248 , C0 , RI1754c610_2);
or ( n48075 , n17247 , n17248 );
buf ( n48076 , n48075 );
buf ( n48077 , RI174c29e8_805);
not ( n48078 , n46791 );
and ( n48079 , n48078 , n46934 );
xor ( n48080 , n39348 , n48079 );
not ( n17249 , n29614 );
and ( n17250 , n17249 , RI173c46f0_1798);
and ( n17251 , n48080 , n29614 );
or ( n48081 , n17250 , n17251 );
not ( n17252 , RI1754c610_2);
and ( n17253 , n17252 , n48081 );
and ( n17254 , C0 , RI1754c610_2);
or ( n48082 , n17253 , n17254 );
buf ( n48083 , n48082 );
not ( n48084 , n47160 );
and ( n48085 , n48084 , n43035 );
xor ( n48086 , n47157 , n48085 );
not ( n17255 , n29614 );
and ( n17256 , n17255 , RI17411c10_1421);
and ( n17257 , n48086 , n29614 );
or ( n48087 , n17256 , n17257 );
not ( n17258 , RI1754c610_2);
and ( n17259 , n17258 , n48087 );
and ( n17260 , C0 , RI1754c610_2);
or ( n48088 , n17259 , n17260 );
buf ( n48089 , n48088 );
buf ( n48090 , RI174944d0_1013);
xor ( n48091 , n30584 , n38167 );
xor ( n48092 , n48091 , n33728 );
not ( n48093 , n48092 );
and ( n48094 , n48093 , n37351 );
xor ( n48095 , n43888 , n48094 );
not ( n17261 , n29614 );
and ( n17262 , n17261 , RI173e81f8_1624);
and ( n17263 , n48095 , n29614 );
or ( n48096 , n17262 , n17263 );
not ( n17264 , RI1754c610_2);
and ( n17265 , n17264 , n48096 );
and ( n17266 , C0 , RI1754c610_2);
or ( n48097 , n17265 , n17266 );
buf ( n48098 , n48097 );
not ( n48099 , n45164 );
and ( n48100 , n48099 , n44963 );
xor ( n48101 , n38838 , n48100 );
not ( n17267 , n29614 );
and ( n17268 , n17267 , RI174713b8_1184);
and ( n17269 , n48101 , n29614 );
or ( n48102 , n17268 , n17269 );
not ( n17270 , RI1754c610_2);
and ( n17271 , n17270 , n48102 );
and ( n17272 , C0 , RI1754c610_2);
or ( n48103 , n17271 , n17272 );
buf ( n48104 , n48103 );
not ( n17273 , n27683 );
and ( n17274 , n17273 , RI19abeda8_2342);
and ( n17275 , RI19ac7d90_2271 , n27683 );
or ( n48105 , n17274 , n17275 );
not ( n17276 , RI1754c610_2);
and ( n17277 , n17276 , n48105 );
and ( n17278 , C0 , RI1754c610_2);
or ( n48106 , n17277 , n17278 );
buf ( n48107 , n48106 );
not ( n17279 , n27683 );
and ( n17280 , n17279 , RI19a99d28_2613);
and ( n17281 , RI19aa3418_2543 , n27683 );
or ( n48108 , n17280 , n17281 );
not ( n17282 , RI1754c610_2);
and ( n17283 , n17282 , n48108 );
and ( n17284 , C0 , RI1754c610_2);
or ( n48109 , n17283 , n17284 );
buf ( n48110 , n48109 );
xor ( n48111 , n36456 , n37104 );
xor ( n48112 , n48111 , n35986 );
xor ( n48113 , n31663 , n30604 );
xor ( n48114 , n48113 , n30741 );
not ( n48115 , n48114 );
xor ( n48116 , n41577 , n39065 );
xor ( n48117 , n48116 , n37331 );
and ( n48118 , n48115 , n48117 );
xor ( n48119 , n48112 , n48118 );
not ( n17285 , n29614 );
and ( n17286 , n17285 , RI173fc040_1527);
and ( n17287 , n48119 , n29614 );
or ( n48120 , n17286 , n17287 );
not ( n17288 , RI1754c610_2);
and ( n17289 , n17288 , n48120 );
and ( n17290 , C0 , RI1754c610_2);
or ( n48121 , n17289 , n17290 );
buf ( n48122 , n48121 );
not ( n48123 , n45473 );
and ( n48124 , n48123 , n45475 );
xor ( n48125 , n42449 , n48124 );
not ( n17291 , n29614 );
and ( n17292 , n17291 , RI17473b18_1172);
and ( n17293 , n48125 , n29614 );
or ( n48126 , n17292 , n17293 );
not ( n17294 , RI1754c610_2);
and ( n17295 , n17294 , n48126 );
and ( n17296 , C0 , RI1754c610_2);
or ( n48127 , n17295 , n17296 );
buf ( n48128 , n48127 );
not ( n48129 , n44850 );
xor ( n48130 , n33054 , n36227 );
xor ( n48131 , n48130 , n40743 );
and ( n48132 , n48129 , n48131 );
xor ( n48133 , n44847 , n48132 );
not ( n17297 , n29614 );
and ( n17298 , n17297 , RI173ce7b8_1749);
and ( n17299 , n48133 , n29614 );
or ( n48134 , n17298 , n17299 );
not ( n17300 , RI1754c610_2);
and ( n17301 , n17300 , n48134 );
and ( n17302 , C0 , RI1754c610_2);
or ( n48135 , n17301 , n17302 );
buf ( n48136 , n48135 );
not ( n48137 , n44072 );
and ( n48138 , n48137 , n42158 );
xor ( n48139 , n44069 , n48138 );
not ( n17303 , n29614 );
and ( n17304 , n17303 , RI173d5df0_1713);
and ( n17305 , n48139 , n29614 );
or ( n48140 , n17304 , n17305 );
not ( n17306 , RI1754c610_2);
and ( n17307 , n17306 , n48140 );
and ( n17308 , C0 , RI1754c610_2);
or ( n48141 , n17307 , n17308 );
buf ( n48142 , n48141 );
not ( n48143 , n47126 );
and ( n48144 , n48143 , n47128 );
xor ( n48145 , n46396 , n48144 );
not ( n17309 , n29614 );
and ( n17310 , n17309 , RI174aadc0_903);
and ( n17311 , n48145 , n29614 );
or ( n48146 , n17310 , n17311 );
not ( n17312 , RI1754c610_2);
and ( n17313 , n17312 , n48146 );
and ( n17314 , C0 , RI1754c610_2);
or ( n48147 , n17313 , n17314 );
buf ( n48148 , n48147 );
not ( n48149 , n41330 );
and ( n48150 , n48149 , n39960 );
xor ( n48151 , n41327 , n48150 );
not ( n17315 , n29614 );
and ( n17316 , n17315 , RI1744a448_1374);
and ( n17317 , n48151 , n29614 );
or ( n48152 , n17316 , n17317 );
not ( n17318 , RI1754c610_2);
and ( n17319 , n17318 , n48152 );
and ( n17320 , C0 , RI1754c610_2);
or ( n48153 , n17319 , n17320 );
buf ( n48154 , n48153 );
not ( n48155 , n41905 );
and ( n48156 , n48155 , n41907 );
xor ( n48157 , n43383 , n48156 );
not ( n17321 , n29614 );
and ( n17322 , n17321 , RI173e2618_1652);
and ( n17323 , n48157 , n29614 );
or ( n48158 , n17322 , n17323 );
not ( n17324 , RI1754c610_2);
and ( n17325 , n17324 , n48158 );
and ( n17326 , C0 , RI1754c610_2);
or ( n48159 , n17325 , n17326 );
buf ( n48160 , n48159 );
not ( n48161 , n37652 );
and ( n48162 , n48161 , n44600 );
xor ( n48163 , n37580 , n48162 );
not ( n17327 , n29614 );
and ( n17328 , n17327 , RI174bae28_829);
and ( n17329 , n48163 , n29614 );
or ( n48164 , n17328 , n17329 );
not ( n17330 , RI1754c610_2);
and ( n17331 , n17330 , n48164 );
and ( n17332 , C0 , RI1754c610_2);
or ( n48165 , n17331 , n17332 );
buf ( n48166 , n48165 );
xor ( n48167 , n36332 , n40718 );
xor ( n48168 , n48167 , n38676 );
xor ( n48169 , n41145 , n34087 );
xor ( n48170 , n48169 , n34127 );
not ( n48171 , n48170 );
xor ( n48172 , n38578 , n29109 );
xor ( n48173 , n48172 , n40463 );
and ( n48174 , n48171 , n48173 );
xor ( n48175 , n48168 , n48174 );
not ( n17333 , n29614 );
and ( n17334 , n17333 , RI17523be8_655);
and ( n17335 , n48175 , n29614 );
or ( n48176 , n17334 , n17335 );
not ( n17336 , RI1754c610_2);
and ( n17337 , n17336 , n48176 );
and ( n17338 , C0 , RI1754c610_2);
or ( n48177 , n17337 , n17338 );
buf ( n48178 , n48177 );
xor ( n48179 , n40423 , n39816 );
xor ( n48180 , n48179 , n35052 );
xor ( n48181 , n36049 , n34475 );
xor ( n48182 , n48181 , n37371 );
not ( n48183 , n48182 );
and ( n48184 , n48183 , n47306 );
xor ( n48185 , n48180 , n48184 );
not ( n17339 , n29614 );
and ( n17340 , n17339 , RI1744e5e8_1354);
and ( n17341 , n48185 , n29614 );
or ( n48186 , n17340 , n17341 );
not ( n17342 , RI1754c610_2);
and ( n17343 , n17342 , n48186 );
and ( n17344 , C0 , RI1754c610_2);
or ( n48187 , n17343 , n17344 );
buf ( n48188 , n48187 );
not ( n48189 , n42010 );
and ( n48190 , n48189 , n42761 );
xor ( n48191 , n42004 , n48190 );
not ( n17345 , n29614 );
and ( n17346 , n17345 , RI17456298_1316);
and ( n17347 , n48191 , n29614 );
or ( n48192 , n17346 , n17347 );
not ( n17348 , RI1754c610_2);
and ( n17349 , n17348 , n48192 );
and ( n17350 , C0 , RI1754c610_2);
or ( n48193 , n17349 , n17350 );
buf ( n48194 , n48193 );
not ( n17351 , n27683 );
and ( n17352 , n17351 , RI19a86fc0_2745);
and ( n17353 , RI19a887a8_2735 , n27683 );
or ( n48195 , n17352 , n17353 );
not ( n17354 , RI1754c610_2);
and ( n17355 , n17354 , n48195 );
and ( n17356 , C0 , RI1754c610_2);
or ( n48196 , n17355 , n17356 );
buf ( n48197 , n48196 );
buf ( n48198 , RI1750f710_718);
xor ( n48199 , n35973 , n37744 );
xor ( n48200 , n48199 , n35438 );
not ( n48201 , n48200 );
and ( n48202 , n48201 , n46721 );
xor ( n48203 , n47390 , n48202 );
not ( n17357 , n29614 );
and ( n17358 , n17357 , RI17393d48_2035);
and ( n17359 , n48203 , n29614 );
or ( n48204 , n17358 , n17359 );
not ( n17360 , RI1754c610_2);
and ( n17361 , n17360 , n48204 );
and ( n17362 , C0 , RI1754c610_2);
or ( n48205 , n17361 , n17362 );
buf ( n48206 , n48205 );
buf ( n48207 , RI174c0af8_811);
xor ( n48208 , n40033 , n40855 );
xor ( n48209 , n48208 , n38574 );
not ( n48210 , n48024 );
and ( n48211 , n48210 , n48026 );
xor ( n48212 , n48209 , n48211 );
not ( n17363 , n29614 );
and ( n17364 , n17363 , RI173c0550_1818);
and ( n17365 , n48212 , n29614 );
or ( n48213 , n17364 , n17365 );
not ( n17366 , RI1754c610_2);
and ( n17367 , n17366 , n48213 );
and ( n17368 , C0 , RI1754c610_2);
or ( n48214 , n17367 , n17368 );
buf ( n48215 , n48214 );
not ( n48216 , n40544 );
and ( n48217 , n48216 , n40565 );
xor ( n48218 , n45679 , n48217 );
not ( n17369 , n29614 );
and ( n17370 , n17369 , RI174972c0_999);
and ( n17371 , n48218 , n29614 );
or ( n48219 , n17370 , n17371 );
not ( n17372 , RI1754c610_2);
and ( n17373 , n17372 , n48219 );
and ( n17374 , C0 , RI1754c610_2);
or ( n48220 , n17373 , n17374 );
buf ( n48221 , n48220 );
not ( n48222 , n44585 );
and ( n48223 , n48222 , n40255 );
xor ( n48224 , n44582 , n48223 );
not ( n17375 , n29614 );
and ( n17376 , n17375 , RI173d3690_1725);
and ( n17377 , n48224 , n29614 );
or ( n48225 , n17376 , n17377 );
not ( n17378 , RI1754c610_2);
and ( n17379 , n17378 , n48225 );
and ( n17380 , C0 , RI1754c610_2);
or ( n48226 , n17379 , n17380 );
buf ( n48227 , n48226 );
not ( n17381 , n27683 );
and ( n17382 , n17381 , RI19a89888_2727);
and ( n17383 , RI19a93ba8_2656 , n27683 );
or ( n48228 , n17382 , n17383 );
not ( n17384 , RI1754c610_2);
and ( n17385 , n17384 , n48228 );
and ( n17386 , C0 , RI1754c610_2);
or ( n48229 , n17385 , n17386 );
buf ( n48230 , n48229 );
not ( n48231 , n40120 );
xor ( n48232 , n35621 , n41543 );
xor ( n48233 , n48232 , n34669 );
and ( n48234 , n48231 , n48233 );
xor ( n48235 , n40117 , n48234 );
not ( n17387 , n29614 );
and ( n17388 , n17387 , RI17485548_1086);
and ( n17389 , n48235 , n29614 );
or ( n48236 , n17388 , n17389 );
not ( n17390 , RI1754c610_2);
and ( n17391 , n17390 , n48236 );
and ( n17392 , C0 , RI1754c610_2);
or ( n48237 , n17391 , n17392 );
buf ( n48238 , n48237 );
not ( n17393 , n27683 );
and ( n17394 , n17393 , RI19ac0338_2330);
and ( n17395 , RI19ac9500_2260 , n27683 );
or ( n48239 , n17394 , n17395 );
not ( n17396 , RI1754c610_2);
and ( n17397 , n17396 , n48239 );
and ( n17398 , C0 , RI1754c610_2);
or ( n48240 , n17397 , n17398 );
buf ( n48241 , n48240 );
not ( n17399 , n27683 );
and ( n17400 , n17399 , RI19a9ff20_2569);
and ( n17401 , RI19aa9bb0_2498 , n27683 );
or ( n48242 , n17400 , n17401 );
not ( n17402 , RI1754c610_2);
and ( n17403 , n17402 , n48242 );
and ( n17404 , C0 , RI1754c610_2);
or ( n48243 , n17403 , n17404 );
buf ( n48244 , n48243 );
buf ( n48245 , RI17499048_990);
not ( n48246 , n42532 );
and ( n48247 , n48246 , n42534 );
xor ( n48248 , n43113 , n48247 );
not ( n17405 , n29614 );
and ( n17406 , n17405 , RI174c1020_810);
and ( n17407 , n48248 , n29614 );
or ( n48249 , n17406 , n17407 );
not ( n17408 , RI1754c610_2);
and ( n17409 , n17408 , n48249 );
and ( n17410 , C0 , RI1754c610_2);
or ( n48250 , n17409 , n17410 );
buf ( n48251 , n48250 );
buf ( n48252 , RI17482410_1101);
xor ( n48253 , n36236 , n41370 );
xor ( n48254 , n48253 , n37898 );
not ( n48255 , n43195 );
and ( n48256 , n48255 , n43197 );
xor ( n48257 , n48254 , n48256 );
not ( n17411 , n29614 );
and ( n17412 , n17411 , RI17347650_2093);
and ( n17413 , n48257 , n29614 );
or ( n48258 , n17412 , n17413 );
not ( n17414 , RI1754c610_2);
and ( n17415 , n17414 , n48258 );
and ( n17416 , C0 , RI1754c610_2);
or ( n48259 , n17415 , n17416 );
buf ( n48260 , n48259 );
buf ( n48261 , RI174b8a10_836);
buf ( n48262 , RI174c5850_796);
buf ( n48263 , RI17492748_1022);
buf ( n48264 , RI1749a740_983);
xor ( n48265 , n41658 , n40692 );
xor ( n48266 , n48265 , n43994 );
not ( n48267 , n40177 );
and ( n48268 , n48267 , n40211 );
xor ( n48269 , n48266 , n48268 );
not ( n17417 , n29614 );
and ( n17418 , n17417 , RI174a7fd0_917);
and ( n17419 , n48269 , n29614 );
or ( n48270 , n17418 , n17419 );
not ( n17420 , RI1754c610_2);
and ( n17421 , n17420 , n48270 );
and ( n17422 , C0 , RI1754c610_2);
or ( n48271 , n17421 , n17422 );
buf ( n48272 , n48271 );
not ( n17423 , n27683 );
and ( n17424 , n17423 , RI19ab8430_2393);
and ( n17425 , RI19ac1148_2322 , n27683 );
or ( n48273 , n17424 , n17425 );
not ( n17426 , RI1754c610_2);
and ( n17427 , n17426 , n48273 );
and ( n17428 , C0 , RI1754c610_2);
or ( n48274 , n17427 , n17428 );
buf ( n48275 , n48274 );
not ( n17429 , n27683 );
and ( n17430 , n17429 , RI19a9f728_2573);
and ( n17431 , RI19aa9430_2501 , n27683 );
or ( n48276 , n17430 , n17431 );
not ( n17432 , RI1754c610_2);
and ( n17433 , n17432 , n48276 );
and ( n17434 , C0 , RI1754c610_2);
or ( n48277 , n17433 , n17434 );
buf ( n48278 , n48277 );
not ( n17435 , n27683 );
and ( n17436 , n17435 , RI19aad300_2474);
and ( n17437 , RI19ab7008_2402 , n27683 );
or ( n48279 , n17436 , n17437 );
not ( n17438 , RI1754c610_2);
and ( n17439 , n17438 , n48279 );
and ( n17440 , C0 , RI1754c610_2);
or ( n48280 , n17439 , n17440 );
buf ( n48281 , n48280 );
buf ( n48282 , RI174cde60_770);
xor ( n48283 , n43273 , n41099 );
xor ( n48284 , n48283 , n30604 );
xor ( n48285 , n35215 , n43492 );
xor ( n48286 , n48285 , n38634 );
not ( n48287 , n48286 );
xor ( n48288 , n30260 , n35311 );
xor ( n48289 , n48288 , n35361 );
and ( n48290 , n48287 , n48289 );
xor ( n48291 , n48284 , n48290 );
not ( n17441 , n29614 );
and ( n17442 , n17441 , RI1752c720_628);
and ( n17443 , n48291 , n29614 );
or ( n48292 , n17442 , n17443 );
not ( n17444 , RI1754c610_2);
and ( n17445 , n17444 , n48292 );
and ( n17446 , C0 , RI1754c610_2);
or ( n48293 , n17445 , n17446 );
buf ( n48294 , n48293 );
xor ( n48295 , n34095 , n42377 );
xor ( n48296 , n48295 , n33991 );
not ( n48297 , n48296 );
and ( n48298 , n48297 , n47694 );
xor ( n48299 , n46983 , n48298 );
not ( n17447 , n29614 );
and ( n17448 , n17447 , RI1752ffd8_617);
and ( n17449 , n48299 , n29614 );
or ( n48300 , n17448 , n17449 );
not ( n17450 , RI1754c610_2);
and ( n17451 , n17450 , n48300 );
and ( n17452 , C0 , RI1754c610_2);
or ( n48301 , n17451 , n17452 );
buf ( n48302 , n48301 );
buf ( n48303 , RI174b5518_852);
xor ( n48304 , n41918 , n42033 );
xor ( n48305 , n48304 , n37987 );
xor ( n48306 , n38225 , n39450 );
xor ( n48307 , n48306 , n39467 );
not ( n48308 , n48307 );
xor ( n48309 , n36934 , n32620 );
xor ( n48310 , n48309 , n33337 );
and ( n48311 , n48308 , n48310 );
xor ( n48312 , n48305 , n48311 );
not ( n17453 , n29614 );
and ( n17454 , n17453 , RI174abe28_898);
and ( n17455 , n48312 , n29614 );
or ( n48313 , n17454 , n17455 );
not ( n17456 , RI1754c610_2);
and ( n17457 , n17456 , n48313 );
and ( n17458 , C0 , RI1754c610_2);
or ( n48314 , n17457 , n17458 );
buf ( n48315 , n48314 );
buf ( n48316 , RI1749dbc0_967);
buf ( n48317 , RI1748ceb0_1049);
xor ( n48318 , n36905 , n32560 );
xor ( n48319 , n48318 , n32620 );
not ( n48320 , n47824 );
and ( n48321 , n48320 , n47826 );
xor ( n48322 , n48319 , n48321 );
not ( n17459 , n29614 );
and ( n17460 , n17459 , RI1744f998_1348);
and ( n17461 , n48322 , n29614 );
or ( n48323 , n17460 , n17461 );
not ( n17462 , RI1754c610_2);
and ( n17463 , n17462 , n48323 );
and ( n17464 , C0 , RI1754c610_2);
or ( n48324 , n17463 , n17464 );
buf ( n48325 , n48324 );
not ( n17465 , n27683 );
and ( n17466 , n17465 , RI19aa2248_2551);
and ( n17467 , RI19aac838_2479 , n27683 );
or ( n48326 , n17466 , n17467 );
not ( n17468 , RI1754c610_2);
and ( n17469 , n17468 , n48326 );
and ( n17470 , C0 , RI1754c610_2);
or ( n48327 , n17469 , n17470 );
buf ( n48328 , n48327 );
not ( n48329 , n43099 );
and ( n48330 , n48329 , n45912 );
xor ( n48331 , n43096 , n48330 );
not ( n17471 , n29614 );
and ( n17472 , n17471 , RI17359698_2089);
and ( n17473 , n48331 , n29614 );
or ( n48332 , n17472 , n17473 );
not ( n17474 , RI1754c610_2);
and ( n17475 , n17474 , n48332 );
and ( n17476 , C0 , RI1754c610_2);
or ( n48333 , n17475 , n17476 );
buf ( n48334 , n48333 );
not ( n17477 , n27683 );
and ( n17478 , n17477 , RI19ab11d0_2445);
and ( n17479 , RI19abaf50_2374 , n27683 );
or ( n48335 , n17478 , n17479 );
not ( n17480 , RI1754c610_2);
and ( n17481 , n17480 , n48335 );
and ( n17482 , C0 , RI1754c610_2);
or ( n48336 , n17481 , n17482 );
buf ( n48337 , n48336 );
not ( n17483 , n27683 );
and ( n17484 , n17483 , RI19ab0528_2451);
and ( n17485 , RI19aba398_2379 , n27683 );
or ( n48338 , n17484 , n17485 );
not ( n17486 , RI1754c610_2);
and ( n17487 , n17486 , n48338 );
and ( n17488 , C0 , RI1754c610_2);
or ( n48339 , n17487 , n17488 );
buf ( n48340 , n48339 );
xor ( n48341 , n38941 , n36917 );
xor ( n48342 , n48341 , n36947 );
not ( n48343 , n48342 );
xor ( n48344 , n41786 , n35955 );
xor ( n48345 , n48344 , n42554 );
and ( n48346 , n48343 , n48345 );
xor ( n48347 , n47607 , n48346 );
not ( n17489 , n29614 );
and ( n17490 , n17489 , RI17409f60_1459);
and ( n17491 , n48347 , n29614 );
or ( n48348 , n17490 , n17491 );
not ( n17492 , RI1754c610_2);
and ( n17493 , n17492 , n48348 );
and ( n17494 , C0 , RI1754c610_2);
or ( n48349 , n17493 , n17494 );
buf ( n48350 , n48349 );
not ( n48351 , n41564 );
xor ( n48352 , n40396 , n32973 );
xor ( n48353 , n48352 , n39816 );
and ( n48354 , n48351 , n48353 );
xor ( n48355 , n41561 , n48354 );
not ( n17495 , n29614 );
and ( n17496 , n17495 , RI173a88b0_1934);
and ( n17497 , n48355 , n29614 );
or ( n48356 , n17496 , n17497 );
not ( n17498 , RI1754c610_2);
and ( n17499 , n17498 , n48356 );
and ( n17500 , C0 , RI1754c610_2);
or ( n48357 , n17499 , n17500 );
buf ( n48358 , n48357 );
not ( n48359 , n40839 );
and ( n48360 , n48359 , n40857 );
xor ( n48361 , n44647 , n48360 );
not ( n17501 , n29614 );
and ( n17502 , n17501 , RI1749add0_981);
and ( n17503 , n48361 , n29614 );
or ( n48362 , n17502 , n17503 );
not ( n17504 , RI1754c610_2);
and ( n17505 , n17504 , n48362 );
and ( n17506 , C0 , RI1754c610_2);
or ( n48363 , n17505 , n17506 );
buf ( n48364 , n48363 );
not ( n17507 , n27683 );
and ( n17508 , n17507 , RI19ac2a98_2309);
and ( n17509 , RI19acba08_2242 , n27683 );
or ( n48365 , n17508 , n17509 );
not ( n17510 , RI1754c610_2);
and ( n17511 , n17510 , n48365 );
and ( n17512 , C0 , RI1754c610_2);
or ( n48366 , n17511 , n17512 );
buf ( n48367 , n48366 );
not ( n48368 , n44452 );
and ( n48369 , n48368 , n46695 );
xor ( n48370 , n44449 , n48369 );
not ( n17513 , n29614 );
and ( n17514 , n17513 , RI174afc80_879);
and ( n17515 , n48370 , n29614 );
or ( n48371 , n17514 , n17515 );
not ( n17516 , RI1754c610_2);
and ( n17517 , n17516 , n48371 );
and ( n17518 , C0 , RI1754c610_2);
or ( n48372 , n17517 , n17518 );
buf ( n48373 , n48372 );
xor ( n48374 , n38879 , n31506 );
xor ( n48375 , n48374 , n31621 );
xor ( n48376 , n30695 , n33728 );
xor ( n48377 , n48376 , n33778 );
not ( n48378 , n48377 );
xor ( n48379 , n41425 , n43464 );
xor ( n48380 , n48379 , n44146 );
and ( n48381 , n48378 , n48380 );
xor ( n48382 , n48375 , n48381 );
not ( n17519 , n29614 );
and ( n17520 , n17519 , RI1744be88_1366);
and ( n17521 , n48382 , n29614 );
or ( n48383 , n17520 , n17521 );
not ( n17522 , RI1754c610_2);
and ( n17523 , n17522 , n48383 );
and ( n17524 , C0 , RI1754c610_2);
or ( n48384 , n17523 , n17524 );
buf ( n48385 , n48384 );
not ( n17525 , n27683 );
and ( n17526 , n17525 , RI19a9eaf8_2579);
and ( n17527 , RI19aa81e8_2508 , n27683 );
or ( n48386 , n17526 , n17527 );
not ( n17528 , RI1754c610_2);
and ( n17529 , n17528 , n48386 );
and ( n17530 , C0 , RI1754c610_2);
or ( n48387 , n17529 , n17530 );
buf ( n48388 , n48387 );
xor ( n48389 , n38801 , n39621 );
xor ( n48390 , n48389 , n40855 );
not ( n48391 , n42266 );
and ( n48392 , n48391 , n42268 );
xor ( n48393 , n48390 , n48392 );
not ( n17531 , n29614 );
and ( n17532 , n17531 , RI174b16c0_871);
and ( n17533 , n48393 , n29614 );
or ( n48394 , n17532 , n17533 );
not ( n17534 , RI1754c610_2);
and ( n17535 , n17534 , n48394 );
and ( n17536 , C0 , RI1754c610_2);
or ( n48395 , n17535 , n17536 );
buf ( n48396 , n48395 );
xor ( n48397 , n31254 , n42049 );
xor ( n48398 , n48397 , n37849 );
not ( n48399 , n48398 );
and ( n48400 , n48399 , n42369 );
xor ( n48401 , n45839 , n48400 );
not ( n17537 , n29614 );
and ( n17538 , n17537 , RI174b5ba8_850);
and ( n17539 , n48401 , n29614 );
or ( n48402 , n17538 , n17539 );
not ( n17540 , RI1754c610_2);
and ( n17541 , n17540 , n48402 );
and ( n17542 , C0 , RI1754c610_2);
or ( n48403 , n17541 , n17542 );
buf ( n48404 , n48403 );
not ( n48405 , n43745 );
and ( n48406 , n48405 , n43747 );
xor ( n48407 , n43850 , n48406 );
not ( n17543 , n29614 );
and ( n17544 , n17543 , RI1733fce8_2130);
and ( n17545 , n48407 , n29614 );
or ( n48408 , n17544 , n17545 );
not ( n17546 , RI1754c610_2);
and ( n17547 , n17546 , n48408 );
and ( n17548 , C0 , RI1754c610_2);
or ( n48409 , n17547 , n17548 );
buf ( n48410 , n48409 );
xor ( n48411 , n39177 , n40166 );
xor ( n48412 , n48411 , n41590 );
not ( n48413 , n48266 );
and ( n48414 , n48413 , n40177 );
xor ( n48415 , n48412 , n48414 );
not ( n17549 , n29614 );
and ( n17550 , n17549 , RI17499390_989);
and ( n17551 , n48415 , n29614 );
or ( n48416 , n17550 , n17551 );
not ( n17552 , RI1754c610_2);
and ( n17553 , n17552 , n48416 );
and ( n17554 , C0 , RI1754c610_2);
or ( n48417 , n17553 , n17554 );
buf ( n48418 , n48417 );
not ( n48419 , n47362 );
and ( n48420 , n48419 , n41936 );
xor ( n48421 , n41898 , n48420 );
not ( n17555 , n29614 );
and ( n17556 , n17555 , RI1744aad8_1372);
and ( n17557 , n48421 , n29614 );
or ( n48422 , n17556 , n17557 );
not ( n17558 , RI1754c610_2);
and ( n17559 , n17558 , n48422 );
and ( n17560 , C0 , RI1754c610_2);
or ( n48423 , n17559 , n17560 );
buf ( n48424 , n48423 );
not ( n17561 , n27683 );
and ( n17562 , n17561 , RI19a946e8_2651);
and ( n17563 , RI19a9eaf8_2579 , n27683 );
or ( n48425 , n17562 , n17563 );
not ( n17564 , RI1754c610_2);
and ( n17565 , n17564 , n48425 );
and ( n17566 , C0 , RI1754c610_2);
or ( n48426 , n17565 , n17566 );
buf ( n48427 , n48426 );
xor ( n48428 , n30671 , n33728 );
xor ( n48429 , n48428 , n33778 );
not ( n48430 , n46197 );
and ( n48431 , n48430 , n46199 );
xor ( n48432 , n48429 , n48431 );
not ( n17567 , n29614 );
and ( n17568 , n17567 , RI174c0af8_811);
and ( n17569 , n48432 , n29614 );
or ( n48433 , n17568 , n17569 );
not ( n17570 , RI1754c610_2);
and ( n17571 , n17570 , n48433 );
and ( n17572 , C0 , RI1754c610_2);
or ( n48434 , n17571 , n17572 );
buf ( n48435 , n48434 );
not ( n48436 , n41076 );
and ( n48437 , n48436 , n41078 );
xor ( n48438 , n41829 , n48437 );
not ( n17573 , n29614 );
and ( n17574 , n17573 , RI173e50c0_1639);
and ( n17575 , n48438 , n29614 );
or ( n48439 , n17574 , n17575 );
not ( n17576 , RI1754c610_2);
and ( n17577 , n17576 , n48439 );
and ( n17578 , C0 , RI1754c610_2);
or ( n48440 , n17577 , n17578 );
buf ( n48441 , n48440 );
not ( n17579 , n27683 );
and ( n17580 , n17579 , RI19a9f188_2576);
and ( n17581 , RI19aa8bc0_2505 , n27683 );
or ( n48442 , n17580 , n17581 );
not ( n17582 , RI1754c610_2);
and ( n17583 , n17582 , n48442 );
and ( n17584 , C0 , RI1754c610_2);
or ( n48443 , n17583 , n17584 );
buf ( n48444 , n48443 );
xor ( n48445 , n38643 , n34300 );
xor ( n48446 , n48445 , n34340 );
xor ( n48447 , n28467 , n41799 );
xor ( n48448 , n48447 , n40381 );
not ( n48449 , n48448 );
xor ( n48450 , n35720 , n39563 );
xor ( n48451 , n48450 , n35416 );
and ( n48452 , n48449 , n48451 );
xor ( n48453 , n48446 , n48452 );
not ( n17585 , n29614 );
and ( n17586 , n17585 , RI17512aa0_708);
and ( n17587 , n48453 , n29614 );
or ( n48454 , n17586 , n17587 );
not ( n17588 , RI1754c610_2);
and ( n17589 , n17588 , n48454 );
and ( n17590 , C0 , RI1754c610_2);
or ( n48455 , n17589 , n17590 );
buf ( n48456 , n48455 );
not ( n17591 , n27683 );
and ( n17592 , n17591 , RI19ab1518_2444);
and ( n17593 , RI19abb298_2373 , n27683 );
or ( n48457 , n17592 , n17593 );
not ( n17594 , RI1754c610_2);
and ( n17595 , n17594 , n48457 );
and ( n17596 , C0 , RI1754c610_2);
or ( n48458 , n17595 , n17596 );
buf ( n48459 , n48458 );
not ( n48460 , n38496 );
and ( n48461 , n48460 , n34128 );
xor ( n48462 , n46343 , n48461 );
not ( n17597 , n29614 );
and ( n17598 , n17597 , RI173bc6f8_1837);
and ( n17599 , n48462 , n29614 );
or ( n48463 , n17598 , n17599 );
not ( n17600 , RI1754c610_2);
and ( n17601 , n17600 , n48463 );
and ( n17602 , C0 , RI1754c610_2);
or ( n48464 , n17601 , n17602 );
buf ( n48465 , n48464 );
xor ( n48466 , n34484 , n29610 );
xor ( n48467 , n48466 , n31380 );
not ( n48468 , n46826 );
and ( n48469 , n48468 , n46828 );
xor ( n48470 , n48467 , n48469 );
not ( n17603 , n29614 );
and ( n17604 , n17603 , RI173ccd78_1757);
and ( n17605 , n48470 , n29614 );
or ( n48471 , n17604 , n17605 );
not ( n17606 , RI1754c610_2);
and ( n17607 , n17606 , n48471 );
and ( n17608 , C0 , RI1754c610_2);
or ( n48472 , n17607 , n17608 );
buf ( n48473 , n48472 );
not ( n17609 , n27683 );
and ( n17610 , n17609 , RI19abddb8_2351);
and ( n17611 , RI19ac6bc0_2279 , n27683 );
or ( n48474 , n17610 , n17611 );
not ( n17612 , RI1754c610_2);
and ( n17613 , n17612 , n48474 );
and ( n17614 , C0 , RI1754c610_2);
or ( n48475 , n17613 , n17614 );
buf ( n48476 , n48475 );
not ( n17615 , n27683 );
and ( n17616 , n17615 , RI19abb5e0_2372);
and ( n17617 , RI19ac3d58_2300 , n27683 );
or ( n48477 , n17616 , n17617 );
not ( n17618 , RI1754c610_2);
and ( n17619 , n17618 , n48477 );
and ( n17620 , C0 , RI1754c610_2);
or ( n48478 , n17619 , n17620 );
buf ( n48479 , n48478 );
xor ( n48480 , n29065 , n34517 );
xor ( n48481 , n48480 , n35911 );
not ( n48482 , n48481 );
and ( n48483 , n48482 , n43534 );
xor ( n48484 , n46469 , n48483 );
not ( n17621 , n29614 );
and ( n17622 , n17621 , RI173ed0b8_1600);
and ( n17623 , n48484 , n29614 );
or ( n48485 , n17622 , n17623 );
not ( n17624 , RI1754c610_2);
and ( n17625 , n17624 , n48485 );
and ( n17626 , C0 , RI1754c610_2);
or ( n48486 , n17625 , n17626 );
buf ( n48487 , n48486 );
xor ( n48488 , n41929 , n42033 );
xor ( n48489 , n48488 , n37987 );
not ( n48490 , n47984 );
and ( n48491 , n48490 , n47986 );
xor ( n48492 , n48489 , n48491 );
not ( n17627 , n29614 );
and ( n17628 , n17627 , RI17490678_1032);
and ( n17629 , n48492 , n29614 );
or ( n48493 , n17628 , n17629 );
not ( n17630 , RI1754c610_2);
and ( n17631 , n17630 , n48493 );
and ( n17632 , C0 , RI1754c610_2);
or ( n48494 , n17631 , n17632 );
buf ( n48495 , n48494 );
and ( n48496 , RI1754af18_51 , n34844 );
buf ( n48497 , n48496 );
not ( n17633 , n34859 );
and ( n17634 , n17633 , n48497 );
and ( n17635 , RI1754af18_51 , n34859 );
or ( n48498 , n17634 , n17635 );
not ( n17636 , RI19a22f70_2797);
and ( n17637 , n17636 , n48498 );
and ( n17638 , C0 , RI19a22f70_2797);
or ( n48499 , n17637 , n17638 );
not ( n17639 , n27683 );
and ( n17640 , n17639 , RI19a23330_2795);
and ( n17641 , n48499 , n27683 );
or ( n48500 , n17640 , n17641 );
not ( n17642 , RI1754c610_2);
and ( n17643 , n17642 , n48500 );
and ( n17644 , C0 , RI1754c610_2);
or ( n48501 , n17643 , n17644 );
buf ( n48502 , n48501 );
xor ( n48503 , n39642 , n35216 );
xor ( n48504 , n48503 , n41241 );
not ( n48505 , n47168 );
and ( n48506 , n48505 , n47170 );
xor ( n48507 , n48504 , n48506 );
not ( n17645 , n29614 );
and ( n17646 , n17645 , RI1744b7f8_1368);
and ( n17647 , n48507 , n29614 );
or ( n48508 , n17646 , n17647 );
not ( n17648 , RI1754c610_2);
and ( n17649 , n17648 , n48508 );
and ( n17650 , C0 , RI1754c610_2);
or ( n48509 , n17649 , n17650 );
buf ( n48510 , n48509 );
not ( n48511 , n40390 );
and ( n48512 , n48511 , n40392 );
xor ( n48513 , n45143 , n48512 );
not ( n17651 , n29614 );
and ( n17652 , n17651 , RI174bb350_828);
and ( n17653 , n48513 , n29614 );
or ( n48514 , n17652 , n17653 );
not ( n17654 , RI1754c610_2);
and ( n17655 , n17654 , n48514 );
and ( n17656 , C0 , RI1754c610_2);
or ( n48515 , n17655 , n17656 );
buf ( n48516 , n48515 );
not ( n17657 , n27683 );
and ( n17658 , n17657 , RI19acda60_2227);
and ( n17659 , RI19a90368_2681 , n27683 );
or ( n48517 , n17658 , n17659 );
not ( n17660 , RI1754c610_2);
and ( n17661 , n17660 , n48517 );
and ( n17662 , C0 , RI1754c610_2);
or ( n48518 , n17661 , n17662 );
buf ( n48519 , n48518 );
not ( n48520 , n28469 );
and ( n48521 , n48520 , n29110 );
xor ( n48522 , n44559 , n48521 );
not ( n17663 , n29614 );
and ( n17664 , n17663 , RI1749f948_958);
and ( n17665 , n48522 , n29614 );
or ( n48523 , n17664 , n17665 );
not ( n17666 , RI1754c610_2);
and ( n17667 , n17666 , n48523 );
and ( n17668 , C0 , RI1754c610_2);
or ( n48524 , n17667 , n17668 );
buf ( n48525 , n48524 );
buf ( n48526 , RI174b23e0_867);
buf ( n48527 , RI174a0cf8_952);
not ( n48528 , n38116 );
and ( n48529 , n48528 , n38168 );
xor ( n48530 , n45500 , n48529 );
not ( n17669 , n29614 );
and ( n17670 , n17669 , RI1744b168_1370);
and ( n17671 , n48530 , n29614 );
or ( n48531 , n17670 , n17671 );
not ( n17672 , RI1754c610_2);
and ( n17673 , n17672 , n48531 );
and ( n17674 , C0 , RI1754c610_2);
or ( n48532 , n17673 , n17674 );
buf ( n48533 , n48532 );
xor ( n48534 , n42296 , n40769 );
xor ( n48535 , n48534 , n40949 );
not ( n48536 , n46246 );
and ( n48537 , n48536 , n44459 );
xor ( n48538 , n48535 , n48537 );
not ( n17675 , n29614 );
and ( n17676 , n17675 , RI17446fc8_1390);
and ( n17677 , n48538 , n29614 );
or ( n48539 , n17676 , n17677 );
not ( n17678 , RI1754c610_2);
and ( n17679 , n17678 , n48539 );
and ( n17680 , C0 , RI1754c610_2);
or ( n48540 , n17679 , n17680 );
buf ( n48541 , n48540 );
not ( n17681 , n27683 );
and ( n17682 , n17681 , RI19ab52f8_2415);
and ( n17683 , RI19abe9e8_2344 , n27683 );
or ( n48542 , n17682 , n17683 );
not ( n17684 , RI1754c610_2);
and ( n17685 , n17684 , n48542 );
and ( n17686 , C0 , RI1754c610_2);
or ( n48543 , n17685 , n17686 );
buf ( n48544 , n48543 );
xor ( n48545 , n33688 , n41854 );
xor ( n48546 , n48545 , n40283 );
not ( n48547 , n48546 );
xor ( n48548 , n39130 , n28111 );
xor ( n48549 , n48548 , n28468 );
and ( n48550 , n48547 , n48549 );
xor ( n48551 , n47435 , n48550 );
not ( n17687 , n29614 );
and ( n17688 , n17687 , RI17399298_2009);
and ( n17689 , n48551 , n29614 );
or ( n48552 , n17688 , n17689 );
not ( n17690 , RI1754c610_2);
and ( n17691 , n17690 , n48552 );
and ( n17692 , C0 , RI1754c610_2);
or ( n48553 , n17691 , n17692 );
buf ( n48554 , n48553 );
and ( n48555 , RI1754b080_48 , n34844 );
and ( n48556 , RI1754b080_48 , n34847 );
or ( n48557 , n48555 , n48556 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n17693 , n34859 );
and ( n17694 , n17693 , n48557 );
and ( n17695 , RI1754b080_48 , n34859 );
or ( n48558 , n17694 , n17695 );
not ( n17696 , RI19a22f70_2797);
and ( n17697 , n17696 , n48558 );
and ( n17698 , C0 , RI19a22f70_2797);
or ( n48559 , n17697 , n17698 );
not ( n17699 , n27683 );
and ( n17700 , n17699 , RI19ac36c8_2303);
and ( n17701 , n48559 , n27683 );
or ( n48560 , n17700 , n17701 );
not ( n17702 , RI1754c610_2);
and ( n17703 , n17702 , n48560 );
and ( n17704 , C0 , RI1754c610_2);
or ( n48561 , n17703 , n17704 );
buf ( n48562 , n48561 );
not ( n48563 , n45141 );
and ( n48564 , n48563 , n45143 );
xor ( n48565 , n40438 , n48564 );
not ( n17705 , n29614 );
and ( n17706 , n17705 , RI17530a28_615);
and ( n17707 , n48565 , n29614 );
or ( n48566 , n17706 , n17707 );
not ( n17708 , RI1754c610_2);
and ( n17709 , n17708 , n48566 );
and ( n17710 , C0 , RI1754c610_2);
or ( n48567 , n17709 , n17710 );
buf ( n48568 , n48567 );
not ( n48569 , n40632 );
and ( n48570 , n48569 , n45856 );
xor ( n48571 , n40626 , n48570 );
not ( n17711 , n29614 );
and ( n17712 , n17711 , RI17415a68_1402);
and ( n17713 , n48571 , n29614 );
or ( n48572 , n17712 , n17713 );
not ( n17714 , RI1754c610_2);
and ( n17715 , n17714 , n48572 );
and ( n17716 , C0 , RI1754c610_2);
or ( n48573 , n17715 , n17716 );
buf ( n48574 , n48573 );
not ( n48575 , n47602 );
and ( n48576 , n48575 , n47604 );
xor ( n48577 , n48345 , n48576 );
not ( n17717 , n29614 );
and ( n17718 , n17717 , RI173de478_1672);
and ( n17719 , n48577 , n29614 );
or ( n48578 , n17718 , n17719 );
not ( n17720 , RI1754c610_2);
and ( n17721 , n17720 , n48578 );
and ( n17722 , C0 , RI1754c610_2);
or ( n48579 , n17721 , n17722 );
buf ( n48580 , n48579 );
xor ( n48581 , n33222 , n31317 );
xor ( n48582 , n48581 , n40302 );
xor ( n48583 , n36070 , n37371 );
xor ( n48584 , n48583 , n36682 );
not ( n48585 , n48584 );
and ( n48586 , n48585 , n44874 );
xor ( n48587 , n48582 , n48586 );
not ( n17723 , n29614 );
and ( n17724 , n17723 , RI173c2968_1807);
and ( n17725 , n48587 , n29614 );
or ( n48588 , n17724 , n17725 );
not ( n17726 , RI1754c610_2);
and ( n17727 , n17726 , n48588 );
and ( n17728 , C0 , RI1754c610_2);
or ( n48589 , n17727 , n17728 );
buf ( n48590 , n48589 );
xor ( n48591 , n39943 , n38724 );
xor ( n48592 , n48591 , n29425 );
not ( n48593 , n47063 );
and ( n48594 , n48593 , n47065 );
xor ( n48595 , n48592 , n48594 );
not ( n17729 , n29614 );
and ( n17730 , n17729 , RI17514eb8_701);
and ( n17731 , n48595 , n29614 );
or ( n48596 , n17730 , n17731 );
not ( n17732 , RI1754c610_2);
and ( n17733 , n17732 , n48596 );
and ( n17734 , C0 , RI1754c610_2);
or ( n48597 , n17733 , n17734 );
buf ( n48598 , n48597 );
not ( n17735 , n27683 );
and ( n17736 , n17735 , RI19abf4b0_2338);
and ( n17737 , RI19ac8510_2267 , n27683 );
or ( n48599 , n17736 , n17737 );
not ( n17738 , RI1754c610_2);
and ( n17739 , n17738 , n48599 );
and ( n17740 , C0 , RI1754c610_2);
or ( n48600 , n17739 , n17740 );
buf ( n48601 , n48600 );
not ( n17741 , n27683 );
and ( n17742 , n17741 , RI19ab16f8_2443);
and ( n17743 , RI19abb5e0_2372 , n27683 );
or ( n48602 , n17742 , n17743 );
not ( n17744 , RI1754c610_2);
and ( n17745 , n17744 , n48602 );
and ( n17746 , C0 , RI1754c610_2);
or ( n48603 , n17745 , n17746 );
buf ( n48604 , n48603 );
not ( n48605 , n46942 );
and ( n48606 , n48605 , n35362 );
xor ( n48607 , n47682 , n48606 );
not ( n17747 , n29614 );
and ( n17748 , n17747 , RI17470350_1189);
and ( n17749 , n48607 , n29614 );
or ( n48608 , n17748 , n17749 );
not ( n17750 , RI1754c610_2);
and ( n17751 , n17750 , n48608 );
and ( n17752 , C0 , RI1754c610_2);
or ( n48609 , n17751 , n17752 );
buf ( n48610 , n48609 );
xor ( n48611 , n39064 , n39702 );
xor ( n48612 , n48611 , n39914 );
not ( n48613 , n46812 );
and ( n48614 , n48613 , n46814 );
xor ( n48615 , n48612 , n48614 );
not ( n17753 , n29614 );
and ( n17754 , n17753 , RI17403cf0_1489);
and ( n17755 , n48615 , n29614 );
or ( n48616 , n17754 , n17755 );
not ( n17756 , RI1754c610_2);
and ( n17757 , n17756 , n48616 );
and ( n17758 , C0 , RI1754c610_2);
or ( n48617 , n17757 , n17758 );
buf ( n48618 , n48617 );
not ( n48619 , n47337 );
and ( n48620 , n48619 , n47370 );
xor ( n48621 , n47334 , n48620 );
not ( n17759 , n29614 );
and ( n17760 , n17759 , RI173aca50_1914);
and ( n17761 , n48621 , n29614 );
or ( n48622 , n17760 , n17761 );
not ( n17762 , RI1754c610_2);
and ( n17763 , n17762 , n48622 );
and ( n17764 , C0 , RI1754c610_2);
or ( n48623 , n17763 , n17764 );
buf ( n48624 , n48623 );
not ( n17765 , RI1754a720_68);
and ( n17766 , n17765 , RI19a22f70_2797);
and ( n17767 , C1 , RI1754a720_68);
or ( n48625 , n17766 , n17767 );
not ( n48626 , RI1754c610_2);
and ( n48627 , n48625 , n48626 );
buf ( n48628 , n48627 );
xor ( n48629 , n39770 , n33125 );
xor ( n48630 , n48629 , n33175 );
not ( n48631 , n48630 );
xor ( n48632 , n36966 , n41818 );
xor ( n48633 , n48632 , n40662 );
and ( n48634 , n48631 , n48633 );
xor ( n48635 , n44935 , n48634 );
not ( n17768 , n29614 );
and ( n17769 , n17768 , RI17532918_609);
and ( n17770 , n48635 , n29614 );
or ( n48636 , n17769 , n17770 );
not ( n17771 , RI1754c610_2);
and ( n17772 , n17771 , n48636 );
and ( n17773 , C0 , RI1754c610_2);
or ( n48637 , n17772 , n17773 );
buf ( n48638 , n48637 );
xor ( n48639 , n39256 , n35361 );
xor ( n48640 , n48639 , n38445 );
not ( n48641 , n48640 );
xor ( n48642 , n32298 , n36003 );
xor ( n48643 , n48642 , n38553 );
and ( n48644 , n48641 , n48643 );
xor ( n48645 , n36160 , n48644 );
not ( n17774 , n29614 );
and ( n17775 , n17774 , RI174c05d0_812);
and ( n17776 , n48645 , n29614 );
or ( n48646 , n17775 , n17776 );
not ( n17777 , RI1754c610_2);
and ( n17778 , n17777 , n48646 );
and ( n17779 , C0 , RI1754c610_2);
or ( n48647 , n17778 , n17779 );
buf ( n48648 , n48647 );
buf ( n48649 , RI1746d218_1204);
not ( n17780 , RI1754c610_2);
and ( n17781 , n17780 , RI17539830_589);
and ( n17782 , C0 , RI1754c610_2);
or ( n48650 , n17781 , n17782 );
buf ( n48651 , n48650 );
not ( n48652 , n47435 );
and ( n48653 , n48652 , n48546 );
xor ( n48654 , n47432 , n48653 );
not ( n17783 , n29614 );
and ( n17784 , n17783 , RI1738ace8_2079);
and ( n17785 , n48654 , n29614 );
or ( n48655 , n17784 , n17785 );
not ( n17786 , RI1754c610_2);
and ( n17787 , n17786 , n48655 );
and ( n17788 , C0 , RI1754c610_2);
or ( n48656 , n17787 , n17788 );
buf ( n48657 , n48656 );
xor ( n48658 , n37116 , n40237 );
xor ( n48659 , n48658 , n40254 );
not ( n48660 , n48659 );
and ( n48661 , n48660 , n45603 );
xor ( n48662 , n43571 , n48661 );
not ( n17789 , n29614 );
and ( n17790 , n17789 , RI1733d588_2142);
and ( n17791 , n48662 , n29614 );
or ( n48663 , n17790 , n17791 );
not ( n17792 , RI1754c610_2);
and ( n17793 , n17792 , n48663 );
and ( n17794 , C0 , RI1754c610_2);
or ( n48664 , n17793 , n17794 );
buf ( n48665 , n48664 );
not ( n48666 , n40260 );
and ( n48667 , n48666 , n44582 );
xor ( n48668 , n40257 , n48667 );
not ( n17795 , n29614 );
and ( n17796 , n17795 , RI173ff178_1512);
and ( n17797 , n48668 , n29614 );
or ( n48669 , n17796 , n17797 );
not ( n17798 , RI1754c610_2);
and ( n17799 , n17798 , n48669 );
and ( n17800 , C0 , RI1754c610_2);
or ( n48670 , n17799 , n17800 );
buf ( n48671 , n48670 );
not ( n17801 , n27683 );
and ( n17802 , n17801 , RI19ab0870_2450);
and ( n17803 , RI19aba578_2378 , n27683 );
or ( n48672 , n17802 , n17803 );
not ( n17804 , RI1754c610_2);
and ( n17805 , n17804 , n48672 );
and ( n17806 , C0 , RI1754c610_2);
or ( n48673 , n17805 , n17806 );
buf ( n48674 , n48673 );
not ( n48675 , n44183 );
and ( n48676 , n48675 , n44185 );
xor ( n48677 , n40891 , n48676 );
not ( n17807 , n29614 );
and ( n17808 , n17807 , RI17472df8_1176);
and ( n17809 , n48677 , n29614 );
or ( n48678 , n17808 , n17809 );
not ( n17810 , RI1754c610_2);
and ( n17811 , n17810 , n48678 );
and ( n17812 , C0 , RI1754c610_2);
or ( n48679 , n17811 , n17812 );
buf ( n48680 , n48679 );
not ( n17813 , n27683 );
and ( n17814 , n17813 , RI19acf8d8_2214);
and ( n17815 , RI19aa4318_2536 , n27683 );
or ( n48681 , n17814 , n17815 );
not ( n17816 , RI1754c610_2);
and ( n17817 , n17816 , n48681 );
and ( n17818 , C0 , RI1754c610_2);
or ( n48682 , n17817 , n17818 );
buf ( n48683 , n48682 );
xor ( n48684 , n41798 , n35955 );
xor ( n48685 , n48684 , n42554 );
xor ( n48686 , n32231 , n36003 );
xor ( n48687 , n48686 , n38553 );
not ( n48688 , n48687 );
xor ( n48689 , n33633 , n35069 );
xor ( n48690 , n48689 , n41854 );
and ( n48691 , n48688 , n48690 );
xor ( n48692 , n48685 , n48691 );
not ( n17819 , n29614 );
and ( n17820 , n17819 , RI173b67d0_1866);
and ( n17821 , n48692 , n29614 );
or ( n48693 , n17820 , n17821 );
not ( n17822 , RI1754c610_2);
and ( n17823 , n17822 , n48693 );
and ( n17824 , C0 , RI1754c610_2);
or ( n48694 , n17823 , n17824 );
buf ( n48695 , n48694 );
not ( n48696 , n44447 );
and ( n48697 , n48696 , n44449 );
xor ( n48698 , n46698 , n48697 );
not ( n17825 , n29614 );
and ( n17826 , n17825 , RI17520330_666);
and ( n17827 , n48698 , n29614 );
or ( n48699 , n17826 , n17827 );
not ( n17828 , RI1754c610_2);
and ( n17829 , n17828 , n48699 );
and ( n17830 , C0 , RI1754c610_2);
or ( n48700 , n17829 , n17830 );
buf ( n48701 , n48700 );
not ( n17831 , n27683 );
and ( n17832 , n17831 , RI19acb828_2243);
and ( n17833 , RI19a87218_2744 , n27683 );
or ( n48702 , n17832 , n17833 );
not ( n17834 , RI1754c610_2);
and ( n17835 , n17834 , n48702 );
and ( n17836 , C0 , RI1754c610_2);
or ( n48703 , n17835 , n17836 );
buf ( n48704 , n48703 );
not ( n17837 , n27683 );
and ( n17838 , n17837 , RI19aa90e8_2502);
and ( n17839 , RI19ab2f58_2432 , n27683 );
or ( n48705 , n17838 , n17839 );
not ( n17840 , RI1754c610_2);
and ( n17841 , n17840 , n48705 );
and ( n17842 , C0 , RI1754c610_2);
or ( n48706 , n17841 , n17842 );
buf ( n48707 , n48706 );
not ( n48708 , n40130 );
and ( n48709 , n48708 , n40167 );
xor ( n48710 , n45466 , n48709 );
not ( n17843 , n29614 );
and ( n17844 , n17843 , RI174a23f0_945);
and ( n17845 , n48710 , n29614 );
or ( n48711 , n17844 , n17845 );
not ( n17846 , RI1754c610_2);
and ( n17847 , n17846 , n48711 );
and ( n17848 , C0 , RI1754c610_2);
or ( n48712 , n17847 , n17848 );
buf ( n48713 , n48712 );
not ( n17849 , n27683 );
and ( n17850 , n17849 , RI19a8acb0_2719);
and ( n17851 , RI19a94b98_2649 , n27683 );
or ( n48714 , n17850 , n17851 );
not ( n17852 , RI1754c610_2);
and ( n17853 , n17852 , n48714 );
and ( n17854 , C0 , RI1754c610_2);
or ( n48715 , n17853 , n17854 );
buf ( n48716 , n48715 );
xor ( n48717 , n39082 , n36377 );
xor ( n48718 , n48717 , n39131 );
not ( n48719 , n48718 );
and ( n48720 , n48719 , n46311 );
xor ( n48721 , n45075 , n48720 );
not ( n17855 , n29614 );
and ( n17856 , n17855 , RI17454ba0_1323);
and ( n17857 , n48721 , n29614 );
or ( n48722 , n17856 , n17857 );
not ( n17858 , RI1754c610_2);
and ( n17859 , n17858 , n48722 );
and ( n17860 , C0 , RI1754c610_2);
or ( n48723 , n17859 , n17860 );
buf ( n48724 , n48723 );
not ( n48725 , n45319 );
and ( n48726 , n48725 , n45321 );
xor ( n48727 , n46951 , n48726 );
not ( n17861 , n29614 );
and ( n17862 , n17861 , RI173915e8_2047);
and ( n17863 , n48727 , n29614 );
or ( n48728 , n17862 , n17863 );
not ( n17864 , RI1754c610_2);
and ( n17865 , n17864 , n48728 );
and ( n17866 , C0 , RI1754c610_2);
or ( n48729 , n17865 , n17866 );
buf ( n48730 , n48729 );
xor ( n48731 , n39851 , n36742 );
xor ( n48732 , n48731 , n42504 );
xor ( n48733 , n37168 , n40254 );
xor ( n48734 , n48733 , n40718 );
not ( n48735 , n48734 );
xor ( n48736 , n38175 , n32220 );
xor ( n48737 , n48736 , n32309 );
and ( n48738 , n48735 , n48737 );
xor ( n48739 , n48732 , n48738 );
not ( n17867 , n29614 );
and ( n17868 , n17867 , RI1748d1f8_1048);
and ( n17869 , n48739 , n29614 );
or ( n48740 , n17868 , n17869 );
not ( n17870 , RI1754c610_2);
and ( n17871 , n17870 , n48740 );
and ( n17872 , C0 , RI1754c610_2);
or ( n48741 , n17871 , n17872 );
buf ( n48742 , n48741 );
buf ( n48743 , RI174ad868_890);
xor ( n48744 , n36536 , n37438 );
xor ( n48745 , n48744 , n30247 );
not ( n48746 , n48745 );
xor ( n48747 , n41762 , n38188 );
xor ( n48748 , n48747 , n36195 );
and ( n48749 , n48746 , n48748 );
xor ( n48750 , n45617 , n48749 );
not ( n17873 , n29614 );
and ( n17874 , n17873 , RI174a0320_955);
and ( n17875 , n48750 , n29614 );
or ( n48751 , n17874 , n17875 );
not ( n17876 , RI1754c610_2);
and ( n17877 , n17876 , n48751 );
and ( n17878 , C0 , RI1754c610_2);
or ( n48752 , n17877 , n17878 );
buf ( n48753 , n48752 );
buf ( n48754 , RI174b5860_851);
buf ( n48755 , RI1749d878_968);
buf ( n48756 , RI174a5bb8_928);
not ( n48757 , n41592 );
and ( n48758 , n48757 , n45239 );
xor ( n48759 , n41573 , n48758 );
not ( n17879 , n29614 );
and ( n17880 , n17879 , RI173b50d8_1873);
and ( n17881 , n48759 , n29614 );
or ( n48760 , n17880 , n17881 );
not ( n17882 , RI1754c610_2);
and ( n17883 , n17882 , n48760 );
and ( n17884 , C0 , RI1754c610_2);
or ( n48761 , n17883 , n17884 );
buf ( n48762 , n48761 );
not ( n17885 , n27683 );
and ( n17886 , n17885 , RI19ab1860_2442);
and ( n17887 , RI19abb748_2371 , n27683 );
or ( n48763 , n17886 , n17887 );
not ( n17888 , RI1754c610_2);
and ( n17889 , n17888 , n48763 );
and ( n17890 , C0 , RI1754c610_2);
or ( n48764 , n17889 , n17890 );
buf ( n48765 , n48764 );
not ( n17891 , n27683 );
and ( n17892 , n17891 , RI19a94b98_2649);
and ( n17893 , RI19a9efa8_2577 , n27683 );
or ( n48766 , n17892 , n17893 );
not ( n17894 , RI1754c610_2);
and ( n17895 , n17894 , n48766 );
and ( n17896 , C0 , RI1754c610_2);
or ( n48767 , n17895 , n17896 );
buf ( n48768 , n48767 );
xor ( n48769 , n40854 , n35009 );
xor ( n48770 , n48769 , n28816 );
not ( n48771 , n48770 );
and ( n48772 , n48771 , n39415 );
xor ( n48773 , n47731 , n48772 );
not ( n17897 , n29614 );
and ( n17898 , n17897 , RI17497c98_996);
and ( n17899 , n48773 , n29614 );
or ( n48774 , n17898 , n17899 );
not ( n17900 , RI1754c610_2);
and ( n17901 , n17900 , n48774 );
and ( n17902 , C0 , RI1754c610_2);
or ( n48775 , n17901 , n17902 );
buf ( n48776 , n48775 );
not ( n48777 , n44784 );
xor ( n48778 , n36586 , n39791 );
xor ( n48779 , n48778 , n40915 );
and ( n48780 , n48777 , n48779 );
xor ( n48781 , n44781 , n48780 );
not ( n17903 , n29614 );
and ( n17904 , n17903 , RI17531478_613);
and ( n17905 , n48781 , n29614 );
or ( n48782 , n17904 , n17905 );
not ( n17906 , RI1754c610_2);
and ( n17907 , n17906 , n48782 );
and ( n17908 , C0 , RI1754c610_2);
or ( n48783 , n17907 , n17908 );
buf ( n48784 , n48783 );
buf ( n48785 , RI17467980_1231);
not ( n48786 , n40383 );
and ( n48787 , n48786 , n40978 );
xor ( n48788 , n40361 , n48787 );
not ( n17909 , n29614 );
and ( n17910 , n17909 , RI17339dc0_2159);
and ( n17911 , n48788 , n29614 );
or ( n48789 , n17910 , n17911 );
not ( n17912 , RI1754c610_2);
and ( n17913 , n17912 , n48789 );
and ( n17914 , C0 , RI1754c610_2);
or ( n48790 , n17913 , n17914 );
buf ( n48791 , n48790 );
not ( n48792 , n39508 );
and ( n48793 , n48792 , n39526 );
xor ( n48794 , n46708 , n48793 );
not ( n17915 , n29614 );
and ( n17916 , n17915 , RI17531ec8_611);
and ( n17917 , n48794 , n29614 );
or ( n48795 , n17916 , n17917 );
not ( n17918 , RI1754c610_2);
and ( n17919 , n17918 , n48795 );
and ( n17920 , C0 , RI1754c610_2);
or ( n48796 , n17919 , n17920 );
buf ( n48797 , n48796 );
xor ( n48798 , n35153 , n37915 );
xor ( n48799 , n48798 , n43492 );
xor ( n48800 , n37226 , n39467 );
xor ( n48801 , n48800 , n41391 );
not ( n48802 , n48801 );
xor ( n48803 , n36280 , n37311 );
xor ( n48804 , n48803 , n37942 );
and ( n48805 , n48802 , n48804 );
xor ( n48806 , n48799 , n48805 );
not ( n17921 , n29614 );
and ( n17922 , n17921 , RI173d7ec0_1703);
and ( n17923 , n48806 , n29614 );
or ( n48807 , n17922 , n17923 );
not ( n17924 , RI1754c610_2);
and ( n17925 , n17924 , n48807 );
and ( n17926 , C0 , RI1754c610_2);
or ( n48808 , n17925 , n17926 );
buf ( n48809 , n48808 );
not ( n48810 , n44290 );
and ( n48811 , n48810 , n42968 );
xor ( n48812 , n44287 , n48811 );
not ( n17927 , n29614 );
and ( n17928 , n17927 , RI173d6e58_1708);
and ( n17929 , n48812 , n29614 );
or ( n48813 , n17928 , n17929 );
not ( n17930 , RI1754c610_2);
and ( n17931 , n17930 , n48813 );
and ( n17932 , C0 , RI1754c610_2);
or ( n48814 , n17931 , n17932 );
buf ( n48815 , n48814 );
not ( n48816 , n44698 );
xor ( n48817 , n39396 , n35594 );
xor ( n48818 , n48817 , n32403 );
and ( n48819 , n48816 , n48818 );
xor ( n48820 , n37341 , n48819 );
not ( n17933 , n29614 );
and ( n17934 , n17933 , RI17485f20_1083);
and ( n17935 , n48820 , n29614 );
or ( n48821 , n17934 , n17935 );
not ( n17936 , RI1754c610_2);
and ( n17937 , n17936 , n48821 );
and ( n17938 , C0 , RI1754c610_2);
or ( n48822 , n17937 , n17938 );
buf ( n48823 , n48822 );
not ( n17939 , n27683 );
and ( n17940 , n17939 , RI19abfc30_2334);
and ( n17941 , RI19ac8c18_2264 , n27683 );
or ( n48824 , n17940 , n17941 );
not ( n17942 , RI1754c610_2);
and ( n17943 , n17942 , n48824 );
and ( n17944 , C0 , RI1754c610_2);
or ( n48825 , n17943 , n17944 );
buf ( n48826 , n48825 );
xor ( n48827 , n38133 , n31053 );
xor ( n48828 , n48827 , n35494 );
xor ( n48829 , n39873 , n42504 );
xor ( n48830 , n48829 , n41818 );
not ( n48831 , n48830 );
and ( n48832 , n48831 , n45624 );
xor ( n48833 , n48828 , n48832 );
not ( n17945 , n29614 );
and ( n17946 , n17945 , RI174c00a8_813);
and ( n17947 , n48833 , n29614 );
or ( n48834 , n17946 , n17947 );
not ( n17948 , RI1754c610_2);
and ( n17949 , n17948 , n48834 );
and ( n17950 , C0 , RI1754c610_2);
or ( n48835 , n17949 , n17950 );
buf ( n48836 , n48835 );
xor ( n48837 , n32077 , n36702 );
xor ( n48838 , n48837 , n38872 );
not ( n48839 , n48838 );
and ( n48840 , n48839 , n47716 );
xor ( n48841 , n44575 , n48840 );
not ( n17951 , n29614 );
and ( n17952 , n17951 , RI174cba48_777);
and ( n17953 , n48841 , n29614 );
or ( n48842 , n17952 , n17953 );
not ( n17954 , RI1754c610_2);
and ( n17955 , n17954 , n48842 );
and ( n17956 , C0 , RI1754c610_2);
or ( n48843 , n17955 , n17956 );
buf ( n48844 , n48843 );
not ( n17957 , n27683 );
and ( n17958 , n17957 , RI19ab2328_2438);
and ( n17959 , RI19abc378_2366 , n27683 );
or ( n48845 , n17958 , n17959 );
not ( n17960 , RI1754c610_2);
and ( n17961 , n17960 , n48845 );
and ( n17962 , C0 , RI1754c610_2);
or ( n48846 , n17961 , n17962 );
buf ( n48847 , n48846 );
not ( n17963 , n27683 );
and ( n17964 , n17963 , RI19ab1ba8_2441);
and ( n17965 , RI19abbc70_2369 , n27683 );
or ( n48848 , n17964 , n17965 );
not ( n17966 , RI1754c610_2);
and ( n17967 , n17966 , n48848 );
and ( n17968 , C0 , RI1754c610_2);
or ( n48849 , n17967 , n17968 );
buf ( n48850 , n48849 );
not ( n17969 , n27683 );
and ( n17970 , n17969 , RI19aaa150_2495);
and ( n17971 , RI19ab4038_2423 , n27683 );
or ( n48851 , n17970 , n17971 );
not ( n17972 , RI1754c610_2);
and ( n17973 , n17972 , n48851 );
and ( n17974 , C0 , RI1754c610_2);
or ( n48852 , n17973 , n17974 );
buf ( n48853 , n48852 );
not ( n17975 , n27683 );
and ( n17976 , n17975 , RI19ab2148_2439);
and ( n17977 , RI19abc198_2367 , n27683 );
or ( n48854 , n17976 , n17977 );
not ( n17978 , RI1754c610_2);
and ( n17979 , n17978 , n48854 );
and ( n17980 , C0 , RI1754c610_2);
or ( n48855 , n17979 , n17980 );
buf ( n48856 , n48855 );
not ( n17981 , n27683 );
and ( n17982 , n17981 , RI19ab1ef0_2440);
and ( n17983 , RI19abbe50_2368 , n27683 );
or ( n48857 , n17982 , n17983 );
not ( n17984 , RI1754c610_2);
and ( n17985 , n17984 , n48857 );
and ( n17986 , C0 , RI1754c610_2);
or ( n48858 , n17985 , n17986 );
buf ( n48859 , n48858 );
not ( n48860 , n33779 );
and ( n48861 , n48860 , n44625 );
xor ( n48862 , n33698 , n48861 );
not ( n17987 , n29614 );
and ( n17988 , n17987 , RI17402c88_1494);
and ( n17989 , n48862 , n29614 );
or ( n48863 , n17988 , n17989 );
not ( n17990 , RI1754c610_2);
and ( n17991 , n17990 , n48863 );
and ( n17992 , C0 , RI1754c610_2);
or ( n48864 , n17991 , n17992 );
buf ( n48865 , n48864 );
not ( n48866 , n43122 );
xor ( n48867 , n36265 , n37311 );
xor ( n48868 , n48867 , n37942 );
and ( n48869 , n48866 , n48868 );
xor ( n48870 , n42100 , n48869 );
not ( n17993 , n29614 );
and ( n17994 , n17993 , RI17346930_2097);
and ( n17995 , n48870 , n29614 );
or ( n48871 , n17994 , n17995 );
not ( n17996 , RI1754c610_2);
and ( n17997 , n17996 , n48871 );
and ( n17998 , C0 , RI1754c610_2);
or ( n48872 , n17997 , n17998 );
buf ( n48873 , n48872 );
not ( n48874 , n48804 );
xor ( n48875 , n39181 , n40166 );
xor ( n48876 , n48875 , n41590 );
and ( n48877 , n48874 , n48876 );
xor ( n48878 , n48801 , n48877 );
not ( n17999 , n29614 );
and ( n18000 , n17999 , RI173e67b8_1632);
and ( n18001 , n48878 , n29614 );
or ( n48879 , n18000 , n18001 );
not ( n18002 , RI1754c610_2);
and ( n18003 , n18002 , n48879 );
and ( n18004 , C0 , RI1754c610_2);
or ( n48880 , n18003 , n18004 );
buf ( n48881 , n48880 );
xor ( n48882 , n34551 , n40563 );
xor ( n48883 , n48882 , n35544 );
not ( n48884 , n48883 );
and ( n48885 , n48884 , n47202 );
xor ( n48886 , n31381 , n48885 );
not ( n18005 , n29614 );
and ( n18006 , n18005 , RI174c7c68_789);
and ( n18007 , n48886 , n29614 );
or ( n48887 , n18006 , n18007 );
not ( n18008 , RI1754c610_2);
and ( n18009 , n18008 , n48887 );
and ( n18010 , C0 , RI1754c610_2);
or ( n48888 , n18009 , n18010 );
buf ( n48889 , n48888 );
buf ( n48890 , RI17512050_710);
xor ( n48891 , n37629 , n40149 );
xor ( n48892 , n48891 , n40166 );
xor ( n48893 , n35729 , n39563 );
xor ( n48894 , n48893 , n35416 );
not ( n48895 , n48894 );
and ( n48896 , n48895 , n46111 );
xor ( n48897 , n48892 , n48896 );
not ( n18011 , n29614 );
and ( n18012 , n18011 , RI1733dc18_2140);
and ( n18013 , n48897 , n29614 );
or ( n48898 , n18012 , n18013 );
not ( n18014 , RI1754c610_2);
and ( n18015 , n18014 , n48898 );
and ( n18016 , C0 , RI1754c610_2);
or ( n48899 , n18015 , n18016 );
buf ( n48900 , n48899 );
not ( n48901 , n48310 );
xor ( n48902 , n36247 , n41370 );
xor ( n48903 , n48902 , n37898 );
and ( n48904 , n48901 , n48903 );
xor ( n48905 , n48307 , n48904 );
not ( n18017 , n29614 );
and ( n18018 , n18017 , RI174bb878_827);
and ( n18019 , n48905 , n29614 );
or ( n48906 , n18018 , n18019 );
not ( n18020 , RI1754c610_2);
and ( n18021 , n18020 , n48906 );
and ( n18022 , C0 , RI1754c610_2);
or ( n48907 , n18021 , n18022 );
buf ( n48908 , n48907 );
buf ( n48909 , RI17480688_1110);
xor ( n48910 , n36677 , n39635 );
xor ( n48911 , n48910 , n39655 );
xor ( n48912 , n33879 , n41146 );
xor ( n48913 , n48912 , n37291 );
not ( n48914 , n48913 );
xor ( n48915 , n36199 , n32923 );
xor ( n48916 , n48915 , n32973 );
and ( n48917 , n48914 , n48916 );
xor ( n48918 , n48911 , n48917 );
not ( n18023 , n29614 );
and ( n18024 , n18023 , RI173f9c28_1538);
and ( n18025 , n48918 , n29614 );
or ( n48919 , n18024 , n18025 );
not ( n18026 , RI1754c610_2);
and ( n18027 , n18026 , n48919 );
and ( n18028 , C0 , RI1754c610_2);
or ( n48920 , n18027 , n18028 );
buf ( n48921 , n48920 );
not ( n48922 , n37312 );
and ( n48923 , n48922 , n37333 );
xor ( n48924 , n48818 , n48923 );
not ( n18029 , n29614 );
and ( n18030 , n18029 , RI174a3110_941);
and ( n18031 , n48924 , n29614 );
or ( n48925 , n18030 , n18031 );
not ( n18032 , RI1754c610_2);
and ( n18033 , n18032 , n48925 );
and ( n18034 , C0 , RI1754c610_2);
or ( n48926 , n18033 , n18034 );
buf ( n48927 , n48926 );
not ( n18035 , n27683 );
and ( n18036 , n18035 , RI19aa1438_2558);
and ( n18037 , RI19aab410_2487 , n27683 );
or ( n48928 , n18036 , n18037 );
not ( n18038 , RI1754c610_2);
and ( n18039 , n18038 , n48928 );
and ( n18040 , C0 , RI1754c610_2);
or ( n48929 , n18039 , n18040 );
buf ( n48930 , n48929 );
xor ( n48931 , n35509 , n38532 );
xor ( n48932 , n48931 , n38933 );
xor ( n48933 , n36147 , n39151 );
xor ( n48934 , n48933 , n38267 );
not ( n48935 , n48934 );
xor ( n48936 , n33465 , n40360 );
xor ( n48937 , n48936 , n35176 );
and ( n48938 , n48935 , n48937 );
xor ( n48939 , n48932 , n48938 );
not ( n18041 , n29614 );
and ( n18042 , n18041 , RI173f6e38_1552);
and ( n18043 , n48939 , n29614 );
or ( n48940 , n18042 , n18043 );
not ( n18044 , RI1754c610_2);
and ( n18045 , n18044 , n48940 );
and ( n18046 , C0 , RI1754c610_2);
or ( n48941 , n18045 , n18046 );
buf ( n48942 , n48941 );
not ( n48943 , n47771 );
and ( n48944 , n48943 , n43280 );
xor ( n48945 , n47768 , n48944 );
not ( n18047 , n29614 );
and ( n18048 , n18047 , RI1750fc38_717);
and ( n18049 , n48945 , n29614 );
or ( n48946 , n18048 , n18049 );
not ( n18050 , RI1754c610_2);
and ( n18051 , n18050 , n48946 );
and ( n18052 , C0 , RI1754c610_2);
or ( n48947 , n18051 , n18052 );
buf ( n48948 , n48947 );
xor ( n48949 , n41817 , n39262 );
xor ( n48950 , n48949 , n39282 );
xor ( n48951 , n40365 , n42554 );
xor ( n48952 , n48951 , n34725 );
not ( n48953 , n48952 );
xor ( n48954 , n33356 , n39005 );
xor ( n48955 , n48954 , n39543 );
and ( n48956 , n48953 , n48955 );
xor ( n48957 , n48950 , n48956 );
not ( n18053 , n29614 );
and ( n18054 , n18053 , RI173f8f08_1542);
and ( n18055 , n48957 , n29614 );
or ( n48958 , n18054 , n18055 );
not ( n18056 , RI1754c610_2);
and ( n18057 , n18056 , n48958 );
and ( n18058 , C0 , RI1754c610_2);
or ( n48959 , n18057 , n18058 );
buf ( n48960 , n48959 );
xor ( n48961 , n32413 , n35622 );
xor ( n48962 , n48961 , n35639 );
xor ( n48963 , n33709 , n35514 );
xor ( n48964 , n48963 , n40486 );
not ( n48965 , n48964 );
and ( n48966 , n48965 , n43621 );
xor ( n48967 , n48962 , n48966 );
not ( n18059 , n29614 );
and ( n18060 , n18059 , RI174486c0_1383);
and ( n18061 , n48967 , n29614 );
or ( n48968 , n18060 , n18061 );
not ( n18062 , RI1754c610_2);
and ( n18063 , n18062 , n48968 );
and ( n18064 , C0 , RI1754c610_2);
or ( n48969 , n18063 , n18064 );
buf ( n48970 , n48969 );
buf ( n48971 , RI174be6e0_818);
buf ( n48972 , RI17496f78_1000);
xor ( n48973 , n34742 , n42619 );
xor ( n48974 , n48973 , n41990 );
not ( n48975 , n48974 );
xor ( n48976 , n37097 , n37716 );
xor ( n48977 , n48976 , n37744 );
and ( n48978 , n48975 , n48977 );
xor ( n48979 , n41320 , n48978 );
not ( n18065 , n29614 );
and ( n18066 , n18065 , RI174bfb80_814);
and ( n18067 , n48979 , n29614 );
or ( n48980 , n18066 , n18067 );
not ( n18068 , RI1754c610_2);
and ( n18069 , n18068 , n48980 );
and ( n18070 , C0 , RI1754c610_2);
or ( n48981 , n18069 , n18070 );
buf ( n48982 , n48981 );
buf ( n48983 , RI174737d0_1173);
not ( n48984 , n33176 );
xor ( n48985 , n38792 , n40516 );
xor ( n48986 , n48985 , n40966 );
and ( n48987 , n48984 , n48986 );
xor ( n48988 , n33070 , n48987 );
not ( n18071 , n29614 );
and ( n18072 , n18071 , RI175110d8_713);
and ( n18073 , n48988 , n29614 );
or ( n48989 , n18072 , n18073 );
not ( n18074 , RI1754c610_2);
and ( n18075 , n18074 , n48989 );
and ( n18076 , C0 , RI1754c610_2);
or ( n48990 , n18075 , n18076 );
buf ( n48991 , n48990 );
not ( n48992 , n44739 );
and ( n48993 , n48992 , n35129 );
xor ( n48994 , n46235 , n48993 );
not ( n18077 , n29614 );
and ( n18078 , n18077 , RI173a5ac0_1948);
and ( n18079 , n48994 , n29614 );
or ( n48995 , n18078 , n18079 );
not ( n18080 , RI1754c610_2);
and ( n18081 , n18080 , n48995 );
and ( n18082 , C0 , RI1754c610_2);
or ( n48996 , n18081 , n18082 );
buf ( n48997 , n48996 );
not ( n48998 , n48582 );
and ( n48999 , n48998 , n48584 );
xor ( n49000 , n44879 , n48999 );
not ( n18083 , n29614 );
and ( n18084 , n18083 , RI173b3d28_1879);
and ( n18085 , n49000 , n29614 );
or ( n49001 , n18084 , n18085 );
not ( n18086 , RI1754c610_2);
and ( n18087 , n18086 , n49001 );
and ( n18088 , C0 , RI1754c610_2);
or ( n49002 , n18087 , n18088 );
buf ( n49003 , n49002 );
not ( n18089 , n27683 );
and ( n18090 , n18089 , RI19ac69e0_2280);
and ( n18091 , RI19acf428_2216 , n27683 );
or ( n49004 , n18090 , n18091 );
not ( n18092 , RI1754c610_2);
and ( n18093 , n18092 , n49004 );
and ( n18094 , C0 , RI1754c610_2);
or ( n49005 , n18093 , n18094 );
buf ( n49006 , n49005 );
not ( n18095 , n27683 );
and ( n18096 , n18095 , RI19ac30b0_2306);
and ( n18097 , RI19acc020_2239 , n27683 );
or ( n49007 , n18096 , n18097 );
not ( n18098 , RI1754c610_2);
and ( n18099 , n18098 , n49007 );
and ( n18100 , C0 , RI1754c610_2);
or ( n49008 , n18099 , n18100 );
buf ( n49009 , n49008 );
not ( n18101 , n27683 );
and ( n18102 , n18101 , RI19abcbe8_2361);
and ( n18103 , RI19ac5540_2289 , n27683 );
or ( n49010 , n18102 , n18103 );
not ( n18104 , RI1754c610_2);
and ( n18105 , n18104 , n49010 );
and ( n18106 , C0 , RI1754c610_2);
or ( n49011 , n18105 , n18106 );
buf ( n49012 , n49011 );
not ( n49013 , n45182 );
and ( n49014 , n49013 , n45184 );
xor ( n49015 , n44100 , n49014 );
not ( n18107 , n29614 );
and ( n18108 , n18107 , RI17404d58_1484);
and ( n18109 , n49015 , n29614 );
or ( n49016 , n18108 , n18109 );
not ( n18110 , RI1754c610_2);
and ( n18111 , n18110 , n49016 );
and ( n18112 , C0 , RI1754c610_2);
or ( n49017 , n18111 , n18112 );
buf ( n49018 , n49017 );
not ( n49019 , n47050 );
xor ( n49020 , n38808 , n39621 );
xor ( n49021 , n49020 , n40855 );
and ( n49022 , n49019 , n49021 );
xor ( n49023 , n41436 , n49022 );
not ( n18113 , n29614 );
and ( n18114 , n18113 , RI173437f8_2112);
and ( n18115 , n49023 , n29614 );
or ( n49024 , n18114 , n18115 );
not ( n18116 , RI1754c610_2);
and ( n18117 , n18116 , n49024 );
and ( n18118 , C0 , RI1754c610_2);
or ( n49025 , n18117 , n18118 );
buf ( n49026 , n49025 );
xor ( n49027 , n35199 , n43492 );
xor ( n49028 , n49027 , n38634 );
not ( n49029 , n47778 );
and ( n49030 , n49029 , n47780 );
xor ( n49031 , n49028 , n49030 );
not ( n18119 , n29614 );
and ( n18120 , n18119 , RI174816f0_1105);
and ( n18121 , n49031 , n29614 );
or ( n49032 , n18120 , n18121 );
not ( n18122 , RI1754c610_2);
and ( n18123 , n18122 , n49032 );
and ( n18124 , C0 , RI1754c610_2);
or ( n49033 , n18123 , n18124 );
buf ( n49034 , n49033 );
not ( n49035 , n48916 );
xor ( n49036 , n38972 , n41590 );
xor ( n49037 , n49036 , n35804 );
and ( n49038 , n49035 , n49037 );
xor ( n49039 , n48913 , n49038 );
not ( n18125 , n29614 );
and ( n18126 , n18125 , RI17408520_1467);
and ( n18127 , n49039 , n29614 );
or ( n49040 , n18126 , n18127 );
not ( n18128 , RI1754c610_2);
and ( n18129 , n18128 , n49040 );
and ( n18130 , C0 , RI1754c610_2);
or ( n49041 , n18129 , n18130 );
buf ( n49042 , n49041 );
not ( n49043 , n43650 );
and ( n49044 , n49043 , n43652 );
xor ( n49045 , n46071 , n49044 );
not ( n18131 , n29614 );
and ( n18132 , n18131 , RI174bf658_815);
and ( n18133 , n49045 , n29614 );
or ( n49046 , n18132 , n18133 );
not ( n18134 , RI1754c610_2);
and ( n18135 , n18134 , n49046 );
and ( n18136 , C0 , RI1754c610_2);
or ( n49047 , n18135 , n18136 );
buf ( n49048 , n49047 );
not ( n18137 , n27683 );
and ( n18138 , n18137 , RI19a99698_2616);
and ( n18139 , RI19aa3058_2545 , n27683 );
or ( n49049 , n18138 , n18139 );
not ( n18140 , RI1754c610_2);
and ( n18141 , n18140 , n49049 );
and ( n18142 , C0 , RI1754c610_2);
or ( n49050 , n18141 , n18142 );
buf ( n49051 , n49050 );
xor ( n49052 , n41783 , n35955 );
xor ( n49053 , n49052 , n42554 );
not ( n49054 , n43207 );
and ( n49055 , n49054 , n43209 );
xor ( n49056 , n49053 , n49055 );
not ( n18143 , n29614 );
and ( n18144 , n18143 , RI17465bf8_1240);
and ( n18145 , n49056 , n29614 );
or ( n49057 , n18144 , n18145 );
not ( n18146 , RI1754c610_2);
and ( n18147 , n18146 , n49057 );
and ( n18148 , C0 , RI1754c610_2);
or ( n49058 , n18147 , n18148 );
buf ( n49059 , n49058 );
not ( n18149 , n27683 );
and ( n18150 , n18149 , RI19ab0a50_2449);
and ( n18151 , RI19aba8c0_2377 , n27683 );
or ( n49060 , n18150 , n18151 );
not ( n18152 , RI1754c610_2);
and ( n18153 , n18152 , n49060 );
and ( n18154 , C0 , RI1754c610_2);
or ( n49061 , n18153 , n18154 );
buf ( n49062 , n49061 );
buf ( n49063 , RI174aa0a0_907);
xor ( n49064 , n39323 , n35416 );
xor ( n49065 , n49064 , n29843 );
xor ( n49066 , n40572 , n37048 );
xor ( n49067 , n49066 , n36772 );
not ( n49068 , n49067 );
xor ( n49069 , n34508 , n31380 );
xor ( n49070 , n49069 , n36463 );
and ( n49071 , n49068 , n49070 );
xor ( n49072 , n49065 , n49071 );
not ( n18155 , n29614 );
and ( n18156 , n18155 , RI173d1278_1736);
and ( n18157 , n49072 , n29614 );
or ( n49073 , n18156 , n18157 );
not ( n18158 , RI1754c610_2);
and ( n18159 , n18158 , n49073 );
and ( n18160 , C0 , RI1754c610_2);
or ( n49074 , n18159 , n18160 );
buf ( n49075 , n49074 );
buf ( n49076 , RI174a9380_911);
xor ( n49077 , n34137 , n33069 );
xor ( n49078 , n49077 , n42264 );
xor ( n49079 , n37808 , n31213 );
xor ( n49080 , n49079 , n31317 );
not ( n49081 , n49080 );
and ( n49082 , n49081 , n43584 );
xor ( n49083 , n49078 , n49082 );
not ( n18161 , n29614 );
and ( n18162 , n18161 , RI173950f8_2029);
and ( n18163 , n49083 , n29614 );
or ( n49084 , n18162 , n18163 );
not ( n18164 , RI1754c610_2);
and ( n18165 , n18164 , n49084 );
and ( n18166 , C0 , RI1754c610_2);
or ( n49085 , n18165 , n18166 );
buf ( n49086 , n49085 );
not ( n18167 , n27683 );
and ( n18168 , n18167 , RI19a919e8_2671);
and ( n18169 , RI19a9bd80_2599 , n27683 );
or ( n49087 , n18168 , n18169 );
not ( n18170 , RI1754c610_2);
and ( n18171 , n18170 , n49087 );
and ( n18172 , C0 , RI1754c610_2);
or ( n49088 , n18171 , n18172 );
buf ( n49089 , n49088 );
not ( n18173 , n27683 );
and ( n18174 , n18173 , RI19a9ce60_2591);
and ( n18175 , RI19aa6640_2520 , n27683 );
or ( n49090 , n18174 , n18175 );
not ( n18176 , RI1754c610_2);
and ( n18177 , n18176 , n49090 );
and ( n18178 , C0 , RI1754c610_2);
or ( n49091 , n18177 , n18178 );
buf ( n49092 , n49091 );
not ( n49093 , n47639 );
xor ( n49094 , n37743 , n41772 );
xor ( n49095 , n49094 , n32663 );
and ( n49096 , n49093 , n49095 );
xor ( n49097 , n47636 , n49096 );
not ( n18179 , n29614 );
and ( n18180 , n18179 , RI174d1208_760);
and ( n18181 , n49097 , n29614 );
or ( n49098 , n18180 , n18181 );
not ( n18182 , RI1754c610_2);
and ( n18183 , n18182 , n49098 );
and ( n18184 , C0 , RI1754c610_2);
or ( n49099 , n18183 , n18184 );
buf ( n49100 , n49099 );
not ( n49101 , n48643 );
and ( n49102 , n49101 , n36149 );
xor ( n49103 , n48640 , n49102 );
not ( n18185 , n29614 );
and ( n18186 , n18185 , RI17508078_741);
and ( n18187 , n49103 , n29614 );
or ( n49104 , n18186 , n18187 );
not ( n18188 , RI1754c610_2);
and ( n18189 , n18188 , n49104 );
and ( n18190 , C0 , RI1754c610_2);
or ( n49105 , n18189 , n18190 );
buf ( n49106 , n49105 );
not ( n18191 , n27683 );
and ( n18192 , n18191 , RI19acd5b0_2229);
and ( n18193 , RI19a8d230_2703 , n27683 );
or ( n49107 , n18192 , n18193 );
not ( n18194 , RI1754c610_2);
and ( n18195 , n18194 , n49107 );
and ( n18196 , C0 , RI1754c610_2);
or ( n49108 , n18195 , n18196 );
buf ( n49109 , n49108 );
not ( n18197 , n27683 );
and ( n18198 , n18197 , RI19ac9de8_2256);
and ( n18199 , RI19a85058_2759 , n27683 );
or ( n49110 , n18198 , n18199 );
not ( n18200 , RI1754c610_2);
and ( n18201 , n18200 , n49110 );
and ( n18202 , C0 , RI1754c610_2);
or ( n49111 , n18201 , n18202 );
buf ( n49112 , n49111 );
not ( n18203 , n27683 );
and ( n18204 , n18203 , RI19a8b4a8_2716);
and ( n18205 , RI19a95750_2644 , n27683 );
or ( n49113 , n18204 , n18205 );
not ( n18206 , RI1754c610_2);
and ( n18207 , n18206 , n49113 );
and ( n18208 , C0 , RI1754c610_2);
or ( n49114 , n18207 , n18208 );
buf ( n49115 , n49114 );
not ( n18209 , n27683 );
and ( n18210 , n18209 , RI19abd4d0_2356);
and ( n18211 , RI19ac5e28_2285 , n27683 );
or ( n49116 , n18210 , n18211 );
not ( n18212 , RI1754c610_2);
and ( n18213 , n18212 , n49116 );
and ( n18214 , C0 , RI1754c610_2);
or ( n49117 , n18213 , n18214 );
buf ( n49118 , n49117 );
xor ( n49119 , n39122 , n28111 );
xor ( n49120 , n49119 , n28468 );
not ( n49121 , n49120 );
and ( n49122 , n49121 , n44791 );
xor ( n49123 , n43468 , n49122 );
not ( n18215 , n29614 );
and ( n18216 , n18215 , RI174be6e0_818);
and ( n18217 , n49123 , n29614 );
or ( n49124 , n18216 , n18217 );
not ( n18218 , RI1754c610_2);
and ( n18219 , n18218 , n49124 );
and ( n18220 , C0 , RI1754c610_2);
or ( n49125 , n18219 , n18220 );
buf ( n49126 , n49125 );
not ( n49127 , n42866 );
and ( n49128 , n49127 , n46480 );
xor ( n49129 , n42754 , n49128 );
not ( n18221 , n29614 );
and ( n18222 , n18221 , RI174bf130_816);
and ( n18223 , n49129 , n29614 );
or ( n49130 , n18222 , n18223 );
not ( n18224 , RI1754c610_2);
and ( n18225 , n18224 , n49130 );
and ( n18226 , C0 , RI1754c610_2);
or ( n49131 , n18225 , n18226 );
buf ( n49132 , n49131 );
xor ( n49133 , n42308 , n40769 );
xor ( n49134 , n49133 , n40949 );
not ( n49135 , n32621 );
and ( n49136 , n49135 , n32716 );
xor ( n49137 , n49134 , n49136 );
not ( n18227 , n29614 );
and ( n18228 , n18227 , RI173379a8_2170);
and ( n18229 , n49137 , n29614 );
or ( n49138 , n18228 , n18229 );
not ( n18230 , RI1754c610_2);
and ( n18231 , n18230 , n49138 );
and ( n18232 , C0 , RI1754c610_2);
or ( n49139 , n18231 , n18232 );
buf ( n49140 , n49139 );
not ( n18233 , n27683 );
and ( n18234 , n18233 , RI19ac4b68_2294);
and ( n18235 , RI19acd808_2228 , n27683 );
or ( n49141 , n18234 , n18235 );
not ( n18236 , RI1754c610_2);
and ( n18237 , n18236 , n49141 );
and ( n18238 , C0 , RI1754c610_2);
or ( n49142 , n18237 , n18238 );
buf ( n49143 , n49142 );
xor ( n49144 , n39970 , n41934 );
xor ( n49145 , n49144 , n40341 );
xor ( n49146 , n41790 , n35955 );
xor ( n49147 , n49146 , n42554 );
not ( n49148 , n49147 );
xor ( n49149 , n29350 , n40034 );
xor ( n49150 , n49149 , n40051 );
and ( n49151 , n49148 , n49150 );
xor ( n49152 , n49145 , n49151 );
not ( n18239 , n29614 );
and ( n18240 , n18239 , RI174bec08_817);
and ( n18241 , n49152 , n29614 );
or ( n49153 , n18240 , n18241 );
not ( n18242 , RI1754c610_2);
and ( n18243 , n18242 , n49153 );
and ( n18244 , C0 , RI1754c610_2);
or ( n49154 , n18243 , n18244 );
buf ( n49155 , n49154 );
buf ( n49156 , RI17474ec8_1166);
not ( n18245 , n27683 );
and ( n18246 , n18245 , RI19a90a70_2678);
and ( n18247 , RI19a9aac0_2607 , n27683 );
or ( n49157 , n18246 , n18247 );
not ( n18248 , RI1754c610_2);
and ( n18249 , n18248 , n49157 );
and ( n18250 , C0 , RI1754c610_2);
or ( n49158 , n18249 , n18250 );
buf ( n49159 , n49158 );
and ( n49160 , RI1754af90_50 , n34844 );
and ( n49161 , RI1754af90_50 , n34847 );
buf ( n49162 , n34850 );
or ( n49163 , n49160 , n49161 , n49162 , C0 , C0 , C0 , C0 , C0 );
not ( n18251 , n34859 );
and ( n18252 , n18251 , n49163 );
and ( n18253 , RI1754af90_50 , n34859 );
or ( n49164 , n18252 , n18253 );
not ( n18254 , RI19a22f70_2797);
and ( n18255 , n18254 , n49164 );
and ( n18256 , C0 , RI19a22f70_2797);
or ( n49165 , n18255 , n18256 );
not ( n18257 , n27683 );
and ( n18258 , n18257 , RI19ac6878_2281);
and ( n18259 , n49165 , n27683 );
or ( n49166 , n18258 , n18259 );
not ( n18260 , RI1754c610_2);
and ( n18261 , n18260 , n49166 );
and ( n18262 , C0 , RI1754c610_2);
or ( n49167 , n18261 , n18262 );
buf ( n49168 , n49167 );
not ( n49169 , n47731 );
and ( n49170 , n49169 , n48770 );
xor ( n49171 , n39420 , n49170 );
not ( n18263 , n29614 );
and ( n18264 , n18263 , RI17489058_1068);
and ( n18265 , n49171 , n29614 );
or ( n49172 , n18264 , n18265 );
not ( n18266 , RI1754c610_2);
and ( n18267 , n18266 , n49172 );
and ( n18268 , C0 , RI1754c610_2);
or ( n49173 , n18267 , n18268 );
buf ( n49174 , n49173 );
not ( n18269 , n27683 );
and ( n18270 , n18269 , RI19aa7090_2516);
and ( n18271 , RI19ab11d0_2445 , n27683 );
or ( n49175 , n18270 , n18271 );
not ( n18272 , RI1754c610_2);
and ( n18273 , n18272 , n49175 );
and ( n18274 , C0 , RI1754c610_2);
or ( n49176 , n18273 , n18274 );
buf ( n49177 , n49176 );
buf ( n49178 , RI174c3e88_801);
buf ( n49179 , RI174937b0_1017);
buf ( n49180 , RI17479a40_1143);
not ( n49181 , n45488 );
xor ( n49182 , n35191 , n43492 );
xor ( n49183 , n49182 , n38634 );
and ( n49184 , n49181 , n49183 );
xor ( n49185 , n45485 , n49184 );
not ( n18275 , n29614 );
and ( n18276 , n18275 , RI173c1c48_1811);
and ( n18277 , n49185 , n29614 );
or ( n49186 , n18276 , n18277 );
not ( n18278 , RI1754c610_2);
and ( n18279 , n18278 , n49186 );
and ( n18280 , C0 , RI1754c610_2);
or ( n49187 , n18279 , n18280 );
buf ( n49188 , n49187 );
xor ( n49189 , n37695 , n37579 );
xor ( n49190 , n49189 , n38495 );
not ( n49191 , n46733 );
and ( n49192 , n49191 , n46735 );
xor ( n49193 , n49190 , n49192 );
not ( n18281 , n29614 );
and ( n18282 , n18281 , RI173ffe98_1508);
and ( n18283 , n49193 , n29614 );
or ( n49194 , n18282 , n18283 );
not ( n18284 , RI1754c610_2);
and ( n18285 , n18284 , n49194 );
and ( n18286 , C0 , RI1754c610_2);
or ( n49195 , n18285 , n18286 );
buf ( n49196 , n49195 );
not ( n18287 , n27683 );
and ( n18288 , n18287 , RI19ac5108_2291);
and ( n18289 , RI19acdcb8_2226 , n27683 );
or ( n49197 , n18288 , n18289 );
not ( n18290 , RI1754c610_2);
and ( n18291 , n18290 , n49197 );
and ( n18292 , C0 , RI1754c610_2);
or ( n49198 , n18291 , n18292 );
buf ( n49199 , n49198 );
xor ( n49200 , n35626 , n34669 );
xor ( n49201 , n49200 , n31831 );
not ( n49202 , n49201 );
and ( n49203 , n49202 , n48429 );
xor ( n49204 , n46202 , n49203 );
not ( n18293 , n29614 );
and ( n18294 , n18293 , RI17535ca8_599);
and ( n18295 , n49204 , n29614 );
or ( n49205 , n18294 , n18295 );
not ( n18296 , RI1754c610_2);
and ( n18297 , n18296 , n49205 );
and ( n18298 , C0 , RI1754c610_2);
or ( n49206 , n18297 , n18298 );
buf ( n49207 , n49206 );
not ( n49208 , n44164 );
xor ( n49209 , n35699 , n39543 );
xor ( n49210 , n49209 , n39563 );
and ( n49211 , n49208 , n49210 );
xor ( n49212 , n44161 , n49211 );
not ( n18299 , n29614 );
and ( n18300 , n18299 , RI17453b38_1328);
and ( n18301 , n49212 , n29614 );
or ( n49213 , n18300 , n18301 );
not ( n18302 , RI1754c610_2);
and ( n18303 , n18302 , n49213 );
and ( n18304 , C0 , RI1754c610_2);
or ( n49214 , n18303 , n18304 );
buf ( n49215 , n49214 );
xor ( n49216 , n41681 , n41885 );
xor ( n49217 , n49216 , n30923 );
not ( n49218 , n48168 );
and ( n49219 , n49218 , n48170 );
xor ( n49220 , n49217 , n49219 );
not ( n18305 , n29614 );
and ( n18306 , n18305 , RI1750cdd0_726);
and ( n18307 , n49220 , n29614 );
or ( n49221 , n18306 , n18307 );
not ( n18308 , RI1754c610_2);
and ( n18309 , n18308 , n49221 );
and ( n18310 , C0 , RI1754c610_2);
or ( n49222 , n18309 , n18310 );
buf ( n49223 , n49222 );
not ( n18311 , n27683 );
and ( n18312 , n18311 , RI19a82b50_2775);
and ( n18313 , RI19aaf448_2459 , n27683 );
or ( n49224 , n18312 , n18313 );
not ( n18314 , RI1754c610_2);
and ( n18315 , n18314 , n49224 );
and ( n18316 , C0 , RI1754c610_2);
or ( n49225 , n18315 , n18316 );
buf ( n49226 , n49225 );
not ( n49227 , n43237 );
and ( n49228 , n49227 , n43239 );
xor ( n49229 , n45269 , n49228 );
not ( n18317 , n29614 );
and ( n18318 , n18317 , RI1747b7c8_1134);
and ( n18319 , n49229 , n29614 );
or ( n49230 , n18318 , n18319 );
not ( n18320 , RI1754c610_2);
and ( n18321 , n18320 , n49230 );
and ( n18322 , C0 , RI1754c610_2);
or ( n49231 , n18321 , n18322 );
buf ( n49232 , n49231 );
xor ( n49233 , n38871 , n41125 );
xor ( n49234 , n49233 , n31506 );
not ( n49235 , n49234 );
xor ( n49236 , n33417 , n36252 );
xor ( n49237 , n49236 , n40360 );
and ( n49238 , n49235 , n49237 );
xor ( n49239 , n46432 , n49238 );
not ( n18323 , n29614 );
and ( n18324 , n18323 , RI173b2630_1886);
and ( n18325 , n49239 , n29614 );
or ( n49240 , n18324 , n18325 );
not ( n18326 , RI1754c610_2);
and ( n18327 , n18326 , n49240 );
and ( n18328 , C0 , RI1754c610_2);
or ( n49241 , n18327 , n18328 );
buf ( n49242 , n49241 );
not ( n18329 , n27683 );
and ( n18330 , n18329 , RI19acbc60_2241);
and ( n18331 , RI19a876c8_2742 , n27683 );
or ( n49243 , n18330 , n18331 );
not ( n18332 , RI1754c610_2);
and ( n18333 , n18332 , n49243 );
and ( n18334 , C0 , RI1754c610_2);
or ( n49244 , n18333 , n18334 );
buf ( n49245 , n49244 );
not ( n18335 , n27683 );
and ( n18336 , n18335 , RI19ac7f70_2270);
and ( n18337 , RI19a82d30_2774 , n27683 );
or ( n49246 , n18336 , n18337 );
not ( n18338 , RI1754c610_2);
and ( n18339 , n18338 , n49246 );
and ( n18340 , C0 , RI1754c610_2);
or ( n49247 , n18339 , n18340 );
buf ( n49248 , n49247 );
buf ( n49249 , RI174b5ba8_850);
not ( n18341 , n27683 );
and ( n18342 , n18341 , RI19aa3ee0_2538);
and ( n18343 , RI19aae458_2466 , n27683 );
or ( n49250 , n18342 , n18343 );
not ( n18344 , RI1754c610_2);
and ( n18345 , n18344 , n49250 );
and ( n18346 , C0 , RI1754c610_2);
or ( n49251 , n18345 , n18346 );
buf ( n49252 , n49251 );
buf ( n49253 , RI1749d530_969);
not ( n49254 , n41320 );
and ( n49255 , n49254 , n48974 );
xor ( n49256 , n41317 , n49255 );
not ( n18347 , n29614 );
and ( n18348 , n18347 , RI174ae8d0_885);
and ( n18349 , n49256 , n29614 );
or ( n49257 , n18348 , n18349 );
not ( n18350 , RI1754c610_2);
and ( n18351 , n18350 , n49257 );
and ( n18352 , C0 , RI1754c610_2);
or ( n49258 , n18351 , n18352 );
buf ( n49259 , n49258 );
not ( n49260 , n42655 );
and ( n49261 , n49260 , n40464 );
xor ( n49262 , n47873 , n49261 );
not ( n18353 , n29614 );
and ( n18354 , n18353 , RI173e39c8_1646);
and ( n18355 , n49262 , n29614 );
or ( n49263 , n18354 , n18355 );
not ( n18356 , RI1754c610_2);
and ( n18357 , n18356 , n49263 );
and ( n18358 , C0 , RI1754c610_2);
or ( n49264 , n18357 , n18358 );
buf ( n49265 , n49264 );
not ( n49266 , n47906 );
and ( n49267 , n49266 , n47908 );
xor ( n49268 , n47024 , n49267 );
not ( n18359 , n29614 );
and ( n18360 , n18359 , RI1744df58_1356);
and ( n18361 , n49268 , n29614 );
or ( n49269 , n18360 , n18361 );
not ( n18362 , RI1754c610_2);
and ( n18363 , n18362 , n49269 );
and ( n18364 , C0 , RI1754c610_2);
or ( n49270 , n18363 , n18364 );
buf ( n49271 , n49270 );
xor ( n49272 , n38978 , n41590 );
xor ( n49273 , n49272 , n35804 );
not ( n49274 , n49273 );
and ( n49275 , n49274 , n44779 );
xor ( n49276 , n48779 , n49275 );
not ( n18365 , n29614 );
and ( n18366 , n18365 , RI174bbda0_826);
and ( n18367 , n49276 , n29614 );
or ( n49277 , n18366 , n18367 );
not ( n18368 , RI1754c610_2);
and ( n18369 , n18368 , n49277 );
and ( n18370 , C0 , RI1754c610_2);
or ( n49278 , n18369 , n18370 );
buf ( n49279 , n49278 );
not ( n49280 , n48006 );
and ( n49281 , n49280 , n43079 );
xor ( n49282 , n41345 , n49281 );
not ( n18371 , n29614 );
and ( n18372 , n18371 , RI17334870_2185);
and ( n18373 , n49282 , n29614 );
or ( n49283 , n18372 , n18373 );
not ( n18374 , RI1754c610_2);
and ( n18375 , n18374 , n49283 );
and ( n18376 , C0 , RI1754c610_2);
or ( n49284 , n18375 , n18376 );
buf ( n49285 , n49284 );
buf ( n49286 , RI1747df28_1122);
buf ( n49287 , RI17465bf8_1240);
not ( n18377 , n27683 );
and ( n18378 , n18377 , RI19a843b0_2764);
and ( n18379 , RI19abe2e0_2348 , n27683 );
or ( n49288 , n18378 , n18379 );
not ( n18380 , RI1754c610_2);
and ( n18381 , n18380 , n49288 );
and ( n18382 , C0 , RI1754c610_2);
or ( n49289 , n18381 , n18382 );
buf ( n49290 , n49289 );
xor ( n49291 , n36909 , n32560 );
xor ( n49292 , n49291 , n32620 );
xor ( n49293 , n41239 , n38634 );
xor ( n49294 , n49293 , n38648 );
not ( n49295 , n49294 );
xor ( n49296 , n32714 , n36209 );
xor ( n49297 , n49296 , n40412 );
and ( n49298 , n49295 , n49297 );
xor ( n49299 , n49292 , n49298 );
not ( n18383 , n29614 );
and ( n18384 , n18383 , RI173a4710_1954);
and ( n18385 , n49299 , n29614 );
or ( n49300 , n18384 , n18385 );
not ( n18386 , RI1754c610_2);
and ( n18387 , n18386 , n49300 );
and ( n18388 , C0 , RI1754c610_2);
or ( n49301 , n18387 , n18388 );
buf ( n49302 , n49301 );
and ( n49303 , RI1754bda0_20 , n34844 );
and ( n49304 , RI1754bda0_20 , n34847 );
and ( n49305 , RI1754bda0_20 , n34850 );
and ( n49306 , RI1754bda0_20 , n34852 );
and ( n49307 , RI1754bda0_20 , n34854 );
or ( n49308 , n49303 , n49304 , n49305 , n49306 , n49307 , C0 , C0 , C0 );
not ( n18389 , n34859 );
and ( n18390 , n18389 , n49308 );
and ( n18391 , RI1754bda0_20 , n34859 );
or ( n49309 , n18390 , n18391 );
not ( n18392 , RI19a22f70_2797);
and ( n18393 , n18392 , n49309 );
and ( n18394 , C0 , RI19a22f70_2797);
or ( n49310 , n18393 , n18394 );
not ( n18395 , n27683 );
and ( n18396 , n18395 , RI19a99ad0_2614);
and ( n18397 , n49310 , n27683 );
or ( n49311 , n18396 , n18397 );
not ( n18398 , RI1754c610_2);
and ( n18399 , n18398 , n49311 );
and ( n18400 , C0 , RI1754c610_2);
or ( n49312 , n18399 , n18400 );
buf ( n49313 , n49312 );
not ( n18401 , n27683 );
and ( n18402 , n18401 , RI19a92bb8_2663);
and ( n18403 , RI19a9ce60_2591 , n27683 );
or ( n49314 , n18402 , n18403 );
not ( n18404 , RI1754c610_2);
and ( n18405 , n18404 , n49314 );
and ( n18406 , C0 , RI1754c610_2);
or ( n49315 , n18405 , n18406 );
buf ( n49316 , n49315 );
not ( n49317 , n44389 );
and ( n49318 , n49317 , n44391 );
xor ( n49319 , n45765 , n49318 );
not ( n18407 , n29614 );
and ( n18408 , n18407 , RI175212a8_663);
and ( n18409 , n49319 , n29614 );
or ( n49320 , n18408 , n18409 );
not ( n18410 , RI1754c610_2);
and ( n18411 , n18410 , n49320 );
and ( n18412 , C0 , RI1754c610_2);
or ( n49321 , n18411 , n18412 );
buf ( n49322 , n49321 );
not ( n49323 , n34042 );
and ( n49324 , n49323 , n39622 );
xor ( n49325 , n33936 , n49324 );
not ( n18413 , n29614 );
and ( n18414 , n18413 , RI1749c180_975);
and ( n18415 , n49325 , n29614 );
or ( n49326 , n18414 , n18415 );
not ( n18416 , RI1754c610_2);
and ( n18417 , n18416 , n49326 );
and ( n18418 , C0 , RI1754c610_2);
or ( n49327 , n18417 , n18418 );
buf ( n49328 , n49327 );
not ( n18419 , n27683 );
and ( n18420 , n18419 , RI19ac1b98_2316);
and ( n18421 , RI19acb120_2247 , n27683 );
or ( n49329 , n18420 , n18421 );
not ( n18422 , RI1754c610_2);
and ( n18423 , n18422 , n49329 );
and ( n18424 , C0 , RI1754c610_2);
or ( n49330 , n18423 , n18424 );
buf ( n49331 , n49330 );
not ( n49332 , n41773 );
and ( n49333 , n49332 , n42922 );
xor ( n49334 , n41754 , n49333 );
not ( n18425 , n29614 );
and ( n18426 , n18425 , RI174ce8b0_768);
and ( n18427 , n49334 , n29614 );
or ( n49335 , n18426 , n18427 );
not ( n18428 , RI1754c610_2);
and ( n18429 , n18428 , n49335 );
and ( n18430 , C0 , RI1754c610_2);
or ( n49336 , n18429 , n18430 );
buf ( n49337 , n49336 );
not ( n49338 , n44988 );
xor ( n49339 , n35505 , n38532 );
xor ( n49340 , n49339 , n38933 );
and ( n49341 , n49338 , n49340 );
xor ( n49342 , n44985 , n49341 );
or ( n49343 , n31331 , RI17537fd0_593);
or ( n49344 , n49343 , RI175379b8_594);
or ( n49345 , n49344 , RI175373a0_595);
or ( n49346 , n49345 , RI17536d88_596);
or ( n49347 , n49346 , RI17536770_597);
or ( n49348 , n49347 , RI17539e48_588);
xor ( n49349 , n49342 , n49348 );
not ( n18431 , n29614 );
and ( n18432 , n18431 , RI174613c8_1262);
and ( n18433 , n49349 , n29614 );
or ( n49350 , n18432 , n18433 );
not ( n18434 , RI1754c610_2);
and ( n18435 , n18434 , n49350 );
and ( n18436 , C0 , RI1754c610_2);
or ( n49351 , n18435 , n18436 );
buf ( n49352 , n49351 );
buf ( n49353 , RI174bd240_822);
not ( n49354 , n42761 );
and ( n49355 , n49354 , n42763 );
xor ( n49356 , n42010 , n49355 );
not ( n18437 , n29614 );
and ( n18438 , n18437 , RI17487960_1075);
and ( n18439 , n49356 , n29614 );
or ( n49357 , n18438 , n18439 );
not ( n18440 , RI1754c610_2);
and ( n18441 , n18440 , n49357 );
and ( n18442 , C0 , RI1754c610_2);
or ( n49358 , n18441 , n18442 );
buf ( n49359 , n49358 );
buf ( n49360 , RI1749b118_980);
xor ( n49361 , n36499 , n40381 );
xor ( n49362 , n49361 , n37438 );
xor ( n49363 , n41650 , n40692 );
xor ( n49364 , n49363 , n43994 );
not ( n49365 , n49364 );
and ( n49366 , n49365 , n46887 );
xor ( n49367 , n49362 , n49366 );
not ( n18443 , n29614 );
and ( n18444 , n18443 , RI17451db0_1337);
and ( n18445 , n49367 , n29614 );
or ( n49368 , n18444 , n18445 );
not ( n18446 , RI1754c610_2);
and ( n18447 , n18446 , n49368 );
and ( n18448 , C0 , RI1754c610_2);
or ( n49369 , n18447 , n18448 );
buf ( n49370 , n49369 );
buf ( n49371 , RI1748a408_1062);
buf ( n49372 , RI17500f80_757);
not ( n18449 , n27683 );
and ( n18450 , n18449 , RI19aa2e78_2546);
and ( n18451 , RI19aad120_2475 , n27683 );
or ( n49373 , n18450 , n18451 );
not ( n18452 , RI1754c610_2);
and ( n18453 , n18452 , n49373 );
and ( n18454 , C0 , RI1754c610_2);
or ( n49374 , n18453 , n18454 );
buf ( n49375 , n49374 );
xor ( n49376 , n37152 , n40254 );
xor ( n49377 , n49376 , n40718 );
not ( n49378 , n46523 );
and ( n49379 , n49378 , n46525 );
xor ( n49380 , n49377 , n49379 );
not ( n18455 , n29614 );
and ( n18456 , n18455 , RI17475558_1164);
and ( n18457 , n49380 , n29614 );
or ( n49381 , n18456 , n18457 );
not ( n18458 , RI1754c610_2);
and ( n18459 , n18458 , n49381 );
and ( n18460 , C0 , RI1754c610_2);
or ( n49382 , n18459 , n18460 );
buf ( n49383 , n49382 );
not ( n18461 , n27683 );
and ( n18462 , n18461 , RI19a864f8_2750);
and ( n18463 , RI19a23150_2796 , n27683 );
or ( n49384 , n18462 , n18463 );
not ( n18464 , RI1754c610_2);
and ( n18465 , n18464 , n49384 );
and ( n18466 , C0 , RI1754c610_2);
or ( n49385 , n18465 , n18466 );
buf ( n49386 , n49385 );
not ( n49387 , n48353 );
and ( n49388 , n49387 , n42803 );
xor ( n49389 , n41564 , n49388 );
not ( n18467 , n29614 );
and ( n18468 , n18467 , RI173b74f0_1862);
and ( n18469 , n49389 , n29614 );
or ( n49390 , n18468 , n18469 );
not ( n18470 , RI1754c610_2);
and ( n18471 , n18470 , n49390 );
and ( n18472 , C0 , RI1754c610_2);
or ( n49391 , n18471 , n18472 );
buf ( n49392 , n49391 );
xor ( n49393 , n37593 , n40319 );
xor ( n49394 , n49393 , n40149 );
not ( n49395 , n44755 );
and ( n49396 , n49395 , n44757 );
xor ( n49397 , n49394 , n49396 );
not ( n18473 , n29614 );
and ( n18474 , n18473 , RI173cf820_1744);
and ( n18475 , n49397 , n29614 );
or ( n49398 , n18474 , n18475 );
not ( n18476 , RI1754c610_2);
and ( n18477 , n18476 , n49398 );
and ( n18478 , C0 , RI1754c610_2);
or ( n49399 , n18477 , n18478 );
buf ( n49400 , n49399 );
not ( n18479 , n27683 );
and ( n18480 , n18479 , RI19a9a868_2608);
and ( n18481 , RI19aa3ee0_2538 , n27683 );
or ( n49401 , n18480 , n18481 );
not ( n18482 , RI1754c610_2);
and ( n18483 , n18482 , n49401 );
and ( n18484 , C0 , RI1754c610_2);
or ( n49402 , n18483 , n18484 );
buf ( n49403 , n49402 );
not ( n18485 , n27683 );
and ( n18486 , n18485 , RI19a87218_2744);
and ( n18487 , RI19a94df0_2648 , n27683 );
or ( n49404 , n18486 , n18487 );
not ( n18488 , RI1754c610_2);
and ( n18489 , n18488 , n49404 );
and ( n18490 , C0 , RI1754c610_2);
or ( n49405 , n18489 , n18490 );
buf ( n49406 , n49405 );
not ( n49407 , n36875 );
xor ( n49408 , n38237 , n39450 );
xor ( n49409 , n49408 , n39467 );
and ( n49410 , n49407 , n49409 );
xor ( n49411 , n36803 , n49410 );
not ( n18491 , n29614 );
and ( n18492 , n18491 , RI1738f518_2057);
and ( n18493 , n49411 , n29614 );
or ( n49412 , n18492 , n18493 );
not ( n18494 , RI1754c610_2);
and ( n18495 , n18494 , n49412 );
and ( n18496 , C0 , RI1754c610_2);
or ( n49413 , n18495 , n18496 );
buf ( n49414 , n49413 );
not ( n49415 , n31926 );
and ( n49416 , n49415 , n42715 );
xor ( n49417 , n31726 , n49416 );
not ( n18497 , n29614 );
and ( n18498 , n18497 , RI173af4f8_1901);
and ( n18499 , n49417 , n29614 );
or ( n49418 , n18498 , n18499 );
not ( n18500 , RI1754c610_2);
and ( n18501 , n18500 , n49418 );
and ( n18502 , C0 , RI1754c610_2);
or ( n49419 , n18501 , n18502 );
buf ( n49420 , n49419 );
xor ( n49421 , n36276 , n37311 );
xor ( n49422 , n49421 , n37942 );
xor ( n49423 , n39058 , n39702 );
xor ( n49424 , n49423 , n39914 );
not ( n49425 , n49424 );
xor ( n49426 , n40807 , n40437 );
xor ( n49427 , n49426 , n42635 );
and ( n49428 , n49425 , n49427 );
xor ( n49429 , n49422 , n49428 );
not ( n18503 , n29614 );
and ( n18504 , n18503 , RI1748ade0_1059);
and ( n18505 , n49429 , n29614 );
or ( n49430 , n18504 , n18505 );
not ( n18506 , RI1754c610_2);
and ( n18507 , n18506 , n49430 );
and ( n18508 , C0 , RI1754c610_2);
or ( n49431 , n18507 , n18508 );
buf ( n49432 , n49431 );
not ( n49433 , n34476 );
and ( n49434 , n49433 , n39162 );
xor ( n49435 , n34446 , n49434 );
not ( n18509 , n29614 );
and ( n18510 , n18509 , RI1752ad58_633);
and ( n18511 , n49435 , n29614 );
or ( n49436 , n18510 , n18511 );
not ( n18512 , RI1754c610_2);
and ( n18513 , n18512 , n49436 );
and ( n18514 , C0 , RI1754c610_2);
or ( n49437 , n18513 , n18514 );
buf ( n49438 , n49437 );
not ( n49439 , n42925 );
and ( n49440 , n49439 , n41752 );
xor ( n49441 , n42922 , n49440 );
not ( n18515 , n29614 );
and ( n18516 , n18515 , RI1752d170_626);
and ( n18517 , n49441 , n29614 );
or ( n49442 , n18516 , n18517 );
not ( n18518 , RI1754c610_2);
and ( n18519 , n18518 , n49442 );
and ( n18520 , C0 , RI1754c610_2);
or ( n49443 , n18519 , n18520 );
buf ( n49444 , n49443 );
not ( n49445 , n48955 );
xor ( n49446 , n40846 , n35009 );
xor ( n49447 , n49446 , n28816 );
and ( n49448 , n49445 , n49447 );
xor ( n49449 , n48952 , n49448 );
not ( n18521 , n29614 );
and ( n18522 , n18521 , RI17412fc0_1415);
and ( n18523 , n49449 , n29614 );
or ( n49450 , n18522 , n18523 );
not ( n18524 , RI1754c610_2);
and ( n18525 , n18524 , n49450 );
and ( n18526 , C0 , RI1754c610_2);
or ( n49451 , n18525 , n18526 );
buf ( n49452 , n49451 );
xor ( n49453 , n41677 , n41885 );
xor ( n49454 , n49453 , n30923 );
xor ( n49455 , n33320 , n38991 );
xor ( n49456 , n49455 , n39005 );
not ( n49457 , n49456 );
and ( n49458 , n49457 , n42345 );
xor ( n49459 , n49454 , n49458 );
not ( n18527 , n29614 );
and ( n18528 , n18527 , RI173d4068_1722);
and ( n18529 , n49459 , n29614 );
or ( n49460 , n18528 , n18529 );
not ( n18530 , RI1754c610_2);
and ( n18531 , n18530 , n49460 );
and ( n18532 , C0 , RI1754c610_2);
or ( n49461 , n18531 , n18532 );
buf ( n49462 , n49461 );
xor ( n49463 , n34323 , n39604 );
xor ( n49464 , n49463 , n39621 );
not ( n49465 , n48112 );
and ( n49466 , n49465 , n48114 );
xor ( n49467 , n49464 , n49466 );
not ( n18533 , n29614 );
and ( n18534 , n18533 , RI173ed400_1599);
and ( n18535 , n49467 , n29614 );
or ( n49468 , n18534 , n18535 );
not ( n18536 , RI1754c610_2);
and ( n18537 , n18536 , n49468 );
and ( n18538 , C0 , RI1754c610_2);
or ( n49469 , n18537 , n18538 );
buf ( n49470 , n49469 );
not ( n49471 , n49150 );
xor ( n49472 , n39004 , n35804 );
xor ( n49473 , n49472 , n35842 );
and ( n49474 , n49471 , n49473 );
xor ( n49475 , n49147 , n49474 );
not ( n18539 , n29614 );
and ( n18540 , n18539 , RI17506188_747);
and ( n18541 , n49475 , n29614 );
or ( n49476 , n18540 , n18541 );
not ( n18542 , RI1754c610_2);
and ( n18543 , n18542 , n49476 );
and ( n18544 , C0 , RI1754c610_2);
or ( n49477 , n18543 , n18544 );
buf ( n49478 , n49477 );
not ( n18545 , n27683 );
and ( n18546 , n18545 , RI19a97b68_2628);
and ( n18547 , RI19aa1618_2557 , n27683 );
or ( n49479 , n18546 , n18547 );
not ( n18548 , RI1754c610_2);
and ( n18549 , n18548 , n49479 );
and ( n18550 , C0 , RI1754c610_2);
or ( n49480 , n18549 , n18550 );
buf ( n49481 , n49480 );
not ( n49482 , n42997 );
and ( n49483 , n49482 , n46350 );
xor ( n49484 , n42994 , n49483 );
not ( n18551 , n29614 );
and ( n18552 , n18551 , RI17465f40_1239);
and ( n18553 , n49484 , n29614 );
or ( n49485 , n18552 , n18553 );
not ( n18554 , RI1754c610_2);
and ( n18555 , n18554 , n49485 );
and ( n18556 , C0 , RI1754c610_2);
or ( n49486 , n18555 , n18556 );
buf ( n49487 , n49486 );
not ( n18557 , n27683 );
and ( n18558 , n18557 , RI19ab5118_2416);
and ( n18559 , RI19abe808_2345 , n27683 );
or ( n49488 , n18558 , n18559 );
not ( n18560 , RI1754c610_2);
and ( n18561 , n18560 , n49488 );
and ( n18562 , C0 , RI1754c610_2);
or ( n49489 , n18561 , n18562 );
buf ( n49490 , n49489 );
xor ( n49491 , n29879 , n36128 );
xor ( n49492 , n49491 , n36148 );
xor ( n49493 , n41495 , n34445 );
xor ( n49494 , n49493 , n41885 );
not ( n49495 , n49494 );
xor ( n49496 , n38262 , n36530 );
xor ( n49497 , n49496 , n36568 );
and ( n49498 , n49495 , n49497 );
xor ( n49499 , n49492 , n49498 );
not ( n18563 , n29614 );
and ( n18564 , n18563 , RI1738d790_2066);
and ( n18565 , n49499 , n29614 );
or ( n49500 , n18564 , n18565 );
not ( n18566 , RI1754c610_2);
and ( n18567 , n18566 , n49500 );
and ( n18568 , C0 , RI1754c610_2);
or ( n49501 , n18567 , n18568 );
buf ( n49502 , n49501 );
not ( n49503 , n49297 );
xor ( n49504 , n32812 , n37203 );
xor ( n49505 , n49504 , n34150 );
and ( n49506 , n49503 , n49505 );
xor ( n49507 , n49294 , n49506 );
not ( n18569 , n29614 );
and ( n18570 , n18569 , RI173b3008_1883);
and ( n18571 , n49507 , n29614 );
or ( n49508 , n18570 , n18571 );
not ( n18572 , RI1754c610_2);
and ( n18573 , n18572 , n49508 );
and ( n18574 , C0 , RI1754c610_2);
or ( n49509 , n18573 , n18574 );
buf ( n49510 , n49509 );
xor ( n49511 , n35531 , n37460 );
xor ( n49512 , n49511 , n37490 );
xor ( n49513 , n34145 , n33069 );
xor ( n49514 , n49513 , n42264 );
not ( n49515 , n49514 );
xor ( n49516 , n39449 , n38495 );
xor ( n49517 , n49516 , n36611 );
and ( n49518 , n49515 , n49517 );
xor ( n49519 , n49512 , n49518 );
not ( n18575 , n29614 );
and ( n18576 , n18575 , RI173ea610_1613);
and ( n18577 , n49519 , n29614 );
or ( n49520 , n18576 , n18577 );
not ( n18578 , RI1754c610_2);
and ( n18579 , n18578 , n49520 );
and ( n18580 , C0 , RI1754c610_2);
or ( n49521 , n18579 , n18580 );
buf ( n49522 , n49521 );
xor ( n49523 , n40133 , n38948 );
xor ( n49524 , n49523 , n39039 );
not ( n49525 , n49524 );
xor ( n49526 , n36077 , n37371 );
xor ( n49527 , n49526 , n36682 );
and ( n49528 , n49525 , n49527 );
xor ( n49529 , n41745 , n49528 );
not ( n18581 , n29614 );
and ( n18582 , n18581 , RI1749dbc0_967);
and ( n18583 , n49529 , n29614 );
or ( n49530 , n18582 , n18583 );
not ( n18584 , RI1754c610_2);
and ( n18585 , n18584 , n49530 );
and ( n18586 , C0 , RI1754c610_2);
or ( n49531 , n18585 , n18586 );
buf ( n49532 , n49531 );
not ( n49533 , n44437 );
and ( n49534 , n49533 , n46439 );
xor ( n49535 , n44434 , n49534 );
not ( n18587 , n29614 );
and ( n18588 , n18587 , RI174a4808_934);
and ( n18589 , n49535 , n29614 );
or ( n49536 , n18588 , n18589 );
not ( n18590 , RI1754c610_2);
and ( n18591 , n18590 , n49536 );
and ( n18592 , C0 , RI1754c610_2);
or ( n49537 , n18591 , n18592 );
buf ( n49538 , n49537 );
not ( n18593 , n27683 );
and ( n18594 , n18593 , RI19aa5560_2527);
and ( n18595 , RI19aafad8_2456 , n27683 );
or ( n49539 , n18594 , n18595 );
not ( n18596 , RI1754c610_2);
and ( n18597 , n18596 , n49539 );
and ( n18598 , C0 , RI1754c610_2);
or ( n49540 , n18597 , n18598 );
buf ( n49541 , n49540 );
not ( n18599 , n27683 );
and ( n18600 , n18599 , RI19aad468_2473);
and ( n18601 , RI19ab71e8_2401 , n27683 );
or ( n49542 , n18600 , n18601 );
not ( n18602 , RI1754c610_2);
and ( n18603 , n18602 , n49542 );
and ( n18604 , C0 , RI1754c610_2);
or ( n49543 , n18603 , n18604 );
buf ( n49544 , n49543 );
not ( n18605 , n27683 );
and ( n18606 , n18605 , RI19acd100_2231);
and ( n18607 , RI19a89e28_2725 , n27683 );
or ( n49545 , n18606 , n18607 );
not ( n18608 , RI1754c610_2);
and ( n18609 , n18608 , n49545 );
and ( n18610 , C0 , RI1754c610_2);
or ( n49546 , n18609 , n18610 );
buf ( n49547 , n49546 );
xor ( n49548 , n40418 , n39816 );
xor ( n49549 , n49548 , n35052 );
xor ( n49550 , n40842 , n35009 );
xor ( n49551 , n49550 , n28816 );
not ( n49552 , n49551 );
xor ( n49553 , n41421 , n43464 );
xor ( n49554 , n49553 , n44146 );
and ( n49555 , n49552 , n49554 );
xor ( n49556 , n49549 , n49555 );
not ( n18611 , n29614 );
and ( n18612 , n18611 , RI174b3790_861);
and ( n18613 , n49556 , n29614 );
or ( n49557 , n18612 , n18613 );
not ( n18614 , RI1754c610_2);
and ( n18615 , n18614 , n49557 );
and ( n18616 , C0 , RI1754c610_2);
or ( n49558 , n18615 , n18616 );
buf ( n49559 , n49558 );
xor ( n49560 , n34774 , n37255 );
xor ( n49561 , n49560 , n41478 );
xor ( n49562 , n37322 , n39914 );
xor ( n49563 , n49562 , n40237 );
not ( n49564 , n49563 );
xor ( n49565 , n39633 , n35176 );
xor ( n49566 , n49565 , n35216 );
and ( n49567 , n49564 , n49566 );
xor ( n49568 , n49561 , n49567 );
not ( n18617 , n29614 );
and ( n18618 , n18617 , RI174bc2c8_825);
and ( n18619 , n49568 , n29614 );
or ( n49569 , n18618 , n18619 );
not ( n18620 , RI1754c610_2);
and ( n18621 , n18620 , n49569 );
and ( n18622 , C0 , RI1754c610_2);
or ( n49570 , n18621 , n18622 );
buf ( n49571 , n49570 );
xor ( n49572 , n33807 , n39414 );
xor ( n49573 , n49572 , n37186 );
xor ( n49574 , n37547 , n34918 );
xor ( n49575 , n49574 , n34968 );
not ( n49576 , n49575 );
xor ( n49577 , n35954 , n36148 );
xor ( n49578 , n49577 , n37421 );
and ( n49579 , n49576 , n49578 );
xor ( n49580 , n49573 , n49579 );
not ( n18623 , n29614 );
and ( n18624 , n18623 , RI1747f968_1114);
and ( n18625 , n49580 , n29614 );
or ( n49581 , n18624 , n18625 );
not ( n18626 , RI1754c610_2);
and ( n18627 , n18626 , n49581 );
and ( n18628 , C0 , RI1754c610_2);
or ( n49582 , n18627 , n18628 );
buf ( n49583 , n49582 );
xor ( n49584 , n37058 , n38594 );
xor ( n49585 , n49584 , n37716 );
not ( n49586 , n49585 );
xor ( n49587 , n37839 , n33697 );
xor ( n49588 , n49587 , n35128 );
and ( n49589 , n49586 , n49588 );
xor ( n49590 , n49517 , n49589 );
not ( n18629 , n29614 );
and ( n18630 , n18629 , RI17407800_1471);
and ( n18631 , n49590 , n29614 );
or ( n49591 , n18630 , n18631 );
not ( n18632 , RI1754c610_2);
and ( n18633 , n18632 , n49591 );
and ( n18634 , C0 , RI1754c610_2);
or ( n49592 , n18633 , n18634 );
buf ( n49593 , n49592 );
not ( n49594 , n42473 );
xor ( n49595 , n35161 , n37915 );
xor ( n49596 , n49595 , n43492 );
and ( n49597 , n49594 , n49596 );
xor ( n49598 , n42470 , n49597 );
not ( n18635 , n29614 );
and ( n18636 , n18635 , RI174b5ef0_849);
and ( n18637 , n49598 , n29614 );
or ( n49599 , n18636 , n18637 );
not ( n18638 , RI1754c610_2);
and ( n18639 , n18638 , n49599 );
and ( n18640 , C0 , RI1754c610_2);
or ( n49600 , n18639 , n18640 );
buf ( n49601 , n49600 );
not ( n49602 , n49210 );
xor ( n49603 , n30922 , n38115 );
xor ( n49604 , n49603 , n41622 );
and ( n49605 , n49602 , n49604 );
xor ( n49606 , n44164 , n49605 );
not ( n18641 , n29614 );
and ( n18642 , n18641 , RI1746e910_1197);
and ( n18643 , n49606 , n29614 );
or ( n49607 , n18642 , n18643 );
not ( n18644 , RI1754c610_2);
and ( n18645 , n18644 , n49607 );
and ( n18646 , C0 , RI1754c610_2);
or ( n49608 , n18645 , n18646 );
buf ( n49609 , n49608 );
not ( n18647 , n27683 );
and ( n18648 , n18647 , RI19acc020_2239);
and ( n18649 , RI19a87b78_2740 , n27683 );
or ( n49610 , n18648 , n18649 );
not ( n18650 , RI1754c610_2);
and ( n18651 , n18650 , n49610 );
and ( n18652 , C0 , RI1754c610_2);
or ( n49611 , n18651 , n18652 );
buf ( n49612 , n49611 );
buf ( n49613 , RI174abe28_898);
not ( n18653 , n27683 );
and ( n18654 , n18653 , RI19ac74a8_2275);
and ( n18655 , RI19acffe0_2211 , n27683 );
or ( n49614 , n18654 , n18655 );
not ( n18656 , RI1754c610_2);
and ( n18657 , n18656 , n49614 );
and ( n18658 , C0 , RI1754c610_2);
or ( n49615 , n18657 , n18658 );
buf ( n49616 , n49615 );
not ( n49617 , n44809 );
and ( n49618 , n49617 , n44811 );
xor ( n49619 , n38649 , n49618 );
not ( n18659 , n29614 );
and ( n18660 , n18659 , RI174a5870_929);
and ( n18661 , n49619 , n29614 );
or ( n49620 , n18660 , n18661 );
not ( n18662 , RI1754c610_2);
and ( n18663 , n18662 , n49620 );
and ( n18664 , C0 , RI1754c610_2);
or ( n49621 , n18663 , n18664 );
buf ( n49622 , n49621 );
not ( n18665 , n27683 );
and ( n18666 , n18665 , RI19aa3580_2542);
and ( n18667 , RI19aad828_2471 , n27683 );
or ( n49623 , n18666 , n18667 );
not ( n18668 , RI1754c610_2);
and ( n18669 , n18668 , n49623 );
and ( n18670 , C0 , RI1754c610_2);
or ( n49624 , n18669 , n18670 );
buf ( n49625 , n49624 );
buf ( n49626 , RI174a72b0_921);
buf ( n49627 , RI1747c1a0_1131);
not ( n49628 , n45672 );
xor ( n49629 , n37219 , n39467 );
xor ( n49630 , n49629 , n41391 );
and ( n49631 , n49628 , n49630 );
xor ( n49632 , n45669 , n49631 );
not ( n18671 , n29614 );
and ( n18672 , n18671 , RI173ae490_1906);
and ( n18673 , n49632 , n29614 );
or ( n49633 , n18672 , n18673 );
not ( n18674 , RI1754c610_2);
and ( n18675 , n18674 , n49633 );
and ( n18676 , C0 , RI1754c610_2);
or ( n49634 , n18675 , n18676 );
buf ( n49635 , n49634 );
xor ( n49636 , n33426 , n36252 );
xor ( n49637 , n49636 , n40360 );
not ( n49638 , n49637 );
xor ( n49639 , n41848 , n33282 );
xor ( n49640 , n49639 , n37623 );
and ( n49641 , n49638 , n49640 );
xor ( n49642 , n32482 , n49641 );
not ( n18677 , n29614 );
and ( n18678 , n18677 , RI173462a0_2099);
and ( n18679 , n49642 , n29614 );
or ( n49643 , n18678 , n18679 );
not ( n18680 , RI1754c610_2);
and ( n18681 , n18680 , n49643 );
and ( n18682 , C0 , RI1754c610_2);
or ( n49644 , n18681 , n18682 );
buf ( n49645 , n49644 );
not ( n49646 , n41705 );
and ( n49647 , n49646 , n45154 );
xor ( n49648 , n41702 , n49647 );
not ( n18683 , n29614 );
and ( n18684 , n18683 , RI1738c728_2071);
and ( n18685 , n49648 , n29614 );
or ( n49649 , n18684 , n18685 );
not ( n18686 , RI1754c610_2);
and ( n18687 , n18686 , n49649 );
and ( n18688 , C0 , RI1754c610_2);
or ( n49650 , n18687 , n18688 );
buf ( n49651 , n49650 );
not ( n49652 , n41752 );
and ( n49653 , n49652 , n41754 );
xor ( n49654 , n42925 , n49653 );
not ( n18689 , n29614 );
and ( n18690 , n18689 , RI1733ae28_2154);
and ( n18691 , n49654 , n29614 );
or ( n49655 , n18690 , n18691 );
not ( n18692 , RI1754c610_2);
and ( n18693 , n18692 , n49655 );
and ( n18694 , C0 , RI1754c610_2);
or ( n49656 , n18693 , n18694 );
buf ( n49657 , n49656 );
not ( n49658 , n42163 );
and ( n49659 , n49658 , n44069 );
xor ( n49660 , n42160 , n49659 );
not ( n18695 , n29614 );
and ( n18696 , n18695 , RI174018d8_1500);
and ( n18697 , n49660 , n29614 );
or ( n49661 , n18696 , n18697 );
not ( n18698 , RI1754c610_2);
and ( n18699 , n18698 , n49661 );
and ( n18700 , C0 , RI1754c610_2);
or ( n49662 , n18699 , n18700 );
buf ( n49663 , n49662 );
xor ( n49664 , n37555 , n34968 );
xor ( n49665 , n49664 , n39771 );
not ( n49666 , n49665 );
and ( n49667 , n49666 , n45415 );
xor ( n49668 , n45886 , n49667 );
not ( n18701 , n29614 );
and ( n18702 , n18701 , RI174a1a18_948);
and ( n18703 , n49668 , n29614 );
or ( n49669 , n18702 , n18703 );
not ( n18704 , RI1754c610_2);
and ( n18705 , n18704 , n49669 );
and ( n18706 , C0 , RI1754c610_2);
or ( n49670 , n18705 , n18706 );
buf ( n49671 , n49670 );
not ( n49672 , n49362 );
and ( n49673 , n49672 , n49364 );
xor ( n49674 , n46892 , n49673 );
not ( n18707 , n29614 );
and ( n18708 , n18707 , RI17414a00_1407);
and ( n18709 , n49674 , n29614 );
or ( n49675 , n18708 , n18709 );
not ( n18710 , RI1754c610_2);
and ( n18711 , n18710 , n49675 );
and ( n18712 , C0 , RI1754c610_2);
or ( n49676 , n18711 , n18712 );
buf ( n49677 , n49676 );
not ( n18713 , n27683 );
and ( n18714 , n18713 , RI19aab938_2485);
and ( n18715 , RI19ab5640_2413 , n27683 );
or ( n49678 , n18714 , n18715 );
not ( n18716 , RI1754c610_2);
and ( n18717 , n18716 , n49678 );
and ( n18718 , C0 , RI1754c610_2);
or ( n49679 , n18717 , n18718 );
buf ( n49680 , n49679 );
and ( n49681 , RI1754aea0_52 , n34844 );
buf ( n49682 , n49681 );
not ( n18719 , n34859 );
and ( n18720 , n18719 , n49682 );
and ( n18721 , RI1754aea0_52 , n34859 );
or ( n49683 , n18720 , n18721 );
not ( n18722 , RI19a22f70_2797);
and ( n18723 , n18722 , n49683 );
and ( n18724 , C0 , RI19a22f70_2797);
or ( n49684 , n18723 , n18724 );
not ( n18725 , n27683 );
and ( n18726 , n18725 , RI19a23510_2794);
and ( n18727 , n49684 , n27683 );
or ( n49685 , n18726 , n18727 );
not ( n18728 , RI1754c610_2);
and ( n18729 , n18728 , n49685 );
and ( n18730 , C0 , RI1754c610_2);
or ( n49686 , n18729 , n18730 );
buf ( n49687 , n49686 );
not ( n49688 , n39210 );
and ( n49689 , n49688 , n39215 );
xor ( n49690 , n43937 , n49689 );
not ( n18731 , n29614 );
and ( n18732 , n18731 , RI173d74e8_1706);
and ( n18733 , n49690 , n29614 );
or ( n49691 , n18732 , n18733 );
not ( n18734 , RI1754c610_2);
and ( n18735 , n18734 , n49691 );
and ( n18736 , C0 , RI1754c610_2);
or ( n49692 , n18735 , n18736 );
buf ( n49693 , n49692 );
not ( n49694 , n41257 );
xor ( n49695 , n38910 , n42309 );
xor ( n49696 , n49695 , n43464 );
and ( n49697 , n49694 , n49696 );
xor ( n49698 , n41254 , n49697 );
not ( n18737 , n29614 );
and ( n18738 , n18737 , RI17512578_709);
and ( n18739 , n49698 , n29614 );
or ( n49699 , n18738 , n18739 );
not ( n18740 , RI1754c610_2);
and ( n18741 , n18740 , n49699 );
and ( n18742 , C0 , RI1754c610_2);
or ( n49700 , n18741 , n18742 );
buf ( n49701 , n49700 );
buf ( n49702 , RI174889c8_1070);
buf ( n49703 , RI1750aee0_732);
xor ( n49704 , n37120 , n40237 );
xor ( n49705 , n49704 , n40254 );
not ( n49706 , n49705 );
xor ( n49707 , n39650 , n35216 );
xor ( n49708 , n49707 , n41241 );
and ( n49709 , n49706 , n49708 );
xor ( n49710 , n41069 , n49709 );
not ( n18743 , n29614 );
and ( n18744 , n18743 , RI17478000_1151);
and ( n18745 , n49710 , n29614 );
or ( n49711 , n18744 , n18745 );
not ( n18746 , RI1754c610_2);
and ( n18747 , n18746 , n49711 );
and ( n18748 , C0 , RI1754c610_2);
or ( n49712 , n18747 , n18748 );
buf ( n49713 , n49712 );
not ( n49714 , n45087 );
xor ( n49715 , n41841 , n33282 );
xor ( n49716 , n49715 , n37623 );
and ( n49717 , n49714 , n49716 );
xor ( n49718 , n45084 , n49717 );
not ( n18749 , n29614 );
and ( n18750 , n18749 , RI17526f78_645);
and ( n18751 , n49718 , n29614 );
or ( n49719 , n18750 , n18751 );
not ( n18752 , RI1754c610_2);
and ( n18753 , n18752 , n49719 );
and ( n18754 , C0 , RI1754c610_2);
or ( n49720 , n18753 , n18754 );
buf ( n49721 , n49720 );
not ( n18755 , n27683 );
and ( n18756 , n18755 , RI19a8e220_2696);
and ( n18757 , RI19a983d8_2624 , n27683 );
or ( n49722 , n18756 , n18757 );
not ( n18758 , RI1754c610_2);
and ( n18759 , n18758 , n49722 );
and ( n18760 , C0 , RI1754c610_2);
or ( n49723 , n18759 , n18760 );
buf ( n49724 , n49723 );
not ( n49725 , n43621 );
and ( n49726 , n49725 , n43623 );
xor ( n49727 , n48964 , n49726 );
not ( n18761 , n29614 );
and ( n18762 , n18761 , RI17456c70_1313);
and ( n18763 , n49727 , n29614 );
or ( n49728 , n18762 , n18763 );
not ( n18764 , RI1754c610_2);
and ( n18765 , n18764 , n49728 );
and ( n18766 , C0 , RI1754c610_2);
or ( n49729 , n18765 , n18766 );
buf ( n49730 , n49729 );
and ( n49731 , RI1754b260_44 , n34844 );
and ( n49732 , RI1754b260_44 , n34847 );
or ( n49733 , n49731 , n49732 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n18767 , n34859 );
and ( n18768 , n18767 , n49733 );
and ( n18769 , RI1754b260_44 , n34859 );
or ( n49734 , n18768 , n18769 );
not ( n18770 , RI19a22f70_2797);
and ( n18771 , n18770 , n49734 );
and ( n18772 , C0 , RI19a22f70_2797);
or ( n49735 , n18771 , n18772 );
not ( n18773 , n27683 );
and ( n18774 , n18773 , RI19abe2e0_2348);
and ( n18775 , n49735 , n27683 );
or ( n49736 , n18774 , n18775 );
not ( n18776 , RI1754c610_2);
and ( n18777 , n18776 , n49736 );
and ( n18778 , C0 , RI1754c610_2);
or ( n49737 , n18777 , n18778 );
buf ( n49738 , n49737 );
not ( n49739 , n39283 );
and ( n49740 , n49739 , n39285 );
xor ( n49741 , n42227 , n49740 );
not ( n18779 , n29614 );
and ( n18780 , n18779 , RI173bbd20_1840);
and ( n18781 , n49741 , n29614 );
or ( n49742 , n18780 , n18781 );
not ( n18782 , RI1754c610_2);
and ( n18783 , n18782 , n49742 );
and ( n18784 , C0 , RI1754c610_2);
or ( n49743 , n18783 , n18784 );
buf ( n49744 , n49743 );
not ( n18785 , n27683 );
and ( n18786 , n18785 , RI19aa62f8_2521);
and ( n18787 , RI19ab0528_2451 , n27683 );
or ( n49745 , n18786 , n18787 );
not ( n18788 , RI1754c610_2);
and ( n18789 , n18788 , n49745 );
and ( n18790 , C0 , RI1754c610_2);
or ( n49746 , n18789 , n18790 );
buf ( n49747 , n49746 );
xor ( n49748 , n35609 , n41543 );
xor ( n49749 , n49748 , n34669 );
not ( n49750 , n49573 );
and ( n49751 , n49750 , n49575 );
xor ( n49752 , n49749 , n49751 );
not ( n18791 , n29614 );
and ( n18792 , n18791 , RI17471070_1185);
and ( n18793 , n49752 , n29614 );
or ( n49753 , n18792 , n18793 );
not ( n18794 , RI1754c610_2);
and ( n18795 , n18794 , n49753 );
and ( n18796 , C0 , RI1754c610_2);
or ( n49754 , n18795 , n18796 );
buf ( n49755 , n49754 );
not ( n49756 , n48535 );
and ( n49757 , n49756 , n46246 );
xor ( n49758 , n44464 , n49757 );
not ( n18797 , n29614 );
and ( n18798 , n18797 , RI1745c508_1286);
and ( n18799 , n49758 , n29614 );
or ( n49759 , n18798 , n18799 );
not ( n18800 , RI1754c610_2);
and ( n18801 , n18800 , n49759 );
and ( n18802 , C0 , RI1754c610_2);
or ( n49760 , n18801 , n18802 );
buf ( n49761 , n49760 );
not ( n18803 , n27683 );
and ( n18804 , n18803 , RI19aa8080_2509);
and ( n18805 , RI19ab2148_2439 , n27683 );
or ( n49762 , n18804 , n18805 );
not ( n18806 , RI1754c610_2);
and ( n18807 , n18806 , n49762 );
and ( n18808 , C0 , RI1754c610_2);
or ( n49763 , n18807 , n18808 );
buf ( n49764 , n49763 );
buf ( n49765 , RI174b2728_866);
buf ( n49766 , RI174a4178_936);
not ( n18809 , RI1754c610_2);
and ( n18810 , n18809 , RI17537fd0_593);
and ( n18811 , C0 , RI1754c610_2);
or ( n49767 , n18810 , n18811 );
buf ( n49768 , n49767 );
xor ( n49769 , n41844 , n33282 );
xor ( n49770 , n49769 , n37623 );
xor ( n49771 , n36693 , n39655 );
xor ( n49772 , n49771 , n41125 );
not ( n49773 , n49772 );
and ( n49774 , n49773 , n48446 );
xor ( n49775 , n49770 , n49774 );
not ( n18812 , n29614 );
and ( n18813 , n18812 , RI1744f308_1350);
and ( n18814 , n49775 , n29614 );
or ( n49776 , n18813 , n18814 );
not ( n18815 , RI1754c610_2);
and ( n18816 , n18815 , n49776 );
and ( n18817 , C0 , RI1754c610_2);
or ( n49777 , n18816 , n18817 );
buf ( n49778 , n49777 );
not ( n18818 , n27683 );
and ( n18819 , n18818 , RI19aba398_2379);
and ( n18820 , RI19ac2cf0_2308 , n27683 );
or ( n49779 , n18819 , n18820 );
not ( n18821 , RI1754c610_2);
and ( n18822 , n18821 , n49779 );
and ( n18823 , C0 , RI1754c610_2);
or ( n49780 , n18822 , n18823 );
buf ( n49781 , n49780 );
buf ( n49782 , RI17476f98_1156);
buf ( n49783 , RI17468d30_1225);
not ( n49784 , n41971 );
and ( n49785 , n49784 , n41992 );
xor ( n49786 , n46269 , n49785 );
not ( n18824 , n29614 );
and ( n18825 , n18824 , RI17509a40_736);
and ( n18826 , n49786 , n29614 );
or ( n49787 , n18825 , n18826 );
not ( n18827 , RI1754c610_2);
and ( n18828 , n18827 , n49787 );
and ( n18829 , C0 , RI1754c610_2);
or ( n49788 , n18828 , n18829 );
buf ( n49789 , n49788 );
not ( n49790 , n45399 );
xor ( n49791 , n36778 , n38214 );
xor ( n49792 , n49791 , n38244 );
and ( n49793 , n49790 , n49792 );
xor ( n49794 , n44280 , n49793 );
not ( n18830 , n29614 );
and ( n18831 , n18830 , RI175172d0_694);
and ( n18832 , n49794 , n29614 );
or ( n49795 , n18831 , n18832 );
not ( n18833 , RI1754c610_2);
and ( n18834 , n18833 , n49795 );
and ( n18835 , C0 , RI1754c610_2);
or ( n49796 , n18834 , n18835 );
buf ( n49797 , n49796 );
not ( n18836 , n27683 );
and ( n18837 , n18836 , RI19accc50_2233);
and ( n18838 , RI19a88be0_2733 , n27683 );
or ( n49798 , n18837 , n18838 );
not ( n18839 , RI1754c610_2);
and ( n18840 , n18839 , n49798 );
and ( n18841 , C0 , RI1754c610_2);
or ( n49799 , n18840 , n18841 );
buf ( n49800 , n49799 );
buf ( n49801 , RI174b5ef0_849);
buf ( n49802 , RI1749d1e8_970);
not ( n49803 , n39564 );
and ( n49804 , n49803 , n46705 );
xor ( n49805 , n39526 , n49804 );
not ( n18842 , n29614 );
and ( n18843 , n18842 , RI174bc7f0_824);
and ( n18844 , n49805 , n29614 );
or ( n49806 , n18843 , n18844 );
not ( n18845 , RI1754c610_2);
and ( n18846 , n18845 , n49806 );
and ( n18847 , C0 , RI1754c610_2);
or ( n49807 , n18846 , n18847 );
buf ( n49808 , n49807 );
not ( n49809 , n48748 );
and ( n49810 , n49809 , n45612 );
xor ( n49811 , n48745 , n49810 );
not ( n18848 , n29614 );
and ( n18849 , n18848 , RI17466288_1238);
and ( n18850 , n49811 , n29614 );
or ( n49812 , n18849 , n18850 );
not ( n18851 , RI1754c610_2);
and ( n18852 , n18851 , n49812 );
and ( n18853 , C0 , RI1754c610_2);
or ( n49813 , n18852 , n18853 );
buf ( n49814 , n49813 );
not ( n18854 , n27683 );
and ( n18855 , n18854 , RI19acc3e0_2237);
and ( n18856 , RI19a88028_2738 , n27683 );
or ( n49815 , n18855 , n18856 );
not ( n18857 , RI1754c610_2);
and ( n18858 , n18857 , n49815 );
and ( n18859 , C0 , RI1754c610_2);
or ( n49816 , n18858 , n18859 );
buf ( n49817 , n49816 );
xor ( n49818 , n39266 , n38445 );
xor ( n49819 , n49818 , n37549 );
xor ( n49820 , n42337 , n29981 );
xor ( n49821 , n49820 , n35955 );
not ( n49822 , n49821 );
and ( n49823 , n49822 , n43809 );
xor ( n49824 , n49819 , n49823 );
not ( n18860 , n29614 );
and ( n18861 , n18860 , RI17414028_1410);
and ( n18862 , n49824 , n29614 );
or ( n49825 , n18861 , n18862 );
not ( n18863 , RI1754c610_2);
and ( n18864 , n18863 , n49825 );
and ( n18865 , C0 , RI1754c610_2);
or ( n49826 , n18864 , n18865 );
buf ( n49827 , n49826 );
not ( n18866 , n27683 );
and ( n18867 , n18866 , RI19ab9498_2386);
and ( n18868 , RI19ac1b98_2316 , n27683 );
or ( n49828 , n18867 , n18868 );
not ( n18869 , RI1754c610_2);
and ( n18870 , n18869 , n49828 );
and ( n18871 , C0 , RI1754c610_2);
or ( n49829 , n18870 , n18871 );
buf ( n49830 , n49829 );
not ( n49831 , n44891 );
and ( n49832 , n49831 , n45846 );
xor ( n49833 , n44888 , n49832 );
not ( n18872 , n29614 );
and ( n18873 , n18872 , RI17411238_1424);
and ( n18874 , n49833 , n29614 );
or ( n49834 , n18873 , n18874 );
not ( n18875 , RI1754c610_2);
and ( n18876 , n18875 , n49834 );
and ( n18877 , C0 , RI1754c610_2);
or ( n49835 , n18876 , n18877 );
buf ( n49836 , n49835 );
not ( n18878 , n27683 );
and ( n18879 , n18878 , RI19ac4460_2297);
and ( n18880 , RI19acd100_2231 , n27683 );
or ( n49837 , n18879 , n18880 );
not ( n18881 , RI1754c610_2);
and ( n18882 , n18881 , n49837 );
and ( n18883 , C0 , RI1754c610_2);
or ( n49838 , n18882 , n18883 );
buf ( n49839 , n49838 );
not ( n49840 , n46343 );
and ( n49841 , n49840 , n38496 );
xor ( n49842 , n34252 , n49841 );
not ( n18884 , n29614 );
and ( n18885 , n18884 , RI173adab8_1909);
and ( n18886 , n49842 , n29614 );
or ( n49843 , n18885 , n18886 );
not ( n18887 , RI1754c610_2);
and ( n18888 , n18887 , n49843 );
and ( n18889 , C0 , RI1754c610_2);
or ( n49844 , n18888 , n18889 );
buf ( n49845 , n49844 );
not ( n18890 , n27683 );
and ( n18891 , n18890 , RI19acc818_2235);
and ( n18892 , RI19a88460_2736 , n27683 );
or ( n49846 , n18891 , n18892 );
not ( n18893 , RI1754c610_2);
and ( n18894 , n18893 , n49846 );
and ( n18895 , C0 , RI1754c610_2);
or ( n49847 , n18894 , n18895 );
buf ( n49848 , n49847 );
not ( n18896 , n27683 );
and ( n18897 , n18896 , RI19ac0f68_2323);
and ( n18898 , RI19aca298_2254 , n27683 );
or ( n49849 , n18897 , n18898 );
not ( n18899 , RI1754c610_2);
and ( n18900 , n18899 , n49849 );
and ( n18901 , C0 , RI1754c610_2);
or ( n49850 , n18900 , n18901 );
buf ( n49851 , n49850 );
xor ( n49852 , n40000 , n40341 );
xor ( n49853 , n49852 , n40091 );
not ( n49854 , n48932 );
and ( n49855 , n49854 , n48934 );
xor ( n49856 , n49853 , n49855 );
not ( n18902 , n29614 );
and ( n18903 , n18902 , RI173e8540_1623);
and ( n18904 , n49856 , n29614 );
or ( n49857 , n18903 , n18904 );
not ( n18905 , RI1754c610_2);
and ( n18906 , n18905 , n49857 );
and ( n18907 , C0 , RI1754c610_2);
or ( n49858 , n18906 , n18907 );
buf ( n49859 , n49858 );
not ( n49860 , n43534 );
and ( n49861 , n49860 , n43536 );
xor ( n49862 , n48481 , n49861 );
not ( n18908 , n29614 );
and ( n18909 , n18908 , RI173fbcf8_1528);
and ( n18910 , n49862 , n29614 );
or ( n49863 , n18909 , n18910 );
not ( n18911 , RI1754c610_2);
and ( n18912 , n18911 , n49863 );
and ( n18913 , C0 , RI1754c610_2);
or ( n49864 , n18912 , n18913 );
buf ( n49865 , n49864 );
buf ( n49866 , RI174cbf70_776);
not ( n49867 , n45299 );
and ( n49868 , n49867 , n39468 );
xor ( n49869 , n45262 , n49868 );
not ( n18914 , n29614 );
and ( n18915 , n18914 , RI17448d50_1381);
and ( n18916 , n49869 , n29614 );
or ( n49870 , n18915 , n18916 );
not ( n18917 , RI1754c610_2);
and ( n18918 , n18917 , n49870 );
and ( n18919 , C0 , RI1754c610_2);
or ( n49871 , n18918 , n18919 );
buf ( n49872 , n49871 );
buf ( n49873 , RI17491d70_1025);
buf ( n49874 , RI1746b7d8_1212);
not ( n49875 , n38649 );
and ( n49876 , n49875 , n44809 );
xor ( n49877 , n38604 , n49876 );
not ( n18920 , n29614 );
and ( n18921 , n18920 , RI17496c30_1001);
and ( n18922 , n49877 , n29614 );
or ( n49878 , n18921 , n18922 );
not ( n18923 , RI1754c610_2);
and ( n18924 , n18923 , n49878 );
and ( n18925 , C0 , RI1754c610_2);
or ( n49879 , n18924 , n18925 );
buf ( n49880 , n49879 );
not ( n49881 , n49554 );
xor ( n49882 , n30196 , n34755 );
xor ( n49883 , n49882 , n35311 );
and ( n49884 , n49881 , n49883 );
xor ( n49885 , n49551 , n49884 );
not ( n18926 , n29614 );
and ( n18927 , n18926 , RI174c7740_790);
and ( n18928 , n49885 , n29614 );
or ( n49886 , n18927 , n18928 );
not ( n18929 , RI1754c610_2);
and ( n18930 , n18929 , n49886 );
and ( n18931 , C0 , RI1754c610_2);
or ( n49887 , n18930 , n18931 );
buf ( n49888 , n49887 );
xor ( n49889 , n37471 , n42188 );
xor ( n49890 , n49889 , n41526 );
not ( n49891 , n40524 );
and ( n49892 , n49891 , n40526 );
xor ( n49893 , n49890 , n49892 );
not ( n18932 , n29614 );
and ( n18933 , n18932 , RI17394090_2034);
and ( n18934 , n49893 , n29614 );
or ( n49894 , n18933 , n18934 );
not ( n18935 , RI1754c610_2);
and ( n18936 , n18935 , n49894 );
and ( n18937 , C0 , RI1754c610_2);
or ( n49895 , n18936 , n18937 );
buf ( n49896 , n49895 );
xor ( n49897 , n36186 , n32309 );
xor ( n49898 , n49897 , n32923 );
not ( n49899 , n49898 );
xor ( n49900 , n40947 , n38793 );
xor ( n49901 , n49900 , n40563 );
and ( n49902 , n49899 , n49901 );
xor ( n49903 , n45197 , n49902 );
not ( n18938 , n29614 );
and ( n18939 , n18938 , RI17474ec8_1166);
and ( n18940 , n49903 , n29614 );
or ( n49904 , n18939 , n18940 );
not ( n18941 , RI1754c610_2);
and ( n18942 , n18941 , n49904 );
and ( n18943 , C0 , RI1754c610_2);
or ( n49905 , n18942 , n18943 );
buf ( n49906 , n49905 );
xor ( n49907 , n39815 , n37800 );
xor ( n49908 , n49907 , n37814 );
not ( n49909 , n49908 );
and ( n49910 , n49909 , n48305 );
xor ( n49911 , n48903 , n49910 );
not ( n18944 , n29614 );
and ( n18945 , n18944 , RI1751a660_684);
and ( n18946 , n49911 , n29614 );
or ( n49912 , n18945 , n18946 );
not ( n18947 , RI1754c610_2);
and ( n18948 , n18947 , n49912 );
and ( n18949 , C0 , RI1754c610_2);
or ( n49913 , n18948 , n18949 );
buf ( n49914 , n49913 );
xor ( n49915 , n40965 , n36844 );
xor ( n49916 , n49915 , n36874 );
not ( n49917 , n49065 );
and ( n49918 , n49917 , n49067 );
xor ( n49919 , n49916 , n49918 );
not ( n18950 , n29614 );
and ( n18951 , n18950 , RI1740b658_1452);
and ( n18952 , n49919 , n29614 );
or ( n49920 , n18951 , n18952 );
not ( n18953 , RI1754c610_2);
and ( n18954 , n18953 , n49920 );
and ( n18955 , C0 , RI1754c610_2);
or ( n49921 , n18954 , n18955 );
buf ( n49922 , n49921 );
not ( n18956 , n27683 );
and ( n18957 , n18956 , RI19ac63c8_2283);
and ( n18958 , RI19acef78_2218 , n27683 );
or ( n49923 , n18957 , n18958 );
not ( n18959 , RI1754c610_2);
and ( n18960 , n18959 , n49923 );
and ( n18961 , C0 , RI1754c610_2);
or ( n49924 , n18960 , n18961 );
buf ( n49925 , n49924 );
not ( n18962 , n27683 );
and ( n18963 , n18962 , RI19ab82c8_2394);
and ( n18964 , RI19ac0f68_2323 , n27683 );
or ( n49926 , n18963 , n18964 );
not ( n18965 , RI1754c610_2);
and ( n18966 , n18965 , n49926 );
and ( n18967 , C0 , RI1754c610_2);
or ( n49927 , n18966 , n18967 );
buf ( n49928 , n49927 );
not ( n49929 , n44419 );
and ( n49930 , n49929 , n45572 );
xor ( n49931 , n42683 , n49930 );
not ( n18968 , n29614 );
and ( n18969 , n18968 , RI17409240_1463);
and ( n18970 , n49931 , n29614 );
or ( n49932 , n18969 , n18970 );
not ( n18971 , RI1754c610_2);
and ( n18972 , n18971 , n49932 );
and ( n18973 , C0 , RI1754c610_2);
or ( n49933 , n18972 , n18973 );
buf ( n49934 , n49933 );
buf ( n49935 , RI174ca5a8_781);
buf ( n49936 , RI1748f610_1037);
not ( n18974 , n27683 );
and ( n18975 , n18974 , RI19a9c1b8_2597);
and ( n18976 , RI19aa5740_2526 , n27683 );
or ( n49937 , n18975 , n18976 );
not ( n18977 , RI1754c610_2);
and ( n18978 , n18977 , n49937 );
and ( n18979 , C0 , RI1754c610_2);
or ( n49938 , n18978 , n18979 );
buf ( n49939 , n49938 );
buf ( n49940 , RI17484198_1092);
buf ( n49941 , RI1750c8a8_727);
not ( n49942 , n43923 );
and ( n49943 , n49942 , n43925 );
xor ( n49944 , n45204 , n49943 );
not ( n18980 , n29614 );
and ( n18981 , n18980 , RI174bcd18_823);
and ( n18982 , n49944 , n29614 );
or ( n49945 , n18981 , n18982 );
not ( n18983 , RI1754c610_2);
and ( n18984 , n18983 , n49945 );
and ( n18985 , C0 , RI1754c610_2);
or ( n49946 , n18984 , n18985 );
buf ( n49947 , n49946 );
not ( n49948 , n44898 );
and ( n49949 , n49948 , n44900 );
xor ( n49950 , n46804 , n49949 );
not ( n18986 , n29614 );
and ( n18987 , n18986 , RI17389fc8_2083);
and ( n18988 , n49950 , n29614 );
or ( n49951 , n18987 , n18988 );
not ( n18989 , RI1754c610_2);
and ( n18990 , n18989 , n49951 );
and ( n18991 , C0 , RI1754c610_2);
or ( n49952 , n18990 , n18991 );
buf ( n49953 , n49952 );
not ( n49954 , n47744 );
and ( n49955 , n49954 , n45108 );
xor ( n49956 , n47816 , n49955 );
not ( n18992 , n29614 );
and ( n18993 , n18992 , RI17489d78_1064);
and ( n18994 , n49956 , n29614 );
or ( n49957 , n18993 , n18994 );
not ( n18995 , RI1754c610_2);
and ( n18996 , n18995 , n49957 );
and ( n18997 , C0 , RI1754c610_2);
or ( n49958 , n18996 , n18997 );
buf ( n49959 , n49958 );
xor ( n49960 , n33643 , n35069 );
xor ( n49961 , n49960 , n41854 );
xor ( n49962 , n41525 , n33824 );
xor ( n49963 , n49962 , n32786 );
not ( n49964 , n49963 );
xor ( n49965 , n35923 , n36148 );
xor ( n49966 , n49965 , n37421 );
and ( n49967 , n49964 , n49966 );
xor ( n49968 , n49961 , n49967 );
not ( n18998 , n29614 );
and ( n18999 , n18998 , RI173fd738_1520);
and ( n19000 , n49968 , n29614 );
or ( n49969 , n18999 , n19000 );
not ( n19001 , RI1754c610_2);
and ( n19002 , n19001 , n49969 );
and ( n19003 , C0 , RI1754c610_2);
or ( n49970 , n19002 , n19003 );
buf ( n49971 , n49970 );
xor ( n49972 , n36816 , n44146 );
xor ( n49973 , n49972 , n41198 );
not ( n49974 , n40112 );
and ( n49975 , n49974 , n40117 );
xor ( n49976 , n49973 , n49975 );
not ( n19004 , n29614 );
and ( n19005 , n19004 , RI17447658_1388);
and ( n19006 , n49976 , n29614 );
or ( n49977 , n19005 , n19006 );
not ( n19007 , RI1754c610_2);
and ( n19008 , n19007 , n49977 );
and ( n19009 , C0 , RI1754c610_2);
or ( n49978 , n19008 , n19009 );
buf ( n49979 , n49978 );
not ( n49980 , n46442 );
and ( n49981 , n49980 , n44432 );
xor ( n49982 , n46439 , n49981 );
not ( n19010 , n29614 );
and ( n19011 , n19010 , RI17479068_1146);
and ( n19012 , n49982 , n29614 );
or ( n49983 , n19011 , n19012 );
not ( n19013 , RI1754c610_2);
and ( n19014 , n19013 , n49983 );
and ( n19015 , C0 , RI1754c610_2);
or ( n49984 , n19014 , n19015 );
buf ( n49985 , n49984 );
not ( n49986 , n45629 );
and ( n49987 , n49986 , n48828 );
xor ( n49988 , n45626 , n49987 );
not ( n19016 , n29614 );
and ( n19017 , n19016 , RI17535258_601);
and ( n19018 , n49988 , n29614 );
or ( n49989 , n19017 , n19018 );
not ( n19019 , RI1754c610_2);
and ( n19020 , n19019 , n49989 );
and ( n19021 , C0 , RI1754c610_2);
or ( n49990 , n19020 , n19021 );
buf ( n49991 , n49990 );
not ( n49992 , n42803 );
and ( n49993 , n49992 , n41559 );
xor ( n49994 , n48353 , n49993 );
not ( n19022 , n29614 );
and ( n19023 , n19022 , RI1733c520_2147);
and ( n19024 , n49994 , n29614 );
or ( n49995 , n19023 , n19024 );
not ( n19025 , RI1754c610_2);
and ( n19026 , n19025 , n49995 );
and ( n19027 , C0 , RI1754c610_2);
or ( n49996 , n19026 , n19027 );
buf ( n49997 , n49996 );
not ( n49998 , n46202 );
and ( n49999 , n49998 , n49201 );
xor ( n50000 , n46199 , n49999 );
not ( n19028 , n29614 );
and ( n19029 , n19028 , RI1751f3b8_669);
and ( n19030 , n50000 , n29614 );
or ( n50001 , n19029 , n19030 );
not ( n19031 , RI1754c610_2);
and ( n19032 , n19031 , n50001 );
and ( n19033 , C0 , RI1754c610_2);
or ( n50002 , n19032 , n19033 );
buf ( n50003 , n50002 );
xor ( n50004 , n33098 , n38244 );
xor ( n50005 , n50004 , n37235 );
xor ( n50006 , n32278 , n36003 );
xor ( n50007 , n50006 , n38553 );
not ( n50008 , n50007 );
and ( n50009 , n50008 , n49961 );
xor ( n50010 , n50005 , n50009 );
not ( n19034 , n29614 );
and ( n19035 , n19034 , RI173e0548_1662);
and ( n19036 , n50010 , n29614 );
or ( n50011 , n19035 , n19036 );
not ( n19037 , RI1754c610_2);
and ( n19038 , n19037 , n50011 );
and ( n19039 , C0 , RI1754c610_2);
or ( n50012 , n19038 , n19039 );
buf ( n50013 , n50012 );
not ( n19040 , n27683 );
and ( n19041 , n19040 , RI19ac8e70_2263);
and ( n19042 , RI19a83f78_2766 , n27683 );
or ( n50014 , n19041 , n19042 );
not ( n19043 , RI1754c610_2);
and ( n19044 , n19043 , n50014 );
and ( n19045 , C0 , RI1754c610_2);
or ( n50015 , n19044 , n19045 );
buf ( n50016 , n50015 );
xor ( n50017 , n32259 , n36003 );
xor ( n50018 , n50017 , n38553 );
not ( n50019 , n50018 );
xor ( n50020 , n37733 , n41772 );
xor ( n50021 , n50020 , n32663 );
and ( n50022 , n50019 , n50021 );
xor ( n50023 , n45009 , n50022 );
not ( n19046 , n29614 );
and ( n19047 , n19046 , RI174665d0_1237);
and ( n19048 , n50023 , n29614 );
or ( n50024 , n19047 , n19048 );
not ( n19049 , RI1754c610_2);
and ( n19050 , n19049 , n50024 );
and ( n19051 , C0 , RI1754c610_2);
or ( n50025 , n19050 , n19051 );
buf ( n50026 , n50025 );
xor ( n50027 , n44136 , n34572 );
xor ( n50028 , n50027 , n34622 );
xor ( n50029 , n38772 , n40516 );
xor ( n50030 , n50029 , n40966 );
not ( n50031 , n50030 );
and ( n50032 , n50031 , n48732 );
xor ( n50033 , n50028 , n50032 );
not ( n19052 , n29614 );
and ( n19053 , n19052 , RI17470008_1190);
and ( n19054 , n50033 , n29614 );
or ( n50034 , n19053 , n19054 );
not ( n19055 , RI1754c610_2);
and ( n19056 , n19055 , n50034 );
and ( n19057 , C0 , RI1754c610_2);
or ( n50035 , n19056 , n19057 );
buf ( n50036 , n50035 );
not ( n50037 , n43722 );
and ( n50038 , n50037 , n43724 );
xor ( n50039 , n45782 , n50038 );
not ( n19058 , n29614 );
and ( n19059 , n19058 , RI1744d8c8_1358);
and ( n19060 , n50039 , n29614 );
or ( n50040 , n19059 , n19060 );
not ( n19061 , RI1754c610_2);
and ( n19062 , n19061 , n50040 );
and ( n19063 , C0 , RI1754c610_2);
or ( n50041 , n19062 , n19063 );
buf ( n50042 , n50041 );
xor ( n50043 , n40090 , n38037 );
xor ( n50044 , n50043 , n39740 );
not ( n50045 , n49549 );
and ( n50046 , n50045 , n49551 );
xor ( n50047 , n50044 , n50046 );
not ( n19064 , n29614 );
and ( n19065 , n19064 , RI173365f8_2176);
and ( n19066 , n50047 , n29614 );
or ( n50048 , n19065 , n19066 );
not ( n19067 , RI1754c610_2);
and ( n19068 , n19067 , n50048 );
and ( n19069 , C0 , RI1754c610_2);
or ( n50049 , n19068 , n19069 );
buf ( n50050 , n50049 );
xor ( n50051 , n34331 , n39604 );
xor ( n50052 , n50051 , n39621 );
xor ( n50053 , n40165 , n39039 );
xor ( n50054 , n50053 , n39065 );
not ( n50055 , n50054 );
xor ( n50056 , n33704 , n35514 );
xor ( n50057 , n50056 , n40486 );
and ( n50058 , n50055 , n50057 );
xor ( n50059 , n50052 , n50058 );
not ( n19070 , n29614 );
and ( n19071 , n19070 , RI1751c550_678);
and ( n19072 , n50059 , n29614 );
or ( n50060 , n19071 , n19072 );
not ( n19073 , RI1754c610_2);
and ( n19074 , n19073 , n50060 );
and ( n19075 , C0 , RI1754c610_2);
or ( n50061 , n19074 , n19075 );
buf ( n50062 , n50061 );
not ( n50063 , n48048 );
xor ( n50064 , n41282 , n38648 );
xor ( n50065 , n50064 , n40890 );
and ( n50066 , n50063 , n50065 );
xor ( n50067 , n43950 , n50066 );
not ( n19076 , n29614 );
and ( n19077 , n19076 , RI174bd240_822);
and ( n19078 , n50067 , n29614 );
or ( n50068 , n19077 , n19078 );
not ( n19079 , RI1754c610_2);
and ( n19080 , n19079 , n50068 );
and ( n19081 , C0 , RI1754c610_2);
or ( n50069 , n19080 , n19081 );
buf ( n50070 , n50069 );
xor ( n50071 , n41538 , n32786 );
xor ( n50072 , n50071 , n32863 );
not ( n50073 , n50072 );
and ( n50074 , n50073 , n42278 );
xor ( n50075 , n44953 , n50074 );
not ( n19082 , n29614 );
and ( n19083 , n19082 , RI1745bb30_1289);
and ( n19084 , n50075 , n29614 );
or ( n50076 , n19083 , n19084 );
not ( n19085 , RI1754c610_2);
and ( n19086 , n19085 , n50076 );
and ( n19087 , C0 , RI1754c610_2);
or ( n50077 , n19086 , n19087 );
buf ( n50078 , n50077 );
xor ( n50079 , n41124 , n41241 );
xor ( n50080 , n50079 , n41287 );
not ( n50081 , n50080 );
and ( n50082 , n50081 , n45728 );
xor ( n50083 , n46320 , n50082 );
not ( n19088 , n29614 );
and ( n19089 , n19088 , RI173b0bf0_1894);
and ( n19090 , n50083 , n29614 );
or ( n50084 , n19089 , n19090 );
not ( n19091 , RI1754c610_2);
and ( n19092 , n19091 , n50084 );
and ( n19093 , C0 , RI1754c610_2);
or ( n50085 , n19092 , n19093 );
buf ( n50086 , n50085 );
not ( n19094 , n27683 );
and ( n19095 , n19094 , RI19ac3d58_2300);
and ( n19096 , RI19acc9f8_2234 , n27683 );
or ( n50087 , n19095 , n19096 );
not ( n19097 , RI1754c610_2);
and ( n19098 , n19097 , n50087 );
and ( n19099 , C0 , RI1754c610_2);
or ( n50088 , n19098 , n19099 );
buf ( n50089 , n50088 );
not ( n19100 , RI1754c610_2);
and ( n19101 , n19100 , RI19ad0bb0_2206);
and ( n19102 , C0 , RI1754c610_2);
or ( n50090 , n19101 , n19102 );
buf ( n50091 , n50090 );
not ( n50092 , n45017 );
and ( n50093 , n50092 , n41148 );
xor ( n50094 , n47659 , n50093 );
not ( n19103 , n29614 );
and ( n19104 , n19103 , RI17453160_1331);
and ( n19105 , n50094 , n29614 );
or ( n50095 , n19104 , n19105 );
not ( n19106 , RI1754c610_2);
and ( n19107 , n19106 , n50095 );
and ( n19108 , C0 , RI1754c610_2);
or ( n50096 , n19107 , n19108 );
buf ( n50097 , n50096 );
not ( n50098 , n43040 );
and ( n50099 , n50098 , n47157 );
xor ( n50100 , n43037 , n50099 );
not ( n19109 , n29614 );
and ( n19110 , n19109 , RI17516358_697);
and ( n19111 , n50100 , n29614 );
or ( n50101 , n19110 , n19111 );
not ( n19112 , RI1754c610_2);
and ( n19113 , n19112 , n50101 );
and ( n19114 , C0 , RI1754c610_2);
or ( n50102 , n19113 , n19114 );
buf ( n50103 , n50102 );
not ( n50104 , n46708 );
and ( n50105 , n50104 , n39508 );
xor ( n50106 , n46705 , n50105 );
not ( n19115 , n29614 );
and ( n19116 , n19115 , RI1751b5d8_681);
and ( n19117 , n50106 , n29614 );
or ( n50107 , n19116 , n19117 );
not ( n19118 , RI1754c610_2);
and ( n19119 , n19118 , n50107 );
and ( n19120 , C0 , RI1754c610_2);
or ( n50108 , n19119 , n19120 );
buf ( n50109 , n50108 );
not ( n50110 , n45565 );
and ( n50111 , n50110 , n44922 );
xor ( n50112 , n42117 , n50111 );
not ( n19121 , n29614 );
and ( n19122 , n19121 , RI173cc6e8_1759);
and ( n19123 , n50112 , n29614 );
or ( n50113 , n19122 , n19123 );
not ( n19124 , RI1754c610_2);
and ( n19125 , n19124 , n50113 );
and ( n19126 , C0 , RI1754c610_2);
or ( n50114 , n19125 , n19126 );
buf ( n50115 , n50114 );
not ( n50116 , n44976 );
and ( n50117 , n50116 , n47586 );
xor ( n50118 , n44973 , n50117 );
not ( n19127 , n29614 );
and ( n19128 , n19127 , RI174a1040_951);
and ( n19129 , n50118 , n29614 );
or ( n50119 , n19128 , n19129 );
not ( n19130 , RI1754c610_2);
and ( n19131 , n19130 , n50119 );
and ( n19132 , C0 , RI1754c610_2);
or ( n50120 , n19131 , n19132 );
buf ( n50121 , n50120 );
xor ( n50122 , n35241 , n39952 );
xor ( n50123 , n50122 , n42945 );
xor ( n50124 , n40884 , n34340 );
xor ( n50125 , n50124 , n38817 );
not ( n50126 , n50125 );
xor ( n50127 , n41499 , n34445 );
xor ( n50128 , n50127 , n41885 );
and ( n50129 , n50126 , n50128 );
xor ( n50130 , n50123 , n50129 );
not ( n19133 , n29614 );
and ( n19134 , n19133 , RI174737d0_1173);
and ( n19135 , n50130 , n29614 );
or ( n50131 , n19134 , n19135 );
not ( n19136 , RI1754c610_2);
and ( n19137 , n19136 , n50131 );
and ( n19138 , C0 , RI1754c610_2);
or ( n50132 , n19137 , n19138 );
buf ( n50133 , n50132 );
xor ( n50134 , n40914 , n34797 );
xor ( n50135 , n50134 , n34837 );
not ( n50136 , n50135 );
xor ( n50137 , n35774 , n37331 );
xor ( n50138 , n50137 , n37129 );
and ( n50139 , n50136 , n50138 );
xor ( n50140 , n49497 , n50139 );
not ( n19139 , n29614 );
and ( n19140 , n19139 , RI173aa980_1924);
and ( n19141 , n50140 , n29614 );
or ( n50141 , n19140 , n19141 );
not ( n19142 , RI1754c610_2);
and ( n19143 , n19142 , n50141 );
and ( n19144 , C0 , RI1754c610_2);
or ( n50142 , n19143 , n19144 );
buf ( n50143 , n50142 );
buf ( n50144 , RI174837c0_1095);
buf ( n50145 , RI17469a50_1221);
buf ( n50146 , RI17513a18_705);
not ( n50147 , n43317 );
and ( n50148 , n50147 , n46277 );
xor ( n50149 , n43314 , n50148 );
not ( n19145 , n29614 );
and ( n19146 , n19145 , RI173ed748_1598);
and ( n19147 , n50149 , n29614 );
or ( n50150 , n19146 , n19147 );
not ( n19148 , RI1754c610_2);
and ( n19149 , n19148 , n50150 );
and ( n19150 , C0 , RI1754c610_2);
or ( n50151 , n19149 , n19150 );
buf ( n50152 , n50151 );
not ( n50153 , n38285 );
and ( n50154 , n50153 , n43735 );
xor ( n50155 , n38250 , n50154 );
not ( n19151 , n29614 );
and ( n19152 , n19151 , RI173a8568_1935);
and ( n19153 , n50155 , n29614 );
or ( n50156 , n19152 , n19153 );
not ( n19154 , RI1754c610_2);
and ( n19155 , n19154 , n50156 );
and ( n19156 , C0 , RI1754c610_2);
or ( n50157 , n19155 , n19156 );
buf ( n50158 , n50157 );
not ( n19157 , n27683 );
and ( n19158 , n19157 , RI19acf428_2216);
and ( n19159 , RI19aa12d0_2559 , n27683 );
or ( n50159 , n19158 , n19159 );
not ( n19160 , RI1754c610_2);
and ( n19161 , n19160 , n50159 );
and ( n19162 , C0 , RI1754c610_2);
or ( n50160 , n19161 , n19162 );
buf ( n50161 , n50160 );
xor ( n50162 , n35175 , n37915 );
xor ( n50163 , n50162 , n43492 );
not ( n50164 , n41692 );
and ( n50165 , n50164 , n40950 );
xor ( n50166 , n50163 , n50165 );
not ( n19163 , n29614 );
and ( n19164 , n19163 , RI173bee58_1825);
and ( n19165 , n50166 , n29614 );
or ( n50167 , n19164 , n19165 );
not ( n19166 , RI1754c610_2);
and ( n19167 , n19166 , n50167 );
and ( n19168 , C0 , RI1754c610_2);
or ( n50168 , n19167 , n19168 );
buf ( n50169 , n50168 );
xor ( n50170 , n30872 , n38115 );
xor ( n50171 , n50170 , n41622 );
not ( n50172 , n50171 );
and ( n50173 , n50172 , n47194 );
xor ( n50174 , n47036 , n50173 );
not ( n19169 , n29614 );
and ( n19170 , n19169 , RI173da2d8_1692);
and ( n19171 , n50174 , n29614 );
or ( n50175 , n19170 , n19171 );
not ( n19172 , RI1754c610_2);
and ( n19173 , n19172 , n50175 );
and ( n19174 , C0 , RI1754c610_2);
or ( n50176 , n19173 , n19174 );
buf ( n50177 , n50176 );
not ( n50178 , n43714 );
xor ( n50179 , n31924 , n36401 );
xor ( n50180 , n50179 , n33453 );
and ( n50181 , n50178 , n50180 );
xor ( n50182 , n43711 , n50181 );
not ( n19175 , n29614 );
and ( n19176 , n19175 , RI1748c190_1053);
and ( n19177 , n50182 , n29614 );
or ( n50183 , n19176 , n19177 );
not ( n19178 , RI1754c610_2);
and ( n19179 , n19178 , n50183 );
and ( n19180 , C0 , RI1754c610_2);
or ( n50184 , n19179 , n19180 );
buf ( n50185 , n50184 );
xor ( n50186 , n33616 , n41740 );
xor ( n50187 , n50186 , n38371 );
not ( n50188 , n50187 );
xor ( n50189 , n35425 , n32663 );
xor ( n50190 , n50189 , n32715 );
and ( n50191 , n50188 , n50190 );
xor ( n50192 , n47533 , n50191 );
not ( n19181 , n29614 );
and ( n19182 , n19181 , RI173f98e0_1539);
and ( n19183 , n50192 , n29614 );
or ( n50193 , n19182 , n19183 );
not ( n19184 , RI1754c610_2);
and ( n19185 , n19184 , n50193 );
and ( n19186 , C0 , RI1754c610_2);
or ( n50194 , n19185 , n19186 );
buf ( n50195 , n50194 );
not ( n50196 , n47390 );
and ( n50197 , n50196 , n48200 );
xor ( n50198 , n46726 , n50197 );
not ( n19187 , n29614 );
and ( n19188 , n19187 , RI17344ba8_2106);
and ( n19189 , n50198 , n29614 );
or ( n50199 , n19188 , n19189 );
not ( n19190 , RI1754c610_2);
and ( n19191 , n19190 , n50199 );
and ( n19192 , C0 , RI1754c610_2);
or ( n50200 , n19191 , n19192 );
buf ( n50201 , n50200 );
not ( n50202 , n44802 );
and ( n50203 , n50202 , n39302 );
xor ( n50204 , n44799 , n50203 );
not ( n19193 , n29614 );
and ( n19194 , n19193 , RI17342e20_2115);
and ( n19195 , n50204 , n29614 );
or ( n50205 , n19194 , n19195 );
not ( n19196 , RI1754c610_2);
and ( n19197 , n19196 , n50205 );
and ( n19198 , C0 , RI1754c610_2);
or ( n50206 , n19197 , n19198 );
buf ( n50207 , n50206 );
not ( n50208 , n47716 );
and ( n50209 , n50208 , n44570 );
xor ( n50210 , n48838 , n50209 );
not ( n19199 , n29614 );
and ( n19200 , n19199 , RI17513a18_705);
and ( n19201 , n50210 , n29614 );
or ( n50211 , n19200 , n19201 );
not ( n19202 , RI1754c610_2);
and ( n19203 , n19202 , n50211 );
and ( n19204 , C0 , RI1754c610_2);
or ( n50212 , n19203 , n19204 );
buf ( n50213 , n50212 );
xor ( n50214 , n39951 , n38724 );
xor ( n50215 , n50214 , n29425 );
not ( n50216 , n43148 );
and ( n50217 , n50216 , n43150 );
xor ( n50218 , n50215 , n50217 );
not ( n19205 , n29614 );
and ( n19206 , n19205 , RI173bfec0_1820);
and ( n19207 , n50218 , n29614 );
or ( n50219 , n19206 , n19207 );
not ( n19208 , RI1754c610_2);
and ( n19209 , n19208 , n50219 );
and ( n19210 , C0 , RI1754c610_2);
or ( n50220 , n19209 , n19210 );
buf ( n50221 , n50220 );
not ( n50222 , n44886 );
and ( n50223 , n50222 , n44888 );
xor ( n50224 , n45848 , n50223 );
not ( n19211 , n29614 );
and ( n19212 , n19211 , RI1750b408_731);
and ( n19213 , n50224 , n29614 );
or ( n50225 , n19212 , n19213 );
not ( n19214 , RI1754c610_2);
and ( n19215 , n19214 , n50225 );
and ( n19216 , C0 , RI1754c610_2);
or ( n50226 , n19215 , n19216 );
buf ( n50227 , n50226 );
xor ( n50228 , n33964 , n34221 );
xor ( n50229 , n50228 , n34251 );
xor ( n50230 , n29727 , n39091 );
xor ( n50231 , n50230 , n36128 );
not ( n50232 , n50231 );
and ( n50233 , n50232 , n50052 );
xor ( n50234 , n50229 , n50233 );
not ( n19217 , n29614 );
and ( n19218 , n19217 , RI174bd768_821);
and ( n19219 , n50234 , n29614 );
or ( n50235 , n19218 , n19219 );
not ( n19220 , RI1754c610_2);
and ( n19221 , n19220 , n50235 );
and ( n19222 , C0 , RI1754c610_2);
or ( n50236 , n19221 , n19222 );
buf ( n50237 , n50236 );
not ( n50238 , n49596 );
xor ( n50239 , n36426 , n33935 );
xor ( n50240 , n50239 , n36287 );
and ( n50241 , n50238 , n50240 );
xor ( n50242 , n42473 , n50241 );
not ( n19223 , n29614 );
and ( n19224 , n19223 , RI174cb520_778);
and ( n19225 , n50242 , n29614 );
or ( n50243 , n19224 , n19225 );
not ( n19226 , RI1754c610_2);
and ( n19227 , n19226 , n50243 );
and ( n19228 , C0 , RI1754c610_2);
or ( n50244 , n19227 , n19228 );
buf ( n50245 , n50244 );
not ( n19229 , n27683 );
and ( n19230 , n19229 , RI19ab4dd0_2417);
and ( n19231 , RI19abe6a0_2346 , n27683 );
or ( n50246 , n19230 , n19231 );
not ( n19232 , RI1754c610_2);
and ( n19233 , n19232 , n50246 );
and ( n19234 , C0 , RI1754c610_2);
or ( n50247 , n19233 , n19234 );
buf ( n50248 , n50247 );
not ( n50249 , n41288 );
xor ( n50250 , n36127 , n39131 );
xor ( n50251 , n50250 , n39151 );
and ( n50252 , n50249 , n50251 );
xor ( n50253 , n41269 , n50252 );
not ( n19235 , n29614 );
and ( n19236 , n19235 , RI1745d8b8_1280);
and ( n19237 , n50253 , n29614 );
or ( n50254 , n19236 , n19237 );
not ( n19238 , RI1754c610_2);
and ( n19239 , n19238 , n50254 );
and ( n19240 , C0 , RI1754c610_2);
or ( n50255 , n19239 , n19240 );
buf ( n50256 , n50255 );
not ( n50257 , n50128 );
xor ( n50258 , n34796 , n37255 );
xor ( n50259 , n50258 , n41478 );
and ( n50260 , n50257 , n50259 );
xor ( n50261 , n50125 , n50260 );
not ( n19241 , n29614 );
and ( n19242 , n19241 , RI174820c8_1102);
and ( n19243 , n50261 , n29614 );
or ( n50262 , n19242 , n19243 );
not ( n19244 , RI1754c610_2);
and ( n19245 , n19244 , n50262 );
and ( n19246 , C0 , RI1754c610_2);
or ( n50263 , n19245 , n19246 );
buf ( n50264 , n50263 );
and ( n50265 , RI19a24c80_2783 , n43086 );
not ( n19247 , n43088 );
and ( n19248 , n19247 , RI19a24a28_2784);
and ( n19249 , n50265 , n43088 );
or ( n50266 , n19248 , n19249 );
not ( n19250 , RI1754c610_2);
and ( n19251 , n19250 , n50266 );
and ( n19252 , C0 , RI1754c610_2);
or ( n50267 , n19251 , n19252 );
buf ( n50268 , n50267 );
not ( n50269 , n42002 );
and ( n50270 , n50269 , n42004 );
xor ( n50271 , n42763 , n50270 );
not ( n19253 , n29614 );
and ( n19254 , n19253 , RI17477970_1153);
and ( n19255 , n50271 , n29614 );
or ( n50272 , n19254 , n19255 );
not ( n19256 , RI1754c610_2);
and ( n19257 , n19256 , n50272 );
and ( n19258 , C0 , RI1754c610_2);
or ( n50273 , n19257 , n19258 );
buf ( n50274 , n50273 );
xor ( n50275 , n35998 , n35438 );
xor ( n50276 , n50275 , n35458 );
not ( n50277 , n49190 );
and ( n50278 , n50277 , n46733 );
xor ( n50279 , n50276 , n50278 );
not ( n19259 , n29614 );
and ( n19260 , n19259 , RI1752f060_620);
and ( n19261 , n50279 , n29614 );
or ( n50280 , n19260 , n19261 );
not ( n19262 , RI1754c610_2);
and ( n19263 , n19262 , n50280 );
and ( n19264 , C0 , RI1754c610_2);
or ( n50281 , n19263 , n19264 );
buf ( n50282 , n50281 );
not ( n50283 , n40062 );
and ( n50284 , n50283 , n40064 );
xor ( n50285 , n44665 , n50284 );
not ( n19265 , n29614 );
and ( n19266 , n19265 , RI174b1a08_870);
and ( n19267 , n50285 , n29614 );
or ( n50286 , n19266 , n19267 );
not ( n19268 , RI1754c610_2);
and ( n19269 , n19268 , n50286 );
and ( n19270 , C0 , RI1754c610_2);
or ( n50287 , n19269 , n19270 );
buf ( n50288 , n50287 );
not ( n50289 , n37351 );
and ( n50290 , n50289 , n37372 );
xor ( n50291 , n48092 , n50290 );
not ( n19271 , n29614 );
and ( n19272 , n19271 , RI173f67a8_1554);
and ( n19273 , n50291 , n29614 );
or ( n50292 , n19272 , n19273 );
not ( n19274 , RI1754c610_2);
and ( n19275 , n19274 , n50292 );
and ( n19276 , C0 , RI1754c610_2);
or ( n50293 , n19275 , n19276 );
buf ( n50294 , n50293 );
buf ( n50295 , RI174adbb0_889);
buf ( n50296 , RI174b6238_848);
not ( n50297 , n44275 );
and ( n50298 , n50297 , n44277 );
xor ( n50299 , n49792 , n50298 );
not ( n19277 , n29614 );
and ( n19278 , n19277 , RI174aa0a0_907);
and ( n19279 , n50299 , n29614 );
or ( n50300 , n19278 , n19279 );
not ( n19280 , RI1754c610_2);
and ( n19281 , n19280 , n50300 );
and ( n19282 , C0 , RI1754c610_2);
or ( n50301 , n19281 , n19282 );
buf ( n50302 , n50301 );
buf ( n50303 , RI174a0668_954);
buf ( n50304 , RI174a5870_929);
not ( n50305 , n39706 );
and ( n50306 , n50305 , n44037 );
xor ( n50307 , n39703 , n50306 );
not ( n19283 , n29614 );
and ( n19284 , n19283 , RI17476c50_1157);
and ( n19285 , n50307 , n29614 );
or ( n50308 , n19284 , n19285 );
not ( n19286 , RI1754c610_2);
and ( n19287 , n19286 , n50308 );
and ( n19288 , C0 , RI1754c610_2);
or ( n50309 , n19287 , n19288 );
buf ( n50310 , n50309 );
not ( n19289 , n27683 );
and ( n19290 , n19289 , RI19abe4c0_2347);
and ( n19291 , RI19ac7250_2276 , n27683 );
or ( n50311 , n19290 , n19291 );
not ( n19292 , RI1754c610_2);
and ( n19293 , n19292 , n50311 );
and ( n19294 , C0 , RI1754c610_2);
or ( n50312 , n19293 , n19294 );
buf ( n50313 , n50312 );
not ( n50314 , n42968 );
and ( n50315 , n50314 , n42970 );
xor ( n50316 , n44290 , n50315 );
not ( n19295 , n29614 );
and ( n19296 , n19295 , RI1740f4b0_1433);
and ( n19297 , n50316 , n29614 );
or ( n50317 , n19296 , n19297 );
not ( n19298 , RI1754c610_2);
and ( n19299 , n19298 , n50317 );
and ( n19300 , C0 , RI1754c610_2);
or ( n50318 , n19299 , n19300 );
buf ( n50319 , n50318 );
not ( n50320 , n49792 );
and ( n50321 , n50320 , n44275 );
xor ( n50322 , n45399 , n50321 );
not ( n19301 , n29614 );
and ( n19302 , n19301 , RI1752dbc0_624);
and ( n19303 , n50322 , n29614 );
or ( n50323 , n19302 , n19303 );
not ( n19304 , RI1754c610_2);
and ( n19305 , n19304 , n50323 );
and ( n19306 , C0 , RI1754c610_2);
or ( n50324 , n19305 , n19306 );
buf ( n50325 , n50324 );
not ( n50326 , n47528 );
and ( n50327 , n50326 , n47530 );
xor ( n50328 , n50190 , n50327 );
not ( n19307 , n29614 );
and ( n19308 , n19307 , RI173ce128_1751);
and ( n19309 , n50328 , n29614 );
or ( n50329 , n19308 , n19309 );
not ( n19310 , RI1754c610_2);
and ( n19311 , n19310 , n50329 );
and ( n19312 , C0 , RI1754c610_2);
or ( n50330 , n19311 , n19312 );
buf ( n50331 , n50330 );
not ( n19313 , n27683 );
and ( n19314 , n19313 , RI19aa0d30_2562);
and ( n19315 , RI19aaac18_2490 , n27683 );
or ( n50332 , n19314 , n19315 );
not ( n19316 , RI1754c610_2);
and ( n19317 , n19316 , n50332 );
and ( n19318 , C0 , RI1754c610_2);
or ( n50333 , n19317 , n19318 );
buf ( n50334 , n50333 );
not ( n50335 , n45197 );
and ( n50336 , n50335 , n49898 );
xor ( n50337 , n45194 , n50336 );
not ( n19319 , n29614 );
and ( n19320 , n19319 , RI17466918_1236);
and ( n19321 , n50337 , n29614 );
or ( n50338 , n19320 , n19321 );
not ( n19322 , RI1754c610_2);
and ( n19323 , n19322 , n50338 );
and ( n19324 , C0 , RI1754c610_2);
or ( n50339 , n19323 , n19324 );
buf ( n50340 , n50339 );
not ( n50341 , n42793 );
and ( n50342 , n50341 , n44729 );
xor ( n50343 , n42790 , n50342 );
not ( n19325 , n29614 );
and ( n19326 , n19325 , RI17400528_1506);
and ( n19327 , n50343 , n29614 );
or ( n50344 , n19326 , n19327 );
not ( n19328 , RI1754c610_2);
and ( n19329 , n19328 , n50344 );
and ( n19330 , C0 , RI1754c610_2);
or ( n50345 , n19329 , n19330 );
buf ( n50346 , n50345 );
not ( n50347 , n44879 );
and ( n50348 , n50347 , n48582 );
xor ( n50349 , n44876 , n50348 );
not ( n19331 , n29614 );
and ( n19332 , n19331 , RI173a5778_1949);
and ( n19333 , n50349 , n29614 );
or ( n50350 , n19332 , n19333 );
not ( n19334 , RI1754c610_2);
and ( n19335 , n19334 , n50350 );
and ( n19336 , C0 , RI1754c610_2);
or ( n50351 , n19335 , n19336 );
buf ( n50352 , n50351 );
buf ( n50353 , RI174868f8_1080);
buf ( n50354 , RI17476908_1158);
buf ( n50355 , RI17508ac8_739);
not ( n50356 , n33283 );
and ( n50357 , n50356 , n33398 );
xor ( n50358 , n41010 , n50357 );
not ( n19337 , n29614 );
and ( n19338 , n19337 , RI173e15b0_1657);
and ( n19339 , n50358 , n29614 );
or ( n50359 , n19338 , n19339 );
not ( n19340 , RI1754c610_2);
and ( n19341 , n19340 , n50359 );
and ( n19342 , C0 , RI1754c610_2);
or ( n50360 , n19341 , n19342 );
buf ( n50361 , n50360 );
buf ( n50362 , RI174bfb80_814);
not ( n50363 , n41022 );
xor ( n50364 , n32675 , n36209 );
xor ( n50365 , n50364 , n40412 );
and ( n50366 , n50363 , n50365 );
xor ( n50367 , n41019 , n50366 );
not ( n19343 , n29614 );
and ( n19344 , n19343 , RI1748d888_1046);
and ( n19345 , n50367 , n29614 );
or ( n50368 , n19344 , n19345 );
not ( n19346 , RI1754c610_2);
and ( n19347 , n19346 , n50368 );
and ( n19348 , C0 , RI1754c610_2);
or ( n50369 , n19347 , n19348 );
buf ( n50370 , n50369 );
not ( n19349 , n27683 );
and ( n19350 , n19349 , RI19a90188_2682);
and ( n19351 , RI19a9a3b8_2610 , n27683 );
or ( n50371 , n19350 , n19351 );
not ( n19352 , RI1754c610_2);
and ( n19353 , n19352 , n50371 );
and ( n19354 , C0 , RI1754c610_2);
or ( n50372 , n19353 , n19354 );
buf ( n50373 , n50372 );
not ( n50374 , n46220 );
and ( n50375 , n50374 , n43312 );
xor ( n50376 , n46277 , n50375 );
not ( n19355 , n29614 );
and ( n19356 , n19355 , RI1740a938_1456);
and ( n19357 , n50376 , n29614 );
or ( n50377 , n19356 , n19357 );
not ( n19358 , RI1754c610_2);
and ( n19359 , n19358 , n50377 );
and ( n19360 , C0 , RI1754c610_2);
or ( n50378 , n19359 , n19360 );
buf ( n50379 , n50378 );
not ( n50380 , n44347 );
and ( n50381 , n50380 , n44349 );
xor ( n50382 , n47576 , n50381 );
not ( n19361 , n29614 );
and ( n19362 , n19361 , RI173c2ff8_1805);
and ( n19363 , n50382 , n29614 );
or ( n50383 , n19362 , n19363 );
not ( n19364 , RI1754c610_2);
and ( n19365 , n19364 , n50383 );
and ( n19366 , C0 , RI1754c610_2);
or ( n50384 , n19365 , n19366 );
buf ( n50385 , n50384 );
buf ( n50386 , RI174ab798_900);
buf ( n50387 , RI1748df18_1044);
buf ( n50388 , RI17496258_1004);
not ( n19367 , n27683 );
and ( n19368 , n19367 , RI19abc198_2367);
and ( n19369 , RI19ac46b8_2296 , n27683 );
or ( n50389 , n19368 , n19369 );
not ( n19370 , RI1754c610_2);
and ( n19371 , n19370 , n50389 );
and ( n19372 , C0 , RI1754c610_2);
or ( n50390 , n19371 , n19372 );
buf ( n50391 , n50390 );
not ( n50392 , n45856 );
and ( n50393 , n50392 , n43304 );
xor ( n50394 , n40632 , n50393 );
not ( n19373 , n29614 );
and ( n19374 , n19373 , RI17452e18_1332);
and ( n19375 , n50394 , n29614 );
or ( n50395 , n19374 , n19375 );
not ( n19376 , RI1754c610_2);
and ( n19377 , n19376 , n50395 );
and ( n19378 , C0 , RI1754c610_2);
or ( n50396 , n19377 , n19378 );
buf ( n50397 , n50396 );
buf ( n50398 , RI17485200_1087);
buf ( n50399 , RI17470008_1190);
buf ( n50400 , RI17510688_715);
xor ( n50401 , n40310 , n37869 );
xor ( n50402 , n50401 , n38948 );
xor ( n50403 , n36697 , n39655 );
xor ( n50404 , n50403 , n41125 );
not ( n50405 , n50404 );
and ( n50406 , n50405 , n46966 );
xor ( n50407 , n50402 , n50406 );
not ( n19379 , n29614 );
and ( n19380 , n19379 , RI173a43c8_1955);
and ( n19381 , n50407 , n29614 );
or ( n50408 , n19380 , n19381 );
not ( n19382 , RI1754c610_2);
and ( n19383 , n19382 , n50408 );
and ( n19384 , C0 , RI1754c610_2);
or ( n50409 , n19383 , n19384 );
buf ( n50410 , n50409 );
not ( n50411 , n44464 );
and ( n50412 , n50411 , n48535 );
xor ( n50413 , n44461 , n50412 );
not ( n19385 , n29614 );
and ( n19386 , n19385 , RI1739b9f8_1997);
and ( n19387 , n50413 , n29614 );
or ( n50414 , n19386 , n19387 );
not ( n19388 , RI1754c610_2);
and ( n19389 , n19388 , n50414 );
and ( n19390 , C0 , RI1754c610_2);
or ( n50415 , n19389 , n19390 );
buf ( n50416 , n50415 );
buf ( n50417 , RI17470698_1188);
not ( n50418 , n49492 );
and ( n50419 , n50418 , n49494 );
xor ( n50420 , n50138 , n50419 );
not ( n19391 , n29614 );
and ( n19392 , n19391 , RI1733e5f0_2137);
and ( n19393 , n50420 , n29614 );
or ( n50421 , n19392 , n19393 );
not ( n19394 , RI1754c610_2);
and ( n19395 , n19394 , n50421 );
and ( n19396 , C0 , RI1754c610_2);
or ( n50422 , n19395 , n19396 );
buf ( n50423 , n50422 );
xor ( n50424 , n42300 , n40769 );
xor ( n50425 , n50424 , n40949 );
xor ( n50426 , n34714 , n42605 );
xor ( n50427 , n50426 , n42619 );
not ( n50428 , n50427 );
xor ( n50429 , n39542 , n35842 );
xor ( n50430 , n50429 , n38401 );
and ( n50431 , n50428 , n50430 );
xor ( n50432 , n50425 , n50431 );
not ( n19397 , n29614 );
and ( n19398 , n19397 , RI1747e5b8_1120);
and ( n19399 , n50432 , n29614 );
or ( n50433 , n19398 , n19399 );
not ( n19400 , RI1754c610_2);
and ( n19401 , n19400 , n50433 );
and ( n19402 , C0 , RI1754c610_2);
or ( n50434 , n19401 , n19402 );
buf ( n50435 , n50434 );
not ( n50436 , n42133 );
and ( n50437 , n50436 , n42135 );
xor ( n50438 , n48013 , n50437 );
not ( n19403 , n29614 );
and ( n19404 , n19403 , RI17405a78_1480);
and ( n19405 , n50438 , n29614 );
or ( n50439 , n19404 , n19405 );
not ( n19406 , RI1754c610_2);
and ( n19407 , n19406 , n50439 );
and ( n19408 , C0 , RI1754c610_2);
or ( n50440 , n19407 , n19408 );
buf ( n50441 , n50440 );
xor ( n50442 , n28881 , n34517 );
xor ( n50443 , n50442 , n35911 );
not ( n50444 , n50443 );
and ( n50445 , n50444 , n48504 );
xor ( n50446 , n47173 , n50445 );
not ( n19409 , n29614 );
and ( n19410 , n19409 , RI173c9268_1775);
and ( n19411 , n50446 , n29614 );
or ( n50447 , n19410 , n19411 );
not ( n19412 , RI1754c610_2);
and ( n19413 , n19412 , n50447 );
and ( n19414 , C0 , RI1754c610_2);
or ( n50448 , n19413 , n19414 );
buf ( n50449 , n50448 );
not ( n19415 , n27683 );
and ( n19416 , n19415 , RI19a93068_2661);
and ( n19417 , RI19a9d400_2589 , n27683 );
or ( n50450 , n19416 , n19417 );
not ( n19418 , RI1754c610_2);
and ( n19419 , n19418 , n50450 );
and ( n19420 , C0 , RI1754c610_2);
or ( n50451 , n19419 , n19420 );
buf ( n50452 , n50451 );
xor ( n50453 , n33924 , n37291 );
xor ( n50454 , n50453 , n37311 );
xor ( n50455 , n41286 , n38648 );
xor ( n50456 , n50455 , n40890 );
not ( n50457 , n50456 );
and ( n50458 , n50457 , n42643 );
xor ( n50459 , n50454 , n50458 );
not ( n19421 , n29614 );
and ( n19422 , n19421 , RI173b4a48_1875);
and ( n19423 , n50459 , n29614 );
or ( n50460 , n19422 , n19423 );
not ( n19424 , RI1754c610_2);
and ( n19425 , n19424 , n50460 );
and ( n19426 , C0 , RI1754c610_2);
or ( n50461 , n19425 , n19426 );
buf ( n50462 , n50461 );
xor ( n50463 , n37700 , n40463 );
xor ( n50464 , n50463 , n41772 );
xor ( n50465 , n40497 , n41430 );
xor ( n50466 , n50465 , n36844 );
not ( n50467 , n50466 );
and ( n50468 , n50467 , n50425 );
xor ( n50469 , n50464 , n50468 );
not ( n19427 , n29614 );
and ( n19428 , n19427 , RI17461710_1261);
and ( n19429 , n50469 , n29614 );
or ( n50470 , n19428 , n19429 );
not ( n19430 , RI1754c610_2);
and ( n19431 , n19430 , n50470 );
and ( n19432 , C0 , RI1754c610_2);
or ( n50471 , n19431 , n19432 );
buf ( n50472 , n50471 );
not ( n50473 , n42278 );
and ( n50474 , n50473 , n42280 );
xor ( n50475 , n50072 , n50474 );
not ( n19433 , n29614 );
and ( n19434 , n19433 , RI174c1a70_808);
and ( n19435 , n50475 , n29614 );
or ( n50476 , n19434 , n19435 );
not ( n19436 , RI1754c610_2);
and ( n19437 , n19436 , n50476 );
and ( n19438 , C0 , RI1754c610_2);
or ( n50477 , n19437 , n19438 );
buf ( n50478 , n50477 );
xor ( n50479 , n37773 , n43994 );
xor ( n50480 , n50479 , n31213 );
xor ( n50481 , n36637 , n40412 );
xor ( n50482 , n50481 , n40437 );
not ( n50483 , n50482 );
xor ( n50484 , n41193 , n34622 );
xor ( n50485 , n50484 , n39397 );
and ( n50486 , n50483 , n50485 );
xor ( n50487 , n50480 , n50486 );
not ( n19439 , n29614 );
and ( n19440 , n19439 , RI174758a0_1163);
and ( n19441 , n50487 , n29614 );
or ( n50488 , n19440 , n19441 );
not ( n19442 , RI1754c610_2);
and ( n19443 , n19442 , n50488 );
and ( n19444 , C0 , RI1754c610_2);
or ( n50489 , n19443 , n19444 );
buf ( n50490 , n50489 );
not ( n50491 , n44945 );
and ( n50492 , n50491 , n44471 );
xor ( n50493 , n44942 , n50492 );
not ( n19445 , n29614 );
and ( n19446 , n19445 , RI17528940_640);
and ( n19447 , n50493 , n29614 );
or ( n50494 , n19446 , n19447 );
not ( n19448 , RI1754c610_2);
and ( n19449 , n19448 , n50494 );
and ( n19450 , C0 , RI1754c610_2);
or ( n50495 , n19449 , n19450 );
buf ( n50496 , n50495 );
not ( n19451 , n27683 );
and ( n19452 , n19451 , RI19a9d658_2588);
and ( n19453 , RI19aa6d48_2517 , n27683 );
or ( n50497 , n19452 , n19453 );
not ( n19454 , RI1754c610_2);
and ( n19455 , n19454 , n50497 );
and ( n19456 , C0 , RI1754c610_2);
or ( n50498 , n19455 , n19456 );
buf ( n50499 , n50498 );
not ( n19457 , n27683 );
and ( n19458 , n19457 , RI19ab6ae0_2404);
and ( n19459 , RI19abfd98_2333 , n27683 );
or ( n50500 , n19458 , n19459 );
not ( n19460 , RI1754c610_2);
and ( n19461 , n19460 , n50500 );
and ( n19462 , C0 , RI1754c610_2);
or ( n50501 , n19461 , n19462 );
buf ( n50502 , n50501 );
not ( n19463 , n27683 );
and ( n19464 , n19463 , RI19a87470_2743);
and ( n19465 , RI19aa40c0_2537 , n27683 );
or ( n50503 , n19464 , n19465 );
not ( n19466 , RI1754c610_2);
and ( n19467 , n19466 , n50503 );
and ( n19468 , C0 , RI1754c610_2);
or ( n50504 , n19467 , n19468 );
buf ( n50505 , n50504 );
not ( n50506 , n38449 );
and ( n50507 , n50506 , n46414 );
xor ( n50508 , n38446 , n50507 );
not ( n19469 , n29614 );
and ( n19470 , n19469 , RI173b7ec8_1859);
and ( n19471 , n50508 , n29614 );
or ( n50509 , n19470 , n19471 );
not ( n19472 , RI1754c610_2);
and ( n19473 , n19472 , n50509 );
and ( n19474 , C0 , RI1754c610_2);
or ( n50510 , n19473 , n19474 );
buf ( n50511 , n50510 );
not ( n50512 , n44159 );
and ( n50513 , n50512 , n44161 );
xor ( n50514 , n49604 , n50513 );
not ( n19475 , n29614 );
and ( n19476 , n19475 , RI1744a100_1375);
and ( n19477 , n50514 , n29614 );
or ( n50515 , n19476 , n19477 );
not ( n19478 , RI1754c610_2);
and ( n19479 , n19478 , n50515 );
and ( n19480 , C0 , RI1754c610_2);
or ( n50516 , n19479 , n19480 );
buf ( n50517 , n50516 );
buf ( n50518 , RI1746f978_1192);
not ( n19481 , n27683 );
and ( n19482 , n19481 , RI19a976b8_2630);
and ( n19483 , RI19aa10f0_2560 , n27683 );
or ( n50519 , n19482 , n19483 );
not ( n19484 , RI1754c610_2);
and ( n19485 , n19484 , n50519 );
and ( n19486 , C0 , RI1754c610_2);
or ( n50520 , n19485 , n19486 );
buf ( n50521 , n50520 );
buf ( n50522 , RI1746ec58_1196);
not ( n50523 , n46267 );
and ( n50524 , n50523 , n46269 );
xor ( n50525 , n41995 , n50524 );
not ( n19487 , n29614 );
and ( n19488 , n19487 , RI174affc8_878);
and ( n19489 , n50525 , n29614 );
or ( n50526 , n19488 , n19489 );
not ( n19490 , RI1754c610_2);
and ( n19491 , n19490 , n50526 );
and ( n19492 , C0 , RI1754c610_2);
or ( n50527 , n19491 , n19492 );
buf ( n50528 , n50527 );
xor ( n50529 , n42549 , n37421 );
xor ( n50530 , n50529 , n42605 );
not ( n50531 , n50530 );
xor ( n50532 , n42032 , n41049 );
xor ( n50533 , n50532 , n41504 );
and ( n50534 , n50531 , n50533 );
xor ( n50535 , n46140 , n50534 );
not ( n19493 , n29614 );
and ( n19494 , n19493 , RI1750e270_722);
and ( n19495 , n50535 , n29614 );
or ( n50536 , n19494 , n19495 );
not ( n19496 , RI1754c610_2);
and ( n19497 , n19496 , n50536 );
and ( n19498 , C0 , RI1754c610_2);
or ( n50537 , n19497 , n19498 );
buf ( n50538 , n50537 );
not ( n50539 , n45794 );
xor ( n50540 , n38478 , n39771 );
xor ( n50541 , n50540 , n39791 );
and ( n50542 , n50539 , n50541 );
xor ( n50543 , n45791 , n50542 );
not ( n19499 , n29614 );
and ( n19500 , n19499 , RI173bb690_1842);
and ( n19501 , n50543 , n29614 );
or ( n50544 , n19500 , n19501 );
not ( n19502 , RI1754c610_2);
and ( n19503 , n19502 , n50544 );
and ( n19504 , C0 , RI1754c610_2);
or ( n50545 , n19503 , n19504 );
buf ( n50546 , n50545 );
not ( n50547 , n39415 );
and ( n50548 , n50547 , n39417 );
xor ( n50549 , n48770 , n50548 );
not ( n19505 , n29614 );
and ( n19506 , n19505 , RI174a6590_925);
and ( n19507 , n50549 , n29614 );
or ( n50550 , n19506 , n19507 );
not ( n19508 , RI1754c610_2);
and ( n19509 , n19508 , n50550 );
and ( n19510 , C0 , RI1754c610_2);
or ( n50551 , n19509 , n19510 );
buf ( n50552 , n50551 );
not ( n50553 , n47586 );
and ( n50554 , n50553 , n45954 );
xor ( n50555 , n44976 , n50554 );
not ( n19511 , n29614 );
and ( n19512 , n19511 , RI17466c60_1235);
and ( n19513 , n50555 , n29614 );
or ( n50556 , n19512 , n19513 );
not ( n19514 , RI1754c610_2);
and ( n19515 , n19514 , n50556 );
and ( n19516 , C0 , RI1754c610_2);
or ( n50557 , n19515 , n19516 );
buf ( n50558 , n50557 );
not ( n50559 , n45360 );
xor ( n50560 , n33494 , n40360 );
xor ( n50561 , n50560 , n35176 );
and ( n50562 , n50559 , n50561 );
xor ( n50563 , n44338 , n50562 );
not ( n19517 , n29614 );
and ( n19518 , n19517 , RI17395440_2028);
and ( n19519 , n50563 , n29614 );
or ( n50564 , n19518 , n19519 );
not ( n19520 , RI1754c610_2);
and ( n19521 , n19520 , n50564 );
and ( n19522 , C0 , RI1754c610_2);
or ( n50565 , n19521 , n19522 );
buf ( n50566 , n50565 );
not ( n50567 , n50533 );
and ( n50568 , n50567 , n46135 );
xor ( n50569 , n50530 , n50568 );
not ( n19523 , n29614 );
and ( n19524 , n19523 , RI175255b0_650);
and ( n19525 , n50569 , n29614 );
or ( n50570 , n19524 , n19525 );
not ( n19526 , RI1754c610_2);
and ( n19527 , n19526 , n50570 );
and ( n19528 , C0 , RI1754c610_2);
or ( n50571 , n19527 , n19528 );
buf ( n50572 , n50571 );
not ( n19529 , n27683 );
and ( n19530 , n19529 , RI19aca298_2254);
and ( n19531 , RI19a85760_2756 , n27683 );
or ( n50573 , n19530 , n19531 );
not ( n19532 , RI1754c610_2);
and ( n19533 , n19532 , n50573 );
and ( n19534 , C0 , RI1754c610_2);
or ( n50574 , n19533 , n19534 );
buf ( n50575 , n50574 );
buf ( n50576 , RI17471070_1185);
buf ( n50577 , RI17500a58_758);
buf ( n50578 , RI1746aab8_1216);
xor ( n50579 , n38855 , n41125 );
xor ( n50580 , n50579 , n31506 );
not ( n50581 , n49028 );
and ( n50582 , n50581 , n47778 );
xor ( n50583 , n50580 , n50582 );
not ( n19535 , n29614 );
and ( n19536 , n19535 , RI17472ab0_1177);
and ( n19537 , n50583 , n29614 );
or ( n50584 , n19536 , n19537 );
not ( n19538 , RI1754c610_2);
and ( n19539 , n19538 , n50584 );
and ( n19540 , C0 , RI1754c610_2);
or ( n50585 , n19539 , n19540 );
buf ( n50586 , n50585 );
not ( n50587 , n46427 );
and ( n50588 , n50587 , n46429 );
xor ( n50589 , n49237 , n50588 );
not ( n19541 , n29614 );
and ( n19542 , n19541 , RI174493e0_1379);
and ( n19543 , n50589 , n29614 );
or ( n50590 , n19542 , n19543 );
not ( n19544 , RI1754c610_2);
and ( n19545 , n19544 , n50590 );
and ( n19546 , C0 , RI1754c610_2);
or ( n50591 , n19545 , n19546 );
buf ( n50592 , n50591 );
not ( n50593 , n44575 );
and ( n50594 , n50593 , n48838 );
xor ( n50595 , n44572 , n50594 );
not ( n19547 , n29614 );
and ( n19548 , n19547 , RI174b6238_848);
and ( n19549 , n50595 , n29614 );
or ( n50596 , n19548 , n19549 );
not ( n19550 , RI1754c610_2);
and ( n19551 , n19550 , n50596 );
and ( n19552 , C0 , RI1754c610_2);
or ( n50597 , n19551 , n19552 );
buf ( n50598 , n50597 );
not ( n50599 , n46500 );
and ( n50600 , n50599 , n45224 );
xor ( n50601 , n46497 , n50600 );
not ( n19553 , n29614 );
and ( n19554 , n19553 , RI1745ec68_1274);
and ( n19555 , n50601 , n29614 );
or ( n50602 , n19554 , n19555 );
not ( n19556 , RI1754c610_2);
and ( n19557 , n19556 , n50602 );
and ( n19558 , C0 , RI1754c610_2);
or ( n50603 , n19557 , n19558 );
buf ( n50604 , n50603 );
not ( n19559 , n27683 );
and ( n19560 , n19559 , RI19aad648_2472);
and ( n19561 , RI19ab73c8_2400 , n27683 );
or ( n50605 , n19560 , n19561 );
not ( n19562 , RI1754c610_2);
and ( n19563 , n19562 , n50605 );
and ( n19564 , C0 , RI1754c610_2);
or ( n50606 , n19563 , n19564 );
buf ( n50607 , n50606 );
not ( n50608 , n45385 );
and ( n50609 , n50608 , n45387 );
xor ( n50610 , n41717 , n50609 );
not ( n19565 , n29614 );
and ( n19566 , n19565 , RI173bd760_1832);
and ( n19567 , n50610 , n29614 );
or ( n50611 , n19566 , n19567 );
not ( n19568 , RI1754c610_2);
and ( n19569 , n19568 , n50611 );
and ( n19570 , C0 , RI1754c610_2);
or ( n50612 , n19569 , n19570 );
buf ( n50613 , n50612 );
and ( n50614 , RI1754ae28_53 , n34844 );
buf ( n50615 , n50614 );
not ( n19571 , n34859 );
and ( n19572 , n19571 , n50615 );
and ( n19573 , RI1754ae28_53 , n34859 );
or ( n50616 , n19572 , n19573 );
not ( n19574 , RI19a22f70_2797);
and ( n19575 , n19574 , n50616 );
and ( n19576 , C0 , RI19a22f70_2797);
or ( n50617 , n19575 , n19576 );
not ( n19577 , n27683 );
and ( n19578 , n19577 , RI19a23678_2793);
and ( n19579 , n50617 , n27683 );
or ( n50618 , n19578 , n19579 );
not ( n19580 , RI1754c610_2);
and ( n19581 , n19580 , n50618 );
and ( n19582 , C0 , RI1754c610_2);
or ( n50619 , n19581 , n19582 );
buf ( n50620 , n50619 );
not ( n19583 , n27683 );
and ( n19584 , n19583 , RI19a9b678_2602);
and ( n19585 , RI19aa4cf0_2531 , n27683 );
or ( n50621 , n19584 , n19585 );
not ( n19586 , RI1754c610_2);
and ( n19587 , n19586 , n50621 );
and ( n19588 , C0 , RI1754c610_2);
or ( n50622 , n19587 , n19588 );
buf ( n50623 , n50622 );
not ( n19589 , n27683 );
and ( n19590 , n19589 , RI19a86750_2749);
and ( n19591 , RI19a83b40_2768 , n27683 );
or ( n50624 , n19590 , n19591 );
not ( n19592 , RI1754c610_2);
and ( n19593 , n19592 , n50624 );
and ( n19594 , C0 , RI1754c610_2);
or ( n50625 , n19593 , n19594 );
buf ( n50626 , n50625 );
not ( n50627 , n49716 );
and ( n50628 , n50627 , n46678 );
xor ( n50629 , n45087 , n50628 );
not ( n19595 , n29614 );
and ( n19596 , n19595 , RI17337318_2172);
and ( n19597 , n50629 , n29614 );
or ( n50630 , n19596 , n19597 );
not ( n19598 , RI1754c610_2);
and ( n19599 , n19598 , n50630 );
and ( n19600 , C0 , RI1754c610_2);
or ( n50631 , n19599 , n19600 );
buf ( n50632 , n50631 );
not ( n50633 , n43507 );
and ( n50634 , n50633 , n48390 );
xor ( n50635 , n42271 , n50634 );
not ( n19601 , n29614 );
and ( n19602 , n19601 , RI17522c70_658);
and ( n19603 , n50635 , n29614 );
or ( n50636 , n19602 , n19603 );
not ( n19604 , RI1754c610_2);
and ( n19605 , n19604 , n50636 );
and ( n19606 , C0 , RI1754c610_2);
or ( n50637 , n19605 , n19606 );
buf ( n50638 , n50637 );
not ( n50639 , n42086 );
and ( n50640 , n50639 , n40693 );
xor ( n50641 , n42083 , n50640 );
not ( n19607 , n29614 );
and ( n19608 , n19607 , RI173df4e0_1667);
and ( n19609 , n50641 , n29614 );
or ( n50642 , n19608 , n19609 );
not ( n19610 , RI1754c610_2);
and ( n19611 , n19610 , n50642 );
and ( n19612 , C0 , RI1754c610_2);
or ( n50643 , n19611 , n19612 );
buf ( n50644 , n50643 );
buf ( n50645 , RI17498328_994);
buf ( n50646 , RI17461710_1261);
buf ( n50647 , RI174bc2c8_825);
not ( n50648 , n45262 );
and ( n50649 , n50648 , n45299 );
xor ( n50650 , n39479 , n50649 );
not ( n19613 , n29614 );
and ( n19614 , n19613 , RI17332110_2197);
and ( n19615 , n50650 , n29614 );
or ( n50651 , n19614 , n19615 );
not ( n19616 , RI1754c610_2);
and ( n19617 , n19616 , n50651 );
and ( n19618 , C0 , RI1754c610_2);
or ( n50652 , n19617 , n19618 );
buf ( n50653 , n50652 );
xor ( n50654 , n38162 , n35494 );
xor ( n50655 , n50654 , n35514 );
not ( n50656 , n50655 );
and ( n50657 , n50656 , n42702 );
xor ( n50658 , n37105 , n50657 );
not ( n19619 , n29614 );
and ( n19620 , n19619 , RI17515e30_698);
and ( n19621 , n50658 , n29614 );
or ( n50659 , n19620 , n19621 );
not ( n19622 , RI1754c610_2);
and ( n19623 , n19622 , n50659 );
and ( n19624 , C0 , RI1754c610_2);
or ( n50660 , n19623 , n19624 );
buf ( n50661 , n50660 );
buf ( n50662 , RI174c8190_788);
not ( n50663 , n47761 );
and ( n50664 , n50663 , n46372 );
xor ( n50665 , n45284 , n50664 );
not ( n19625 , n29614 );
and ( n19626 , n19625 , RI1740ead8_1436);
and ( n19627 , n50665 , n29614 );
or ( n50666 , n19626 , n19627 );
not ( n19628 , RI1754c610_2);
and ( n19629 , n19628 , n50666 );
and ( n19630 , C0 , RI1754c610_2);
or ( n50667 , n19629 , n19630 );
buf ( n50668 , n50667 );
not ( n50669 , n46069 );
and ( n50670 , n50669 , n46071 );
xor ( n50671 , n43655 , n50670 );
not ( n19631 , n29614 );
and ( n19632 , n19631 , RI17534808_603);
and ( n19633 , n50671 , n29614 );
or ( n50672 , n19632 , n19633 );
not ( n19634 , RI1754c610_2);
and ( n19635 , n19634 , n50672 );
and ( n19636 , C0 , RI1754c610_2);
or ( n50673 , n19635 , n19636 );
buf ( n50674 , n50673 );
not ( n50675 , n50229 );
and ( n50676 , n50675 , n50231 );
xor ( n50677 , n50057 , n50676 );
not ( n19637 , n29614 );
and ( n19638 , n19637 , RI174ad520_891);
and ( n19639 , n50677 , n29614 );
or ( n50678 , n19638 , n19639 );
not ( n19640 , RI1754c610_2);
and ( n19641 , n19640 , n50678 );
and ( n19642 , C0 , RI1754c610_2);
or ( n50679 , n19641 , n19642 );
buf ( n50680 , n50679 );
not ( n50681 , n39792 );
and ( n50682 , n50681 , n39818 );
xor ( n50683 , n47961 , n50682 );
not ( n19643 , n29614 );
and ( n19644 , n19643 , RI173e5408_1638);
and ( n19645 , n50683 , n29614 );
or ( n50684 , n19644 , n19645 );
not ( n19646 , RI1754c610_2);
and ( n19647 , n19646 , n50684 );
and ( n19648 , C0 , RI1754c610_2);
or ( n50685 , n19647 , n19648 );
buf ( n50686 , n50685 );
buf ( n50687 , RI174909c0_1031);
buf ( n50688 , RI1748aa98_1060);
buf ( n50689 , RI17508078_741);
not ( n50690 , n42692 );
xor ( n50691 , n37853 , n35128 );
xor ( n50692 , n50691 , n36917 );
and ( n50693 , n50690 , n50692 );
xor ( n50694 , n36253 , n50693 );
not ( n19649 , n29614 );
and ( n19650 , n19649 , RI174cc498_775);
and ( n19651 , n50694 , n29614 );
or ( n50695 , n19650 , n19651 );
not ( n19652 , RI1754c610_2);
and ( n19653 , n19652 , n50695 );
and ( n19654 , C0 , RI1754c610_2);
or ( n50696 , n19653 , n19654 );
buf ( n50697 , n50696 );
not ( n19655 , n27683 );
and ( n19656 , n19655 , RI19a8f648_2687);
and ( n19657 , RI19a99698_2616 , n27683 );
or ( n50698 , n19656 , n19657 );
not ( n19658 , RI1754c610_2);
and ( n19659 , n19658 , n50698 );
and ( n19660 , C0 , RI1754c610_2);
or ( n50699 , n19659 , n19660 );
buf ( n50700 , n50699 );
not ( n50701 , n49512 );
and ( n50702 , n50701 , n49514 );
xor ( n50703 , n49588 , n50702 );
not ( n19661 , n29614 );
and ( n19662 , n19661 , RI173dbd18_1684);
and ( n19663 , n50703 , n29614 );
or ( n50704 , n19662 , n19663 );
not ( n19664 , RI1754c610_2);
and ( n19665 , n19664 , n50704 );
and ( n19666 , C0 , RI1754c610_2);
or ( n50705 , n19665 , n19666 );
buf ( n50706 , n50705 );
buf ( n50707 , RI1746c1b0_1209);
not ( n19667 , n34859 );
and ( n19668 , n19667 , C0 );
and ( n19669 , RI1754a888_65 , n34859 );
or ( n50708 , n19668 , n19669 );
not ( n19670 , RI19a22f70_2797);
and ( n19671 , n19670 , n50708 );
and ( n19672 , C0 , RI19a22f70_2797);
or ( n50709 , n19671 , n19672 );
not ( n19673 , n27683 );
and ( n19674 , n19673 , RI19ac1d78_2315);
and ( n19675 , n50709 , n27683 );
or ( n50710 , n19674 , n19675 );
not ( n19676 , RI1754c610_2);
and ( n19677 , n19676 , n50710 );
and ( n19678 , C0 , RI1754c610_2);
or ( n50711 , n19677 , n19678 );
buf ( n50712 , n50711 );
xor ( n50713 , n40569 , n37048 );
xor ( n50714 , n50713 , n36772 );
not ( n50715 , n50480 );
and ( n50716 , n50715 , n50482 );
xor ( n50717 , n50714 , n50716 );
not ( n19679 , n29614 );
and ( n19680 , n19679 , RI17466fa8_1234);
and ( n19681 , n50717 , n29614 );
or ( n50718 , n19680 , n19681 );
not ( n19682 , RI1754c610_2);
and ( n19683 , n19682 , n50718 );
and ( n19684 , C0 , RI1754c610_2);
or ( n50719 , n19683 , n19684 );
buf ( n50720 , n50719 );
not ( n50721 , n43589 );
and ( n50722 , n50721 , n49078 );
xor ( n50723 , n43586 , n50722 );
not ( n19685 , n29614 );
and ( n19686 , n19685 , RI173c0be0_1816);
and ( n19687 , n50723 , n29614 );
or ( n50724 , n19686 , n19687 );
not ( n19688 , RI1754c610_2);
and ( n19689 , n19688 , n50724 );
and ( n19690 , C0 , RI1754c610_2);
or ( n50725 , n19689 , n19690 );
buf ( n50726 , n50725 );
xor ( n50727 , n35637 , n34669 );
xor ( n50728 , n50727 , n31831 );
not ( n50729 , n50728 );
and ( n50730 , n50729 , n43439 );
xor ( n50731 , n40320 , n50730 );
not ( n19691 , n29614 );
and ( n19692 , n19691 , RI17484eb8_1088);
and ( n19693 , n50731 , n29614 );
or ( n50732 , n19692 , n19693 );
not ( n19694 , RI1754c610_2);
and ( n19695 , n19694 , n50732 );
and ( n19696 , C0 , RI1754c610_2);
or ( n50733 , n19695 , n19696 );
buf ( n50734 , n50733 );
not ( n50735 , n48504 );
and ( n50736 , n50735 , n47168 );
xor ( n50737 , n50443 , n50736 );
not ( n19697 , n29614 );
and ( n19698 , n19697 , RI1740e100_1439);
and ( n19699 , n50737 , n29614 );
or ( n50738 , n19698 , n19699 );
not ( n19700 , RI1754c610_2);
and ( n19701 , n19700 , n50738 );
and ( n19702 , C0 , RI1754c610_2);
or ( n50739 , n19701 , n19702 );
buf ( n50740 , n50739 );
xor ( n50741 , n40741 , n31925 );
xor ( n50742 , n50741 , n34475 );
not ( n50743 , n50742 );
and ( n50744 , n50743 , n45529 );
xor ( n50745 , n46566 , n50744 );
not ( n19703 , n29614 );
and ( n19704 , n19703 , RI173ea958_1612);
and ( n19705 , n50745 , n29614 );
or ( n50746 , n19704 , n19705 );
not ( n19706 , RI1754c610_2);
and ( n19707 , n19706 , n50746 );
and ( n19708 , C0 , RI1754c610_2);
or ( n50747 , n19707 , n19708 );
buf ( n50748 , n50747 );
not ( n50749 , n40916 );
and ( n50750 , n50749 , n47552 );
xor ( n50751 , n40903 , n50750 );
not ( n19709 , n29614 );
and ( n19710 , n19709 , RI17457648_1310);
and ( n19711 , n50751 , n29614 );
or ( n50752 , n19710 , n19711 );
not ( n19712 , RI1754c610_2);
and ( n19713 , n19712 , n50752 );
and ( n19714 , C0 , RI1754c610_2);
or ( n50753 , n19713 , n19714 );
buf ( n50754 , n50753 );
xor ( n50755 , n35437 , n32663 );
xor ( n50756 , n50755 , n32715 );
not ( n50757 , n50756 );
and ( n50758 , n50757 , n44224 );
xor ( n50759 , n45557 , n50758 );
not ( n19715 , n29614 );
and ( n19716 , n19715 , RI17498d00_991);
and ( n19717 , n50759 , n29614 );
or ( n50760 , n19716 , n19717 );
not ( n19718 , RI1754c610_2);
and ( n19719 , n19718 , n50760 );
and ( n19720 , C0 , RI1754c610_2);
or ( n50761 , n19719 , n19720 );
buf ( n50762 , n50761 );
buf ( n50763 , RI17472ab0_1177);
buf ( n50764 , RI174620e8_1258);
not ( n19721 , n27683 );
and ( n19722 , n19721 , RI19aaa330_2494);
and ( n19723 , RI19ab4380_2422 , n27683 );
or ( n50765 , n19722 , n19723 );
not ( n19724 , RI1754c610_2);
and ( n19725 , n19724 , n50765 );
and ( n19726 , C0 , RI1754c610_2);
or ( n50766 , n19725 , n19726 );
buf ( n50767 , n50766 );
not ( n50768 , n44953 );
and ( n50769 , n50768 , n50072 );
xor ( n50770 , n42283 , n50769 );
not ( n19727 , n29614 );
and ( n19728 , n19727 , RI1744d238_1360);
and ( n19729 , n50770 , n29614 );
or ( n50771 , n19728 , n19729 );
not ( n19730 , RI1754c610_2);
and ( n19731 , n19730 , n50771 );
and ( n19732 , C0 , RI1754c610_2);
or ( n50772 , n19731 , n19732 );
buf ( n50773 , n50772 );
not ( n50774 , n47109 );
and ( n50775 , n50774 , n44193 );
xor ( n50776 , n42206 , n50775 );
not ( n19733 , n29614 );
and ( n19734 , n19733 , RI174c7218_791);
and ( n19735 , n50776 , n29614 );
or ( n50777 , n19734 , n19735 );
not ( n19736 , RI1754c610_2);
and ( n19737 , n19736 , n50777 );
and ( n19738 , C0 , RI1754c610_2);
or ( n50778 , n19737 , n19738 );
buf ( n50779 , n50778 );
not ( n50780 , n49566 );
xor ( n50781 , n33647 , n35069 );
xor ( n50782 , n50781 , n41854 );
and ( n50783 , n50780 , n50782 );
xor ( n50784 , n49563 , n50783 );
not ( n19739 , n29614 );
and ( n19740 , n19739 , RI17501ef8_754);
and ( n19741 , n50784 , n29614 );
or ( n50785 , n19740 , n19741 );
not ( n19742 , RI1754c610_2);
and ( n19743 , n19742 , n50785 );
and ( n19744 , C0 , RI1754c610_2);
or ( n50786 , n19743 , n19744 );
buf ( n50787 , n50786 );
xor ( n50788 , n42023 , n41049 );
xor ( n50789 , n50788 , n41504 );
not ( n50790 , n44831 );
and ( n50791 , n50790 , n42832 );
xor ( n50792 , n50789 , n50791 );
not ( n19745 , n29614 );
and ( n19746 , n19745 , RI17391930_2046);
and ( n19747 , n50792 , n29614 );
or ( n50793 , n19746 , n19747 );
not ( n19748 , RI1754c610_2);
and ( n19749 , n19748 , n50793 );
and ( n19750 , C0 , RI1754c610_2);
or ( n50794 , n19749 , n19750 );
buf ( n50795 , n50794 );
not ( n50796 , n42095 );
and ( n50797 , n50796 , n42097 );
xor ( n50798 , n48868 , n50797 );
not ( n19751 , n29614 );
and ( n19752 , n19751 , RI17444ef8_1400);
and ( n19753 , n50798 , n29614 );
or ( n50799 , n19752 , n19753 );
not ( n19754 , RI1754c610_2);
and ( n19755 , n19754 , n50799 );
and ( n19756 , C0 , RI1754c610_2);
or ( n50800 , n19755 , n19756 );
buf ( n50801 , n50800 );
not ( n50802 , n42345 );
and ( n50803 , n50802 , n42347 );
xor ( n50804 , n49456 , n50803 );
not ( n19757 , n29614 );
and ( n19758 , n19757 , RI173e2960_1651);
and ( n19759 , n50804 , n29614 );
or ( n50805 , n19758 , n19759 );
not ( n19760 , RI1754c610_2);
and ( n19761 , n19760 , n50805 );
and ( n19762 , C0 , RI1754c610_2);
or ( n50806 , n19761 , n19762 );
buf ( n50807 , n50806 );
not ( n19763 , n27683 );
and ( n19764 , n19763 , RI19aa1d20_2554);
and ( n19765 , RI19aabcf8_2483 , n27683 );
or ( n50808 , n19764 , n19765 );
not ( n19766 , RI1754c610_2);
and ( n19767 , n19766 , n50808 );
and ( n19768 , C0 , RI1754c610_2);
or ( n50809 , n19767 , n19768 );
buf ( n50810 , n50809 );
xor ( n50811 , n40205 , n34041 );
xor ( n50812 , n50811 , n41934 );
not ( n50813 , n50812 );
and ( n50814 , n50813 , n48612 );
xor ( n50815 , n46817 , n50814 );
not ( n19769 , n29614 );
and ( n19770 , n19769 , RI173e6b00_1631);
and ( n19771 , n50815 , n29614 );
or ( n50816 , n19770 , n19771 );
not ( n19772 , RI1754c610_2);
and ( n19773 , n19772 , n50816 );
and ( n19774 , C0 , RI1754c610_2);
or ( n50817 , n19773 , n19774 );
buf ( n50818 , n50817 );
buf ( n50819 , RI174ce388_769);
buf ( n50820 , RI174b6580_847);
xor ( n50821 , n37622 , n40319 );
xor ( n50822 , n50821 , n40149 );
not ( n50823 , n41602 );
and ( n50824 , n50823 , n41623 );
xor ( n50825 , n50822 , n50824 );
not ( n19775 , n29614 );
and ( n19776 , n19775 , RI174a9038_912);
and ( n19777 , n50825 , n29614 );
or ( n50826 , n19776 , n19777 );
not ( n19778 , RI1754c610_2);
and ( n19779 , n19778 , n50826 );
and ( n19780 , C0 , RI1754c610_2);
or ( n50827 , n19779 , n19780 );
buf ( n50828 , n50827 );
buf ( n50829 , RI174a0320_955);
buf ( n50830 , RI1748cb68_1050);
not ( n19781 , n27683 );
and ( n19782 , n19781 , RI19abb298_2373);
and ( n19783 , RI19ac3b00_2301 , n27683 );
or ( n50831 , n19782 , n19783 );
not ( n19784 , RI1754c610_2);
and ( n19785 , n19784 , n50831 );
and ( n19786 , C0 , RI1754c610_2);
or ( n50832 , n19785 , n19786 );
buf ( n50833 , n50832 );
buf ( n50834 , RI1748ade0_1059);
buf ( n50835 , RI174d1208_760);
buf ( n50836 , RI1747b138_1136);
buf ( n50837 , RI17464ed8_1244);
not ( n50838 , n44618 );
and ( n50839 , n50838 , n48039 );
xor ( n50840 , n44615 , n50839 );
not ( n19787 , n29614 );
and ( n19788 , n19787 , RI174672f0_1233);
and ( n19789 , n50840 , n29614 );
or ( n50841 , n19788 , n19789 );
not ( n19790 , RI1754c610_2);
and ( n19791 , n19790 , n50841 );
and ( n19792 , C0 , RI1754c610_2);
or ( n50842 , n19791 , n19792 );
buf ( n50843 , n50842 );
buf ( n50844 , RI174b2a70_865);
not ( n19793 , n27683 );
and ( n19794 , n19793 , RI19a89018_2731);
and ( n19795 , RI19a93068_2661 , n27683 );
or ( n50845 , n19794 , n19795 );
not ( n19796 , RI1754c610_2);
and ( n19797 , n19796 , n50845 );
and ( n19798 , C0 , RI1754c610_2);
or ( n50846 , n19797 , n19798 );
buf ( n50847 , n50846 );
buf ( n50848 , RI174a3e30_937);
buf ( n50849 , RI17464500_1247);
not ( n19799 , n27683 );
and ( n19800 , n19799 , RI19aa9430_2501);
and ( n19801 , RI19ab3138_2431 , n27683 );
or ( n50850 , n19800 , n19801 );
not ( n19802 , RI1754c610_2);
and ( n19803 , n19802 , n50850 );
and ( n19804 , C0 , RI1754c610_2);
or ( n50851 , n19803 , n19804 );
buf ( n50852 , n50851 );
xor ( n50853 , n33796 , n39414 );
xor ( n50854 , n50853 , n37186 );
not ( n50855 , n50854 );
and ( n50856 , n50855 , n43709 );
xor ( n50857 , n50180 , n50856 );
not ( n19805 , n29614 );
and ( n19806 , n19805 , RI174a51e0_931);
and ( n19807 , n50857 , n29614 );
or ( n50858 , n19806 , n19807 );
not ( n19808 , RI1754c610_2);
and ( n19809 , n19808 , n50858 );
and ( n19810 , C0 , RI1754c610_2);
or ( n50859 , n19809 , n19810 );
buf ( n50860 , n50859 );
not ( n50861 , n42643 );
and ( n50862 , n50861 , n42645 );
xor ( n50863 , n50456 , n50862 );
not ( n19811 , n29614 );
and ( n19812 , n19811 , RI173b6e60_1864);
and ( n19813 , n50863 , n29614 );
or ( n50864 , n19812 , n19813 );
not ( n19814 , RI1754c610_2);
and ( n19815 , n19814 , n50864 );
and ( n19816 , C0 , RI1754c610_2);
or ( n50865 , n19815 , n19816 );
buf ( n50866 , n50865 );
not ( n50867 , n37916 );
and ( n50868 , n50867 , n40664 );
xor ( n50869 , n37875 , n50868 );
not ( n19817 , n29614 );
and ( n19818 , n19817 , RI173fee30_1513);
and ( n19819 , n50869 , n29614 );
or ( n50870 , n19818 , n19819 );
not ( n19820 , RI1754c610_2);
and ( n19821 , n19820 , n50870 );
and ( n19822 , C0 , RI1754c610_2);
or ( n50871 , n19821 , n19822 );
buf ( n50872 , n50871 );
not ( n50873 , n44214 );
and ( n50874 , n50873 , n45269 );
xor ( n50875 , n43242 , n50874 );
not ( n19823 , n29614 );
and ( n19824 , n19823 , RI174a72b0_921);
and ( n19825 , n50875 , n29614 );
or ( n50876 , n19824 , n19825 );
not ( n19826 , RI1754c610_2);
and ( n19827 , n19826 , n50876 );
and ( n19828 , C0 , RI1754c610_2);
or ( n50877 , n19827 , n19828 );
buf ( n50878 , n50877 );
not ( n50879 , n48732 );
and ( n50880 , n50879 , n48734 );
xor ( n50881 , n50030 , n50880 );
not ( n19829 , n29614 );
and ( n19830 , n19829 , RI1747ec48_1118);
and ( n19831 , n50881 , n29614 );
or ( n50882 , n19830 , n19831 );
not ( n19832 , RI1754c610_2);
and ( n19833 , n19832 , n50882 );
and ( n19834 , C0 , RI1754c610_2);
or ( n50883 , n19833 , n19834 );
buf ( n50884 , n50883 );
and ( n50885 , RI19a240c8_2788 , n43086 );
not ( n19835 , n43088 );
and ( n19836 , n19835 , RI19a23e70_2789);
and ( n19837 , n50885 , n43088 );
or ( n50886 , n19836 , n19837 );
not ( n19838 , RI1754c610_2);
and ( n19839 , n19838 , n50886 );
and ( n19840 , C0 , RI1754c610_2);
or ( n50887 , n19839 , n19840 );
buf ( n50888 , n50887 );
not ( n50889 , n49901 );
and ( n50890 , n50889 , n45192 );
xor ( n50891 , n49898 , n50890 );
not ( n19841 , n29614 );
and ( n19842 , n19841 , RI17483b08_1094);
and ( n19843 , n50891 , n29614 );
or ( n50892 , n19842 , n19843 );
not ( n19844 , RI1754c610_2);
and ( n19845 , n19844 , n50892 );
and ( n19846 , C0 , RI1754c610_2);
or ( n50893 , n19845 , n19846 );
buf ( n50894 , n50893 );
not ( n50895 , n50464 );
and ( n50896 , n50895 , n50466 );
xor ( n50897 , n50430 , n50896 );
not ( n19847 , n29614 );
and ( n19848 , n19847 , RI1749b7a8_978);
and ( n19849 , n50897 , n29614 );
or ( n50898 , n19848 , n19849 );
not ( n19850 , RI1754c610_2);
and ( n19851 , n19850 , n50898 );
and ( n19852 , C0 , RI1754c610_2);
or ( n50899 , n19851 , n19852 );
buf ( n50900 , n50899 );
not ( n50901 , n48633 );
and ( n50902 , n50901 , n44930 );
xor ( n50903 , n48630 , n50902 );
not ( n19853 , n29614 );
and ( n19854 , n19853 , RI174022b0_1497);
and ( n19855 , n50903 , n29614 );
or ( n50904 , n19854 , n19855 );
not ( n19856 , RI1754c610_2);
and ( n19857 , n19856 , n50904 );
and ( n19858 , C0 , RI1754c610_2);
or ( n50905 , n19857 , n19858 );
buf ( n50906 , n50905 );
not ( n19859 , n27683 );
and ( n19860 , n19859 , RI19ac0860_2327);
and ( n19861 , RI19ac9b90_2257 , n27683 );
or ( n50907 , n19860 , n19861 );
not ( n19862 , RI1754c610_2);
and ( n19863 , n19862 , n50907 );
and ( n19864 , C0 , RI1754c610_2);
or ( n50908 , n19863 , n19864 );
buf ( n50909 , n50908 );
not ( n50910 , n45846 );
and ( n50911 , n50910 , n45848 );
xor ( n50912 , n44891 , n50911 );
not ( n19865 , n29614 );
and ( n19866 , n19865 , RI1744ec78_1352);
and ( n19867 , n50912 , n29614 );
or ( n50913 , n19866 , n19867 );
not ( n19868 , RI1754c610_2);
and ( n19869 , n19868 , n50913 );
and ( n19870 , C0 , RI1754c610_2);
or ( n50914 , n19869 , n19870 );
buf ( n50915 , n50914 );
not ( n50916 , n37105 );
and ( n50917 , n50916 , n50655 );
xor ( n50918 , n37054 , n50917 );
not ( n19871 , n29614 );
and ( n19872 , n19871 , RI174ce388_769);
and ( n19873 , n50918 , n29614 );
or ( n50919 , n19872 , n19873 );
not ( n19874 , RI1754c610_2);
and ( n19875 , n19874 , n50919 );
and ( n19876 , C0 , RI1754c610_2);
or ( n50920 , n19875 , n19876 );
buf ( n50921 , n50920 );
not ( n19877 , n27683 );
and ( n19878 , n19877 , RI19ab4bf0_2418);
and ( n19879 , RI19abe4c0_2347 , n27683 );
or ( n50922 , n19878 , n19879 );
not ( n19880 , RI1754c610_2);
and ( n19881 , n19880 , n50922 );
and ( n19882 , C0 , RI1754c610_2);
or ( n50923 , n19881 , n19882 );
buf ( n50924 , n50923 );
not ( n50925 , n45415 );
and ( n50926 , n50925 , n45417 );
xor ( n50927 , n49665 , n50926 );
not ( n19883 , n29614 );
and ( n19884 , n19883 , RI17467638_1232);
and ( n19885 , n50927 , n29614 );
or ( n50928 , n19884 , n19885 );
not ( n19886 , RI1754c610_2);
and ( n19887 , n19886 , n50928 );
and ( n19888 , C0 , RI1754c610_2);
or ( n50929 , n19887 , n19888 );
buf ( n50930 , n50929 );
not ( n50931 , n31381 );
and ( n50932 , n50931 , n48883 );
xor ( n50933 , n31318 , n50932 );
not ( n19889 , n29614 );
and ( n19890 , n19889 , RI174b3ad8_860);
and ( n19891 , n50933 , n29614 );
or ( n50934 , n19890 , n19891 );
not ( n19892 , RI1754c610_2);
and ( n19893 , n19892 , n50934 );
and ( n19894 , C0 , RI1754c610_2);
or ( n50935 , n19893 , n19894 );
buf ( n50936 , n50935 );
not ( n50937 , RI17539e48_588);
and ( n50938 , RI1753aa78_586 , n50937 );
or ( n50939 , n50938 , n27689 );
not ( n50940 , RI1754c610_2);
and ( n50941 , n50939 , n50940 );
buf ( n50942 , n50941 );
not ( n50943 , n45514 );
and ( n50944 , n50943 , n45516 );
xor ( n50945 , n46155 , n50944 );
not ( n19895 , n29614 );
and ( n19896 , n19895 , RI173f6460_1555);
and ( n19897 , n50945 , n29614 );
or ( n50946 , n19896 , n19897 );
not ( n19898 , RI1754c610_2);
and ( n19899 , n19898 , n50946 );
and ( n19900 , C0 , RI1754c610_2);
or ( n50947 , n19899 , n19900 );
buf ( n50948 , n50947 );
not ( n50949 , n42194 );
xor ( n50950 , n32914 , n38553 );
xor ( n50951 , n50950 , n41659 );
and ( n50952 , n50949 , n50951 );
xor ( n50953 , n42191 , n50952 );
not ( n19901 , n29614 );
and ( n19902 , n19901 , RI1747a760_1139);
and ( n19903 , n50953 , n29614 );
or ( n50954 , n19902 , n19903 );
not ( n19904 , RI1754c610_2);
and ( n19905 , n19904 , n50954 );
and ( n19906 , C0 , RI1754c610_2);
or ( n50955 , n19905 , n19906 );
buf ( n50956 , n50955 );
not ( n50957 , n49973 );
and ( n50958 , n50957 , n40112 );
xor ( n50959 , n48233 , n50958 );
not ( n19907 , n29614 );
and ( n19908 , n19907 , RI17460d38_1264);
and ( n19909 , n50959 , n29614 );
or ( n50960 , n19908 , n19909 );
not ( n19910 , RI1754c610_2);
and ( n19911 , n19910 , n50960 );
and ( n19912 , C0 , RI1754c610_2);
or ( n50961 , n19911 , n19912 );
buf ( n50962 , n50961 );
not ( n19913 , n27683 );
and ( n19914 , n19913 , RI19a991e8_2618);
and ( n19915 , RI19aa2c20_2547 , n27683 );
or ( n50963 , n19914 , n19915 );
not ( n19916 , RI1754c610_2);
and ( n19917 , n19916 , n50963 );
and ( n19918 , C0 , RI1754c610_2);
or ( n50964 , n19917 , n19918 );
buf ( n50965 , n50964 );
xor ( n50966 , n43265 , n41099 );
xor ( n50967 , n50966 , n30604 );
not ( n50968 , n47839 );
and ( n50969 , n50968 , n38678 );
xor ( n50970 , n50967 , n50969 );
not ( n19919 , n29614 );
and ( n19920 , n19919 , RI1747d898_1124);
and ( n19921 , n50970 , n29614 );
or ( n50971 , n19920 , n19921 );
not ( n19922 , RI1754c610_2);
and ( n19923 , n19922 , n50971 );
and ( n19924 , C0 , RI1754c610_2);
or ( n50972 , n19923 , n19924 );
buf ( n50973 , n50972 );
not ( n50974 , n44747 );
and ( n50975 , n50974 , n44613 );
xor ( n50976 , n48039 , n50975 );
not ( n19925 , n29614 );
and ( n19926 , n19925 , RI174844e0_1091);
and ( n19927 , n50976 , n29614 );
or ( n50977 , n19926 , n19927 );
not ( n19928 , RI1754c610_2);
and ( n19929 , n19928 , n50977 );
and ( n19930 , C0 , RI1754c610_2);
or ( n50978 , n19929 , n19930 );
buf ( n50979 , n50978 );
not ( n50980 , n43826 );
xor ( n50981 , n38561 , n28816 );
xor ( n50982 , n50981 , n29109 );
and ( n50983 , n50980 , n50982 );
xor ( n50984 , n43823 , n50983 );
not ( n19931 , n29614 );
and ( n19932 , n19931 , RI173b5ab0_1870);
and ( n19933 , n50984 , n29614 );
or ( n50985 , n19932 , n19933 );
not ( n19934 , RI1754c610_2);
and ( n19935 , n19934 , n50985 );
and ( n19936 , C0 , RI1754c610_2);
or ( n50986 , n19935 , n19936 );
buf ( n50987 , n50986 );
not ( n19937 , n27683 );
and ( n19938 , n19937 , RI19a8cb28_2706);
and ( n19939 , RI19a96e48_2634 , n27683 );
or ( n50988 , n19938 , n19939 );
not ( n19940 , RI1754c610_2);
and ( n19941 , n19940 , n50988 );
and ( n19942 , C0 , RI1754c610_2);
or ( n50989 , n19941 , n19942 );
buf ( n50990 , n50989 );
and ( n50991 , RI1754bbc0_24 , n34844 );
and ( n50992 , RI1754bbc0_24 , n34847 );
and ( n50993 , RI1754bbc0_24 , n34850 );
and ( n50994 , RI1754bbc0_24 , n34852 );
and ( n50995 , RI1754bbc0_24 , n34854 );
or ( n50996 , n50991 , n50992 , n50993 , n50994 , n50995 , C0 , C0 , C0 );
not ( n19943 , n34859 );
and ( n19944 , n19943 , n50996 );
and ( n19945 , RI1754bbc0_24 , n34859 );
or ( n50997 , n19944 , n19945 );
not ( n19946 , RI19a22f70_2797);
and ( n19947 , n19946 , n50997 );
and ( n19948 , C0 , RI19a22f70_2797);
or ( n50998 , n19947 , n19948 );
not ( n19949 , n27683 );
and ( n19950 , n19949 , RI19a9fcc8_2570);
and ( n19951 , n50998 , n27683 );
or ( n50999 , n19950 , n19951 );
not ( n19952 , RI1754c610_2);
and ( n19953 , n19952 , n50999 );
and ( n19954 , C0 , RI1754c610_2);
or ( n51000 , n19953 , n19954 );
buf ( n51001 , n51000 );
not ( n51002 , n43814 );
and ( n51003 , n51002 , n49819 );
xor ( n51004 , n43811 , n51003 );
not ( n19955 , n29614 );
and ( n19956 , n19955 , RI17332458_2196);
and ( n19957 , n51004 , n29614 );
or ( n51005 , n19956 , n19957 );
not ( n19958 , RI1754c610_2);
and ( n19959 , n19958 , n51005 );
and ( n19960 , C0 , RI1754c610_2);
or ( n51006 , n19959 , n19960 );
buf ( n51007 , n51006 );
not ( n51008 , n46951 );
and ( n51009 , n51008 , n45319 );
xor ( n51010 , n46550 , n51009 );
not ( n19961 , n29614 );
and ( n19962 , n19961 , RI17342448_2118);
and ( n19963 , n51010 , n29614 );
or ( n51011 , n19962 , n19963 );
not ( n19964 , RI1754c610_2);
and ( n19965 , n19964 , n51011 );
and ( n19966 , C0 , RI1754c610_2);
or ( n51012 , n19965 , n19966 );
buf ( n51013 , n51012 );
not ( n19967 , n27683 );
and ( n19968 , n19967 , RI19a846f8_2763);
and ( n19969 , RI19abf690_2337 , n27683 );
or ( n51014 , n19968 , n19969 );
not ( n19970 , RI1754c610_2);
and ( n19971 , n19970 , n51014 );
and ( n19972 , C0 , RI1754c610_2);
or ( n51015 , n19971 , n19972 );
buf ( n51016 , n51015 );
xor ( n51017 , n41040 , n34395 );
xor ( n51018 , n51017 , n34445 );
not ( n51019 , n41959 );
and ( n51020 , n51019 , n41961 );
xor ( n51021 , n51018 , n51020 );
not ( n19973 , n29614 );
and ( n19974 , n19973 , RI1747cb78_1128);
and ( n19975 , n51021 , n29614 );
or ( n51022 , n19974 , n19975 );
not ( n19976 , RI1754c610_2);
and ( n19977 , n19976 , n51022 );
and ( n19978 , C0 , RI1754c610_2);
or ( n51023 , n19977 , n19978 );
buf ( n51024 , n51023 );
not ( n51025 , n41296 );
and ( n51026 , n51025 , n41317 );
xor ( n51027 , n48977 , n51026 );
not ( n19979 , n29614 );
and ( n19980 , n19979 , RI1751e440_672);
and ( n19981 , n51027 , n29614 );
or ( n51028 , n19980 , n19981 );
not ( n19982 , RI1754c610_2);
and ( n19983 , n19982 , n51028 );
and ( n19984 , C0 , RI1754c610_2);
or ( n51029 , n19983 , n19984 );
buf ( n51030 , n51029 );
not ( n51031 , n41837 );
and ( n51032 , n51031 , n41855 );
xor ( n51033 , n47515 , n51032 );
not ( n19985 , n29614 );
and ( n19986 , n19985 , RI17467980_1231);
and ( n19987 , n51033 , n29614 );
or ( n51034 , n19986 , n19987 );
not ( n19988 , RI1754c610_2);
and ( n19989 , n19988 , n51034 );
and ( n19990 , C0 , RI1754c610_2);
or ( n51035 , n19989 , n19990 );
buf ( n51036 , n51035 );
not ( n51037 , n43421 );
and ( n51038 , n51037 , n43423 );
xor ( n51039 , n46365 , n51038 );
not ( n19991 , n29614 );
and ( n19992 , n19991 , RI17518248_691);
and ( n19993 , n51039 , n29614 );
or ( n51040 , n19992 , n19993 );
not ( n19994 , RI1754c610_2);
and ( n19995 , n19994 , n51040 );
and ( n19996 , C0 , RI1754c610_2);
or ( n51041 , n19995 , n19996 );
buf ( n51042 , n51041 );
not ( n51043 , n46391 );
and ( n51044 , n51043 , n46393 );
xor ( n51045 , n47128 , n51044 );
not ( n19997 , n29614 );
and ( n19998 , n19997 , RI174d0cc8_761);
and ( n19999 , n51045 , n29614 );
or ( n51046 , n19998 , n19999 );
not ( n20000 , RI1754c610_2);
and ( n20001 , n20000 , n51046 );
and ( n20002 , C0 , RI1754c610_2);
or ( n51047 , n20001 , n20002 );
buf ( n51048 , n51047 );
xor ( n51049 , n42595 , n38284 );
xor ( n51050 , n51049 , n39856 );
xor ( n51051 , n31010 , n41622 );
xor ( n51052 , n51051 , n38512 );
not ( n51053 , n51052 );
and ( n51054 , n51053 , n41947 );
xor ( n51055 , n51050 , n51054 );
not ( n20003 , n29614 );
and ( n20004 , n20003 , RI1738e4b0_2062);
and ( n20005 , n51055 , n29614 );
or ( n51056 , n20004 , n20005 );
not ( n20006 , RI1754c610_2);
and ( n20007 , n20006 , n51056 );
and ( n20008 , C0 , RI1754c610_2);
or ( n51057 , n20007 , n20008 );
buf ( n51058 , n51057 );
not ( n20009 , RI1754c610_2);
and ( n20010 , n20009 , RI19ad0e08_2205);
and ( n20011 , C0 , RI1754c610_2);
or ( n51059 , n20010 , n20011 );
buf ( n51060 , n51059 );
xor ( n51061 , n42334 , n29981 );
xor ( n51062 , n51061 , n35955 );
not ( n51063 , n51062 );
and ( n51064 , n51063 , n47318 );
xor ( n51065 , n46040 , n51064 );
not ( n20012 , n29614 );
and ( n20013 , n20012 , RI17339730_2161);
and ( n20014 , n51065 , n29614 );
or ( n51066 , n20013 , n20014 );
not ( n20015 , RI1754c610_2);
and ( n20016 , n20015 , n51066 );
and ( n20017 , C0 , RI1754c610_2);
or ( n51067 , n20016 , n20017 );
buf ( n51068 , n51067 );
not ( n51069 , n47024 );
and ( n51070 , n51069 , n47906 );
xor ( n51071 , n47021 , n51070 );
not ( n20018 , n29614 );
and ( n20019 , n20018 , RI17410860_1427);
and ( n20020 , n51071 , n29614 );
or ( n51072 , n20019 , n20020 );
not ( n20021 , RI1754c610_2);
and ( n20022 , n20021 , n51072 );
and ( n20023 , C0 , RI1754c610_2);
or ( n51073 , n20022 , n20023 );
buf ( n51074 , n51073 );
xor ( n51075 , n40050 , n38574 );
xor ( n51076 , n51075 , n38594 );
xor ( n51077 , n39775 , n33175 );
xor ( n51078 , n51077 , n34797 );
not ( n51079 , n51078 );
and ( n51080 , n51079 , n45716 );
xor ( n51081 , n51076 , n51080 );
not ( n20024 , n29614 );
and ( n20025 , n20024 , RI1752e610_622);
and ( n20026 , n51081 , n29614 );
or ( n51082 , n20025 , n20026 );
not ( n20027 , RI1754c610_2);
and ( n20028 , n20027 , n51082 );
and ( n20029 , C0 , RI1754c610_2);
or ( n51083 , n20028 , n20029 );
buf ( n51084 , n51083 );
xor ( n51085 , n33844 , n41146 );
xor ( n51086 , n51085 , n37291 );
not ( n51087 , n47634 );
and ( n51088 , n51087 , n47636 );
xor ( n51089 , n51086 , n51088 );
not ( n20030 , n29614 );
and ( n20031 , n20030 , RI174ab108_902);
and ( n20032 , n51089 , n29614 );
or ( n51090 , n20031 , n20032 );
not ( n20033 , RI1754c610_2);
and ( n20034 , n20033 , n51090 );
and ( n20035 , C0 , RI1754c610_2);
or ( n51091 , n20034 , n20035 );
buf ( n51092 , n51091 );
not ( n51093 , n43839 );
and ( n51094 , n51093 , n41267 );
xor ( n51095 , n50251 , n51094 );
not ( n20036 , n29614 );
and ( n20037 , n20036 , RI173eb678_1608);
and ( n20038 , n51095 , n29614 );
or ( n51096 , n20037 , n20038 );
not ( n20039 , RI1754c610_2);
and ( n20040 , n20039 , n51096 );
and ( n20041 , C0 , RI1754c610_2);
or ( n51097 , n20040 , n20041 );
buf ( n51098 , n51097 );
not ( n51099 , n44303 );
and ( n51100 , n51099 , n44305 );
xor ( n51101 , n47400 , n51100 );
not ( n20042 , n29614 );
and ( n20043 , n20042 , RI173eddd8_1596);
and ( n20044 , n51101 , n29614 );
or ( n51102 , n20043 , n20044 );
not ( n20045 , RI1754c610_2);
and ( n20046 , n20045 , n51102 );
and ( n20047 , C0 , RI1754c610_2);
or ( n51103 , n20046 , n20047 );
buf ( n51104 , n51103 );
not ( n51105 , n43683 );
and ( n51106 , n51105 , n42735 );
xor ( n51107 , n43680 , n51106 );
not ( n20048 , n29614 );
and ( n20049 , n20048 , RI1745b158_1292);
and ( n20050 , n51107 , n29614 );
or ( n51108 , n20049 , n20050 );
not ( n20051 , RI1754c610_2);
and ( n20052 , n20051 , n51108 );
and ( n20053 , C0 , RI1754c610_2);
or ( n51109 , n20052 , n20053 );
buf ( n51110 , n51109 );
not ( n51111 , n43212 );
xor ( n51112 , n37290 , n34127 );
xor ( n51113 , n51112 , n40190 );
and ( n51114 , n51111 , n51113 );
xor ( n51115 , n43209 , n51114 );
not ( n20054 , n29614 );
and ( n20055 , n20054 , RI17482aa0_1099);
and ( n20056 , n51115 , n29614 );
or ( n51116 , n20055 , n20056 );
not ( n20057 , RI1754c610_2);
and ( n20058 , n20057 , n51116 );
and ( n20059 , C0 , RI1754c610_2);
or ( n51117 , n20058 , n20059 );
buf ( n51118 , n51117 );
buf ( n51119 , RI17478690_1149);
xor ( n51120 , n40340 , n37987 );
xor ( n51121 , n51120 , n38037 );
xor ( n51122 , n42538 , n37421 );
xor ( n51123 , n51122 , n42605 );
not ( n51124 , n51123 );
and ( n51125 , n51124 , n46778 );
xor ( n51126 , n51121 , n51125 );
not ( n20060 , n29614 );
and ( n20061 , n20060 , RI173bacb8_1845);
and ( n20062 , n51126 , n29614 );
or ( n51127 , n20061 , n20062 );
not ( n20063 , RI1754c610_2);
and ( n20064 , n20063 , n51127 );
and ( n20065 , C0 , RI1754c610_2);
or ( n51128 , n20064 , n20065 );
buf ( n51129 , n51128 );
not ( n51130 , n47173 );
and ( n51131 , n51130 , n50443 );
xor ( n51132 , n47170 , n51131 );
not ( n20066 , n29614 );
and ( n20067 , n20066 , RI174ae588_886);
and ( n20068 , n51132 , n29614 );
or ( n51133 , n20067 , n20068 );
not ( n20069 , RI1754c610_2);
and ( n20070 , n20069 , n51133 );
and ( n20071 , C0 , RI1754c610_2);
or ( n51134 , n20070 , n20071 );
buf ( n51135 , n51134 );
not ( n51136 , n49966 );
and ( n51137 , n51136 , n50005 );
xor ( n51138 , n49963 , n51137 );
not ( n20072 , n29614 );
and ( n20073 , n20072 , RI1740c030_1449);
and ( n20074 , n51138 , n29614 );
or ( n51139 , n20073 , n20074 );
not ( n20075 , RI1754c610_2);
and ( n20076 , n20075 , n51139 );
and ( n20077 , C0 , RI1754c610_2);
or ( n51140 , n20076 , n20077 );
buf ( n51141 , n51140 );
xor ( n51142 , n42634 , n35052 );
xor ( n51143 , n51142 , n35069 );
not ( n51144 , n48254 );
and ( n51145 , n51144 , n43195 );
xor ( n51146 , n51143 , n51145 );
not ( n20078 , n29614 );
and ( n20079 , n20078 , RI173c22d8_1809);
and ( n20080 , n51146 , n29614 );
or ( n51147 , n20079 , n20080 );
not ( n20081 , RI1754c610_2);
and ( n20082 , n20081 , n51147 );
and ( n20083 , C0 , RI1754c610_2);
or ( n51148 , n20082 , n20083 );
buf ( n51149 , n51148 );
buf ( n51150 , RI174aa3e8_906);
xor ( n51151 , n31342 , n37074 );
xor ( n51152 , n51151 , n37104 );
not ( n51153 , n51152 );
and ( n51154 , n51153 , n49853 );
xor ( n51155 , n48937 , n51154 );
not ( n20084 , n29614 );
and ( n20085 , n20084 , RI173caff0_1766);
and ( n20086 , n51155 , n29614 );
or ( n51156 , n20085 , n20086 );
not ( n20087 , RI1754c610_2);
and ( n20088 , n20087 , n51156 );
and ( n20089 , C0 , RI1754c610_2);
or ( n51157 , n20088 , n20089 );
buf ( n51158 , n51157 );
not ( n51159 , n49604 );
and ( n51160 , n51159 , n44159 );
xor ( n51161 , n49210 , n51160 );
not ( n20090 , n29614 );
and ( n20091 , n20090 , RI17389938_2085);
and ( n20092 , n51161 , n29614 );
or ( n51162 , n20091 , n20092 );
not ( n20093 , RI1754c610_2);
and ( n20094 , n20093 , n51162 );
and ( n20095 , C0 , RI1754c610_2);
or ( n51163 , n20094 , n20095 );
buf ( n51164 , n51163 );
not ( n51165 , n44368 );
and ( n51166 , n51165 , n42017 );
xor ( n51167 , n45643 , n51166 );
not ( n20096 , n29614 );
and ( n20097 , n20096 , RI173dd758_1676);
and ( n20098 , n51167 , n29614 );
or ( n51168 , n20097 , n20098 );
not ( n20099 , RI1754c610_2);
and ( n20100 , n20099 , n51168 );
and ( n20101 , C0 , RI1754c610_2);
or ( n51169 , n20100 , n20101 );
buf ( n51170 , n51169 );
not ( n51171 , n33826 );
and ( n51172 , n51171 , n33936 );
xor ( n51173 , n39656 , n51172 );
not ( n20102 , n29614 );
and ( n20103 , n20102 , RI17449a70_1377);
and ( n20104 , n51173 , n29614 );
or ( n51174 , n20103 , n20104 );
not ( n20105 , RI1754c610_2);
and ( n20106 , n20105 , n51174 );
and ( n20107 , C0 , RI1754c610_2);
or ( n51175 , n20106 , n20107 );
buf ( n51176 , n51175 );
buf ( n51177 , RI174a9038_912);
buf ( n51178 , RI17472420_1179);
buf ( n51179 , RI19a23e70_2789);
not ( n51180 , n41372 );
and ( n51181 , n51180 , n41374 );
xor ( n51182 , n43373 , n51181 );
not ( n20108 , n29614 );
and ( n20109 , n20108 , RI174637e0_1251);
and ( n20110 , n51182 , n29614 );
or ( n51183 , n20109 , n20110 );
not ( n20111 , RI1754c610_2);
and ( n20112 , n20111 , n51183 );
and ( n20113 , C0 , RI1754c610_2);
or ( n51184 , n20112 , n20113 );
buf ( n51185 , n51184 );
not ( n51186 , n46135 );
and ( n51187 , n51186 , n46137 );
xor ( n51188 , n50533 , n51187 );
not ( n20114 , n29614 );
and ( n20115 , n20114 , RI17335f68_2178);
and ( n20116 , n51188 , n29614 );
or ( n51189 , n20115 , n20116 );
not ( n20117 , RI1754c610_2);
and ( n20118 , n20117 , n51189 );
and ( n20119 , C0 , RI1754c610_2);
or ( n51190 , n20118 , n20119 );
buf ( n51191 , n51190 );
not ( n51192 , n45962 );
and ( n51193 , n51192 , n36743 );
xor ( n51194 , n49409 , n51193 );
not ( n20120 , n29614 );
and ( n20121 , n20120 , RI173ac708_1915);
and ( n20122 , n51194 , n29614 );
or ( n51195 , n20121 , n20122 );
not ( n20123 , RI1754c610_2);
and ( n20124 , n20123 , n51195 );
and ( n20125 , C0 , RI1754c610_2);
or ( n51196 , n20124 , n20125 );
buf ( n51197 , n51196 );
xor ( n51198 , n31814 , n34644 );
xor ( n51199 , n51198 , n36401 );
not ( n51200 , n48209 );
and ( n51201 , n51200 , n48024 );
xor ( n51202 , n51199 , n51201 );
not ( n20126 , n29614 );
and ( n20127 , n20126 , RI173b1910_1890);
and ( n20128 , n51202 , n29614 );
or ( n51203 , n20127 , n20128 );
not ( n20129 , RI1754c610_2);
and ( n20130 , n20129 , n51203 );
and ( n20131 , C0 , RI1754c610_2);
or ( n51204 , n20130 , n20131 );
buf ( n51205 , n51204 );
not ( n51206 , n42574 );
and ( n51207 , n51206 , n42576 );
xor ( n51208 , n42888 , n51207 );
not ( n20132 , n29614 );
and ( n20133 , n20132 , RI17406798_1476);
and ( n20134 , n51208 , n29614 );
or ( n51209 , n20133 , n20134 );
not ( n20135 , RI1754c610_2);
and ( n20136 , n20135 , n51209 );
and ( n20137 , C0 , RI1754c610_2);
or ( n51210 , n20136 , n20137 );
buf ( n51211 , n51210 );
not ( n20138 , n27683 );
and ( n20139 , n20138 , RI19aabb90_2484);
and ( n20140 , RI19ab5820_2412 , n27683 );
or ( n51212 , n20139 , n20140 );
not ( n20141 , RI1754c610_2);
and ( n20142 , n20141 , n51212 );
and ( n20143 , C0 , RI1754c610_2);
or ( n51213 , n20142 , n20143 );
buf ( n51214 , n51213 );
buf ( n51215 , RI17462ac0_1255);
buf ( n51216 , RI17466fa8_1234);
not ( n51217 , n48390 );
and ( n51218 , n51217 , n42266 );
xor ( n51219 , n43507 , n51218 );
not ( n20144 , n29614 );
and ( n20145 , n20144 , RI17334528_2186);
and ( n20146 , n51219 , n29614 );
or ( n51220 , n20145 , n20146 );
not ( n20147 , RI1754c610_2);
and ( n20148 , n20147 , n51220 );
and ( n20149 , C0 , RI1754c610_2);
or ( n51221 , n20148 , n20149 );
buf ( n51222 , n51221 );
not ( n51223 , n46311 );
and ( n51224 , n51223 , n45070 );
xor ( n51225 , n48718 , n51224 );
not ( n20150 , n29614 );
and ( n20151 , n20150 , RI1747a0d0_1141);
and ( n20152 , n51225 , n29614 );
or ( n51226 , n20151 , n20152 );
not ( n20153 , RI1754c610_2);
and ( n20154 , n20153 , n51226 );
and ( n20155 , C0 , RI1754c610_2);
or ( n51227 , n20154 , n20155 );
buf ( n51228 , n51227 );
xor ( n51229 , n40930 , n38793 );
xor ( n51230 , n51229 , n40563 );
not ( n51231 , n51230 );
and ( n51232 , n51231 , n49145 );
xor ( n51233 , n49473 , n51232 );
not ( n20156 , n29614 );
and ( n20157 , n20156 , RI17533db8_605);
and ( n20158 , n51233 , n29614 );
or ( n51234 , n20157 , n20158 );
not ( n20159 , RI1754c610_2);
and ( n20160 , n20159 , n51234 );
and ( n20161 , C0 , RI1754c610_2);
or ( n51235 , n20160 , n20161 );
buf ( n51236 , n51235 );
xor ( n51237 , n32842 , n37203 );
xor ( n51238 , n51237 , n34150 );
not ( n51239 , n51238 );
and ( n51240 , n51239 , n48911 );
xor ( n51241 , n49037 , n51240 );
not ( n20162 , n29614 );
and ( n20163 , n20162 , RI173dca38_1680);
and ( n20164 , n51241 , n29614 );
or ( n51242 , n20163 , n20164 );
not ( n20165 , RI1754c610_2);
and ( n20166 , n20165 , n51242 );
and ( n20167 , C0 , RI1754c610_2);
or ( n51243 , n20166 , n20167 );
buf ( n51244 , n51243 );
xor ( n51245 , n35409 , n41068 );
xor ( n51246 , n51245 , n39091 );
not ( n51247 , n50822 );
and ( n51248 , n51247 , n41602 );
xor ( n51249 , n51246 , n51248 );
not ( n20168 , n29614 );
and ( n20169 , n20168 , RI1749a740_983);
and ( n20170 , n51249 , n29614 );
or ( n51250 , n20169 , n20170 );
not ( n20171 , RI1754c610_2);
and ( n20172 , n20171 , n51250 );
and ( n20173 , C0 , RI1754c610_2);
or ( n51251 , n20172 , n20173 );
buf ( n51252 , n51251 );
not ( n20174 , n27683 );
and ( n20175 , n20174 , RI19aa4cf0_2531);
and ( n20176 , RI19aaf088_2461 , n27683 );
or ( n51253 , n20175 , n20176 );
not ( n20177 , RI1754c610_2);
and ( n20178 , n20177 , n51253 );
and ( n20179 , C0 , RI1754c610_2);
or ( n51254 , n20178 , n20179 );
buf ( n51255 , n51254 );
not ( n51256 , n47646 );
and ( n51257 , n51256 , n47648 );
xor ( n51258 , n46921 , n51257 );
not ( n20180 , n29614 );
and ( n20181 , n20180 , RI17450a00_1343);
and ( n20182 , n51258 , n29614 );
or ( n51259 , n20181 , n20182 );
not ( n20183 , RI1754c610_2);
and ( n20184 , n20183 , n51259 );
and ( n20185 , C0 , RI1754c610_2);
or ( n51260 , n20184 , n20185 );
buf ( n51261 , n51260 );
buf ( n51262 , RI1748b470_1057);
buf ( n51263 , RI174d07a0_762);
not ( n51264 , n48892 );
and ( n51265 , n51264 , n48894 );
xor ( n51266 , n46116 , n51265 );
not ( n20186 , n29614 );
and ( n20187 , n20186 , RI173b88a0_1856);
and ( n20188 , n51266 , n29614 );
or ( n51267 , n20187 , n20188 );
not ( n20189 , RI1754c610_2);
and ( n20190 , n20189 , n51267 );
and ( n20191 , C0 , RI1754c610_2);
or ( n51268 , n20190 , n20191 );
buf ( n51269 , n51268 );
xor ( n51270 , n37914 , n32048 );
xor ( n51271 , n51270 , n32108 );
not ( n51272 , n51271 );
and ( n51273 , n51272 , n45942 );
xor ( n51274 , n47012 , n51273 );
not ( n20192 , n29614 );
and ( n20193 , n20192 , RI174965a0_1003);
and ( n20194 , n51274 , n29614 );
or ( n51275 , n20193 , n20194 );
not ( n20195 , RI1754c610_2);
and ( n20196 , n20195 , n51275 );
and ( n20197 , C0 , RI1754c610_2);
or ( n51276 , n20196 , n20197 );
buf ( n51277 , n51276 );
not ( n20198 , n27683 );
and ( n20199 , n20198 , RI19a8db18_2699);
and ( n20200 , RI19a97b68_2628 , n27683 );
or ( n51278 , n20199 , n20200 );
not ( n20201 , RI1754c610_2);
and ( n20202 , n20201 , n51278 );
and ( n20203 , C0 , RI1754c610_2);
or ( n51279 , n20202 , n20203 );
buf ( n51280 , n51279 );
xor ( n51281 , n34986 , n42945 );
xor ( n51282 , n51281 , n34497 );
xor ( n51283 , n40554 , n40966 );
xor ( n51284 , n51283 , n37460 );
not ( n51285 , n51284 );
and ( n51286 , n51285 , n44171 );
xor ( n51287 , n51282 , n51286 );
not ( n20204 , n29614 );
and ( n20205 , n20204 , RI1744cba8_1362);
and ( n20206 , n51287 , n29614 );
or ( n51288 , n20205 , n20206 );
not ( n20207 , RI1754c610_2);
and ( n20208 , n20207 , n51288 );
and ( n20209 , C0 , RI1754c610_2);
or ( n51289 , n20208 , n20209 );
buf ( n51290 , n51289 );
not ( n51291 , n47829 );
xor ( n51292 , n38660 , n39347 );
xor ( n51293 , n51292 , n42344 );
and ( n51294 , n51291 , n51293 );
xor ( n51295 , n47826 , n51294 );
not ( n20210 , n29614 );
and ( n20211 , n20210 , RI17519c10_686);
and ( n20212 , n51295 , n29614 );
or ( n51296 , n20211 , n20212 );
not ( n20213 , RI1754c610_2);
and ( n20214 , n20213 , n51296 );
and ( n20215 , C0 , RI1754c610_2);
or ( n51297 , n20214 , n20215 );
buf ( n51298 , n51297 );
not ( n20216 , n27683 );
and ( n20217 , n20216 , RI19a96740_2637);
and ( n20218 , RI19aa05b0_2566 , n27683 );
or ( n51299 , n20217 , n20218 );
not ( n20219 , RI1754c610_2);
and ( n20220 , n20219 , n51299 );
and ( n20221 , C0 , RI1754c610_2);
or ( n51300 , n20220 , n20221 );
buf ( n51301 , n51300 );
not ( n20222 , n27683 );
and ( n20223 , n20222 , RI19a90f20_2676);
and ( n20224 , RI19a9af70_2605 , n27683 );
or ( n51302 , n20223 , n20224 );
not ( n20225 , RI1754c610_2);
and ( n20226 , n20225 , n51302 );
and ( n20227 , C0 , RI1754c610_2);
or ( n51303 , n20226 , n20227 );
buf ( n51304 , n51303 );
not ( n51305 , n50005 );
and ( n51306 , n51305 , n50007 );
xor ( n51307 , n49966 , n51306 );
not ( n20228 , n29614 );
and ( n20229 , n20228 , RI173d1c50_1733);
and ( n20230 , n51307 , n29614 );
or ( n51308 , n20229 , n20230 );
not ( n20231 , RI1754c610_2);
and ( n20232 , n20231 , n51308 );
and ( n20233 , C0 , RI1754c610_2);
or ( n51309 , n20232 , n20233 );
buf ( n51310 , n51309 );
xor ( n51311 , n36669 , n39635 );
xor ( n51312 , n51311 , n39655 );
not ( n51313 , n51312 );
and ( n51314 , n51313 , n49292 );
xor ( n51315 , n49505 , n51314 );
not ( n20234 , n29614 );
and ( n20235 , n20234 , RI17346c78_2096);
and ( n20236 , n51315 , n29614 );
or ( n51316 , n20235 , n20236 );
not ( n20237 , RI1754c610_2);
and ( n20238 , n20237 , n51316 );
and ( n20239 , C0 , RI1754c610_2);
or ( n51317 , n20238 , n20239 );
buf ( n51318 , n51317 );
not ( n20240 , n27683 );
and ( n20241 , n20240 , RI19a82d30_2774);
and ( n20242 , RI19ab0c30_2448 , n27683 );
or ( n51319 , n20241 , n20242 );
not ( n20243 , RI1754c610_2);
and ( n20244 , n20243 , n51319 );
and ( n20245 , C0 , RI1754c610_2);
or ( n51320 , n20244 , n20245 );
buf ( n51321 , n51320 );
buf ( n51322 , n34844 );
buf ( n51323 , n51322 );
not ( n20246 , n34859 );
and ( n20247 , n20246 , n51323 );
and ( n20248 , RI1754a810_66 , n34859 );
or ( n51324 , n20247 , n20248 );
not ( n20249 , RI19a22f70_2797);
and ( n20250 , n20249 , n51324 );
and ( n20251 , C0 , RI19a22f70_2797);
or ( n51325 , n20250 , n20251 );
not ( n20252 , n27683 );
and ( n20253 , n20252 , RI19ad0238_2210);
and ( n20254 , n51325 , n27683 );
or ( n51326 , n20253 , n20254 );
not ( n20255 , RI1754c610_2);
and ( n20256 , n20255 , n51326 );
and ( n20257 , C0 , RI1754c610_2);
or ( n51327 , n20256 , n20257 );
buf ( n51328 , n51327 );
not ( n51329 , n50425 );
and ( n51330 , n51329 , n50427 );
xor ( n51331 , n50466 , n51330 );
not ( n20258 , n29614 );
and ( n20259 , n20258 , RI1746fcc0_1191);
and ( n20260 , n51331 , n29614 );
or ( n51332 , n20259 , n20260 );
not ( n20261 , RI1754c610_2);
and ( n20262 , n20261 , n51332 );
and ( n20263 , C0 , RI1754c610_2);
or ( n51333 , n20262 , n20263 );
buf ( n51334 , n51333 );
buf ( n51335 , RI174ac4b8_896);
buf ( n51336 , RI174a6f68_922);
not ( n20264 , n27683 );
and ( n20265 , n20264 , RI19ab7f80_2395);
and ( n20266 , RI19ac0d88_2324 , n27683 );
or ( n51337 , n20265 , n20266 );
not ( n20267 , RI1754c610_2);
and ( n20268 , n20267 , n51337 );
and ( n20269 , C0 , RI1754c610_2);
or ( n51338 , n20268 , n20269 );
buf ( n51339 , n51338 );
buf ( n51340 , RI17463b28_1250);
not ( n51341 , n47607 );
and ( n51342 , n51341 , n48342 );
xor ( n51343 , n47604 , n51342 );
not ( n20270 , n29614 );
and ( n20271 , n20270 , RI173fb9b0_1529);
and ( n20272 , n51343 , n29614 );
or ( n51344 , n20271 , n20272 );
not ( n20273 , RI1754c610_2);
and ( n20274 , n20273 , n51344 );
and ( n20275 , C0 , RI1754c610_2);
or ( n51345 , n20274 , n20275 );
buf ( n51346 , n51345 );
not ( n51347 , n46916 );
and ( n51348 , n51347 , n46918 );
xor ( n51349 , n47648 , n51348 );
not ( n20276 , n29614 );
and ( n20277 , n20276 , RI1752b7a8_631);
and ( n20278 , n51349 , n29614 );
or ( n51350 , n20277 , n20278 );
not ( n20279 , RI1754c610_2);
and ( n20280 , n20279 , n51350 );
and ( n20281 , C0 , RI1754c610_2);
or ( n51351 , n20280 , n20281 );
buf ( n51352 , n51351 );
xor ( n51353 , n37254 , n41391 );
xor ( n51354 , n51353 , n39686 );
not ( n51355 , n51354 );
xor ( n51356 , n32155 , n35986 );
xor ( n51357 , n51356 , n36003 );
and ( n51358 , n51355 , n51357 );
xor ( n51359 , n42878 , n51358 );
not ( n20282 , n29614 );
and ( n20283 , n20282 , RI173f9598_1540);
and ( n20284 , n51359 , n29614 );
or ( n51360 , n20283 , n20284 );
not ( n20285 , RI1754c610_2);
and ( n20286 , n20285 , n51360 );
and ( n20287 , C0 , RI1754c610_2);
or ( n51361 , n20286 , n20287 );
buf ( n51362 , n51361 );
not ( n51363 , n50276 );
and ( n51364 , n51363 , n49190 );
xor ( n51365 , n46738 , n51364 );
not ( n20288 , n29614 );
and ( n20289 , n20288 , RI1745f988_1270);
and ( n20290 , n51365 , n29614 );
or ( n51366 , n20289 , n20290 );
not ( n20291 , RI1754c610_2);
and ( n20292 , n20291 , n51366 );
and ( n20293 , C0 , RI1754c610_2);
or ( n51367 , n20292 , n20293 );
buf ( n51368 , n51367 );
not ( n51369 , n45819 );
and ( n51370 , n51369 , n48013 );
xor ( n51371 , n42138 , n51370 );
not ( n20294 , n29614 );
and ( n20295 , n20294 , RI173e8888_1622);
and ( n20296 , n51371 , n29614 );
or ( n51372 , n20295 , n20296 );
not ( n20297 , RI1754c610_2);
and ( n20298 , n20297 , n51372 );
and ( n20299 , C0 , RI1754c610_2);
or ( n51373 , n20298 , n20299 );
buf ( n51374 , n51373 );
not ( n51375 , n50180 );
and ( n51376 , n51375 , n50854 );
xor ( n51377 , n43714 , n51376 );
not ( n20300 , n29614 );
and ( n20301 , n20300 , RI173a71b8_1941);
and ( n20302 , n51377 , n29614 );
or ( n51378 , n20301 , n20302 );
not ( n20303 , RI1754c610_2);
and ( n20304 , n20303 , n51378 );
and ( n20305 , C0 , RI1754c610_2);
or ( n51379 , n20304 , n20305 );
buf ( n51380 , n51379 );
not ( n51381 , n43809 );
and ( n51382 , n51381 , n43811 );
xor ( n51383 , n49821 , n51382 );
not ( n20306 , n29614 );
and ( n20307 , n20306 , RI17451720_1339);
and ( n20308 , n51383 , n29614 );
or ( n51384 , n20307 , n20308 );
not ( n20309 , RI1754c610_2);
and ( n20310 , n20309 , n51384 );
and ( n20311 , C0 , RI1754c610_2);
or ( n51385 , n20310 , n20311 );
buf ( n51386 , n51385 );
not ( n20312 , n27683 );
and ( n20313 , n20312 , RI19a97208_2632);
and ( n20314 , RI19aa0d30_2562 , n27683 );
or ( n51387 , n20313 , n20314 );
not ( n20315 , RI1754c610_2);
and ( n20316 , n20315 , n51387 );
and ( n20317 , C0 , RI1754c610_2);
or ( n51388 , n20316 , n20317 );
buf ( n51389 , n51388 );
not ( n51390 , n32109 );
and ( n51391 , n51390 , n32310 );
xor ( n51392 , n49640 , n51391 );
not ( n20318 , n29614 );
and ( n20319 , n20318 , RI173a4080_1956);
and ( n20320 , n51392 , n29614 );
or ( n51393 , n20319 , n20320 );
not ( n20321 , RI1754c610_2);
and ( n20322 , n20321 , n51393 );
and ( n20323 , C0 , RI1754c610_2);
or ( n51394 , n20322 , n20323 );
buf ( n51395 , n51394 );
buf ( n51396 , RI174b3100_863);
buf ( n51397 , RI1749ffd8_956);
buf ( n51398 , RI17494ea8_1010);
not ( n51399 , n43153 );
xor ( n51400 , n33021 , n35639 );
xor ( n51401 , n51400 , n36227 );
and ( n51402 , n51399 , n51401 );
xor ( n51403 , n43150 , n51402 );
not ( n20324 , n29614 );
and ( n20325 , n20324 , RI173943d8_2033);
and ( n20326 , n51403 , n29614 );
or ( n51404 , n20325 , n20326 );
not ( n20327 , RI1754c610_2);
and ( n20328 , n20327 , n51404 );
and ( n20329 , C0 , RI1754c610_2);
or ( n51405 , n20328 , n20329 );
buf ( n51406 , n51405 );
buf ( n51407 , RI174c1548_809);
xor ( n51408 , n40328 , n37987 );
xor ( n51409 , n51408 , n38037 );
not ( n51410 , n51409 );
and ( n51411 , n51410 , n43249 );
xor ( n51412 , n36402 , n51411 );
not ( n20330 , n29614 );
and ( n20331 , n20330 , RI174a3e30_937);
and ( n20332 , n51412 , n29614 );
or ( n51413 , n20331 , n20332 );
not ( n20333 , RI1754c610_2);
and ( n20334 , n20333 , n51413 );
and ( n20335 , C0 , RI1754c610_2);
or ( n51414 , n20334 , n20335 );
buf ( n51415 , n51414 );
not ( n20336 , n27683 );
and ( n20337 , n20336 , RI19a9de50_2585);
and ( n20338 , RI19aa7888_2513 , n27683 );
or ( n51416 , n20337 , n20338 );
not ( n20339 , RI1754c610_2);
and ( n20340 , n20339 , n51416 );
and ( n20341 , C0 , RI1754c610_2);
or ( n51417 , n20340 , n20341 );
buf ( n51418 , n51417 );
xor ( n51419 , n37799 , n43994 );
xor ( n51420 , n51419 , n31213 );
xor ( n51421 , n37722 , n41772 );
xor ( n51422 , n51421 , n32663 );
not ( n51423 , n51422 );
and ( n51424 , n51423 , n48375 );
xor ( n51425 , n51420 , n51424 );
not ( n20342 , n29614 );
and ( n20343 , n20342 , RI173cdde0_1752);
and ( n20344 , n51425 , n29614 );
or ( n51426 , n20343 , n20344 );
not ( n20345 , RI1754c610_2);
and ( n20346 , n20345 , n51426 );
and ( n20347 , C0 , RI1754c610_2);
or ( n51427 , n20346 , n20347 );
buf ( n51428 , n51427 );
not ( n20348 , n27683 );
and ( n20349 , n20348 , RI19abebc8_2343);
and ( n20350 , RI19ac7b38_2272 , n27683 );
or ( n51429 , n20349 , n20350 );
not ( n20351 , RI1754c610_2);
and ( n20352 , n20351 , n51429 );
and ( n20353 , C0 , RI1754c610_2);
or ( n51430 , n20352 , n20353 );
buf ( n51431 , n51430 );
not ( n20354 , n27683 );
and ( n20355 , n20354 , RI19a876c8_2742);
and ( n20356 , RI19ab3a20_2426 , n27683 );
or ( n51432 , n20355 , n20356 );
not ( n20357 , RI1754c610_2);
and ( n20358 , n20357 , n51432 );
and ( n20359 , C0 , RI1754c610_2);
or ( n51433 , n20358 , n20359 );
buf ( n51434 , n51433 );
not ( n51435 , n50028 );
and ( n51436 , n51435 , n50030 );
xor ( n51437 , n48737 , n51436 );
not ( n20360 , n29614 );
and ( n20361 , n20360 , RI17461a58_1260);
and ( n20362 , n51437 , n29614 );
or ( n51438 , n20361 , n20362 );
not ( n20363 , RI1754c610_2);
and ( n20364 , n20363 , n51438 );
and ( n20365 , C0 , RI1754c610_2);
or ( n51439 , n20364 , n20365 );
buf ( n51440 , n51439 );
xor ( n51441 , n35979 , n37744 );
xor ( n51442 , n51441 , n35438 );
not ( n51443 , n51442 );
xor ( n51444 , n34299 , n38886 );
xor ( n51445 , n51444 , n39604 );
and ( n51446 , n51443 , n51445 );
xor ( n51447 , n44152 , n51446 );
not ( n20366 , n29614 );
and ( n20367 , n20366 , RI17488680_1071);
and ( n20368 , n51447 , n29614 );
or ( n51448 , n20367 , n20368 );
not ( n20369 , RI1754c610_2);
and ( n20370 , n20369 , n51448 );
and ( n20371 , C0 , RI1754c610_2);
or ( n51449 , n20370 , n20371 );
buf ( n51450 , n51449 );
not ( n51451 , n47855 );
xor ( n51452 , n39138 , n28468 );
xor ( n51453 , n51452 , n36530 );
and ( n51454 , n51451 , n51453 );
xor ( n51455 , n47852 , n51454 );
not ( n20372 , n29614 );
and ( n20373 , n20372 , RI173b9908_1851);
and ( n20374 , n51455 , n29614 );
or ( n51456 , n20373 , n20374 );
not ( n20375 , RI1754c610_2);
and ( n20376 , n20375 , n51456 );
and ( n20377 , C0 , RI1754c610_2);
or ( n51457 , n20376 , n20377 );
buf ( n51458 , n51457 );
xor ( n51459 , n40189 , n33991 );
xor ( n51460 , n51459 , n34041 );
not ( n51461 , n29982 );
and ( n51462 , n51461 , n30462 );
xor ( n51463 , n51460 , n51462 );
not ( n20378 , n29614 );
and ( n20379 , n20378 , RI173ba2e0_1848);
and ( n20380 , n51463 , n29614 );
or ( n51464 , n20379 , n20380 );
not ( n20381 , RI1754c610_2);
and ( n20382 , n20381 , n51464 );
and ( n20383 , C0 , RI1754c610_2);
or ( n51465 , n20382 , n20383 );
buf ( n51466 , n51465 );
not ( n51467 , n51050 );
and ( n51468 , n51467 , n51052 );
xor ( n51469 , n41952 , n51468 );
not ( n20384 , n29614 );
and ( n20385 , n20384 , RI1733efc8_2134);
and ( n20386 , n51469 , n29614 );
or ( n51470 , n20385 , n20386 );
not ( n20387 , RI1754c610_2);
and ( n20388 , n20387 , n51470 );
and ( n20389 , C0 , RI1754c610_2);
or ( n51471 , n20388 , n20389 );
buf ( n51472 , n51471 );
not ( n20390 , n27683 );
and ( n20391 , n20390 , RI19acef78_2218);
and ( n20392 , RI19a9e6c0_2581 , n27683 );
or ( n51473 , n20391 , n20392 );
not ( n20393 , RI1754c610_2);
and ( n20394 , n20393 , n51473 );
and ( n20395 , C0 , RI1754c610_2);
or ( n51474 , n20394 , n20395 );
buf ( n51475 , n51474 );
not ( n51476 , n48828 );
and ( n51477 , n51476 , n48830 );
xor ( n51478 , n45629 , n51477 );
not ( n20396 , n29614 );
and ( n20397 , n20396 , RI174aec18_884);
and ( n20398 , n51478 , n29614 );
or ( n51479 , n20397 , n20398 );
not ( n20399 , RI1754c610_2);
and ( n20400 , n20399 , n51479 );
and ( n20401 , C0 , RI1754c610_2);
or ( n51480 , n20400 , n20401 );
buf ( n51481 , n51480 );
not ( n51482 , n48319 );
and ( n51483 , n51482 , n47824 );
xor ( n51484 , n51293 , n51483 );
not ( n20402 , n29614 );
and ( n20403 , n20402 , RI174125e8_1418);
and ( n20404 , n51484 , n29614 );
or ( n51485 , n20403 , n20404 );
not ( n20405 , RI1754c610_2);
and ( n20406 , n20405 , n51485 );
and ( n20407 , C0 , RI1754c610_2);
or ( n51486 , n20406 , n20407 );
buf ( n51487 , n51486 );
not ( n20408 , n27683 );
and ( n20409 , n20408 , RI19abdbd8_2352);
and ( n20410 , RI19ac69e0_2280 , n27683 );
or ( n51488 , n20409 , n20410 );
not ( n20411 , RI1754c610_2);
and ( n20412 , n20411 , n51488 );
and ( n20413 , C0 , RI1754c610_2);
or ( n51489 , n20412 , n20413 );
buf ( n51490 , n51489 );
not ( n51491 , n42369 );
and ( n51492 , n51491 , n42378 );
xor ( n51493 , n48398 , n51492 );
not ( n20414 , n29614 );
and ( n20415 , n20414 , RI174caff8_779);
and ( n20416 , n51493 , n29614 );
or ( n51494 , n20415 , n20416 );
not ( n20417 , RI1754c610_2);
and ( n20418 , n20417 , n51494 );
and ( n20419 , C0 , RI1754c610_2);
or ( n51495 , n20418 , n20419 );
buf ( n51496 , n51495 );
not ( n20420 , n27683 );
and ( n20421 , n20420 , RI19ab92b8_2387);
and ( n20422 , RI19ac1a30_2317 , n27683 );
or ( n51497 , n20421 , n20422 );
not ( n20423 , RI1754c610_2);
and ( n20424 , n20423 , n51497 );
and ( n20425 , C0 , RI1754c610_2);
or ( n51498 , n20424 , n20425 );
buf ( n51499 , n51498 );
and ( n51500 , RI1754b440_40 , n34844 );
and ( n51501 , RI1754b440_40 , n34847 );
and ( n51502 , RI1754b440_40 , n34850 );
or ( n51503 , n51500 , n51501 , n51502 , C0 , C0 , C0 , C0 , C0 );
not ( n20426 , n34859 );
and ( n20427 , n20426 , n51503 );
and ( n20428 , RI1754b440_40 , n34859 );
or ( n51504 , n20427 , n20428 );
not ( n20429 , RI19a22f70_2797);
and ( n20430 , n20429 , n51504 );
and ( n20431 , C0 , RI19a22f70_2797);
or ( n51505 , n20430 , n20431 );
not ( n20432 , n27683 );
and ( n20433 , n20432 , RI19ab8778_2392);
and ( n20434 , n51505 , n27683 );
or ( n51506 , n20433 , n20434 );
not ( n20435 , RI1754c610_2);
and ( n20436 , n20435 , n51506 );
and ( n20437 , C0 , RI1754c610_2);
or ( n51507 , n20436 , n20437 );
buf ( n51508 , n51507 );
xor ( n51509 , n38667 , n39347 );
xor ( n51510 , n51509 , n42344 );
not ( n51511 , n45826 );
and ( n51512 , n51511 , n45828 );
xor ( n51513 , n51510 , n51512 );
not ( n20438 , n29614 );
and ( n20439 , n20438 , RI17486f88_1078);
and ( n20440 , n51513 , n29614 );
or ( n51514 , n20439 , n20440 );
not ( n20441 , RI1754c610_2);
and ( n20442 , n20441 , n51514 );
and ( n20443 , C0 , RI1754c610_2);
or ( n51515 , n20442 , n20443 );
buf ( n51516 , n51515 );
not ( n51517 , n41171 );
and ( n51518 , n51517 , n44408 );
xor ( n51519 , n41165 , n51518 );
not ( n20444 , n29614 );
and ( n20445 , n20444 , RI173c8bd8_1777);
and ( n20446 , n51519 , n29614 );
or ( n51520 , n20445 , n20446 );
not ( n20447 , RI1754c610_2);
and ( n20448 , n20447 , n51520 );
and ( n20449 , C0 , RI1754c610_2);
or ( n51521 , n20448 , n20449 );
buf ( n51522 , n51521 );
not ( n51523 , n50057 );
and ( n51524 , n51523 , n50229 );
xor ( n51525 , n50054 , n51524 );
not ( n20450 , n29614 );
and ( n20451 , n20450 , RI17533368_607);
and ( n20452 , n51525 , n29614 );
or ( n51526 , n20451 , n20452 );
not ( n20453 , RI1754c610_2);
and ( n20454 , n20453 , n51526 );
and ( n20455 , C0 , RI1754c610_2);
or ( n51527 , n20454 , n20455 );
buf ( n51528 , n51527 );
not ( n51529 , n42960 );
and ( n51530 , n51529 , n35515 );
xor ( n51531 , n45063 , n51530 );
not ( n20456 , n29614 );
and ( n20457 , n20456 , RI173cc058_1761);
and ( n20458 , n51531 , n29614 );
or ( n51532 , n20457 , n20458 );
not ( n20459 , RI1754c610_2);
and ( n20460 , n20459 , n51532 );
and ( n20461 , C0 , RI1754c610_2);
or ( n51533 , n20460 , n20461 );
buf ( n51534 , n51533 );
not ( n51535 , n43327 );
and ( n51536 , n51535 , n37923 );
xor ( n51537 , n43324 , n51536 );
not ( n20462 , n29614 );
and ( n20463 , n20462 , RI17411f58_1420);
and ( n20464 , n51537 , n29614 );
or ( n51538 , n20463 , n20464 );
not ( n20465 , RI1754c610_2);
and ( n20466 , n20465 , n51538 );
and ( n20467 , C0 , RI1754c610_2);
or ( n51539 , n20466 , n20467 );
buf ( n51540 , n51539 );
not ( n51541 , n43969 );
and ( n51542 , n51541 , n43971 );
xor ( n51543 , n47295 , n51542 );
not ( n20468 , n29614 );
and ( n20469 , n20468 , RI17333e98_2188);
and ( n20470 , n51543 , n29614 );
or ( n51544 , n20469 , n20470 );
not ( n20471 , RI1754c610_2);
and ( n20472 , n20471 , n51544 );
and ( n20473 , C0 , RI1754c610_2);
or ( n51545 , n20472 , n20473 );
buf ( n51546 , n51545 );
not ( n51547 , n43200 );
and ( n51548 , n51547 , n51143 );
xor ( n51549 , n43197 , n51548 );
not ( n20474 , n29614 );
and ( n20475 , n20474 , RI173a5430_1950);
and ( n20476 , n51549 , n29614 );
or ( n51550 , n20475 , n20476 );
not ( n20477 , RI1754c610_2);
and ( n20478 , n20477 , n51550 );
and ( n20479 , C0 , RI1754c610_2);
or ( n51551 , n20478 , n20479 );
buf ( n51552 , n51551 );
and ( n51553 , RI1754adb0_54 , n34844 );
buf ( n51554 , n51553 );
not ( n20480 , n34859 );
and ( n20481 , n20480 , n51554 );
and ( n20482 , RI1754adb0_54 , n34859 );
or ( n51555 , n20481 , n20482 );
not ( n20483 , RI19a22f70_2797);
and ( n20484 , n20483 , n51555 );
and ( n20485 , C0 , RI19a22f70_2797);
or ( n51556 , n20484 , n20485 );
not ( n20486 , n27683 );
and ( n20487 , n20486 , RI19a23858_2792);
and ( n20488 , n51556 , n27683 );
or ( n51557 , n20487 , n20488 );
not ( n20489 , RI1754c610_2);
and ( n20490 , n20489 , n51557 );
and ( n20491 , C0 , RI1754c610_2);
or ( n51558 , n20490 , n20491 );
buf ( n51559 , n51558 );
xor ( n51560 , n36119 , n39131 );
xor ( n51561 , n51560 , n39151 );
not ( n51562 , n42480 );
and ( n51563 , n51562 , n42482 );
xor ( n51564 , n51561 , n51563 );
not ( n20492 , n29614 );
and ( n20493 , n20492 , RI173e3d10_1645);
and ( n20494 , n51564 , n29614 );
or ( n51565 , n20493 , n20494 );
not ( n20495 , RI1754c610_2);
and ( n20496 , n20495 , n51565 );
and ( n20497 , C0 , RI1754c610_2);
or ( n51566 , n20496 , n20497 );
buf ( n51567 , n51566 );
and ( n51568 , RI1754c3b8_7 , n34844 );
and ( n51569 , RI1754c3b8_7 , n34847 );
and ( n51570 , RI1754c3b8_7 , n34850 );
and ( n51571 , RI1754c3b8_7 , n34852 );
and ( n51572 , RI1754c3b8_7 , n34854 );
and ( n51573 , RI1754c3b8_7 , n34856 );
and ( n51574 , RI1754c3b8_7 , n39233 );
or ( n51575 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , C0 );
not ( n20498 , n34859 );
and ( n20499 , n20498 , n51575 );
and ( n20500 , RI1754c3b8_7 , n34859 );
or ( n51576 , n20499 , n20500 );
not ( n20501 , RI19a22f70_2797);
and ( n20502 , n20501 , n51576 );
and ( n20503 , C0 , RI19a22f70_2797);
or ( n51577 , n20502 , n20503 );
not ( n20504 , n27683 );
and ( n20505 , n20504 , RI19a88a00_2734);
and ( n20506 , n51577 , n27683 );
or ( n51578 , n20505 , n20506 );
not ( n20507 , RI1754c610_2);
and ( n20508 , n20507 , n51578 );
and ( n20509 , C0 , RI1754c610_2);
or ( n51579 , n20508 , n20509 );
buf ( n51580 , n51579 );
xor ( n51581 , n36850 , n41198 );
xor ( n51582 , n51581 , n41215 );
not ( n51583 , n51582 );
and ( n51584 , n51583 , n48799 );
xor ( n51585 , n48876 , n51584 );
not ( n20510 , n29614 );
and ( n20511 , n20510 , RI174039a8_1490);
and ( n20512 , n51585 , n29614 );
or ( n51586 , n20511 , n20512 );
not ( n20513 , RI1754c610_2);
and ( n20514 , n20513 , n51586 );
and ( n20515 , C0 , RI1754c610_2);
or ( n51587 , n20514 , n20515 );
buf ( n51588 , n51587 );
not ( n51589 , n44501 );
xor ( n51590 , n42618 , n39856 );
xor ( n51591 , n51590 , n39886 );
and ( n51592 , n51589 , n51591 );
xor ( n51593 , n42825 , n51592 );
not ( n20516 , n29614 );
and ( n20517 , n20516 , RI17480340_1111);
and ( n20518 , n51593 , n29614 );
or ( n51594 , n20517 , n20518 );
not ( n20519 , RI1754c610_2);
and ( n20520 , n20519 , n51594 );
and ( n20521 , C0 , RI1754c610_2);
or ( n51595 , n20520 , n20521 );
buf ( n51596 , n51595 );
not ( n51597 , n47318 );
and ( n51598 , n51597 , n46035 );
xor ( n51599 , n51062 , n51598 );
not ( n20522 , n29614 );
and ( n20523 , n20522 , RI174b6580_847);
and ( n20524 , n51599 , n29614 );
or ( n51600 , n20523 , n20524 );
not ( n20525 , RI1754c610_2);
and ( n20526 , n20525 , n51600 );
and ( n20527 , C0 , RI1754c610_2);
or ( n51601 , n20526 , n20527 );
buf ( n51602 , n51601 );
not ( n20528 , n27683 );
and ( n20529 , n20528 , RI19ab6900_2405);
and ( n20530 , RI19abfc30_2334 , n27683 );
or ( n51603 , n20529 , n20530 );
not ( n20531 , RI1754c610_2);
and ( n20532 , n20531 , n51603 );
and ( n20533 , C0 , RI1754c610_2);
or ( n51604 , n20532 , n20533 );
buf ( n51605 , n51604 );
not ( n51606 , n42648 );
and ( n51607 , n51606 , n50454 );
xor ( n51608 , n42645 , n51607 );
not ( n20534 , n29614 );
and ( n20535 , n20534 , RI17458368_1306);
and ( n20536 , n51608 , n29614 );
or ( n51609 , n20535 , n20536 );
not ( n20537 , RI1754c610_2);
and ( n20538 , n20537 , n51609 );
and ( n20539 , C0 , RI1754c610_2);
or ( n51610 , n20538 , n20539 );
buf ( n51611 , n51610 );
not ( n51612 , n41780 );
and ( n51613 , n51612 , n41801 );
xor ( n51614 , n42402 , n51613 );
not ( n20540 , n29614 );
and ( n20541 , n20540 , RI173c7198_1785);
and ( n20542 , n51614 , n29614 );
or ( n51615 , n20541 , n20542 );
not ( n20543 , RI1754c610_2);
and ( n20544 , n20543 , n51615 );
and ( n20545 , C0 , RI1754c610_2);
or ( n51616 , n20544 , n20545 );
buf ( n51617 , n51616 );
xor ( n51618 , n43984 , n40808 );
xor ( n51619 , n51618 , n40828 );
not ( n51620 , n51619 );
and ( n51621 , n51620 , n49749 );
xor ( n51622 , n49578 , n51621 );
not ( n20546 , n29614 );
and ( n20547 , n20546 , RI1749cb58_972);
and ( n20548 , n51622 , n29614 );
or ( n51623 , n20547 , n20548 );
not ( n20549 , RI1754c610_2);
and ( n20550 , n20549 , n51623 );
and ( n20551 , C0 , RI1754c610_2);
or ( n51624 , n20550 , n20551 );
buf ( n51625 , n51624 );
not ( n20552 , n27683 );
and ( n20553 , n20552 , RI19ac8330_2268);
and ( n20554 , RI19a831e0_2772 , n27683 );
or ( n51626 , n20553 , n20554 );
not ( n20555 , RI1754c610_2);
and ( n20556 , n20555 , n51626 );
and ( n20557 , C0 , RI1754c610_2);
or ( n51627 , n20556 , n20557 );
buf ( n51628 , n51627 );
not ( n20558 , n27683 );
and ( n20559 , n20558 , RI19a8c498_2709);
and ( n20560 , RI19a964e8_2638 , n27683 );
or ( n51629 , n20559 , n20560 );
not ( n20561 , RI1754c610_2);
and ( n20562 , n20561 , n51629 );
and ( n20563 , C0 , RI1754c610_2);
or ( n51630 , n20562 , n20563 );
buf ( n51631 , n51630 );
not ( n20564 , n27683 );
and ( n20565 , n20564 , RI19ac5bd0_2286);
and ( n20566 , RI19ace870_2221 , n27683 );
or ( n51632 , n20565 , n20566 );
not ( n20567 , RI1754c610_2);
and ( n20568 , n20567 , n51632 );
and ( n20569 , C0 , RI1754c610_2);
or ( n51633 , n20568 , n20569 );
buf ( n51634 , n51633 );
xor ( n51635 , n33586 , n41740 );
xor ( n51636 , n51635 , n38371 );
not ( n51637 , n51636 );
and ( n51638 , n51637 , n49377 );
xor ( n51639 , n46528 , n51638 );
not ( n20570 , n29614 );
and ( n20571 , n20570 , RI17445f60_1395);
and ( n20572 , n51639 , n29614 );
or ( n51640 , n20571 , n20572 );
not ( n20573 , RI1754c610_2);
and ( n20574 , n20573 , n51640 );
and ( n20575 , C0 , RI1754c610_2);
or ( n51641 , n20574 , n20575 );
buf ( n51642 , n51641 );
not ( n20576 , n27683 );
and ( n20577 , n20576 , RI19aa0790_2565);
and ( n20578 , RI19aaa330_2494 , n27683 );
or ( n51643 , n20577 , n20578 );
not ( n20579 , RI1754c610_2);
and ( n20580 , n20579 , n51643 );
and ( n20581 , C0 , RI1754c610_2);
or ( n51644 , n20580 , n20581 );
buf ( n51645 , n51644 );
buf ( n51646 , RI17492400_1023);
not ( n51647 , n46140 );
and ( n51648 , n51647 , n50530 );
xor ( n51649 , n46137 , n51648 );
not ( n20582 , n29614 );
and ( n20583 , n20582 , RI174c6cf0_792);
and ( n20584 , n51649 , n29614 );
or ( n51650 , n20583 , n20584 );
not ( n20585 , RI1754c610_2);
and ( n20586 , n20585 , n51650 );
and ( n20587 , C0 , RI1754c610_2);
or ( n51651 , n20586 , n20587 );
buf ( n51652 , n51651 );
buf ( n51653 , RI17485890_1085);
not ( n51654 , n44100 );
and ( n51655 , n51654 , n45182 );
xor ( n51656 , n44097 , n51655 );
not ( n20588 , n29614 );
and ( n20589 , n20588 , RI173f6118_1556);
and ( n20590 , n51656 , n29614 );
or ( n51657 , n20589 , n20590 );
not ( n20591 , RI1754c610_2);
and ( n20592 , n20591 , n51657 );
and ( n20593 , C0 , RI1754c610_2);
or ( n51658 , n20592 , n20593 );
buf ( n51659 , n51658 );
not ( n20594 , n27683 );
and ( n20595 , n20594 , RI19ab48a8_2419);
and ( n20596 , RI19abe100_2349 , n27683 );
or ( n51660 , n20595 , n20596 );
not ( n20597 , RI1754c610_2);
and ( n20598 , n20597 , n51660 );
and ( n20599 , C0 , RI1754c610_2);
or ( n51661 , n20598 , n20599 );
buf ( n51662 , n51661 );
buf ( n51663 , RI1750a490_734);
not ( n51664 , n46887 );
and ( n51665 , n51664 , n46889 );
xor ( n51666 , n49364 , n51665 );
not ( n20600 , n29614 );
and ( n20601 , n20600 , RI174606a8_1266);
and ( n20602 , n51666 , n29614 );
or ( n51667 , n20601 , n20602 );
not ( n20603 , RI1754c610_2);
and ( n20604 , n20603 , n51667 );
and ( n20605 , C0 , RI1754c610_2);
or ( n51668 , n20604 , n20605 );
buf ( n51669 , n51668 );
not ( n51670 , n37267 );
and ( n51671 , n51670 , n44244 );
xor ( n51672 , n37261 , n51671 );
not ( n20606 , n29614 );
and ( n20607 , n20606 , RI17402940_1495);
and ( n20608 , n51672 , n29614 );
or ( n51673 , n20607 , n20608 );
not ( n20609 , RI1754c610_2);
and ( n20610 , n20609 , n51673 );
and ( n20611 , C0 , RI1754c610_2);
or ( n51674 , n20610 , n20611 );
buf ( n51675 , n51674 );
not ( n20612 , n27683 );
and ( n20613 , n20612 , RI19aadd50_2469);
and ( n20614 , RI19ab7878_2398 , n27683 );
or ( n51676 , n20613 , n20614 );
not ( n20615 , RI1754c610_2);
and ( n20616 , n20615 , n51676 );
and ( n20617 , C0 , RI1754c610_2);
or ( n51677 , n20616 , n20617 );
buf ( n51678 , n51677 );
buf ( n51679 , RI174c5d78_795);
not ( n20618 , n27683 );
and ( n20619 , n20618 , RI19abca80_2362);
and ( n20620 , RI19ac52e8_2290 , n27683 );
or ( n51680 , n20619 , n20620 );
not ( n20621 , RI1754c610_2);
and ( n20622 , n20621 , n51680 );
and ( n20623 , C0 , RI1754c610_2);
or ( n51681 , n20622 , n20623 );
buf ( n51682 , n51681 );
xor ( n51683 , n35146 , n37915 );
xor ( n51684 , n51683 , n43492 );
not ( n51685 , n51684 );
xor ( n51686 , n34010 , n34251 );
xor ( n51687 , n51686 , n42033 );
and ( n51688 , n51685 , n51687 );
xor ( n51689 , n49427 , n51688 );
not ( n20624 , n29614 );
and ( n20625 , n20624 , RI174a8318_916);
and ( n20626 , n51689 , n29614 );
or ( n51690 , n20625 , n20626 );
not ( n20627 , RI1754c610_2);
and ( n20628 , n20627 , n51690 );
and ( n20629 , C0 , RI1754c610_2);
or ( n51691 , n20628 , n20629 );
buf ( n51692 , n51691 );
not ( n51693 , n48779 );
and ( n51694 , n51693 , n49273 );
xor ( n51695 , n44784 , n51694 );
not ( n20630 , n29614 );
and ( n20631 , n20630 , RI174ac4b8_896);
and ( n20632 , n51695 , n29614 );
or ( n51696 , n20631 , n20632 );
not ( n20633 , RI1754c610_2);
and ( n20634 , n20633 , n51696 );
and ( n20635 , C0 , RI1754c610_2);
or ( n51697 , n20634 , n20635 );
buf ( n51698 , n51697 );
buf ( n51699 , RI17482aa0_1099);
buf ( n51700 , RI17471d90_1181);
buf ( n51701 , RI1750e798_721);
not ( n20636 , n27683 );
and ( n20637 , n20636 , RI19aad828_2471);
and ( n20638 , RI19ab7530_2399 , n27683 );
or ( n51702 , n20637 , n20638 );
not ( n20639 , RI1754c610_2);
and ( n20640 , n20639 , n51702 );
and ( n20641 , C0 , RI1754c610_2);
or ( n51703 , n20640 , n20641 );
buf ( n51704 , n51703 );
not ( n20642 , n27683 );
and ( n20643 , n20642 , RI19aba050_2380);
and ( n20644 , RI19ac2a98_2309 , n27683 );
or ( n51705 , n20643 , n20644 );
not ( n20645 , RI1754c610_2);
and ( n20646 , n20645 , n51705 );
and ( n20647 , C0 , RI1754c610_2);
or ( n51706 , n20646 , n20647 );
buf ( n51707 , n51706 );
not ( n51708 , n47332 );
and ( n51709 , n51708 , n47334 );
xor ( n51710 , n47372 , n51709 );
not ( n20648 , n29614 );
and ( n20649 , n20648 , RI1738f860_2056);
and ( n20650 , n51710 , n29614 );
or ( n51711 , n20649 , n20650 );
not ( n20651 , RI1754c610_2);
and ( n20652 , n20651 , n51711 );
and ( n20653 , C0 , RI1754c610_2);
or ( n51712 , n20652 , n20653 );
buf ( n51713 , n51712 );
not ( n51714 , n47445 );
and ( n51715 , n51714 , n43292 );
xor ( n51716 , n47442 , n51715 );
not ( n20654 , n29614 );
and ( n20655 , n20654 , RI1748b470_1057);
and ( n20656 , n51716 , n29614 );
or ( n51717 , n20655 , n20656 );
not ( n20657 , RI1754c610_2);
and ( n20658 , n20657 , n51717 );
and ( n20659 , C0 , RI1754c610_2);
or ( n51718 , n20658 , n20659 );
buf ( n51719 , n51718 );
not ( n20660 , n27683 );
and ( n20661 , n20660 , RI19aa71f8_2515);
and ( n20662 , RI19ab1518_2444 , n27683 );
or ( n51720 , n20661 , n20662 );
not ( n20663 , RI1754c610_2);
and ( n20664 , n20663 , n51720 );
and ( n20665 , C0 , RI1754c610_2);
or ( n51721 , n20664 , n20665 );
buf ( n51722 , n51721 );
not ( n51723 , n44791 );
and ( n51724 , n51723 , n43447 );
xor ( n51725 , n49120 , n51724 );
not ( n20666 , n29614 );
and ( n20667 , n20666 , RI17503de8_748);
and ( n20668 , n51725 , n29614 );
or ( n51726 , n20667 , n20668 );
not ( n20669 , RI1754c610_2);
and ( n20670 , n20669 , n51726 );
and ( n20671 , C0 , RI1754c610_2);
or ( n51727 , n20670 , n20671 );
buf ( n51728 , n51727 );
not ( n51729 , n50138 );
and ( n51730 , n51729 , n49492 );
xor ( n51731 , n50135 , n51730 );
not ( n20672 , n29614 );
and ( n20673 , n20672 , RI173b9278_1853);
and ( n20674 , n51731 , n29614 );
or ( n51732 , n20673 , n20674 );
not ( n20675 , RI1754c610_2);
and ( n20676 , n20675 , n51732 );
and ( n20677 , C0 , RI1754c610_2);
or ( n51733 , n20676 , n20677 );
buf ( n51734 , n51733 );
not ( n51735 , n44922 );
and ( n51736 , n51735 , n42112 );
xor ( n51737 , n45565 , n51736 );
not ( n20678 , n29614 );
and ( n20679 , n20678 , RI173daff8_1688);
and ( n20680 , n51737 , n29614 );
or ( n51738 , n20679 , n20680 );
not ( n20681 , RI1754c610_2);
and ( n20682 , n20681 , n51738 );
and ( n20683 , C0 , RI1754c610_2);
or ( n51739 , n20682 , n20683 );
buf ( n51740 , n51739 );
not ( n51741 , n44625 );
and ( n51742 , n51741 , n44627 );
xor ( n51743 , n33779 , n51742 );
not ( n20684 , n29614 );
and ( n20685 , n20684 , RI173c8548_1779);
and ( n20686 , n51743 , n29614 );
or ( n51744 , n20685 , n20686 );
not ( n20687 , RI1754c610_2);
and ( n20688 , n20687 , n51744 );
and ( n20689 , C0 , RI1754c610_2);
or ( n51745 , n20688 , n20689 );
buf ( n51746 , n51745 );
buf ( n51747 , RI174adef8_888);
not ( n51748 , n50454 );
and ( n51749 , n51748 , n50456 );
xor ( n51750 , n42648 , n51749 );
not ( n20690 , n29614 );
and ( n20691 , n20690 , RI17499d68_986);
and ( n20692 , n51750 , n29614 );
or ( n51751 , n20691 , n20692 );
not ( n20693 , RI1754c610_2);
and ( n20694 , n20693 , n51751 );
and ( n20695 , C0 , RI1754c610_2);
or ( n51752 , n20694 , n20695 );
buf ( n51753 , n51752 );
not ( n51754 , n45643 );
and ( n51755 , n51754 , n44368 );
xor ( n51756 , n42051 , n51755 );
not ( n20696 , n29614 );
and ( n20697 , n20696 , RI173cf190_1746);
and ( n20698 , n51756 , n29614 );
or ( n51757 , n20697 , n20698 );
not ( n20699 , RI1754c610_2);
and ( n20700 , n20699 , n51757 );
and ( n20701 , C0 , RI1754c610_2);
or ( n51758 , n20700 , n20701 );
buf ( n51759 , n51758 );
not ( n20702 , n27683 );
and ( n20703 , n20702 , RI19ac21b0_2313);
and ( n20704 , RI19acb300_2246 , n27683 );
or ( n51760 , n20703 , n20704 );
not ( n20705 , RI1754c610_2);
and ( n20706 , n20705 , n51760 );
and ( n20707 , C0 , RI1754c610_2);
or ( n51761 , n20706 , n20707 );
buf ( n51762 , n51761 );
not ( n20708 , n27683 );
and ( n20709 , n20708 , RI19ac1490_2320);
and ( n20710 , RI19aca9a0_2251 , n27683 );
or ( n51763 , n20709 , n20710 );
not ( n20711 , RI1754c610_2);
and ( n20712 , n20711 , n51763 );
and ( n20713 , C0 , RI1754c610_2);
or ( n51764 , n20712 , n20713 );
buf ( n51765 , n51764 );
buf ( n51766 , RI174a4e98_932);
not ( n51767 , n40693 );
and ( n51768 , n51767 , n40700 );
xor ( n51769 , n42086 , n51768 );
not ( n20714 , n29614 );
and ( n20715 , n20714 , RI173ee120_1595);
and ( n20716 , n51769 , n29614 );
or ( n51770 , n20715 , n20716 );
not ( n20717 , RI1754c610_2);
and ( n20718 , n20717 , n51770 );
and ( n20719 , C0 , RI1754c610_2);
or ( n51771 , n20718 , n20719 );
buf ( n51772 , n51771 );
not ( n51773 , n51293 );
and ( n51774 , n51773 , n48319 );
xor ( n51775 , n47829 , n51774 );
not ( n20720 , n29614 );
and ( n20721 , n20720 , RI173f22c0_1575);
and ( n20722 , n51775 , n29614 );
or ( n51776 , n20721 , n20722 );
not ( n20723 , RI1754c610_2);
and ( n20724 , n20723 , n51776 );
and ( n20725 , C0 , RI1754c610_2);
or ( n51777 , n20724 , n20725 );
buf ( n51778 , n51777 );
not ( n20726 , n27683 );
and ( n20727 , n20726 , RI19a9a3b8_2610);
and ( n20728 , RI19aa3aa8_2540 , n27683 );
or ( n51779 , n20727 , n20728 );
not ( n20729 , RI1754c610_2);
and ( n20730 , n20729 , n51779 );
and ( n20731 , C0 , RI1754c610_2);
or ( n51780 , n20730 , n20731 );
buf ( n51781 , n51780 );
buf ( n51782 , RI17476278_1160);
not ( n51783 , n44524 );
and ( n51784 , n51783 , n44526 );
xor ( n51785 , n45690 , n51784 );
not ( n20732 , n29614 );
and ( n20733 , n20732 , RI1745a780_1295);
and ( n20734 , n51785 , n29614 );
or ( n51786 , n20733 , n20734 );
not ( n20735 , RI1754c610_2);
and ( n20736 , n20735 , n51786 );
and ( n20737 , C0 , RI1754c610_2);
or ( n51787 , n20736 , n20737 );
buf ( n51788 , n51787 );
buf ( n51789 , RI1746d560_1203);
not ( n20738 , n27683 );
and ( n20739 , n20738 , RI19a96290_2639);
and ( n20740 , RI19aa0100_2568 , n27683 );
or ( n51790 , n20739 , n20740 );
not ( n20741 , RI1754c610_2);
and ( n20742 , n20741 , n51790 );
and ( n20743 , C0 , RI1754c610_2);
or ( n51791 , n20742 , n20743 );
buf ( n51792 , n51791 );
xor ( n51793 , n35593 , n37490 );
xor ( n51794 , n51793 , n41316 );
not ( n51795 , n51794 );
and ( n51796 , n51795 , n45541 );
xor ( n51797 , n46903 , n51796 );
not ( n20744 , n29614 );
and ( n20745 , n20744 , RI173fd3f0_1521);
and ( n20746 , n51797 , n29614 );
or ( n51798 , n20745 , n20746 );
not ( n20747 , RI1754c610_2);
and ( n20748 , n20747 , n51798 );
and ( n20749 , C0 , RI1754c610_2);
or ( n51799 , n20748 , n20749 );
buf ( n51800 , n51799 );
xor ( n51801 , n40029 , n40855 );
xor ( n51802 , n51801 , n38574 );
not ( n51803 , n51802 );
xor ( n51804 , n30246 , n34755 );
xor ( n51805 , n51804 , n35311 );
and ( n51806 , n51803 , n51805 );
xor ( n51807 , n45809 , n51806 );
not ( n20750 , n29614 );
and ( n20751 , n20750 , RI1745e5d8_1276);
and ( n20752 , n51807 , n29614 );
or ( n51808 , n20751 , n20752 );
not ( n20753 , RI1754c610_2);
and ( n20754 , n20753 , n51808 );
and ( n20755 , C0 , RI1754c610_2);
or ( n51809 , n20754 , n20755 );
buf ( n51810 , n51809 );
xor ( n51811 , n41274 , n38648 );
xor ( n51812 , n51811 , n40890 );
not ( n51813 , n35912 );
and ( n51814 , n51813 , n35956 );
xor ( n51815 , n51812 , n51814 );
not ( n20756 , n29614 );
and ( n20757 , n20756 , RI173599e0_2088);
and ( n20758 , n51815 , n29614 );
or ( n51816 , n20757 , n20758 );
not ( n20759 , RI1754c610_2);
and ( n20760 , n20759 , n51816 );
and ( n20761 , C0 , RI1754c610_2);
or ( n51817 , n20760 , n20761 );
buf ( n51818 , n51817 );
not ( n51819 , n45839 );
and ( n51820 , n51819 , n48398 );
xor ( n51821 , n42381 , n51820 );
not ( n20762 , n29614 );
and ( n20763 , n20762 , RI17338a10_2165);
and ( n20764 , n51821 , n29614 );
or ( n51822 , n20763 , n20764 );
not ( n20765 , RI1754c610_2);
and ( n20766 , n20765 , n51822 );
and ( n20767 , C0 , RI1754c610_2);
or ( n51823 , n20766 , n20767 );
buf ( n51824 , n51823 );
not ( n51825 , n43094 );
and ( n51826 , n51825 , n43096 );
xor ( n51827 , n45914 , n51826 );
not ( n20768 , n29614 );
and ( n20769 , n20768 , RI173b4700_1876);
and ( n20770 , n51827 , n29614 );
or ( n51828 , n20769 , n20770 );
not ( n20771 , RI1754c610_2);
and ( n20772 , n20771 , n51828 );
and ( n20773 , C0 , RI1754c610_2);
or ( n51829 , n20772 , n20773 );
buf ( n51830 , n51829 );
not ( n51831 , n49578 );
and ( n51832 , n51831 , n51619 );
xor ( n51833 , n49575 , n51832 );
not ( n20774 , n29614 );
and ( n20775 , n20774 , RI1748df18_1044);
and ( n20776 , n51833 , n29614 );
or ( n51834 , n20775 , n20776 );
not ( n20777 , RI1754c610_2);
and ( n20778 , n20777 , n51834 );
and ( n20779 , C0 , RI1754c610_2);
or ( n51835 , n20778 , n20779 );
buf ( n51836 , n51835 );
not ( n20780 , n27683 );
and ( n20781 , n20780 , RI19aca748_2252);
and ( n20782 , RI19a85c10_2754 , n27683 );
or ( n51837 , n20781 , n20782 );
not ( n20783 , RI1754c610_2);
and ( n20784 , n20783 , n51837 );
and ( n20785 , C0 , RI1754c610_2);
or ( n51838 , n20784 , n20785 );
buf ( n51839 , n51838 );
buf ( n51840 , RI17494188_1014);
buf ( n51841 , RI1747f620_1115);
not ( n20786 , n27683 );
and ( n20787 , n20786 , RI19a9c848_2594);
and ( n20788 , RI19aa6190_2522 , n27683 );
or ( n51842 , n20787 , n20788 );
not ( n20789 , RI1754c610_2);
and ( n20790 , n20789 , n51842 );
and ( n20791 , C0 , RI1754c610_2);
or ( n51843 , n20790 , n20791 );
buf ( n51844 , n51843 );
not ( n51845 , n46593 );
and ( n51846 , n51845 , n46595 );
xor ( n51847 , n41886 , n51846 );
not ( n20792 , n29614 );
and ( n20793 , n20792 , RI17455c08_1318);
and ( n20794 , n51847 , n29614 );
or ( n51848 , n20793 , n20794 );
not ( n20795 , RI1754c610_2);
and ( n20796 , n20795 , n51848 );
and ( n20797 , C0 , RI1754c610_2);
or ( n51849 , n20796 , n20797 );
buf ( n51850 , n51849 );
buf ( n51851 , RI17514468_703);
buf ( n51852 , RI174c2f10_804);
not ( n51853 , n46870 );
and ( n51854 , n51853 , n45934 );
xor ( n51855 , n41666 , n51854 );
not ( n20798 , n29614 );
and ( n20799 , n20798 , RI173c7828_1783);
and ( n20800 , n51855 , n29614 );
or ( n51856 , n20799 , n20800 );
not ( n20801 , RI1754c610_2);
and ( n20802 , n20801 , n51856 );
and ( n20803 , C0 , RI1754c610_2);
or ( n51857 , n20802 , n20803 );
buf ( n51858 , n51857 );
not ( n51859 , n49377 );
and ( n51860 , n51859 , n46523 );
xor ( n51861 , n51636 , n51860 );
not ( n20804 , n29614 );
and ( n20805 , n20804 , RI17454510_1325);
and ( n20806 , n51861 , n29614 );
or ( n51862 , n20805 , n20806 );
not ( n20807 , RI1754c610_2);
and ( n20808 , n20807 , n51862 );
and ( n20809 , C0 , RI1754c610_2);
or ( n51863 , n20808 , n20809 );
buf ( n51864 , n51863 );
not ( n51865 , n46721 );
and ( n51866 , n51865 , n46723 );
xor ( n51867 , n48200 , n51866 );
not ( n20810 , n29614 );
and ( n20811 , n20810 , RI173a2640_1964);
and ( n20812 , n51867 , n29614 );
or ( n51868 , n20811 , n20812 );
not ( n20813 , RI1754c610_2);
and ( n20814 , n20813 , n51868 );
and ( n20815 , C0 , RI1754c610_2);
or ( n51869 , n20814 , n20815 );
buf ( n51870 , n51869 );
not ( n20816 , n27683 );
and ( n20817 , n20816 , RI19a869a8_2748);
and ( n20818 , RI19a85508_2757 , n27683 );
or ( n51871 , n20817 , n20818 );
not ( n20819 , RI1754c610_2);
and ( n20820 , n20819 , n51871 );
and ( n20821 , C0 , RI1754c610_2);
or ( n51872 , n20820 , n20821 );
buf ( n51873 , n51872 );
not ( n51874 , n44874 );
and ( n51875 , n51874 , n44876 );
xor ( n51876 , n48584 , n51875 );
not ( n20822 , n29614 );
and ( n20823 , n20822 , RI17358cc0_2092);
and ( n20824 , n51876 , n29614 );
or ( n51877 , n20823 , n20824 );
not ( n20825 , RI1754c610_2);
and ( n20826 , n20825 , n51877 );
and ( n20827 , C0 , RI1754c610_2);
or ( n51878 , n20826 , n20827 );
buf ( n51879 , n51878 );
xor ( n51880 , n37541 , n34918 );
xor ( n51881 , n51880 , n34968 );
not ( n51882 , n51881 );
xor ( n51883 , n37614 , n40319 );
xor ( n51884 , n51883 , n40149 );
and ( n51885 , n51882 , n51884 );
xor ( n51886 , n48690 , n51885 );
not ( n20828 , n29614 );
and ( n20829 , n20828 , RI1738b030_2078);
and ( n20830 , n51886 , n29614 );
or ( n51887 , n20829 , n20830 );
not ( n20831 , RI1754c610_2);
and ( n20832 , n20831 , n51887 );
and ( n20833 , C0 , RI1754c610_2);
or ( n51888 , n20832 , n20833 );
buf ( n51889 , n51888 );
not ( n51890 , n42849 );
and ( n51891 , n51890 , n45291 );
xor ( n51892 , n42846 , n51891 );
not ( n20834 , n29614 );
and ( n20835 , n20834 , RI17333808_2190);
and ( n20836 , n51892 , n29614 );
or ( n51893 , n20835 , n20836 );
not ( n20837 , RI1754c610_2);
and ( n20838 , n20837 , n51893 );
and ( n20839 , C0 , RI1754c610_2);
or ( n51894 , n20838 , n20839 );
buf ( n51895 , n51894 );
not ( n51896 , n49134 );
and ( n51897 , n51896 , n32621 );
xor ( n51898 , n42149 , n51897 );
not ( n20840 , n29614 );
and ( n20841 , n20840 , RI175279c8_643);
and ( n20842 , n51898 , n29614 );
or ( n51899 , n20841 , n20842 );
not ( n20843 , RI1754c610_2);
and ( n20844 , n20843 , n51899 );
and ( n20845 , C0 , RI1754c610_2);
or ( n51900 , n20844 , n20845 );
buf ( n51901 , n51900 );
buf ( n51902 , RI1747ec48_1118);
buf ( n51903 , RI1748bb00_1055);
buf ( n51904 , RI174cf828_765);
buf ( n51905 , RI175153e0_700);
not ( n51906 , n47959 );
and ( n51907 , n51906 , n47961 );
xor ( n51908 , n39821 , n51907 );
not ( n20846 , n29614 );
and ( n20847 , n20846 , RI173c7eb8_1781);
and ( n20848 , n51908 , n29614 );
or ( n51909 , n20847 , n20848 );
not ( n20849 , RI1754c610_2);
and ( n20850 , n20849 , n51909 );
and ( n20851 , C0 , RI1754c610_2);
or ( n51910 , n20850 , n20851 );
buf ( n51911 , n51910 );
not ( n20852 , RI1754c610_2);
and ( n20853 , n20852 , RI1753a460_587);
and ( n20854 , C0 , RI1754c610_2);
or ( n51912 , n20853 , n20854 );
buf ( n51913 , n51912 );
not ( n51914 , n49527 );
and ( n51915 , n51914 , n41724 );
xor ( n51916 , n49524 , n51915 );
not ( n20855 , n29614 );
and ( n20856 , n20855 , RI17463b28_1250);
and ( n20857 , n51916 , n29614 );
or ( n51917 , n20856 , n20857 );
not ( n20858 , RI1754c610_2);
and ( n20859 , n20858 , n51917 );
and ( n20860 , C0 , RI1754c610_2);
or ( n51918 , n20859 , n20860 );
buf ( n51919 , n51918 );
not ( n51920 , n49640 );
and ( n51921 , n51920 , n32109 );
xor ( n51922 , n49637 , n51921 );
not ( n20861 , n29614 );
and ( n20862 , n20861 , RI17395788_2027);
and ( n20863 , n51922 , n29614 );
or ( n51923 , n20862 , n20863 );
not ( n20864 , RI1754c610_2);
and ( n20865 , n20864 , n51923 );
and ( n20866 , C0 , RI1754c610_2);
or ( n51924 , n20865 , n20866 );
buf ( n51925 , n51924 );
xor ( n51926 , n39591 , n31621 );
xor ( n51927 , n51926 , n35272 );
not ( n51928 , n39720 );
and ( n51929 , n51928 , n39741 );
xor ( n51930 , n51927 , n51929 );
not ( n20867 , n29614 );
and ( n20868 , n20867 , RI173d8be0_1699);
and ( n20869 , n51930 , n29614 );
or ( n51931 , n20868 , n20869 );
not ( n20870 , RI1754c610_2);
and ( n20871 , n20870 , n51931 );
and ( n20872 , C0 , RI1754c610_2);
or ( n51932 , n20871 , n20872 );
buf ( n51933 , n51932 );
not ( n51934 , n46469 );
and ( n51935 , n51934 , n48481 );
xor ( n51936 , n43539 , n51935 );
not ( n20873 , n29614 );
and ( n20874 , n20873 , RI173de7c0_1671);
and ( n20875 , n51936 , n29614 );
or ( n51937 , n20874 , n20875 );
not ( n20876 , RI1754c610_2);
and ( n20877 , n20876 , n51937 );
and ( n20878 , C0 , RI1754c610_2);
or ( n51938 , n20877 , n20878 );
buf ( n51939 , n51938 );
not ( n51940 , n42444 );
and ( n51941 , n51940 , n42446 );
xor ( n51942 , n45475 , n51941 );
not ( n20879 , n29614 );
and ( n20880 , n20879 , RI17491050_1029);
and ( n20881 , n51942 , n29614 );
or ( n51943 , n20880 , n20881 );
not ( n20882 , RI1754c610_2);
and ( n20883 , n20882 , n51943 );
and ( n20884 , C0 , RI1754c610_2);
or ( n51944 , n20883 , n20884 );
buf ( n51945 , n51944 );
not ( n51946 , n51812 );
and ( n51947 , n51946 , n35912 );
xor ( n51948 , n44316 , n51947 );
not ( n20885 , n29614 );
and ( n20886 , n20885 , RI173c3688_1803);
and ( n20887 , n51948 , n29614 );
or ( n51949 , n20886 , n20887 );
not ( n20888 , RI1754c610_2);
and ( n20889 , n20888 , n51949 );
and ( n20890 , C0 , RI1754c610_2);
or ( n51950 , n20889 , n20890 );
buf ( n51951 , n51950 );
not ( n20891 , n27683 );
and ( n20892 , n20891 , RI19abd2f0_2357);
and ( n20893 , RI19ac5bd0_2286 , n27683 );
or ( n51952 , n20892 , n20893 );
not ( n20894 , RI1754c610_2);
and ( n20895 , n20894 , n51952 );
and ( n20896 , C0 , RI1754c610_2);
or ( n51953 , n20895 , n20896 );
buf ( n51954 , n51953 );
buf ( n51955 , RI1747cec0_1127);
not ( n51956 , n46383 );
and ( n51957 , n51956 , n45667 );
xor ( n51958 , n49630 , n51957 );
not ( n20897 , n29614 );
and ( n20898 , n20897 , RI17341db8_2120);
and ( n20899 , n51958 , n29614 );
or ( n51959 , n20898 , n20899 );
not ( n20900 , RI1754c610_2);
and ( n20901 , n20900 , n51959 );
and ( n20902 , C0 , RI1754c610_2);
or ( n51960 , n20901 , n20902 );
buf ( n51961 , n51960 );
not ( n51962 , n46778 );
and ( n51963 , n51962 , n46780 );
xor ( n51964 , n51123 , n51963 );
not ( n20903 , n29614 );
and ( n20904 , n20903 , RI17340030_2129);
and ( n20905 , n51964 , n29614 );
or ( n51965 , n20904 , n20905 );
not ( n20906 , RI1754c610_2);
and ( n20907 , n20906 , n51965 );
and ( n20908 , C0 , RI1754c610_2);
or ( n51966 , n20907 , n20908 );
buf ( n51967 , n51966 );
not ( n51968 , n36948 );
xor ( n51969 , n38984 , n41590 );
xor ( n51970 , n51969 , n35804 );
and ( n51971 , n51968 , n51970 );
xor ( n51972 , n36892 , n51971 );
not ( n20909 , n29614 );
and ( n20910 , n20909 , RI174534a8_1330);
and ( n20911 , n51972 , n29614 );
or ( n51973 , n20910 , n20911 );
not ( n20912 , RI1754c610_2);
and ( n20913 , n20912 , n51973 );
and ( n20914 , C0 , RI1754c610_2);
or ( n51974 , n20913 , n20914 );
buf ( n51975 , n51974 );
not ( n51976 , n48685 );
and ( n51977 , n51976 , n48687 );
xor ( n51978 , n51884 , n51977 );
not ( n20915 , n29614 );
and ( n20916 , n20915 , RI173a8220_1936);
and ( n20917 , n51978 , n29614 );
or ( n51979 , n20916 , n20917 );
not ( n20918 , RI1754c610_2);
and ( n20919 , n20918 , n51979 );
and ( n20920 , C0 , RI1754c610_2);
or ( n51980 , n20919 , n20920 );
buf ( n51981 , n51980 );
not ( n20921 , n27683 );
and ( n20922 , n20921 , RI19a8be08_2712);
and ( n20923 , RI19a95de0_2641 , n27683 );
or ( n51982 , n20922 , n20923 );
not ( n20924 , RI1754c610_2);
and ( n20925 , n20924 , n51982 );
and ( n20926 , C0 , RI1754c610_2);
or ( n51983 , n20925 , n20926 );
buf ( n51984 , n51983 );
not ( n20927 , n27683 );
and ( n20928 , n20927 , RI19ac0158_2331);
and ( n20929 , RI19ac92a8_2261 , n27683 );
or ( n51985 , n20928 , n20929 );
not ( n20930 , RI1754c610_2);
and ( n20931 , n20930 , n51985 );
and ( n20932 , C0 , RI1754c610_2);
or ( n51986 , n20931 , n20932 );
buf ( n51987 , n51986 );
not ( n20933 , RI1754c610_2);
and ( n20934 , n20933 , RI19ad1060_2204);
and ( n20935 , C0 , RI1754c610_2);
or ( n51988 , n20934 , n20935 );
buf ( n51989 , n51988 );
not ( n51990 , n42878 );
and ( n51991 , n51990 , n51354 );
xor ( n51992 , n42875 , n51991 );
not ( n20936 , n29614 );
and ( n20937 , n20936 , RI173eaca0_1611);
and ( n20938 , n51992 , n29614 );
or ( n51993 , n20937 , n20938 );
not ( n20939 , RI1754c610_2);
and ( n20940 , n20939 , n51993 );
and ( n20941 , C0 , RI1754c610_2);
or ( n51994 , n20940 , n20941 );
buf ( n51995 , n51994 );
xor ( n51996 , n42604 , n38284 );
xor ( n51997 , n51996 , n39856 );
not ( n51998 , n45922 );
and ( n51999 , n51998 , n45924 );
xor ( n52000 , n51997 , n51999 );
not ( n20942 , n29614 );
and ( n20943 , n20942 , RI17332ae8_2194);
and ( n20944 , n52000 , n29614 );
or ( n52001 , n20943 , n20944 );
not ( n20945 , RI1754c610_2);
and ( n20946 , n20945 , n52001 );
and ( n20947 , C0 , RI1754c610_2);
or ( n52002 , n20946 , n20947 );
buf ( n52003 , n52002 );
not ( n20948 , n27683 );
and ( n20949 , n20948 , RI19ac92a8_2261);
and ( n20950 , RI19a843b0_2764 , n27683 );
or ( n52004 , n20949 , n20950 );
not ( n20951 , RI1754c610_2);
and ( n20952 , n20951 , n52004 );
and ( n20953 , C0 , RI1754c610_2);
or ( n52005 , n20952 , n20953 );
buf ( n52006 , n52005 );
not ( n52007 , n41995 );
and ( n52008 , n52007 , n46267 );
xor ( n52009 , n41992 , n52008 );
not ( n20954 , n29614 );
and ( n20955 , n20954 , RI17333178_2192);
and ( n20956 , n52009 , n29614 );
or ( n52010 , n20955 , n20956 );
not ( n20957 , RI1754c610_2);
and ( n20958 , n20957 , n52010 );
and ( n20959 , C0 , RI1754c610_2);
or ( n52011 , n20958 , n20959 );
buf ( n52012 , n52011 );
not ( n52013 , n46983 );
and ( n52014 , n52013 , n48296 );
xor ( n52015 , n46980 , n52014 );
not ( n20960 , n29614 );
and ( n20961 , n20960 , RI175191c0_688);
and ( n20962 , n52015 , n29614 );
or ( n52016 , n20961 , n20962 );
not ( n20963 , RI1754c610_2);
and ( n20964 , n20963 , n52016 );
and ( n20965 , C0 , RI1754c610_2);
or ( n52017 , n20964 , n20965 );
buf ( n52018 , n52017 );
not ( n52019 , n41010 );
and ( n52020 , n52019 , n33283 );
xor ( n52021 , n41007 , n52020 );
not ( n20966 , n29614 );
and ( n20967 , n20966 , RI173d3000_1727);
and ( n20968 , n52021 , n29614 );
or ( n52022 , n20967 , n20968 );
not ( n20969 , RI1754c610_2);
and ( n20970 , n20969 , n52022 );
and ( n20971 , C0 , RI1754c610_2);
or ( n52023 , n20970 , n20971 );
buf ( n52024 , n52023 );
not ( n52025 , n45878 );
xor ( n52026 , n40335 , n37987 );
xor ( n52027 , n52026 , n38037 );
and ( n52028 , n52025 , n52027 );
xor ( n52029 , n45875 , n52028 );
not ( n20972 , n29614 );
and ( n20973 , n20972 , RI174b1d50_869);
and ( n20974 , n52029 , n29614 );
or ( n52030 , n20973 , n20974 );
not ( n20975 , RI1754c610_2);
and ( n20976 , n20975 , n52030 );
and ( n20977 , C0 , RI1754c610_2);
or ( n52031 , n20976 , n20977 );
buf ( n52032 , n52031 );
not ( n52033 , n50021 );
and ( n52034 , n52033 , n45004 );
xor ( n52035 , n50018 , n52034 );
not ( n20978 , n29614 );
and ( n20979 , n20978 , RI17474b80_1167);
and ( n20980 , n52035 , n29614 );
or ( n52036 , n20979 , n20980 );
not ( n20981 , RI1754c610_2);
and ( n20982 , n20981 , n52036 );
and ( n20983 , C0 , RI1754c610_2);
or ( n52037 , n20982 , n20983 );
buf ( n52038 , n52037 );
xor ( n52039 , n33628 , n35069 );
xor ( n52040 , n52039 , n41854 );
not ( n52041 , n41513 );
and ( n52042 , n52041 , n41544 );
xor ( n52043 , n52040 , n52042 );
not ( n20984 , n29614 );
and ( n20985 , n20984 , RI1740fe88_1430);
and ( n20986 , n52043 , n29614 );
or ( n52044 , n20985 , n20986 );
not ( n20987 , RI1754c610_2);
and ( n20988 , n20987 , n52044 );
and ( n20989 , C0 , RI1754c610_2);
or ( n52045 , n20988 , n20989 );
buf ( n52046 , n52045 );
buf ( n52047 , RI174af5f0_881);
buf ( n52048 , RI174a3ae8_938);
buf ( n52049 , RI174793b0_1145);
xor ( n52050 , n31441 , n41287 );
xor ( n52051 , n52050 , n39935 );
not ( n52052 , n52051 );
and ( n52053 , n52052 , n48489 );
xor ( n52054 , n47989 , n52053 );
not ( n20990 , n29614 );
and ( n20991 , n20990 , RI17473488_1174);
and ( n20992 , n52054 , n29614 );
or ( n52055 , n20991 , n20992 );
not ( n20993 , RI1754c610_2);
and ( n20994 , n20993 , n52055 );
and ( n20995 , C0 , RI1754c610_2);
or ( n52056 , n20994 , n20995 );
buf ( n52057 , n52056 );
not ( n52058 , n39960 );
and ( n52059 , n52058 , n40010 );
xor ( n52060 , n41330 , n52059 );
not ( n20996 , n29614 );
and ( n20997 , n20996 , RI17458d40_1303);
and ( n20998 , n52060 , n29614 );
or ( n52061 , n20997 , n20998 );
not ( n20999 , RI1754c610_2);
and ( n21000 , n20999 , n52061 );
and ( n21001 , C0 , RI1754c610_2);
or ( n52062 , n21000 , n21001 );
buf ( n52063 , n52062 );
not ( n52064 , n45905 );
and ( n52065 , n52064 , n47400 );
xor ( n52066 , n44308 , n52065 );
not ( n21002 , n29614 );
and ( n21003 , n21002 , RI173d0bd0_1738);
and ( n21004 , n52066 , n29614 );
or ( n52067 , n21003 , n21004 );
not ( n21005 , RI1754c610_2);
and ( n21006 , n21005 , n52067 );
and ( n21007 , C0 , RI1754c610_2);
or ( n52068 , n21006 , n21007 );
buf ( n52069 , n52068 );
not ( n52070 , n34645 );
xor ( n52071 , n40429 , n39816 );
xor ( n52072 , n52071 , n35052 );
and ( n52073 , n52070 , n52072 );
xor ( n52074 , n34623 , n52073 );
not ( n21008 , n29614 );
and ( n21009 , n21008 , RI173458c8_2102);
and ( n21010 , n52074 , n29614 );
or ( n52075 , n21009 , n21010 );
not ( n21011 , RI1754c610_2);
and ( n21012 , n21011 , n52075 );
and ( n21013 , C0 , RI1754c610_2);
or ( n52076 , n21012 , n21013 );
buf ( n52077 , n52076 );
not ( n21014 , n27683 );
and ( n21015 , n21014 , RI19aa81e8_2508);
and ( n21016 , RI19ab2328_2438 , n27683 );
or ( n52078 , n21015 , n21016 );
not ( n21017 , RI1754c610_2);
and ( n21018 , n21017 , n52078 );
and ( n21019 , C0 , RI1754c610_2);
or ( n52079 , n21018 , n21019 );
buf ( n52080 , n52079 );
buf ( n52081 , RI174b3448_862);
buf ( n52082 , RI1749fc90_957);
buf ( n52083 , RI174996d8_988);
buf ( n52084 , RI174b9eb0_832);
not ( n21020 , n27683 );
and ( n21021 , n21020 , RI19abf2d0_2339);
and ( n21022 , RI19ac8330_2268 , n27683 );
or ( n52085 , n21021 , n21022 );
not ( n21023 , RI1754c610_2);
and ( n21024 , n21023 , n52085 );
and ( n21025 , C0 , RI1754c610_2);
or ( n52086 , n21024 , n21025 );
buf ( n52087 , n52086 );
not ( n52088 , n40595 );
and ( n52089 , n52088 , n40600 );
xor ( n52090 , n39155 , n52089 );
not ( n21026 , n29614 );
and ( n21027 , n21026 , RI173358d8_2180);
and ( n21028 , n52090 , n29614 );
or ( n52091 , n21027 , n21028 );
not ( n21029 , RI1754c610_2);
and ( n21030 , n21029 , n52091 );
and ( n21031 , C0 , RI1754c610_2);
or ( n52092 , n21030 , n21031 );
buf ( n52093 , n52092 );
xor ( n52094 , n33135 , n37235 );
xor ( n52095 , n52094 , n37255 );
not ( n52096 , n46851 );
and ( n52097 , n52096 , n46853 );
xor ( n52098 , n52095 , n52097 );
not ( n21032 , n29614 );
and ( n21033 , n21032 , RI17415090_1405);
and ( n21034 , n52098 , n29614 );
or ( n52099 , n21033 , n21034 );
not ( n21035 , RI1754c610_2);
and ( n21036 , n21035 , n52099 );
and ( n21037 , C0 , RI1754c610_2);
or ( n52100 , n21036 , n21037 );
buf ( n52101 , n52100 );
not ( n52102 , n43888 );
and ( n52103 , n52102 , n48092 );
xor ( n52104 , n37375 , n52103 );
not ( n21038 , n29614 );
and ( n21039 , n21038 , RI173d9900_1695);
and ( n21040 , n52104 , n29614 );
or ( n52105 , n21039 , n21040 );
not ( n21041 , RI1754c610_2);
and ( n21042 , n21041 , n52105 );
and ( n21043 , C0 , RI1754c610_2);
or ( n52106 , n21042 , n21043 );
buf ( n52107 , n52106 );
not ( n21044 , n27683 );
and ( n21045 , n21044 , RI19aa24a0_2550);
and ( n21046 , RI19aaca18_2478 , n27683 );
or ( n52108 , n21045 , n21046 );
not ( n21047 , RI1754c610_2);
and ( n21048 , n21047 , n52108 );
and ( n21049 , C0 , RI1754c610_2);
or ( n52109 , n21048 , n21049 );
buf ( n52110 , n52109 );
xor ( n52111 , n39038 , n36947 );
xor ( n52112 , n52111 , n39702 );
not ( n52113 , n52040 );
and ( n52114 , n52113 , n41513 );
xor ( n52115 , n52112 , n52114 );
not ( n21050 , n29614 );
and ( n21051 , n21050 , RI173db688_1686);
and ( n21052 , n52115 , n29614 );
or ( n52116 , n21051 , n21052 );
not ( n21053 , RI1754c610_2);
and ( n21054 , n21053 , n52116 );
and ( n21055 , C0 , RI1754c610_2);
or ( n52117 , n21054 , n21055 );
buf ( n52118 , n52117 );
not ( n52119 , n51805 );
and ( n52120 , n52119 , n45804 );
xor ( n52121 , n51802 , n52120 );
not ( n21056 , n29614 );
and ( n21057 , n21056 , RI1751d4c8_675);
and ( n21058 , n52121 , n29614 );
or ( n52122 , n21057 , n21058 );
not ( n21059 , RI1754c610_2);
and ( n21060 , n21059 , n52122 );
and ( n21061 , C0 , RI1754c610_2);
or ( n52123 , n21060 , n21061 );
buf ( n52124 , n52123 );
xor ( n52125 , n38068 , n40091 );
xor ( n52126 , n52125 , n40111 );
not ( n52127 , n52126 );
and ( n52128 , n52127 , n47850 );
xor ( n52129 , n51453 , n52128 );
not ( n21062 , n29614 );
and ( n21063 , n21062 , RI1738dad8_2065);
and ( n21064 , n52129 , n29614 );
or ( n52130 , n21063 , n21064 );
not ( n21065 , RI1754c610_2);
and ( n21066 , n21065 , n52130 );
and ( n21067 , C0 , RI1754c610_2);
or ( n52131 , n21066 , n21067 );
buf ( n52132 , n52131 );
xor ( n52133 , n33000 , n35639 );
xor ( n52134 , n52133 , n36227 );
not ( n52135 , n52134 );
and ( n52136 , n52135 , n51927 );
xor ( n52137 , n39747 , n52136 );
not ( n21068 , n29614 );
and ( n21069 , n21068 , RI17404a10_1485);
and ( n21070 , n52137 , n29614 );
or ( n52138 , n21069 , n21070 );
not ( n21071 , RI1754c610_2);
and ( n21072 , n21071 , n52138 );
and ( n21073 , C0 , RI1754c610_2);
or ( n52139 , n21072 , n21073 );
buf ( n52140 , n52139 );
not ( n52141 , n46670 );
and ( n52142 , n52141 , n42429 );
xor ( n52143 , n47139 , n52142 );
not ( n21074 , n29614 );
and ( n21075 , n21074 , RI174896e8_1066);
and ( n21076 , n52143 , n29614 );
or ( n52144 , n21075 , n21076 );
not ( n21077 , RI1754c610_2);
and ( n21078 , n21077 , n52144 );
and ( n21079 , C0 , RI1754c610_2);
or ( n52145 , n21078 , n21079 );
buf ( n52146 , n52145 );
not ( n52147 , n39887 );
and ( n52148 , n52147 , n43981 );
xor ( n52149 , n39833 , n52148 );
not ( n21080 , n29614 );
and ( n21081 , n21080 , RI1740ca08_1446);
and ( n21082 , n52149 , n29614 );
or ( n52150 , n21081 , n21082 );
not ( n21083 , RI1754c610_2);
and ( n21084 , n21083 , n52150 );
and ( n21085 , C0 , RI1754c610_2);
or ( n52151 , n21084 , n21085 );
buf ( n52152 , n52151 );
not ( n21086 , n27683 );
and ( n21087 , n21086 , RI19ac6e18_2278);
and ( n21088 , RI19acf8d8_2214 , n27683 );
or ( n52153 , n21087 , n21088 );
not ( n21089 , RI1754c610_2);
and ( n21090 , n21089 , n52153 );
and ( n21091 , C0 , RI1754c610_2);
or ( n52154 , n21090 , n21091 );
buf ( n52155 , n52154 );
not ( n52156 , n43160 );
and ( n52157 , n52156 , n43162 );
xor ( n52158 , n45591 , n52157 );
not ( n21092 , n29614 );
and ( n21093 , n21092 , RI1745cee0_1283);
and ( n21094 , n52158 , n29614 );
or ( n52159 , n21093 , n21094 );
not ( n21095 , RI1754c610_2);
and ( n21096 , n21095 , n52159 );
and ( n21097 , C0 , RI1754c610_2);
or ( n52160 , n21096 , n21097 );
buf ( n52161 , n52160 );
not ( n21098 , n27683 );
and ( n21099 , n21098 , RI19a95de0_2641);
and ( n21100 , RI19a9fae8_2571 , n27683 );
or ( n52162 , n21099 , n21100 );
not ( n21101 , RI1754c610_2);
and ( n21102 , n21101 , n52162 );
and ( n21103 , C0 , RI1754c610_2);
or ( n52163 , n21102 , n21103 );
buf ( n52164 , n52163 );
not ( n52165 , n42402 );
and ( n52166 , n52165 , n41780 );
xor ( n52167 , n42399 , n52166 );
not ( n21104 , n29614 );
and ( n21105 , n21104 , RI17401590_1501);
and ( n21106 , n52167 , n29614 );
or ( n52168 , n21105 , n21106 );
not ( n21107 , RI1754c610_2);
and ( n21108 , n21107 , n52168 );
and ( n21109 , C0 , RI1754c610_2);
or ( n52169 , n21108 , n21109 );
buf ( n52170 , n52169 );
not ( n52171 , n45519 );
and ( n52172 , n52171 , n46153 );
xor ( n52173 , n45516 , n52172 );
not ( n21110 , n29614 );
and ( n21111 , n21110 , RI173ca960_1768);
and ( n21112 , n52173 , n29614 );
or ( n52174 , n21111 , n21112 );
not ( n21113 , RI1754c610_2);
and ( n21114 , n21113 , n52174 );
and ( n21115 , C0 , RI1754c610_2);
or ( n52175 , n21114 , n21115 );
buf ( n52176 , n52175 );
not ( n21116 , n27683 );
and ( n21117 , n21116 , RI19a9e468_2582);
and ( n21118 , RI19aa7e28_2510 , n27683 );
or ( n52177 , n21117 , n21118 );
not ( n21119 , RI1754c610_2);
and ( n21120 , n21119 , n52177 );
and ( n21121 , C0 , RI1754c610_2);
or ( n52178 , n21120 , n21121 );
buf ( n52179 , n52178 );
xor ( n52180 , n34461 , n33453 );
xor ( n52181 , n52180 , n33505 );
xor ( n52182 , n37974 , n41504 );
xor ( n52183 , n52182 , n41690 );
not ( n52184 , n52183 );
xor ( n52185 , n38108 , n40111 );
xor ( n52186 , n52185 , n43278 );
and ( n52187 , n52184 , n52186 );
xor ( n52188 , n52181 , n52187 );
not ( n21122 , n29614 );
and ( n21123 , n21122 , RI17459718_1300);
and ( n21124 , n52188 , n29614 );
or ( n52189 , n21123 , n21124 );
not ( n21125 , RI1754c610_2);
and ( n21126 , n21125 , n52189 );
and ( n21127 , C0 , RI1754c610_2);
or ( n52190 , n21126 , n21127 );
buf ( n52191 , n52190 );
not ( n52192 , n46414 );
and ( n52193 , n52192 , n44536 );
xor ( n52194 , n38449 , n52193 );
not ( n21128 , n29614 );
and ( n21129 , n21128 , RI1733cef8_2144);
and ( n21130 , n52194 , n29614 );
or ( n52195 , n21129 , n21130 );
not ( n21131 , RI1754c610_2);
and ( n21132 , n21131 , n52195 );
and ( n21133 , C0 , RI1754c610_2);
or ( n52196 , n21132 , n21133 );
buf ( n52197 , n52196 );
and ( n52198 , RI1754ba58_27 , n34844 );
and ( n52199 , RI1754ba58_27 , n34847 );
and ( n52200 , RI1754ba58_27 , n34850 );
and ( n52201 , RI1754ba58_27 , n34852 );
or ( n52202 , n52198 , n52199 , n52200 , n52201 , C0 , C0 , C0 , C0 );
not ( n21134 , n34859 );
and ( n21135 , n21134 , n52202 );
and ( n21136 , RI1754ba58_27 , n34859 );
or ( n52203 , n21135 , n21136 );
not ( n21137 , RI19a22f70_2797);
and ( n21138 , n21137 , n52203 );
and ( n21139 , C0 , RI19a22f70_2797);
or ( n52204 , n21138 , n21139 );
not ( n21140 , n27683 );
and ( n21141 , n21140 , RI19aa4318_2536);
and ( n21142 , n52204 , n27683 );
or ( n52205 , n21141 , n21142 );
not ( n21143 , RI1754c610_2);
and ( n21144 , n21143 , n52205 );
and ( n21145 , C0 , RI1754c610_2);
or ( n52206 , n21144 , n21145 );
buf ( n52207 , n52206 );
xor ( n52208 , n34828 , n41478 );
xor ( n52209 , n52208 , n41146 );
not ( n52210 , n52209 );
and ( n52211 , n52210 , n45307 );
xor ( n52212 , n47226 , n52211 );
not ( n21146 , n29614 );
and ( n21147 , n21146 , RI17512050_710);
and ( n21148 , n52212 , n29614 );
or ( n52213 , n21147 , n21148 );
not ( n21149 , RI1754c610_2);
and ( n21150 , n21149 , n52213 );
and ( n21151 , C0 , RI1754c610_2);
or ( n52214 , n21150 , n21151 );
buf ( n52215 , n52214 );
not ( n52216 , n43050 );
and ( n52217 , n52216 , n42723 );
xor ( n52218 , n43047 , n52217 );
not ( n21152 , n29614 );
and ( n21153 , n21152 , RI17527ef0_642);
and ( n21154 , n52218 , n29614 );
or ( n52219 , n21153 , n21154 );
not ( n21155 , RI1754c610_2);
and ( n21156 , n21155 , n52219 );
and ( n21157 , C0 , RI1754c610_2);
or ( n52220 , n21156 , n21157 );
buf ( n52221 , n52220 );
buf ( n52222 , RI17487618_1076);
buf ( n52223 , RI1747a760_1139);
buf ( n52224 , RI17507100_744);
not ( n52225 , n48289 );
xor ( n52226 , n37144 , n40254 );
xor ( n52227 , n52226 , n40718 );
and ( n52228 , n52225 , n52227 );
xor ( n52229 , n48286 , n52228 );
not ( n21158 , n29614 );
and ( n21159 , n21158 , RI1733a798_2156);
and ( n21160 , n52229 , n29614 );
or ( n52230 , n21159 , n21160 );
not ( n21161 , RI1754c610_2);
and ( n21162 , n21161 , n52230 );
and ( n21163 , C0 , RI1754c610_2);
or ( n52231 , n21162 , n21163 );
buf ( n52232 , n52231 );
not ( n52233 , n46406 );
and ( n52234 , n52233 , n45995 );
xor ( n52235 , n46403 , n52234 );
not ( n21164 , n29614 );
and ( n21165 , n21164 , RI1733d8d0_2141);
and ( n21166 , n52235 , n29614 );
or ( n52236 , n21165 , n21166 );
not ( n21167 , RI1754c610_2);
and ( n21168 , n21167 , n52236 );
and ( n21169 , C0 , RI1754c610_2);
or ( n52237 , n21168 , n21169 );
buf ( n52238 , n52237 );
not ( n52239 , n48962 );
and ( n52240 , n52239 , n48964 );
xor ( n52241 , n43626 , n52240 );
not ( n21170 , n29614 );
and ( n21171 , n21170 , RI174bdc90_820);
and ( n21172 , n52241 , n29614 );
or ( n52242 , n21171 , n21172 );
not ( n21173 , RI1754c610_2);
and ( n21174 , n21173 , n52242 );
and ( n21175 , C0 , RI1754c610_2);
or ( n52243 , n21174 , n21175 );
buf ( n52244 , n52243 );
not ( n21176 , n27683 );
and ( n21177 , n21176 , RI19a96e48_2634);
and ( n21178 , RI19aa0970_2564 , n27683 );
or ( n52245 , n21177 , n21178 );
not ( n21179 , RI1754c610_2);
and ( n21180 , n21179 , n52245 );
and ( n21181 , C0 , RI1754c610_2);
or ( n52246 , n21180 , n21181 );
buf ( n52247 , n52246 );
buf ( n52248 , RI17481a38_1104);
buf ( n52249 , RI17462e08_1254);
xor ( n52250 , n36748 , n39208 );
xor ( n52251 , n52250 , n38214 );
xor ( n52252 , n41730 , n34837 );
xor ( n52253 , n52252 , n33880 );
not ( n52254 , n52253 );
and ( n52255 , n52254 , n46658 );
xor ( n52256 , n52251 , n52255 );
not ( n21182 , n29614 );
and ( n21183 , n21182 , RI173413e0_2123);
and ( n21184 , n52256 , n29614 );
or ( n52257 , n21183 , n21184 );
not ( n21185 , RI1754c610_2);
and ( n21186 , n21185 , n52257 );
and ( n21187 , C0 , RI1754c610_2);
or ( n52258 , n21186 , n21187 );
buf ( n52259 , n52258 );
not ( n52260 , n50541 );
and ( n52261 , n52260 , n47247 );
xor ( n52262 , n45794 , n52261 );
not ( n21188 , n29614 );
and ( n21189 , n21188 , RI17340a08_2126);
and ( n21190 , n52262 , n29614 );
or ( n52263 , n21189 , n21190 );
not ( n21191 , RI1754c610_2);
and ( n21192 , n21191 , n52263 );
and ( n21193 , C0 , RI1754c610_2);
or ( n52264 , n21192 , n21193 );
buf ( n52265 , n52264 );
buf ( n52266 , RI17516880_696);
not ( n52267 , n51113 );
and ( n52268 , n52267 , n49053 );
xor ( n52269 , n43212 , n52268 );
not ( n21194 , n29614 );
and ( n21195 , n21194 , RI174916e0_1027);
and ( n21196 , n52269 , n29614 );
or ( n52270 , n21195 , n21196 );
not ( n21197 , RI1754c610_2);
and ( n21198 , n21197 , n52270 );
and ( n21199 , C0 , RI1754c610_2);
or ( n52271 , n21198 , n21199 );
buf ( n52272 , n52271 );
not ( n52273 , n49819 );
and ( n52274 , n52273 , n49821 );
xor ( n52275 , n43814 , n52274 );
not ( n21200 , n29614 );
and ( n21201 , n21200 , RI174046c8_1486);
and ( n21202 , n52275 , n29614 );
or ( n52276 , n21201 , n21202 );
not ( n21203 , RI1754c610_2);
and ( n21204 , n21203 , n52276 );
and ( n21205 , C0 , RI1754c610_2);
or ( n52277 , n21204 , n21205 );
buf ( n52278 , n52277 );
not ( n52279 , n39747 );
and ( n52280 , n52279 , n52134 );
xor ( n52281 , n39741 , n52280 );
not ( n21206 , n29614 );
and ( n21207 , n21206 , RI173f5dd0_1557);
and ( n21208 , n52281 , n29614 );
or ( n52282 , n21207 , n21208 );
not ( n21209 , RI1754c610_2);
and ( n21210 , n21209 , n52282 );
and ( n21211 , C0 , RI1754c610_2);
or ( n52283 , n21210 , n21211 );
buf ( n52284 , n52283 );
xor ( n52285 , n39466 , n36611 );
xor ( n52286 , n52285 , n33567 );
not ( n52287 , n52286 );
and ( n52288 , n52287 , n44685 );
xor ( n52289 , n46461 , n52288 );
not ( n21212 , n29614 );
and ( n21213 , n21212 , RI173aa638_1925);
and ( n21214 , n52289 , n29614 );
or ( n52290 , n21213 , n21214 );
not ( n21215 , RI1754c610_2);
and ( n21216 , n21215 , n52290 );
and ( n21217 , C0 , RI1754c610_2);
or ( n52291 , n21216 , n21217 );
buf ( n52292 , n52291 );
not ( n52293 , n39307 );
and ( n52294 , n52293 , n44799 );
xor ( n52295 , n39304 , n52294 );
not ( n21218 , n29614 );
and ( n21219 , n21218 , RI173af1b0_1902);
and ( n21220 , n52295 , n29614 );
or ( n52296 , n21219 , n21220 );
not ( n21221 , RI1754c610_2);
and ( n21222 , n21221 , n52296 );
and ( n21223 , C0 , RI1754c610_2);
or ( n52297 , n21222 , n21223 );
buf ( n52298 , n52297 );
not ( n52299 , n49630 );
and ( n52300 , n52299 , n46383 );
xor ( n52301 , n45672 , n52300 );
not ( n21224 , n29614 );
and ( n21225 , n21224 , RI173bcd88_1835);
and ( n21226 , n52301 , n29614 );
or ( n52302 , n21225 , n21226 );
not ( n21227 , RI1754c610_2);
and ( n21228 , n21227 , n52302 );
and ( n21229 , C0 , RI1754c610_2);
or ( n52303 , n21228 , n21229 );
buf ( n52304 , n52303 );
not ( n52305 , n47783 );
and ( n52306 , n52305 , n50580 );
xor ( n52307 , n47780 , n52306 );
not ( n21230 , n29614 );
and ( n21231 , n21230 , RI1749e8e0_963);
and ( n21232 , n52307 , n29614 );
or ( n52308 , n21231 , n21232 );
not ( n21233 , RI1754c610_2);
and ( n21234 , n21233 , n52308 );
and ( n21235 , C0 , RI1754c610_2);
or ( n52309 , n21234 , n21235 );
buf ( n52310 , n52309 );
buf ( n52311 , RI17498d00_991);
not ( n21236 , n27683 );
and ( n21237 , n21236 , RI19ab4740_2420);
and ( n21238 , RI19abdf98_2350 , n27683 );
or ( n52312 , n21237 , n21238 );
not ( n21239 , RI1754c610_2);
and ( n21240 , n21239 , n52312 );
and ( n21241 , C0 , RI1754c610_2);
or ( n52313 , n21240 , n21241 );
buf ( n52314 , n52313 );
xor ( n52315 , n28188 , n41799 );
xor ( n52316 , n52315 , n40381 );
not ( n52317 , n43690 );
and ( n52318 , n52317 , n43692 );
xor ( n52319 , n52316 , n52318 );
not ( n21242 , n29614 );
and ( n21243 , n21242 , RI1733f9a0_2131);
and ( n21244 , n52319 , n29614 );
or ( n52320 , n21243 , n21244 );
not ( n21245 , RI1754c610_2);
and ( n21246 , n21245 , n52320 );
and ( n21247 , C0 , RI1754c610_2);
or ( n52321 , n21246 , n21247 );
buf ( n52322 , n52321 );
buf ( n52323 , RI174bb350_828);
not ( n52324 , n49394 );
and ( n52325 , n52324 , n44755 );
xor ( n52326 , n46516 , n52325 );
not ( n21248 , n29614 );
and ( n21249 , n21248 , RI17409c18_1460);
and ( n21250 , n52326 , n29614 );
or ( n52327 , n21249 , n21250 );
not ( n21251 , RI1754c610_2);
and ( n21252 , n21251 , n52327 );
and ( n21253 , C0 , RI1754c610_2);
or ( n52328 , n21252 , n21253 );
buf ( n52329 , n52328 );
not ( n52330 , n41029 );
and ( n52331 , n52330 , n41050 );
xor ( n52332 , n49708 , n52331 );
not ( n21254 , n29614 );
and ( n21255 , n21254 , RI17494ea8_1010);
and ( n21256 , n52332 , n29614 );
or ( n52333 , n21255 , n21256 );
not ( n21257 , RI1754c610_2);
and ( n21258 , n21257 , n52333 );
and ( n21259 , C0 , RI1754c610_2);
or ( n52334 , n21258 , n21259 );
buf ( n52335 , n52334 );
xor ( n52336 , n39558 , n38401 );
xor ( n52337 , n52336 , n41068 );
not ( n52338 , n52337 );
and ( n52339 , n52338 , n45873 );
xor ( n52340 , n52027 , n52339 );
not ( n21260 , n29614 );
and ( n21261 , n21260 , RI1750c8a8_727);
and ( n21262 , n52340 , n29614 );
or ( n52341 , n21261 , n21262 );
not ( n21263 , RI1754c610_2);
and ( n21264 , n21263 , n52341 );
and ( n21265 , C0 , RI1754c610_2);
or ( n52342 , n21264 , n21265 );
buf ( n52343 , n52342 );
xor ( n52344 , n36673 , n39635 );
xor ( n52345 , n52344 , n39655 );
not ( n52346 , n52345 );
xor ( n52347 , n34118 , n42377 );
xor ( n52348 , n52347 , n33991 );
and ( n52349 , n52346 , n52348 );
xor ( n52350 , n45134 , n52349 );
not ( n21266 , n29614 );
and ( n21267 , n21266 , RI17472768_1178);
and ( n21268 , n52350 , n29614 );
or ( n52351 , n21267 , n21268 );
not ( n21269 , RI1754c610_2);
and ( n21270 , n21269 , n52351 );
and ( n21271 , C0 , RI1754c610_2);
or ( n52352 , n21270 , n21271 );
buf ( n52353 , n52352 );
not ( n52354 , n41443 );
and ( n52355 , n52354 , n41445 );
xor ( n52356 , n43860 , n52355 );
not ( n21272 , n29614 );
and ( n21273 , n21272 , RI173ae148_1907);
and ( n21274 , n52356 , n29614 );
or ( n52357 , n21273 , n21274 );
not ( n21275 , RI1754c610_2);
and ( n21276 , n21275 , n52357 );
and ( n21277 , C0 , RI1754c610_2);
or ( n52358 , n21276 , n21277 );
buf ( n52359 , n52358 );
not ( n52360 , n45307 );
and ( n52361 , n52360 , n45309 );
xor ( n52362 , n52209 , n52361 );
not ( n21278 , n29614 );
and ( n21279 , n21278 , RI17529390_638);
and ( n21280 , n52362 , n29614 );
or ( n52363 , n21279 , n21280 );
not ( n21281 , RI1754c610_2);
and ( n21282 , n21281 , n52363 );
and ( n21283 , C0 , RI1754c610_2);
or ( n52364 , n21282 , n21283 );
buf ( n52365 , n52364 );
not ( n52366 , n43363 );
and ( n52367 , n52366 , n42932 );
xor ( n52368 , n47420 , n52367 );
not ( n21284 , n29614 );
and ( n21285 , n21284 , RI173d4d88_1718);
and ( n21286 , n52368 , n29614 );
or ( n52369 , n21285 , n21286 );
not ( n21287 , RI1754c610_2);
and ( n21288 , n21287 , n52369 );
and ( n21289 , C0 , RI1754c610_2);
or ( n52370 , n21288 , n21289 );
buf ( n52371 , n52370 );
and ( n52372 , RI1754c340_8 , n34844 );
and ( n52373 , RI1754c340_8 , n34847 );
and ( n52374 , RI1754c340_8 , n34850 );
and ( n52375 , RI1754c340_8 , n34852 );
and ( n52376 , RI1754c340_8 , n34854 );
and ( n52377 , RI1754c340_8 , n34856 );
and ( n52378 , RI1754c340_8 , n39233 );
or ( n52379 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , C0 );
not ( n21290 , n34859 );
and ( n21291 , n21290 , n52379 );
and ( n21292 , RI1754c340_8 , n34859 );
or ( n52380 , n21291 , n21292 );
not ( n21293 , RI19a22f70_2797);
and ( n21294 , n21293 , n52380 );
and ( n21295 , C0 , RI19a22f70_2797);
or ( n52381 , n21294 , n21295 );
not ( n21296 , n27683 );
and ( n21297 , n21296 , RI19a88be0_2733);
and ( n21298 , n52381 , n27683 );
or ( n52382 , n21297 , n21298 );
not ( n21299 , RI1754c610_2);
and ( n21300 , n21299 , n52382 );
and ( n21301 , C0 , RI1754c610_2);
or ( n52383 , n21300 , n21301 );
buf ( n52384 , n52383 );
not ( n52385 , n44108 );
and ( n52386 , n52385 , n47295 );
xor ( n52387 , n43974 , n52386 );
not ( n21302 , n29614 );
and ( n21303 , n21302 , RI1750aee0_732);
and ( n21304 , n52387 , n29614 );
or ( n52388 , n21303 , n21304 );
not ( n21305 , RI1754c610_2);
and ( n21306 , n21305 , n52388 );
and ( n21307 , C0 , RI1754c610_2);
or ( n52389 , n21306 , n21307 );
buf ( n52390 , n52389 );
not ( n21308 , n27683 );
and ( n21309 , n21308 , RI19a95930_2643);
and ( n21310 , RI19a9f728_2573 , n27683 );
or ( n52391 , n21309 , n21310 );
not ( n21311 , RI1754c610_2);
and ( n21312 , n21311 , n52391 );
and ( n21313 , C0 , RI1754c610_2);
or ( n52392 , n21312 , n21313 );
buf ( n52393 , n52392 );
not ( n21314 , n27683 );
and ( n21315 , n21314 , RI19ac7958_2273);
and ( n21316 , RI19a82790_2777 , n27683 );
or ( n52394 , n21315 , n21316 );
not ( n21317 , RI1754c610_2);
and ( n21318 , n21317 , n52394 );
and ( n21319 , C0 , RI1754c610_2);
or ( n52395 , n21318 , n21319 );
buf ( n52396 , n52395 );
not ( n52397 , n47202 );
and ( n52398 , n52397 , n31054 );
xor ( n52399 , n48883 , n52398 );
not ( n21320 , n29614 );
and ( n21321 , n21320 , RI1750f710_718);
and ( n21322 , n52399 , n29614 );
or ( n52400 , n21321 , n21322 );
not ( n21323 , RI1754c610_2);
and ( n21324 , n21323 , n52400 );
and ( n21325 , C0 , RI1754c610_2);
or ( n52401 , n21324 , n21325 );
buf ( n52402 , n52401 );
not ( n52403 , n43285 );
and ( n52404 , n52403 , n47768 );
xor ( n52405 , n43282 , n52404 );
not ( n21326 , n29614 );
and ( n21327 , n21326 , RI174b3e20_859);
and ( n21328 , n52405 , n29614 );
or ( n52406 , n21327 , n21328 );
not ( n21329 , RI1754c610_2);
and ( n21330 , n21329 , n52406 );
and ( n21331 , C0 , RI1754c610_2);
or ( n52407 , n21330 , n21331 );
buf ( n52408 , n52407 );
not ( n52409 , n51970 );
xor ( n52410 , n40008 , n40341 );
xor ( n52411 , n52410 , n40091 );
and ( n52412 , n52409 , n52411 );
xor ( n52413 , n36948 , n52412 );
not ( n21332 , n29614 );
and ( n21333 , n21332 , RI1746a0e0_1219);
and ( n21334 , n52413 , n29614 );
or ( n52414 , n21333 , n21334 );
not ( n21335 , RI1754c610_2);
and ( n21336 , n21335 , n52414 );
and ( n21337 , C0 , RI1754c610_2);
or ( n52415 , n21336 , n21337 );
buf ( n52416 , n52415 );
not ( n21338 , n27683 );
and ( n21339 , n21338 , RI19a954f8_2645);
and ( n21340 , RI19a9f368_2575 , n27683 );
or ( n52417 , n21339 , n21340 );
not ( n21341 , RI1754c610_2);
and ( n21342 , n21341 , n52417 );
and ( n21343 , C0 , RI1754c610_2);
or ( n52418 , n21342 , n21343 );
buf ( n52419 , n52418 );
not ( n52420 , n44152 );
and ( n52421 , n52420 , n51442 );
xor ( n52422 , n44149 , n52421 );
not ( n21344 , n29614 );
and ( n21345 , n21344 , RI17479d88_1142);
and ( n21346 , n52422 , n29614 );
or ( n52423 , n21345 , n21346 );
not ( n21347 , RI1754c610_2);
and ( n21348 , n21347 , n52423 );
and ( n21349 , C0 , RI1754c610_2);
or ( n52424 , n21348 , n21349 );
buf ( n52425 , n52424 );
buf ( n52426 , RI174c43b0_800);
buf ( n52427 , RI17471700_1183);
buf ( n52428 , RI17493468_1018);
xor ( n52429 , n40110 , n39740 );
xor ( n52430 , n52429 , n41099 );
not ( n52431 , n52430 );
and ( n52432 , n52431 , n50714 );
xor ( n52433 , n50485 , n52432 );
not ( n21350 , n29614 );
and ( n21351 , n21350 , RI17492a90_1021);
and ( n21352 , n52433 , n29614 );
or ( n52434 , n21351 , n21352 );
not ( n21353 , RI1754c610_2);
and ( n21354 , n21353 , n52434 );
and ( n21355 , C0 , RI1754c610_2);
or ( n52435 , n21354 , n21355 );
buf ( n52436 , n52435 );
not ( n21356 , n27683 );
and ( n21357 , n21356 , RI19abfa50_2335);
and ( n21358 , RI19ac89c0_2265 , n27683 );
or ( n52437 , n21357 , n21358 );
not ( n21359 , RI1754c610_2);
and ( n21360 , n21359 , n52437 );
and ( n21361 , C0 , RI1754c610_2);
or ( n52438 , n21360 , n21361 );
buf ( n52439 , n52438 );
not ( n21362 , n27683 );
and ( n21363 , n21362 , RI19a9af70_2605);
and ( n21364 , RI19aa48b8_2533 , n27683 );
or ( n52440 , n21363 , n21364 );
not ( n21365 , RI1754c610_2);
and ( n21366 , n21365 , n52440 );
and ( n21367 , C0 , RI1754c610_2);
or ( n52441 , n21366 , n21367 );
buf ( n52442 , n52441 );
not ( n21368 , n27683 );
and ( n21369 , n21368 , RI19a8a2d8_2723);
and ( n21370 , RI19a94238_2653 , n27683 );
or ( n52443 , n21369 , n21370 );
not ( n21371 , RI1754c610_2);
and ( n21372 , n21371 , n52443 );
and ( n21373 , C0 , RI1754c610_2);
or ( n52444 , n21372 , n21373 );
buf ( n52445 , n52444 );
not ( n21374 , n34859 );
and ( n21375 , n21374 , C0 );
and ( n21376 , RI1754aa68_61 , n34859 );
or ( n52446 , n21375 , n21376 );
not ( n21377 , RI19a22f70_2797);
and ( n21378 , n21377 , n52446 );
and ( n21379 , C0 , RI19a22f70_2797);
or ( n52447 , n21378 , n21379 );
not ( n21380 , n27683 );
and ( n21381 , n21380 , RI19a887a8_2735);
and ( n21382 , n52447 , n27683 );
or ( n52448 , n21381 , n21382 );
not ( n21383 , RI1754c610_2);
and ( n21384 , n21383 , n52448 );
and ( n21385 , C0 , RI1754c610_2);
or ( n52449 , n21384 , n21385 );
buf ( n52450 , n52449 );
not ( n52451 , n45603 );
and ( n52452 , n52451 , n43566 );
xor ( n52453 , n48659 , n52452 );
not ( n21386 , n29614 );
and ( n21387 , n21386 , RI1738ca70_2070);
and ( n21388 , n52453 , n29614 );
or ( n52454 , n21387 , n21388 );
not ( n21389 , RI1754c610_2);
and ( n21390 , n21389 , n52454 );
and ( n21391 , C0 , RI1754c610_2);
or ( n52455 , n21390 , n21391 );
buf ( n52456 , n52455 );
not ( n52457 , n46921 );
and ( n52458 , n52457 , n47646 );
xor ( n52459 , n46918 , n52458 );
not ( n21392 , n29614 );
and ( n21393 , n21392 , RI17413650_1413);
and ( n21394 , n52459 , n29614 );
or ( n52460 , n21393 , n21394 );
not ( n21395 , RI1754c610_2);
and ( n21396 , n21395 , n52460 );
and ( n21397 , C0 , RI1754c610_2);
or ( n52461 , n21396 , n21397 );
buf ( n52462 , n52461 );
not ( n52463 , n45617 );
and ( n52464 , n52463 , n48745 );
xor ( n52465 , n45614 , n52464 );
not ( n21398 , n29614 );
and ( n21399 , n21398 , RI17491d70_1025);
and ( n21400 , n52465 , n29614 );
or ( n52466 , n21399 , n21400 );
not ( n21401 , RI1754c610_2);
and ( n21402 , n21401 , n52466 );
and ( n21403 , C0 , RI1754c610_2);
or ( n52467 , n21402 , n21403 );
buf ( n52468 , n52467 );
not ( n52469 , n46186 );
and ( n52470 , n52469 , n46254 );
xor ( n52471 , n46183 , n52470 );
not ( n21404 , n29614 );
and ( n21405 , n21404 , RI1747b480_1135);
and ( n21406 , n52471 , n29614 );
or ( n52472 , n21405 , n21406 );
not ( n21407 , RI1754c610_2);
and ( n21408 , n21407 , n52472 );
and ( n21409 , C0 , RI1754c610_2);
or ( n52473 , n21408 , n21409 );
buf ( n52474 , n52473 );
not ( n21410 , n27683 );
and ( n21411 , n21410 , RI19aa6640_2520);
and ( n21412 , RI19ab0870_2450 , n27683 );
or ( n52475 , n21411 , n21412 );
not ( n21413 , RI1754c610_2);
and ( n21414 , n21413 , n52475 );
and ( n21415 , C0 , RI1754c610_2);
or ( n52476 , n21414 , n21415 );
buf ( n52477 , n52476 );
not ( n21416 , n27683 );
and ( n21417 , n21416 , RI19aa5740_2526);
and ( n21418 , RI19aafcb8_2455 , n27683 );
or ( n52478 , n21417 , n21418 );
not ( n21419 , RI1754c610_2);
and ( n21420 , n21419 , n52478 );
and ( n21421 , C0 , RI1754c610_2);
or ( n52479 , n21420 , n21421 );
buf ( n52480 , n52479 );
not ( n21422 , n27683 );
and ( n21423 , n21422 , RI19aa44f8_2535);
and ( n21424 , RI19aae7a0_2465 , n27683 );
or ( n52481 , n21423 , n21424 );
not ( n21425 , RI1754c610_2);
and ( n21426 , n21425 , n52481 );
and ( n21427 , C0 , RI1754c610_2);
or ( n52482 , n21426 , n21427 );
buf ( n52483 , n52482 );
not ( n52484 , n46663 );
and ( n52485 , n52484 , n52251 );
xor ( n52486 , n46660 , n52485 );
not ( n21428 , n29614 );
and ( n21429 , n21428 , RI173ad770_1910);
and ( n21430 , n52486 , n29614 );
or ( n52487 , n21429 , n21430 );
not ( n21431 , RI1754c610_2);
and ( n21432 , n21431 , n52487 );
and ( n21433 , C0 , RI1754c610_2);
or ( n52488 , n21432 , n21433 );
buf ( n52489 , n52488 );
not ( n52490 , n50561 );
and ( n52491 , n52490 , n44333 );
xor ( n52492 , n45360 , n52491 );
not ( n21434 , n29614 );
and ( n21435 , n21434 , RI173a3d38_1957);
and ( n21436 , n52492 , n29614 );
or ( n52493 , n21435 , n21436 );
not ( n21437 , RI1754c610_2);
and ( n21438 , n21437 , n52493 );
and ( n21439 , C0 , RI1754c610_2);
or ( n52494 , n21438 , n21439 );
buf ( n52495 , n52494 );
not ( n52496 , n46698 );
and ( n52497 , n52496 , n44447 );
xor ( n52498 , n46695 , n52497 );
not ( n21440 , n29614 );
and ( n21441 , n21440 , RI17509518_737);
and ( n21442 , n52498 , n29614 );
or ( n52499 , n21441 , n21442 );
not ( n21443 , RI1754c610_2);
and ( n21444 , n21443 , n52499 );
and ( n21445 , C0 , RI1754c610_2);
or ( n52500 , n21444 , n21445 );
buf ( n52501 , n52500 );
xor ( n52502 , n36645 , n40412 );
xor ( n52503 , n52502 , n40437 );
not ( n52504 , n52503 );
and ( n52505 , n52504 , n49916 );
xor ( n52506 , n49070 , n52505 );
not ( n21446 , n29614 );
and ( n21447 , n21446 , RI173ee468_1594);
and ( n21448 , n52506 , n29614 );
or ( n52507 , n21447 , n21448 );
not ( n21449 , RI1754c610_2);
and ( n21450 , n21449 , n52507 );
and ( n21451 , C0 , RI1754c610_2);
or ( n52508 , n21450 , n21451 );
buf ( n52509 , n52508 );
not ( n21452 , n27683 );
and ( n21453 , n21452 , RI19a89720_2728);
and ( n21454 , RI19a93950_2657 , n27683 );
or ( n52510 , n21453 , n21454 );
not ( n21455 , RI1754c610_2);
and ( n21456 , n21455 , n52510 );
and ( n21457 , C0 , RI1754c610_2);
or ( n52511 , n21456 , n21457 );
buf ( n52512 , n52511 );
not ( n52513 , n44051 );
xor ( n52514 , n28421 , n41799 );
xor ( n52515 , n52514 , n40381 );
and ( n52516 , n52513 , n52515 );
xor ( n52517 , n43877 , n52516 );
not ( n21458 , n29614 );
and ( n21459 , n21458 , RI174c67c8_793);
and ( n21460 , n52517 , n29614 );
or ( n52518 , n21459 , n21460 );
not ( n21461 , RI1754c610_2);
and ( n21462 , n21461 , n52518 );
and ( n21463 , C0 , RI1754c610_2);
or ( n52519 , n21462 , n21463 );
buf ( n52520 , n52519 );
not ( n52521 , n42735 );
and ( n52522 , n52521 , n42737 );
xor ( n52523 , n43683 , n52522 );
not ( n21464 , n29614 );
and ( n21465 , n21464 , RI174b75e8_842);
and ( n21466 , n52523 , n29614 );
or ( n52524 , n21465 , n21466 );
not ( n21467 , RI1754c610_2);
and ( n21468 , n21467 , n52524 );
and ( n21469 , C0 , RI1754c610_2);
or ( n52525 , n21468 , n21469 );
buf ( n52526 , n52525 );
not ( n21470 , n27683 );
and ( n21471 , n21470 , RI19a87920_2741);
and ( n21472 , RI19ac1d78_2315 , n27683 );
or ( n52527 , n21471 , n21472 );
not ( n21473 , RI1754c610_2);
and ( n21474 , n21473 , n52527 );
and ( n21475 , C0 , RI1754c610_2);
or ( n52528 , n21474 , n21475 );
buf ( n52529 , n52528 );
not ( n52530 , n45192 );
and ( n52531 , n52530 , n45194 );
xor ( n52532 , n49901 , n52531 );
not ( n21476 , n29614 );
and ( n21477 , n21476 , RI17492400_1023);
and ( n21478 , n52532 , n29614 );
or ( n52533 , n21477 , n21478 );
not ( n21479 , RI1754c610_2);
and ( n21480 , n21479 , n52533 );
and ( n21481 , C0 , RI1754c610_2);
or ( n52534 , n21480 , n21481 );
buf ( n52535 , n52534 );
not ( n52536 , n47682 );
and ( n52537 , n52536 , n46942 );
xor ( n52538 , n35459 , n52537 );
not ( n21482 , n29614 );
and ( n21483 , n21482 , RI17461da0_1259);
and ( n21484 , n52538 , n29614 );
or ( n52539 , n21483 , n21484 );
not ( n21485 , RI1754c610_2);
and ( n21486 , n21485 , n52539 );
and ( n21487 , C0 , RI1754c610_2);
or ( n52540 , n21486 , n21487 );
buf ( n52541 , n52540 );
and ( n52542 , RI1754ad38_55 , n34844 );
buf ( n52543 , n52542 );
not ( n21488 , n34859 );
and ( n21489 , n21488 , n52543 );
and ( n21490 , RI1754ad38_55 , n34859 );
or ( n52544 , n21489 , n21490 );
not ( n21491 , RI19a22f70_2797);
and ( n21492 , n21491 , n52544 );
and ( n21493 , C0 , RI19a22f70_2797);
or ( n52545 , n21492 , n21493 );
not ( n21494 , n27683 );
and ( n21495 , n21494 , RI19a23a38_2791);
and ( n21496 , n52545 , n27683 );
or ( n52546 , n21495 , n21496 );
not ( n21497 , RI1754c610_2);
and ( n21498 , n21497 , n52546 );
and ( n21499 , C0 , RI1754c610_2);
or ( n52547 , n21498 , n21499 );
buf ( n52548 , n52547 );
not ( n52549 , n45224 );
and ( n52550 , n52549 , n45226 );
xor ( n52551 , n46500 , n52550 );
not ( n21500 , n29614 );
and ( n21501 , n21500 , RI17520d80_664);
and ( n21502 , n52551 , n29614 );
or ( n52552 , n21501 , n21502 );
not ( n21503 , RI1754c610_2);
and ( n21504 , n21503 , n52552 );
and ( n21505 , C0 , RI1754c610_2);
or ( n52553 , n21504 , n21505 );
buf ( n52554 , n52553 );
not ( n52555 , n44394 );
and ( n52556 , n52555 , n45762 );
xor ( n52557 , n44391 , n52556 );
not ( n21506 , n29614 );
and ( n21507 , n21506 , RI174b0310_877);
and ( n21508 , n52557 , n29614 );
or ( n52558 , n21507 , n21508 );
not ( n21509 , RI1754c610_2);
and ( n21510 , n21509 , n52558 );
and ( n21511 , C0 , RI1754c610_2);
or ( n52559 , n21510 , n21511 );
buf ( n52560 , n52559 );
not ( n52561 , n44126 );
and ( n52562 , n52561 , n43633 );
xor ( n52563 , n46082 , n52562 );
not ( n21512 , n29614 );
and ( n21513 , n21512 , RI173be480_1828);
and ( n21514 , n52563 , n29614 );
or ( n52564 , n21513 , n21514 );
not ( n21515 , RI1754c610_2);
and ( n21516 , n21515 , n52564 );
and ( n21517 , C0 , RI1754c610_2);
or ( n52565 , n21516 , n21517 );
buf ( n52566 , n52565 );
xor ( n52567 , n31371 , n37074 );
xor ( n52568 , n52567 , n37104 );
not ( n52569 , n48950 );
and ( n52570 , n52569 , n48952 );
xor ( n52571 , n52568 , n52570 );
not ( n21518 , n29614 );
and ( n21519 , n21518 , RI17524638_653);
and ( n21520 , n52571 , n29614 );
or ( n52572 , n21519 , n21520 );
not ( n21521 , RI1754c610_2);
and ( n21522 , n21521 , n52572 );
and ( n21523 , C0 , RI1754c610_2);
or ( n52573 , n21522 , n21523 );
buf ( n52574 , n52573 );
not ( n52575 , n42149 );
and ( n52576 , n52575 , n49134 );
xor ( n52577 , n32864 , n52576 );
not ( n21524 , n29614 );
and ( n21525 , n21524 , RI17510bb0_714);
and ( n21526 , n52577 , n29614 );
or ( n52578 , n21525 , n21526 );
not ( n21527 , RI1754c610_2);
and ( n21528 , n21527 , n52578 );
and ( n21529 , C0 , RI1754c610_2);
or ( n52579 , n21528 , n21529 );
buf ( n52580 , n52579 );
xor ( n52581 , n28687 , n34497 );
xor ( n52582 , n52581 , n34517 );
not ( n52583 , n52582 );
and ( n52584 , n52583 , n48284 );
xor ( n52585 , n52227 , n52584 );
not ( n21530 , n29614 );
and ( n21531 , n21530 , RI174cde60_770);
and ( n21532 , n52585 , n29614 );
or ( n52586 , n21531 , n21532 );
not ( n21533 , RI1754c610_2);
and ( n21534 , n21533 , n52586 );
and ( n21535 , C0 , RI1754c610_2);
or ( n52587 , n21534 , n21535 );
buf ( n52588 , n52587 );
not ( n52589 , n45529 );
and ( n52590 , n52589 , n45531 );
xor ( n52591 , n50742 , n52590 );
not ( n21536 , n29614 );
and ( n21537 , n21536 , RI173f9250_1541);
and ( n21538 , n52591 , n29614 );
or ( n52592 , n21537 , n21538 );
not ( n21539 , RI1754c610_2);
and ( n21540 , n21539 , n52592 );
and ( n21541 , C0 , RI1754c610_2);
or ( n52593 , n21540 , n21541 );
buf ( n52594 , n52593 );
xor ( n52595 , n39625 , n35176 );
xor ( n52596 , n52595 , n35216 );
not ( n52597 , n52596 );
and ( n52598 , n52597 , n41400 );
xor ( n52599 , n46959 , n52598 );
not ( n21542 , n29614 );
and ( n21543 , n21542 , RI17463e70_1249);
and ( n21544 , n52599 , n29614 );
or ( n52600 , n21543 , n21544 );
not ( n21545 , RI1754c610_2);
and ( n21546 , n21545 , n52600 );
and ( n21547 , C0 , RI1754c610_2);
or ( n52601 , n21546 , n21547 );
buf ( n52602 , n52601 );
not ( n52603 , n46289 );
and ( n52604 , n52603 , n43597 );
xor ( n52605 , n41245 , n52604 );
not ( n21548 , n29614 );
and ( n21549 , n21548 , RI173c50c8_1795);
and ( n21550 , n52605 , n29614 );
or ( n52606 , n21549 , n21550 );
not ( n21551 , RI1754c610_2);
and ( n21552 , n21551 , n52606 );
and ( n21553 , C0 , RI1754c610_2);
or ( n52607 , n21552 , n21553 );
buf ( n52608 , n52607 );
not ( n52609 , n45039 );
and ( n52610 , n52609 , n45041 );
xor ( n52611 , n46061 , n52610 );
not ( n21554 , n29614 );
and ( n21555 , n21554 , RI17495f10_1005);
and ( n21556 , n52611 , n29614 );
or ( n52612 , n21555 , n21556 );
not ( n21557 , RI1754c610_2);
and ( n21558 , n21557 , n52612 );
and ( n21559 , C0 , RI1754c610_2);
or ( n52613 , n21558 , n21559 );
buf ( n52614 , n52613 );
buf ( n52615 , RI174caad0_780);
not ( n52616 , n46320 );
and ( n52617 , n52616 , n50080 );
xor ( n52618 , n45733 , n52617 );
not ( n21560 , n29614 );
and ( n21561 , n21560 , RI173a22f8_1965);
and ( n21562 , n52618 , n29614 );
or ( n52619 , n21561 , n21562 );
not ( n21563 , RI1754c610_2);
and ( n21564 , n21563 , n52619 );
and ( n21565 , C0 , RI1754c610_2);
or ( n52620 , n21564 , n21565 );
buf ( n52621 , n52620 );
not ( n52622 , n40343 );
and ( n52623 , n52622 , n40361 );
xor ( n52624 , n40980 , n52623 );
not ( n21566 , n29614 );
and ( n21567 , n21566 , RI17514990_702);
and ( n21568 , n52624 , n29614 );
or ( n52625 , n21567 , n21568 );
not ( n21569 , RI1754c610_2);
and ( n21570 , n21569 , n52625 );
and ( n21571 , C0 , RI1754c610_2);
or ( n52626 , n21570 , n21571 );
buf ( n52627 , n52626 );
buf ( n52628 , RI175038c0_749);
buf ( n52629 , RI1748c4d8_1052);
not ( n52630 , n50251 );
and ( n52631 , n52630 , n43839 );
xor ( n52632 , n41288 , n52631 );
not ( n21572 , n29614 );
and ( n21573 , n21572 , RI1750ecc0_720);
and ( n21574 , n52632 , n29614 );
or ( n52633 , n21573 , n21574 );
not ( n21575 , RI1754c610_2);
and ( n21576 , n21575 , n52633 );
and ( n21577 , C0 , RI1754c610_2);
or ( n52634 , n21576 , n21577 );
buf ( n52635 , n52634 );
buf ( n52636 , RI1748f2c8_1038);
not ( n52637 , n39184 );
and ( n52638 , n52637 , n34341 );
xor ( n52639 , n39162 , n52638 );
not ( n21578 , n29614 );
and ( n21579 , n21578 , RI174b68c8_846);
and ( n21580 , n52639 , n29614 );
or ( n52640 , n21579 , n21580 );
not ( n21581 , RI1754c610_2);
and ( n21582 , n21581 , n52640 );
and ( n21583 , C0 , RI1754c610_2);
or ( n52641 , n21582 , n21583 );
buf ( n52642 , n52641 );
not ( n52643 , n51420 );
and ( n52644 , n52643 , n51422 );
xor ( n52645 , n48380 , n52644 );
not ( n21584 , n29614 );
and ( n21585 , n21584 , RI174b2db8_864);
and ( n21586 , n52645 , n29614 );
or ( n52646 , n21585 , n21586 );
not ( n21587 , RI1754c610_2);
and ( n21588 , n21587 , n52646 );
and ( n21589 , C0 , RI1754c610_2);
or ( n52647 , n21588 , n21589 );
buf ( n52648 , n52647 );
not ( n52649 , n45557 );
and ( n52650 , n52649 , n50756 );
xor ( n52651 , n44229 , n52650 );
not ( n21590 , n29614 );
and ( n21591 , n21590 , RI1748a408_1062);
and ( n21592 , n52651 , n29614 );
or ( n52652 , n21591 , n21592 );
not ( n21593 , RI1754c610_2);
and ( n21594 , n21593 , n52652 );
and ( n21595 , C0 , RI1754c610_2);
or ( n52653 , n21594 , n21595 );
buf ( n52654 , n52653 );
not ( n21596 , n27683 );
and ( n21597 , n21596 , RI19aaa510_2493);
and ( n21598 , RI19ab4560_2421 , n27683 );
or ( n52655 , n21597 , n21598 );
not ( n21599 , RI1754c610_2);
and ( n21600 , n21599 , n52655 );
and ( n21601 , C0 , RI1754c610_2);
or ( n52656 , n21600 , n21601 );
buf ( n52657 , n52656 );
not ( n52658 , n42525 );
and ( n52659 , n52658 , n46645 );
xor ( n52660 , n42522 , n52659 );
not ( n21602 , n29614 );
and ( n21603 , n21602 , RI174001e0_1507);
and ( n21604 , n52660 , n29614 );
or ( n52661 , n21603 , n21604 );
not ( n21605 , RI1754c610_2);
and ( n21606 , n21605 , n52661 );
and ( n21607 , C0 , RI1754c610_2);
or ( n52662 , n21606 , n21607 );
buf ( n52663 , n52662 );
not ( n52664 , n44316 );
and ( n52665 , n52664 , n51812 );
xor ( n52666 , n36004 , n52665 );
not ( n21608 , n29614 );
and ( n21609 , n21608 , RI173b4d90_1874);
and ( n21610 , n52666 , n29614 );
or ( n52667 , n21609 , n21610 );
not ( n21611 , RI1754c610_2);
and ( n21612 , n21611 , n52667 );
and ( n21613 , C0 , RI1754c610_2);
or ( n52668 , n21612 , n21613 );
buf ( n52669 , n52668 );
not ( n52670 , n51591 );
and ( n52671 , n52670 , n42820 );
xor ( n52672 , n44501 , n52671 );
not ( n21614 , n29614 );
and ( n21615 , n21614 , RI1748ef80_1039);
and ( n21616 , n52672 , n29614 );
or ( n52673 , n21615 , n21616 );
not ( n21617 , RI1754c610_2);
and ( n21618 , n21617 , n52673 );
and ( n21619 , C0 , RI1754c610_2);
or ( n52674 , n21618 , n21619 );
buf ( n52675 , n52674 );
not ( n21620 , n27683 );
and ( n21621 , n21620 , RI19aadfa8_2468);
and ( n21622 , RI19ab7a58_2397 , n27683 );
or ( n52676 , n21621 , n21622 );
not ( n21623 , RI1754c610_2);
and ( n21624 , n21623 , n52676 );
and ( n21625 , C0 , RI1754c610_2);
or ( n52677 , n21624 , n21625 );
buf ( n52678 , n52677 );
not ( n52679 , n44247 );
and ( n52680 , n52679 , n37256 );
xor ( n52681 , n44244 , n52680 );
not ( n21626 , n29614 );
and ( n21627 , n21626 , RI173d6b10_1709);
and ( n21628 , n52681 , n29614 );
or ( n52682 , n21627 , n21628 );
not ( n21629 , RI1754c610_2);
and ( n21630 , n21629 , n52682 );
and ( n21631 , C0 , RI1754c610_2);
or ( n52683 , n21630 , n21631 );
buf ( n52684 , n52683 );
not ( n52685 , n49340 );
and ( n52686 , n52685 , n46877 );
xor ( n52687 , n44988 , n52686 );
not ( n21632 , n29614 );
and ( n21633 , n21632 , RI1746f978_1192);
and ( n21634 , n52687 , n29614 );
or ( n52688 , n21633 , n21634 );
not ( n21635 , RI1754c610_2);
and ( n21636 , n21635 , n52688 );
and ( n21637 , C0 , RI1754c610_2);
or ( n52689 , n21636 , n21637 );
buf ( n52690 , n52689 );
not ( n21638 , n27683 );
and ( n21639 , n21638 , RI19aceac8_2220);
and ( n21640 , RI19a9b420_2603 , n27683 );
or ( n52691 , n21639 , n21640 );
not ( n21641 , RI1754c610_2);
and ( n21642 , n21641 , n52691 );
and ( n21643 , C0 , RI1754c610_2);
or ( n52692 , n21642 , n21643 );
buf ( n52693 , n52692 );
not ( n21644 , n27683 );
and ( n21645 , n21644 , RI19aabcf8_2483);
and ( n21646 , RI19ab5a00_2411 , n27683 );
or ( n52694 , n21645 , n21646 );
not ( n21647 , RI1754c610_2);
and ( n21648 , n21647 , n52694 );
and ( n21649 , C0 , RI1754c610_2);
or ( n52695 , n21648 , n21649 );
buf ( n52696 , n52695 );
not ( n21650 , n27683 );
and ( n21651 , n21650 , RI19aa0100_2568);
and ( n21652 , RI19aa9d90_2497 , n27683 );
or ( n52697 , n21651 , n21652 );
not ( n21653 , RI1754c610_2);
and ( n21654 , n21653 , n52697 );
and ( n21655 , C0 , RI1754c610_2);
or ( n52698 , n21654 , n21655 );
buf ( n52699 , n52698 );
not ( n21656 , n27683 );
and ( n21657 , n21656 , RI19a8d410_2702);
and ( n21658 , RI19a97460_2631 , n27683 );
or ( n52700 , n21657 , n21658 );
not ( n21659 , RI1754c610_2);
and ( n21660 , n21659 , n52700 );
and ( n21661 , C0 , RI1754c610_2);
or ( n52701 , n21660 , n21661 );
buf ( n52702 , n52701 );
buf ( n52703 , RI174cc9c0_774);
not ( n52704 , n51143 );
and ( n52705 , n52704 , n48254 );
xor ( n52706 , n43200 , n52705 );
not ( n21662 , n29614 );
and ( n21663 , n21662 , RI173b39e0_1880);
and ( n21664 , n52706 , n29614 );
or ( n52707 , n21663 , n21664 );
not ( n21665 , RI1754c610_2);
and ( n21666 , n21665 , n52707 );
and ( n21667 , C0 , RI1754c610_2);
or ( n52708 , n21666 , n21667 );
buf ( n52709 , n52708 );
buf ( n52710 , RI174b8f38_835);
buf ( n52711 , RI1749a3f8_984);
buf ( n52712 , RI1748dbd0_1045);
not ( n52713 , n40170 );
and ( n52714 , n52713 , n45463 );
xor ( n52715 , n40167 , n52714 );
not ( n21668 , n29614 );
and ( n21669 , n21668 , RI17476908_1158);
and ( n21670 , n52715 , n29614 );
or ( n52716 , n21669 , n21670 );
not ( n21671 , RI1754c610_2);
and ( n21672 , n21671 , n52716 );
and ( n21673 , C0 , RI1754c610_2);
or ( n52717 , n21672 , n21673 );
buf ( n52718 , n52717 );
not ( n21674 , n27683 );
and ( n21675 , n21674 , RI19a84950_2762);
and ( n21676 , RI19ac0a40_2326 , n27683 );
or ( n52719 , n21675 , n21676 );
not ( n21677 , RI1754c610_2);
and ( n21678 , n21677 , n52719 );
and ( n21679 , C0 , RI1754c610_2);
or ( n52720 , n21678 , n21679 );
buf ( n52721 , n52720 );
buf ( n52722 , RI174c6cf0_792);
not ( n52723 , n44058 );
and ( n52724 , n52723 , n38349 );
xor ( n52725 , n44722 , n52724 );
not ( n21680 , n29614 );
and ( n21681 , n21680 , RI17521cf8_661);
and ( n21682 , n52725 , n29614 );
or ( n52726 , n21681 , n21682 );
not ( n21683 , RI1754c610_2);
and ( n21684 , n21683 , n52726 );
and ( n21685 , C0 , RI1754c610_2);
or ( n52727 , n21684 , n21685 );
buf ( n52728 , n52727 );
not ( n52729 , n50190 );
and ( n52730 , n52729 , n47528 );
xor ( n52731 , n50187 , n52730 );
not ( n21686 , n29614 );
and ( n21687 , n21686 , RI174081d8_1468);
and ( n21688 , n52731 , n29614 );
or ( n52732 , n21687 , n21688 );
not ( n21689 , RI1754c610_2);
and ( n21690 , n21689 , n52732 );
and ( n21691 , C0 , RI1754c610_2);
or ( n52733 , n21690 , n21691 );
buf ( n52734 , n52733 );
buf ( n52735 , RI17491a28_1026);
not ( n21692 , n27683 );
and ( n21693 , n21692 , RI19a98d38_2620);
and ( n21694 , RI19aa24a0_2550 , n27683 );
or ( n52736 , n21693 , n21694 );
not ( n21695 , RI1754c610_2);
and ( n21696 , n21695 , n52736 );
and ( n21697 , C0 , RI1754c610_2);
or ( n52737 , n21696 , n21697 );
buf ( n52738 , n52737 );
buf ( n52739 , RI174b3790_861);
not ( n52740 , n40664 );
and ( n52741 , n52740 , n40666 );
xor ( n52742 , n37916 , n52741 );
not ( n21698 , n29614 );
and ( n21699 , n21698 , RI1740d3e0_1443);
and ( n21700 , n52742 , n29614 );
or ( n52743 , n21699 , n21700 );
not ( n21701 , RI1754c610_2);
and ( n21702 , n21701 , n52743 );
and ( n21703 , C0 , RI1754c610_2);
or ( n52744 , n21702 , n21703 );
buf ( n52745 , n52744 );
buf ( n52746 , RI174bec08_817);
not ( n52747 , n41712 );
and ( n52748 , n52747 , n41714 );
xor ( n52749 , n45387 , n52748 );
not ( n21704 , n29614 );
and ( n21705 , n21704 , RI17391c78_2045);
and ( n21706 , n52749 , n29614 );
or ( n52750 , n21705 , n21706 );
not ( n21707 , RI1754c610_2);
and ( n21708 , n21707 , n52750 );
and ( n21709 , C0 , RI1754c610_2);
or ( n52751 , n21708 , n21709 );
buf ( n52752 , n52751 );
not ( n52753 , n38595 );
xor ( n52754 , n31995 , n36682 );
xor ( n52755 , n52754 , n36702 );
and ( n52756 , n52753 , n52755 );
xor ( n52757 , n38554 , n52756 );
not ( n21710 , n29614 );
and ( n21711 , n21710 , RI173c6e50_1786);
and ( n21712 , n52757 , n29614 );
or ( n52758 , n21711 , n21712 );
not ( n21713 , RI1754c610_2);
and ( n21714 , n21713 , n52758 );
and ( n21715 , C0 , RI1754c610_2);
or ( n52759 , n21714 , n21715 );
buf ( n52760 , n52759 );
buf ( n52761 , RI1750be58_729);
buf ( n52762 , RI17468010_1229);
buf ( n52763 , RI1747bb10_1133);
buf ( n52764 , RI17484828_1090);
buf ( n52765 , RI17496c30_1001);
buf ( n52766 , RI1749f948_958);
xor ( n52767 , n41417 , n43464 );
xor ( n52768 , n52767 , n44146 );
not ( n52769 , n51561 );
and ( n52770 , n52769 , n42480 );
xor ( n52771 , n52768 , n52770 );
not ( n21716 , n29614 );
and ( n21717 , n21716 , RI173d5760_1715);
and ( n21718 , n52771 , n29614 );
or ( n52772 , n21717 , n21718 );
not ( n21719 , RI1754c610_2);
and ( n21720 , n21719 , n52772 );
and ( n21721 , C0 , RI1754c610_2);
or ( n52773 , n21720 , n21721 );
buf ( n52774 , n52773 );
not ( n21722 , n27683 );
and ( n21723 , n21722 , RI19ab65b8_2406);
and ( n21724 , RI19abfa50_2335 , n27683 );
or ( n52775 , n21723 , n21724 );
not ( n21725 , RI1754c610_2);
and ( n21726 , n21725 , n52775 );
and ( n21727 , C0 , RI1754c610_2);
or ( n52776 , n21726 , n21727 );
buf ( n52777 , n52776 );
not ( n52778 , n46059 );
and ( n52779 , n52778 , n46061 );
xor ( n52780 , n45044 , n52779 );
not ( n21728 , n29614 );
and ( n21729 , n21728 , RI17478d20_1147);
and ( n21730 , n52780 , n29614 );
or ( n52781 , n21729 , n21730 );
not ( n21731 , RI1754c610_2);
and ( n21732 , n21731 , n52781 );
and ( n21733 , C0 , RI1754c610_2);
or ( n52782 , n21732 , n21733 );
buf ( n52783 , n52782 );
not ( n21734 , n27683 );
and ( n21735 , n21734 , RI19abbe50_2368);
and ( n21736 , RI19ac4460_2297 , n27683 );
or ( n52784 , n21735 , n21736 );
not ( n21737 , RI1754c610_2);
and ( n21738 , n21737 , n52784 );
and ( n21739 , C0 , RI1754c610_2);
or ( n52785 , n21738 , n21739 );
buf ( n52786 , n52785 );
not ( n52787 , n37256 );
and ( n52788 , n52787 , n37261 );
xor ( n52789 , n44247 , n52788 );
not ( n21740 , n29614 );
and ( n21741 , n21740 , RI173e5750_1637);
and ( n21742 , n52789 , n29614 );
or ( n52790 , n21741 , n21742 );
not ( n21743 , RI1754c610_2);
and ( n21744 , n21743 , n52790 );
and ( n21745 , C0 , RI1754c610_2);
or ( n52791 , n21744 , n21745 );
buf ( n52792 , n52791 );
not ( n52793 , n39953 );
and ( n52794 , n52793 , n40829 );
xor ( n52795 , n39915 , n52794 );
not ( n21746 , n29614 );
and ( n21747 , n21746 , RI173a50e8_1951);
and ( n21748 , n52795 , n29614 );
or ( n52796 , n21747 , n21748 );
not ( n21749 , RI1754c610_2);
and ( n21750 , n21749 , n52796 );
and ( n21751 , C0 , RI1754c610_2);
or ( n52797 , n21750 , n21751 );
buf ( n52798 , n52797 );
not ( n52799 , n47226 );
and ( n52800 , n52799 , n52209 );
xor ( n52801 , n45312 , n52800 );
not ( n21752 , n29614 );
and ( n21753 , n21752 , RI174caad0_780);
and ( n21754 , n52801 , n29614 );
or ( n52802 , n21753 , n21754 );
not ( n21755 , RI1754c610_2);
and ( n21756 , n21755 , n52802 );
and ( n21757 , C0 , RI1754c610_2);
or ( n52803 , n21756 , n21757 );
buf ( n52804 , n52803 );
not ( n52805 , n47355 );
xor ( n52806 , n39905 , n33397 );
xor ( n52807 , n52806 , n35710 );
and ( n52808 , n52805 , n52807 );
xor ( n52809 , n44915 , n52808 );
not ( n21758 , n29614 );
and ( n21759 , n21758 , RI17445588_1398);
and ( n21760 , n52809 , n29614 );
or ( n52810 , n21759 , n21760 );
not ( n21761 , RI1754c610_2);
and ( n21762 , n21761 , n52810 );
and ( n21763 , C0 , RI1754c610_2);
or ( n52811 , n21762 , n21763 );
buf ( n52812 , n52811 );
not ( n21764 , n27683 );
and ( n21765 , n21764 , RI19ac2840_2310);
and ( n21766 , RI19acb828_2243 , n27683 );
or ( n52813 , n21765 , n21766 );
not ( n21767 , RI1754c610_2);
and ( n21768 , n21767 , n52813 );
and ( n21769 , C0 , RI1754c610_2);
or ( n52814 , n21768 , n21769 );
buf ( n52815 , n52814 );
buf ( n52816 , RI1750d820_724);
buf ( n52817 , RI17486f88_1078);
not ( n52818 , n46000 );
and ( n52819 , n52818 , n46403 );
xor ( n52820 , n45997 , n52819 );
not ( n21770 , n29614 );
and ( n21771 , n21770 , RI17452788_1334);
and ( n21772 , n52820 , n29614 );
or ( n52821 , n21771 , n21772 );
not ( n21773 , RI1754c610_2);
and ( n21774 , n21773 , n52821 );
and ( n21775 , C0 , RI1754c610_2);
or ( n52822 , n21774 , n21775 );
buf ( n52823 , n52822 );
not ( n52824 , n49708 );
and ( n52825 , n52824 , n41029 );
xor ( n52826 , n49705 , n52825 );
not ( n21776 , n29614 );
and ( n21777 , n21776 , RI174865b0_1081);
and ( n21778 , n52826 , n29614 );
or ( n52827 , n21777 , n21778 );
not ( n21779 , RI1754c610_2);
and ( n21780 , n21779 , n52827 );
and ( n21781 , C0 , RI1754c610_2);
or ( n52828 , n21780 , n21781 );
buf ( n52829 , n52828 );
not ( n21782 , n27683 );
and ( n21783 , n21782 , RI19a9f908_2572);
and ( n21784 , RI19aa9688_2500 , n27683 );
or ( n52830 , n21783 , n21784 );
not ( n21785 , RI1754c610_2);
and ( n21786 , n21785 , n52830 );
and ( n21787 , C0 , RI1754c610_2);
or ( n52831 , n21786 , n21787 );
buf ( n52832 , n52831 );
not ( n21788 , n27683 );
and ( n21789 , n21788 , RI19a920f0_2668);
and ( n21790 , RI19a9c1b8_2597 , n27683 );
or ( n52833 , n21789 , n21790 );
not ( n21791 , RI1754c610_2);
and ( n21792 , n21791 , n52833 );
and ( n21793 , C0 , RI1754c610_2);
or ( n52834 , n21792 , n21793 );
buf ( n52835 , n52834 );
not ( n21794 , RI1754c610_2);
and ( n21795 , n21794 , RI19ad12b8_2203);
and ( n21796 , C0 , RI1754c610_2);
or ( n52836 , n21795 , n21796 );
buf ( n52837 , n52836 );
not ( n52838 , n47430 );
and ( n52839 , n52838 , n47432 );
xor ( n52840 , n48549 , n52839 );
not ( n21797 , n29614 );
and ( n21798 , n21797 , RI173b6488_1867);
and ( n21799 , n52840 , n29614 );
or ( n52841 , n21798 , n21799 );
not ( n21800 , RI1754c610_2);
and ( n21801 , n21800 , n52841 );
and ( n21802 , C0 , RI1754c610_2);
or ( n52842 , n21801 , n21802 );
buf ( n52843 , n52842 );
not ( n52844 , n46257 );
and ( n52845 , n52844 , n46181 );
xor ( n52846 , n46254 , n52845 );
not ( n21803 , n29614 );
and ( n21804 , n21803 , RI17498670_993);
and ( n21805 , n52846 , n29614 );
or ( n52847 , n21804 , n21805 );
not ( n21806 , RI1754c610_2);
and ( n21807 , n21806 , n52847 );
and ( n21808 , C0 , RI1754c610_2);
or ( n52848 , n21807 , n21808 );
buf ( n52849 , n52848 );
not ( n52850 , n45934 );
and ( n52851 , n52850 , n41639 );
xor ( n52852 , n46870 , n52851 );
not ( n21809 , n29614 );
and ( n21810 , n21809 , RI173d6138_1712);
and ( n21811 , n52852 , n29614 );
or ( n52853 , n21810 , n21811 );
not ( n21812 , RI1754c610_2);
and ( n21813 , n21812 , n52853 );
and ( n21814 , C0 , RI1754c610_2);
or ( n52854 , n21813 , n21814 );
buf ( n52855 , n52854 );
not ( n21815 , n27683 );
and ( n21816 , n21815 , RI19ab7da0_2396);
and ( n21817 , RI19ac0ba8_2325 , n27683 );
or ( n52856 , n21816 , n21817 );
not ( n21818 , RI1754c610_2);
and ( n21819 , n21818 , n52856 );
and ( n21820 , C0 , RI1754c610_2);
or ( n52857 , n21819 , n21820 );
buf ( n52858 , n52857 );
not ( n52859 , n42873 );
and ( n52860 , n52859 , n42875 );
xor ( n52861 , n51357 , n52860 );
not ( n21821 , n29614 );
and ( n21822 , n21821 , RI173cd750_1754);
and ( n21823 , n52861 , n29614 );
or ( n52862 , n21822 , n21823 );
not ( n21824 , RI1754c610_2);
and ( n21825 , n21824 , n52862 );
and ( n21826 , C0 , RI1754c610_2);
or ( n52863 , n21825 , n21826 );
buf ( n52864 , n52863 );
not ( n52865 , n47036 );
and ( n52866 , n52865 , n50171 );
xor ( n52867 , n47033 , n52866 );
not ( n21827 , n29614 );
and ( n21828 , n21827 , RI173cb9c8_1763);
and ( n21829 , n52867 , n29614 );
or ( n52868 , n21828 , n21829 );
not ( n21830 , RI1754c610_2);
and ( n21831 , n21830 , n52868 );
and ( n21832 , C0 , RI1754c610_2);
or ( n52869 , n21831 , n21832 );
buf ( n52870 , n52869 );
not ( n52871 , n37170 );
and ( n52872 , n52871 , n37204 );
xor ( n52873 , n47595 , n52872 );
not ( n21833 , n29614 );
and ( n21834 , n21833 , RI173f5a88_1558);
and ( n21835 , n52873 , n29614 );
or ( n52874 , n21834 , n21835 );
not ( n21836 , RI1754c610_2);
and ( n21837 , n21836 , n52874 );
and ( n21838 , C0 , RI1754c610_2);
or ( n52875 , n21837 , n21838 );
buf ( n52876 , n52875 );
not ( n52877 , n48173 );
xor ( n52878 , n37905 , n32048 );
xor ( n52879 , n52878 , n32108 );
and ( n52880 , n52877 , n52879 );
xor ( n52881 , n48170 , n52880 );
not ( n21839 , n29614 );
and ( n21840 , n21839 , RI17335248_2182);
and ( n21841 , n52881 , n29614 );
or ( n52882 , n21840 , n21841 );
not ( n21842 , RI1754c610_2);
and ( n21843 , n21842 , n52882 );
and ( n21844 , C0 , RI1754c610_2);
or ( n52883 , n21843 , n21844 );
buf ( n52884 , n52883 );
not ( n52885 , n44779 );
and ( n52886 , n52885 , n44781 );
xor ( n52887 , n49273 , n52886 );
not ( n21845 , n29614 );
and ( n21846 , n21845 , RI175019d0_755);
and ( n21847 , n52887 , n29614 );
or ( n52888 , n21846 , n21847 );
not ( n21848 , RI1754c610_2);
and ( n21849 , n21848 , n52888 );
and ( n21850 , C0 , RI1754c610_2);
or ( n52889 , n21849 , n21850 );
buf ( n52890 , n52889 );
xor ( n52891 , n37412 , n38267 );
xor ( n52892 , n52891 , n38284 );
not ( n52893 , n46627 );
and ( n52894 , n52893 , n46629 );
xor ( n52895 , n52892 , n52894 );
not ( n21851 , n29614 );
and ( n21852 , n21851 , RI173971c8_2019);
and ( n21853 , n52895 , n29614 );
or ( n52896 , n21852 , n21853 );
not ( n21854 , RI1754c610_2);
and ( n21855 , n21854 , n52896 );
and ( n21856 , C0 , RI1754c610_2);
or ( n52897 , n21855 , n21856 );
buf ( n52898 , n52897 );
not ( n52899 , n46365 );
and ( n52900 , n52899 , n43421 );
xor ( n52901 , n44714 , n52900 );
not ( n21857 , n29614 );
and ( n21858 , n21857 , RI174d07a0_762);
and ( n21859 , n52901 , n29614 );
or ( n52902 , n21858 , n21859 );
not ( n21860 , RI1754c610_2);
and ( n21861 , n21860 , n52902 );
and ( n21862 , C0 , RI1754c610_2);
or ( n52903 , n21861 , n21862 );
buf ( n52904 , n52903 );
not ( n21863 , n27683 );
and ( n21864 , n21863 , RI19acabf8_2250);
and ( n21865 , RI19a860c0_2752 , n27683 );
or ( n52905 , n21864 , n21865 );
not ( n21866 , RI1754c610_2);
and ( n21867 , n21866 , n52905 );
and ( n21868 , C0 , RI1754c610_2);
or ( n52906 , n21867 , n21868 );
buf ( n52907 , n52906 );
not ( n21869 , n27683 );
and ( n21870 , n21869 , RI19ab4560_2421);
and ( n21871 , RI19abddb8_2351 , n27683 );
or ( n52908 , n21870 , n21871 );
not ( n21872 , RI1754c610_2);
and ( n21873 , n21872 , n52908 );
and ( n21874 , C0 , RI1754c610_2);
or ( n52909 , n21873 , n21874 );
buf ( n52910 , n52909 );
buf ( n52911 , RI17511600_712);
buf ( n52912 , RI17481060_1107);
not ( n21875 , n27683 );
and ( n21876 , n21875 , RI19aa3058_2545);
and ( n21877 , RI19aad300_2474 , n27683 );
or ( n52913 , n21876 , n21877 );
not ( n21878 , RI1754c610_2);
and ( n21879 , n21878 , n52913 );
and ( n21880 , C0 , RI1754c610_2);
or ( n52914 , n21879 , n21880 );
buf ( n52915 , n52914 );
not ( n52916 , n33506 );
and ( n52917 , n52916 , n41007 );
xor ( n52918 , n33398 , n52917 );
not ( n21881 , n29614 );
and ( n21882 , n21881 , RI173feae8_1514);
and ( n21883 , n52918 , n29614 );
or ( n52919 , n21882 , n21883 );
not ( n21884 , RI1754c610_2);
and ( n21885 , n21884 , n52919 );
and ( n21886 , C0 , RI1754c610_2);
or ( n52920 , n21885 , n21886 );
buf ( n52921 , n52920 );
not ( n52922 , n36655 );
and ( n52923 , n52922 , n46764 );
xor ( n52924 , n36613 , n52923 );
not ( n21887 , n29614 );
and ( n21888 , n21887 , RI173e0890_1661);
and ( n21889 , n52924 , n29614 );
or ( n52925 , n21888 , n21889 );
not ( n21890 , RI1754c610_2);
and ( n21891 , n21890 , n52925 );
and ( n21892 , C0 , RI1754c610_2);
or ( n52926 , n21891 , n21892 );
buf ( n52927 , n52926 );
not ( n21893 , n27683 );
and ( n21894 , n21893 , RI19aa9688_2500);
and ( n21895 , RI19ab3318_2430 , n27683 );
or ( n52928 , n21894 , n21895 );
not ( n21896 , RI1754c610_2);
and ( n21897 , n21896 , n52928 );
and ( n21898 , C0 , RI1754c610_2);
or ( n52929 , n21897 , n21898 );
buf ( n52930 , n52929 );
not ( n21899 , n27683 );
and ( n21900 , n21899 , RI19aa1618_2557);
and ( n21901 , RI19aab5f0_2486 , n27683 );
or ( n52931 , n21900 , n21901 );
not ( n21902 , RI1754c610_2);
and ( n21903 , n21902 , n52931 );
and ( n21904 , C0 , RI1754c610_2);
or ( n52932 , n21903 , n21904 );
buf ( n52933 , n52932 );
xor ( n52934 , n40705 , n39333 );
xor ( n52935 , n52934 , n39347 );
not ( n52936 , n52935 );
and ( n52937 , n52936 , n50123 );
xor ( n52938 , n50259 , n52937 );
not ( n21905 , n29614 );
and ( n21906 , n21905 , RI1749f2b8_960);
and ( n21907 , n52938 , n29614 );
or ( n52939 , n21906 , n21907 );
not ( n21908 , RI1754c610_2);
and ( n21909 , n21908 , n52939 );
and ( n21910 , C0 , RI1754c610_2);
or ( n52940 , n21909 , n21910 );
buf ( n52941 , n52940 );
not ( n52942 , n51927 );
and ( n52943 , n52942 , n39720 );
xor ( n52944 , n52134 , n52943 );
not ( n21911 , n29614 );
and ( n21912 , n21911 , RI173ca2d0_1770);
and ( n21913 , n52944 , n29614 );
or ( n52945 , n21912 , n21913 );
not ( n21914 , RI1754c610_2);
and ( n21915 , n21914 , n52945 );
and ( n21916 , C0 , RI1754c610_2);
or ( n52946 , n21915 , n21916 );
buf ( n52947 , n52946 );
not ( n52948 , n46966 );
and ( n52949 , n52948 , n46968 );
xor ( n52950 , n50404 , n52949 );
not ( n21917 , n29614 );
and ( n21918 , n21917 , RI173b2cc0_1884);
and ( n21919 , n52950 , n29614 );
or ( n52951 , n21918 , n21919 );
not ( n21920 , RI1754c610_2);
and ( n21921 , n21920 , n52951 );
and ( n21922 , C0 , RI1754c610_2);
or ( n52952 , n21921 , n21922 );
buf ( n52953 , n52952 );
not ( n52954 , n48029 );
and ( n52955 , n52954 , n51199 );
xor ( n52956 , n48026 , n52955 );
not ( n21923 , n29614 );
and ( n21924 , n21923 , RI17394720_2032);
and ( n21925 , n52956 , n29614 );
or ( n52957 , n21924 , n21925 );
not ( n21926 , RI1754c610_2);
and ( n21927 , n21926 , n52957 );
and ( n21928 , C0 , RI1754c610_2);
or ( n52958 , n21927 , n21928 );
buf ( n52959 , n52958 );
buf ( n52960 , RI1747d898_1124);
not ( n52961 , n47194 );
and ( n52962 , n52961 , n47031 );
xor ( n52963 , n50171 , n52962 );
not ( n21929 , n29614 );
and ( n21930 , n21929 , RI173e8bd0_1621);
and ( n21931 , n52963 , n29614 );
or ( n52964 , n21930 , n21931 );
not ( n21932 , RI1754c610_2);
and ( n21933 , n21932 , n52964 );
and ( n21934 , C0 , RI1754c610_2);
or ( n52965 , n21933 , n21934 );
buf ( n52966 , n52965 );
not ( n52967 , n49447 );
and ( n52968 , n52967 , n52568 );
xor ( n52969 , n48955 , n52968 );
not ( n21935 , n29614 );
and ( n21936 , n21935 , RI17450370_1345);
and ( n21937 , n52969 , n29614 );
or ( n52970 , n21936 , n21937 );
not ( n21938 , RI1754c610_2);
and ( n21939 , n21938 , n52970 );
and ( n21940 , C0 , RI1754c610_2);
or ( n52971 , n21939 , n21940 );
buf ( n52972 , n52971 );
not ( n52973 , n32482 );
and ( n52974 , n52973 , n49637 );
xor ( n52975 , n32310 , n52974 );
not ( n21941 , n29614 );
and ( n21942 , n21941 , RI173c1270_1814);
and ( n21943 , n52975 , n29614 );
or ( n52976 , n21942 , n21943 );
not ( n21944 , RI1754c610_2);
and ( n21945 , n21944 , n52976 );
and ( n21946 , C0 , RI1754c610_2);
or ( n52977 , n21945 , n21946 );
buf ( n52978 , n52977 );
not ( n21947 , RI1754c610_2);
and ( n21948 , n21947 , RI175385e8_592);
and ( n21949 , C0 , RI1754c610_2);
or ( n52979 , n21948 , n21949 );
buf ( n52980 , n52979 );
not ( n52981 , n48467 );
and ( n52982 , n52981 , n46826 );
xor ( n52983 , n48056 , n52982 );
not ( n21950 , n29614 );
and ( n21951 , n21950 , RI174074b8_1472);
and ( n21952 , n52983 , n29614 );
or ( n52984 , n21951 , n21952 );
not ( n21953 , RI1754c610_2);
and ( n21954 , n21953 , n52984 );
and ( n21955 , C0 , RI1754c610_2);
or ( n52985 , n21954 , n21955 );
buf ( n52986 , n52985 );
not ( n52987 , n52186 );
xor ( n52988 , n37103 , n37716 );
xor ( n52989 , n52988 , n37744 );
and ( n52990 , n52987 , n52989 );
xor ( n52991 , n52183 , n52990 );
not ( n21956 , n29614 );
and ( n21957 , n21956 , RI174a7940_919);
and ( n21958 , n52991 , n29614 );
or ( n52992 , n21957 , n21958 );
not ( n21959 , RI1754c610_2);
and ( n21960 , n21959 , n52992 );
and ( n21961 , C0 , RI1754c610_2);
or ( n52993 , n21960 , n21961 );
buf ( n52994 , n52993 );
and ( n52995 , RI1754be90_18 , n34844 );
and ( n52996 , RI1754be90_18 , n34847 );
and ( n52997 , RI1754be90_18 , n34850 );
and ( n52998 , RI1754be90_18 , n34852 );
and ( n52999 , RI1754be90_18 , n34854 );
and ( n53000 , RI1754be90_18 , n34856 );
buf ( n53001 , n39233 );
or ( n53002 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , C0 );
not ( n21962 , n34859 );
and ( n21963 , n21962 , n53002 );
and ( n21964 , RI1754be90_18 , n34859 );
or ( n53003 , n21963 , n21964 );
not ( n21965 , RI19a22f70_2797);
and ( n21966 , n21965 , n53003 );
and ( n21967 , C0 , RI19a22f70_2797);
or ( n53004 , n21966 , n21967 );
not ( n21968 , n27683 );
and ( n21969 , n21968 , RI19a96998_2636);
and ( n21970 , n53004 , n27683 );
or ( n53005 , n21969 , n21970 );
not ( n21971 , RI1754c610_2);
and ( n21972 , n21971 , n53005 );
and ( n21973 , C0 , RI1754c610_2);
or ( n53006 , n21972 , n21973 );
buf ( n53007 , n53006 );
and ( n53008 , RI1754c2c8_9 , n34844 );
and ( n53009 , RI1754c2c8_9 , n34847 );
and ( n53010 , RI1754c2c8_9 , n34850 );
and ( n53011 , RI1754c2c8_9 , n34852 );
and ( n53012 , RI1754c2c8_9 , n34854 );
and ( n53013 , RI1754c2c8_9 , n34856 );
and ( n53014 , RI1754c2c8_9 , n39233 );
or ( n53015 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , C0 );
not ( n21974 , n34859 );
and ( n21975 , n21974 , n53015 );
and ( n21976 , RI1754c2c8_9 , n34859 );
or ( n53016 , n21975 , n21976 );
not ( n21977 , RI19a22f70_2797);
and ( n21978 , n21977 , n53016 );
and ( n21979 , C0 , RI19a22f70_2797);
or ( n53017 , n21978 , n21979 );
not ( n21980 , n27683 );
and ( n21981 , n21980 , RI19a88e38_2732);
and ( n21982 , n53017 , n27683 );
or ( n53018 , n21981 , n21982 );
not ( n21983 , RI1754c610_2);
and ( n21984 , n21983 , n53018 );
and ( n21985 , C0 , RI1754c610_2);
or ( n53019 , n21984 , n21985 );
buf ( n53020 , n53019 );
not ( n21986 , n27683 );
and ( n21987 , n21986 , RI19aa38c8_2541);
and ( n21988 , RI19aadd50_2469 , n27683 );
or ( n53021 , n21987 , n21988 );
not ( n21989 , RI1754c610_2);
and ( n21990 , n21989 , n53021 );
and ( n21991 , C0 , RI1754c610_2);
or ( n53022 , n21990 , n21991 );
buf ( n53023 , n53022 );
not ( n21992 , n27683 );
and ( n21993 , n21992 , RI19a8e6d0_2694);
and ( n21994 , RI19a98888_2622 , n27683 );
or ( n53024 , n21993 , n21994 );
not ( n21995 , RI1754c610_2);
and ( n21996 , n21995 , n53024 );
and ( n21997 , C0 , RI1754c610_2);
or ( n53025 , n21996 , n21997 );
buf ( n53026 , n53025 );
not ( n53027 , n39688 );
and ( n53028 , n53027 , n39703 );
xor ( n53029 , n44040 , n53028 );
not ( n21998 , n29614 );
and ( n21999 , n21998 , RI174a2738_944);
and ( n22000 , n53029 , n29614 );
or ( n53030 , n21999 , n22000 );
not ( n22001 , RI1754c610_2);
and ( n22002 , n22001 , n53030 );
and ( n22003 , C0 , RI1754c610_2);
or ( n53031 , n22002 , n22003 );
buf ( n53032 , n53031 );
not ( n53033 , n42980 );
and ( n53034 , n53033 , n42982 );
xor ( n53035 , n45175 , n53034 );
not ( n22004 , n29614 );
and ( n22005 , n22004 , RI1746e5c8_1198);
and ( n22006 , n53035 , n29614 );
or ( n53036 , n22005 , n22006 );
not ( n22007 , RI1754c610_2);
and ( n22008 , n22007 , n53036 );
and ( n22009 , C0 , RI1754c610_2);
or ( n53037 , n22008 , n22009 );
buf ( n53038 , n53037 );
and ( n53039 , RI1754c1d8_11 , n34844 );
and ( n53040 , RI1754c1d8_11 , n34847 );
and ( n53041 , RI1754c1d8_11 , n34850 );
and ( n53042 , RI1754c1d8_11 , n34852 );
and ( n53043 , RI1754c1d8_11 , n34854 );
and ( n53044 , RI1754c1d8_11 , n34856 );
or ( n53045 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , C0 , C0 );
not ( n22010 , n34859 );
and ( n22011 , n22010 , n53045 );
and ( n22012 , RI1754c1d8_11 , n34859 );
or ( n53046 , n22011 , n22012 );
not ( n22013 , RI19a22f70_2797);
and ( n22014 , n22013 , n53046 );
and ( n22015 , C0 , RI19a22f70_2797);
or ( n53047 , n22014 , n22015 );
not ( n22016 , n27683 );
and ( n22017 , n22016 , RI19a8b958_2714);
and ( n22018 , n53047 , n27683 );
or ( n53048 , n22017 , n22018 );
not ( n22019 , RI1754c610_2);
and ( n22020 , n22019 , n53048 );
and ( n22021 , C0 , RI1754c610_2);
or ( n53049 , n22020 , n22021 );
buf ( n53050 , n53049 );
not ( n22022 , n27683 );
and ( n22023 , n22022 , RI19a86c00_2747);
and ( n22024 , RI19a86de0_2746 , n27683 );
or ( n53051 , n22023 , n22024 );
not ( n22025 , RI1754c610_2);
and ( n22026 , n22025 , n53051 );
and ( n22027 , C0 , RI1754c610_2);
or ( n53052 , n22026 , n22027 );
buf ( n53053 , n53052 );
not ( n53054 , n48690 );
and ( n53055 , n53054 , n51881 );
xor ( n53056 , n48687 , n53055 );
not ( n22028 , n29614 );
and ( n22029 , n22028 , RI1733be90_2149);
and ( n22030 , n53056 , n29614 );
or ( n53057 , n22029 , n22030 );
not ( n22031 , RI1754c610_2);
and ( n22032 , n22031 , n53057 );
and ( n22033 , C0 , RI1754c610_2);
or ( n53058 , n22032 , n22033 );
buf ( n53059 , n53058 );
not ( n22034 , n27683 );
and ( n22035 , n22034 , RI19abaf50_2374);
and ( n22036 , RI19ac3920_2302 , n27683 );
or ( n53060 , n22035 , n22036 );
not ( n22037 , RI1754c610_2);
and ( n22038 , n22037 , n53060 );
and ( n22039 , C0 , RI1754c610_2);
or ( n53061 , n22038 , n22039 );
buf ( n53062 , n53061 );
not ( n53063 , n48868 );
and ( n53064 , n53063 , n42095 );
xor ( n53065 , n43122 , n53064 );
not ( n22040 , n29614 );
and ( n22041 , n22040 , RI17447ce8_1386);
and ( n22042 , n53065 , n29614 );
or ( n53066 , n22041 , n22042 );
not ( n22043 , RI1754c610_2);
and ( n22044 , n22043 , n53066 );
and ( n22045 , C0 , RI1754c610_2);
or ( n53067 , n22044 , n22045 );
buf ( n53068 , n53067 );
not ( n53069 , n50044 );
and ( n53070 , n53069 , n49549 );
xor ( n53071 , n49883 , n53070 );
not ( n22046 , n29614 );
and ( n22047 , n22046 , RI17526000_648);
and ( n22048 , n53071 , n29614 );
or ( n53072 , n22047 , n22048 );
not ( n22049 , RI1754c610_2);
and ( n22050 , n22049 , n53072 );
and ( n22051 , C0 , RI1754c610_2);
or ( n53073 , n22050 , n22051 );
buf ( n53074 , n53073 );
not ( n53075 , n45995 );
and ( n53076 , n53075 , n45997 );
xor ( n53077 , n46406 , n53076 );
not ( n22052 , n29614 );
and ( n22053 , n22052 , RI1740fb40_1431);
and ( n22054 , n53077 , n29614 );
or ( n53078 , n22053 , n22054 );
not ( n22055 , RI1754c610_2);
and ( n22056 , n22055 , n53078 );
and ( n22057 , C0 , RI1754c610_2);
or ( n53079 , n22056 , n22057 );
buf ( n53080 , n53079 );
not ( n53081 , n37815 );
and ( n53082 , n53081 , n45248 );
xor ( n53083 , n37745 , n53082 );
not ( n22058 , n29614 );
and ( n22059 , n22058 , RI173ee7b0_1593);
and ( n22060 , n53083 , n29614 );
or ( n53084 , n22059 , n22060 );
not ( n22061 , RI1754c610_2);
and ( n22062 , n22061 , n53084 );
and ( n22063 , C0 , RI1754c610_2);
or ( n53085 , n22062 , n22063 );
buf ( n53086 , n53085 );
not ( n53087 , n37870 );
and ( n53088 , n53087 , n37875 );
xor ( n53089 , n40666 , n53088 );
not ( n22064 , n29614 );
and ( n22065 , n22064 , RI173e18f8_1656);
and ( n22066 , n53089 , n29614 );
or ( n53090 , n22065 , n22066 );
not ( n22067 , RI1754c610_2);
and ( n22068 , n22067 , n53090 );
and ( n22069 , C0 , RI1754c610_2);
or ( n53091 , n22068 , n22069 );
buf ( n53092 , n53091 );
not ( n22070 , n27683 );
and ( n22071 , n22070 , RI19ac5540_2289);
and ( n22072 , RI19ace168_2224 , n27683 );
or ( n53093 , n22071 , n22072 );
not ( n22073 , RI1754c610_2);
and ( n22074 , n22073 , n53093 );
and ( n22075 , C0 , RI1754c610_2);
or ( n53094 , n22074 , n22075 );
buf ( n53095 , n53094 );
not ( n22076 , n27683 );
and ( n22077 , n22076 , RI19a9bd80_2599);
and ( n22078 , RI19aa53f8_2528 , n27683 );
or ( n53096 , n22077 , n22078 );
not ( n22079 , RI1754c610_2);
and ( n22080 , n22079 , n53096 );
and ( n22081 , C0 , RI1754c610_2);
or ( n53097 , n22080 , n22081 );
buf ( n53098 , n53097 );
not ( n53099 , n45728 );
and ( n53100 , n53099 , n45730 );
xor ( n53101 , n50080 , n53100 );
not ( n22082 , n29614 );
and ( n22083 , n22082 , RI173bf4e8_1823);
and ( n22084 , n53101 , n29614 );
or ( n53102 , n22083 , n22084 );
not ( n22085 , RI1754c610_2);
and ( n22086 , n22085 , n53102 );
and ( n22087 , C0 , RI1754c610_2);
or ( n53103 , n22086 , n22087 );
buf ( n53104 , n53103 );
not ( n53105 , n42414 );
and ( n53106 , n53105 , n46008 );
xor ( n53107 , n42411 , n53106 );
not ( n22088 , n29614 );
and ( n22089 , n22088 , RI1748c820_1051);
and ( n22090 , n53107 , n29614 );
or ( n53108 , n22089 , n22090 );
not ( n22091 , RI1754c610_2);
and ( n22092 , n22091 , n53108 );
and ( n22093 , C0 , RI1754c610_2);
or ( n53109 , n22092 , n22093 );
buf ( n53110 , n53109 );
not ( n53111 , n35656 );
and ( n53112 , n53111 , n35761 );
xor ( n53113 , n42564 , n53112 );
not ( n22094 , n29614 );
and ( n22095 , n22094 , RI174a3458_940);
and ( n22096 , n53113 , n29614 );
or ( n53114 , n22095 , n22096 );
not ( n22097 , RI1754c610_2);
and ( n22098 , n22097 , n53114 );
and ( n22099 , C0 , RI1754c610_2);
or ( n53115 , n22098 , n22099 );
buf ( n53116 , n53115 );
not ( n53117 , n46817 );
and ( n53118 , n53117 , n50812 );
xor ( n53119 , n46814 , n53118 );
not ( n22100 , n29614 );
and ( n22101 , n22100 , RI173d8208_1702);
and ( n22102 , n53119 , n29614 );
or ( n53120 , n22101 , n22102 );
not ( n22103 , RI1754c610_2);
and ( n22104 , n22103 , n53120 );
and ( n22105 , C0 , RI1754c610_2);
or ( n53121 , n22104 , n22105 );
buf ( n53122 , n53121 );
not ( n53123 , n48818 );
and ( n53124 , n53123 , n37312 );
xor ( n53125 , n44698 , n53124 );
not ( n22106 , n29614 );
and ( n22107 , n22106 , RI17494818_1012);
and ( n22108 , n53125 , n29614 );
or ( n53126 , n22107 , n22108 );
not ( n22109 , RI1754c610_2);
and ( n22110 , n22109 , n53126 );
and ( n22111 , C0 , RI1754c610_2);
or ( n53127 , n22110 , n22111 );
buf ( n53128 , n53127 );
not ( n53129 , n47533 );
and ( n53130 , n53129 , n50187 );
xor ( n53131 , n47530 , n53130 );
not ( n22112 , n29614 );
and ( n22113 , n22112 , RI173eafe8_1610);
and ( n22114 , n53131 , n29614 );
or ( n53132 , n22113 , n22114 );
not ( n22115 , RI1754c610_2);
and ( n22116 , n22115 , n53132 );
and ( n22117 , C0 , RI1754c610_2);
or ( n53133 , n22116 , n22117 );
buf ( n53134 , n53133 );
not ( n53135 , n43468 );
and ( n53136 , n53135 , n49120 );
xor ( n53137 , n43465 , n53136 );
not ( n22118 , n29614 );
and ( n22119 , n22118 , RI174ad868_890);
and ( n22120 , n53137 , n29614 );
or ( n53138 , n22119 , n22120 );
not ( n22121 , RI1754c610_2);
and ( n22122 , n22121 , n53138 );
and ( n22123 , C0 , RI1754c610_2);
or ( n53139 , n22122 , n22123 );
buf ( n53140 , n53139 );
not ( n22124 , n27683 );
and ( n22125 , n22124 , RI19a9f368_2575);
and ( n22126 , RI19aa8da0_2504 , n27683 );
or ( n53141 , n22125 , n22126 );
not ( n22127 , RI1754c610_2);
and ( n22128 , n22127 , n53141 );
and ( n22129 , C0 , RI1754c610_2);
or ( n53142 , n22128 , n22129 );
buf ( n53143 , n53142 );
not ( n22130 , n27683 );
and ( n22131 , n22130 , RI19a9ed50_2578);
and ( n22132 , RI19aa8530_2507 , n27683 );
or ( n53144 , n22131 , n22132 );
not ( n22133 , RI1754c610_2);
and ( n22134 , n22133 , n53144 );
and ( n22135 , C0 , RI1754c610_2);
or ( n53145 , n22134 , n22135 );
buf ( n53146 , n53145 );
not ( n53147 , n45896 );
and ( n53148 , n53147 , n43821 );
xor ( n53149 , n50982 , n53148 );
not ( n22136 , n29614 );
and ( n22137 , n22136 , RI1738a310_2082);
and ( n22138 , n53149 , n29614 );
or ( n53150 , n22137 , n22138 );
not ( n22139 , RI1754c610_2);
and ( n22140 , n22139 , n53150 );
and ( n22141 , C0 , RI1754c610_2);
or ( n53151 , n22140 , n22141 );
buf ( n53152 , n53151 );
not ( n22142 , n27683 );
and ( n22143 , n22142 , RI19a8aad0_2720);
and ( n22144 , RI19a94940_2650 , n27683 );
or ( n53153 , n22143 , n22144 );
not ( n22145 , RI1754c610_2);
and ( n22146 , n22145 , n53153 );
and ( n22147 , C0 , RI1754c610_2);
or ( n53154 , n22146 , n22147 );
buf ( n53155 , n53154 );
not ( n53156 , n50402 );
and ( n53157 , n53156 , n50404 );
xor ( n53158 , n46971 , n53157 );
not ( n22148 , n29614 );
and ( n22149 , n22148 , RI17395ad0_2026);
and ( n22150 , n53158 , n29614 );
or ( n53159 , n22149 , n22150 );
not ( n22151 , RI1754c610_2);
and ( n22152 , n22151 , n53159 );
and ( n22153 , C0 , RI1754c610_2);
or ( n53160 , n22152 , n22153 );
buf ( n53161 , n53160 );
not ( n53162 , n43079 );
and ( n53163 , n53162 , n41337 );
xor ( n53164 , n48006 , n53163 );
not ( n22154 , n29614 );
and ( n22155 , n22154 , RI17406ae0_1475);
and ( n22156 , n53164 , n29614 );
or ( n53165 , n22155 , n22156 );
not ( n22157 , RI1754c610_2);
and ( n22158 , n22157 , n53165 );
and ( n22159 , C0 , RI1754c610_2);
or ( n53166 , n22158 , n22159 );
buf ( n53167 , n53166 );
buf ( n53168 , RI174af938_880);
not ( n53169 , n42820 );
and ( n53170 , n53169 , n42822 );
xor ( n53171 , n51591 , n53170 );
not ( n22160 , n29614 );
and ( n22161 , n22160 , RI1749d530_969);
and ( n22162 , n53171 , n29614 );
or ( n53172 , n22161 , n22162 );
not ( n22163 , RI1754c610_2);
and ( n22164 , n22163 , n53172 );
and ( n22165 , C0 , RI1754c610_2);
or ( n53173 , n22164 , n22165 );
buf ( n53174 , n53173 );
buf ( n53175 , RI174ac800_895);
not ( n53176 , n43911 );
and ( n53177 , n53176 , n43913 );
xor ( n53178 , n44382 , n53177 );
not ( n22166 , n29614 );
and ( n22167 , n22166 , RI173b08a8_1895);
and ( n22168 , n53178 , n29614 );
or ( n53179 , n22167 , n22168 );
not ( n22169 , RI1754c610_2);
and ( n22170 , n22169 , n53179 );
and ( n22171 , C0 , RI1754c610_2);
or ( n53180 , n22170 , n22171 );
buf ( n53181 , n53180 );
buf ( n53182 , RI1746efa0_1195);
buf ( n53183 , RI1746bb20_1211);
buf ( n53184 , RI17478000_1151);
buf ( n53185 , RI17474838_1168);
buf ( n53186 , RI174a6c20_923);
buf ( n53187 , RI174a37a0_939);
not ( n53188 , n45134 );
and ( n53189 , n53188 , n52345 );
xor ( n53190 , n45131 , n53189 );
not ( n22172 , n29614 );
and ( n22173 , n22172 , RI174641b8_1248);
and ( n22174 , n53190 , n29614 );
or ( n53191 , n22173 , n22174 );
not ( n22175 , RI1754c610_2);
and ( n22176 , n22175 , n53191 );
and ( n22177 , C0 , RI1754c610_2);
or ( n53192 , n22176 , n22177 );
buf ( n53193 , n53192 );
and ( n53194 , RI19a24a28_2784 , n43086 );
not ( n22178 , n43088 );
and ( n22179 , n22178 , RI19a247d0_2785);
and ( n22180 , n53194 , n43088 );
or ( n53195 , n22179 , n22180 );
not ( n22181 , RI1754c610_2);
and ( n22182 , n22181 , n53195 );
and ( n22183 , C0 , RI1754c610_2);
or ( n53196 , n22182 , n22183 );
buf ( n53197 , n53196 );
buf ( n53198 , RI174aa730_905);
buf ( n53199 , RI17469078_1224);
buf ( n53200 , RI174a8cf0_913);
not ( n53201 , n52348 );
and ( n53202 , n53201 , n45129 );
xor ( n53203 , n52345 , n53202 );
not ( n22184 , n29614 );
and ( n22185 , n22184 , RI174813a8_1106);
and ( n22186 , n53203 , n29614 );
or ( n53204 , n22185 , n22186 );
not ( n22187 , RI1754c610_2);
and ( n22188 , n22187 , n53204 );
and ( n22189 , C0 , RI1754c610_2);
or ( n53205 , n22188 , n22189 );
buf ( n53206 , n53205 );
not ( n22190 , n27683 );
and ( n22191 , n22190 , RI19a8efb8_2690);
and ( n22192 , RI19a98f90_2619 , n27683 );
or ( n53207 , n22191 , n22192 );
not ( n22193 , RI1754c610_2);
and ( n22194 , n22193 , n53207 );
and ( n22195 , C0 , RI1754c610_2);
or ( n53208 , n22194 , n22195 );
buf ( n53209 , n53208 );
xor ( n53210 , n39993 , n40341 );
xor ( n53211 , n53210 , n40091 );
xor ( n53212 , n35501 , n38532 );
xor ( n53213 , n53212 , n38933 );
not ( n53214 , n53213 );
xor ( n53215 , n34992 , n42945 );
xor ( n53216 , n53215 , n34497 );
and ( n53217 , n53214 , n53216 );
xor ( n53218 , n53211 , n53217 );
not ( n22196 , n29614 );
and ( n22197 , n22196 , RI17343b40_2111);
and ( n22198 , n53218 , n29614 );
or ( n53219 , n22197 , n22198 );
not ( n22199 , RI1754c610_2);
and ( n22200 , n22199 , n53219 );
and ( n22201 , C0 , RI1754c610_2);
or ( n53220 , n22200 , n22201 );
buf ( n53221 , n53220 );
not ( n53222 , n39115 );
and ( n53223 , n53222 , n39152 );
xor ( n53224 , n40600 , n53223 );
not ( n22202 , n29614 );
and ( n22203 , n22202 , RI174c62a0_794);
and ( n22204 , n53224 , n29614 );
or ( n53225 , n22203 , n22204 );
not ( n22205 , RI1754c610_2);
and ( n22206 , n22205 , n53225 );
and ( n22207 , C0 , RI1754c610_2);
or ( n53226 , n22206 , n22207 );
buf ( n53227 , n53226 );
not ( n53228 , n42325 );
and ( n53229 , n53228 , n43022 );
xor ( n53230 , n42322 , n53229 );
not ( n22208 , n29614 );
and ( n22209 , n22208 , RI174aa3e8_906);
and ( n22210 , n53230 , n29614 );
or ( n53231 , n22209 , n22210 );
not ( n22211 , RI1754c610_2);
and ( n22212 , n22211 , n53231 );
and ( n22213 , C0 , RI1754c610_2);
or ( n53232 , n22212 , n22213 );
buf ( n53233 , n53232 );
not ( n22214 , n27683 );
and ( n22215 , n22214 , RI19acffe0_2211);
and ( n22216 , RI19aa8f80_2503 , n27683 );
or ( n53234 , n22215 , n22216 );
not ( n22217 , RI1754c610_2);
and ( n22218 , n22217 , n53234 );
and ( n22219 , C0 , RI1754c610_2);
or ( n53235 , n22218 , n22219 );
buf ( n53236 , n53235 );
not ( n22220 , n27683 );
and ( n22221 , n22220 , RI19ab8f70_2388);
and ( n22222 , RI19ac1850_2318 , n27683 );
or ( n53237 , n22221 , n22222 );
not ( n22223 , RI1754c610_2);
and ( n22224 , n22223 , n53237 );
and ( n22225 , C0 , RI1754c610_2);
or ( n53238 , n22224 , n22225 );
buf ( n53239 , n53238 );
not ( n22226 , n27683 );
and ( n22227 , n22226 , RI19a936f8_2658);
and ( n22228 , RI19a9d9a0_2587 , n27683 );
or ( n53240 , n22227 , n22228 );
not ( n22229 , RI1754c610_2);
and ( n22230 , n22229 , n53240 );
and ( n22231 , C0 , RI1754c610_2);
or ( n53241 , n22230 , n22231 );
buf ( n53242 , n53241 );
not ( n53243 , n44326 );
and ( n53244 , n53243 , n43662 );
xor ( n53245 , n44323 , n53244 );
not ( n22232 , n29614 );
and ( n22233 , n22232 , RI173c3d18_1801);
and ( n22234 , n53245 , n29614 );
or ( n53246 , n22233 , n22234 );
not ( n22235 , RI1754c610_2);
and ( n22236 , n22235 , n53246 );
and ( n22237 , C0 , RI1754c610_2);
or ( n53247 , n22236 , n22237 );
buf ( n53248 , n53247 );
not ( n53249 , n43004 );
and ( n53250 , n53249 , n42357 );
xor ( n53251 , n44592 , n53250 );
not ( n22238 , n29614 );
and ( n22239 , n22238 , RI1738e168_2063);
and ( n22240 , n53251 , n29614 );
or ( n53252 , n22239 , n22240 );
not ( n22241 , RI1754c610_2);
and ( n22242 , n22241 , n53252 );
and ( n22243 , C0 , RI1754c610_2);
or ( n53253 , n22242 , n22243 );
buf ( n53254 , n53253 );
not ( n53255 , n45075 );
and ( n53256 , n53255 , n48718 );
xor ( n53257 , n45072 , n53256 );
not ( n22244 , n29614 );
and ( n22245 , n22244 , RI174465f0_1393);
and ( n22246 , n53257 , n29614 );
or ( n53258 , n22245 , n22246 );
not ( n22247 , RI1754c610_2);
and ( n22248 , n22247 , n53258 );
and ( n22249 , C0 , RI1754c610_2);
or ( n53259 , n22248 , n22249 );
buf ( n53260 , n53259 );
not ( n53261 , n43597 );
and ( n53262 , n53261 , n41227 );
xor ( n53263 , n46289 , n53262 );
not ( n22250 , n29614 );
and ( n22251 , n22250 , RI173d39d8_1724);
and ( n22252 , n53263 , n29614 );
or ( n53264 , n22251 , n22252 );
not ( n22253 , RI1754c610_2);
and ( n22254 , n22253 , n53264 );
and ( n22255 , C0 , RI1754c610_2);
or ( n53265 , n22254 , n22255 );
buf ( n53266 , n53265 );
not ( n53267 , n47311 );
and ( n53268 , n53267 , n48180 );
xor ( n53269 , n47308 , n53268 );
not ( n22256 , n29614 );
and ( n22257 , n22256 , RI173e6e48_1630);
and ( n22258 , n53269 , n29614 );
or ( n53270 , n22257 , n22258 );
not ( n22259 , RI1754c610_2);
and ( n22260 , n22259 , n53270 );
and ( n22261 , C0 , RI1754c610_2);
or ( n53271 , n22260 , n22261 );
buf ( n53272 , n53271 );
not ( n53273 , n44382 );
and ( n53274 , n53273 , n43911 );
xor ( n53275 , n44379 , n53274 );
not ( n22262 , n29614 );
and ( n22263 , n22262 , RI173a1fb0_1966);
and ( n22264 , n53275 , n29614 );
or ( n53276 , n22263 , n22264 );
not ( n22265 , RI1754c610_2);
and ( n22266 , n22265 , n53276 );
and ( n22267 , C0 , RI1754c610_2);
or ( n53277 , n22266 , n22267 );
buf ( n53278 , n53277 );
not ( n22268 , n27683 );
and ( n22269 , n22268 , RI19a91358_2674);
and ( n22270 , RI19a9b678_2602 , n27683 );
or ( n53279 , n22269 , n22270 );
not ( n22271 , RI1754c610_2);
and ( n22272 , n22271 , n53279 );
and ( n22273 , C0 , RI1754c610_2);
or ( n53280 , n22272 , n22273 );
buf ( n53281 , n53280 );
not ( n53282 , n44147 );
and ( n53283 , n53282 , n44149 );
xor ( n53284 , n51445 , n53283 );
not ( n22274 , n29614 );
and ( n22275 , n22274 , RI174a5bb8_928);
and ( n22276 , n53284 , n29614 );
or ( n53285 , n22275 , n22276 );
not ( n22277 , RI1754c610_2);
and ( n22278 , n22277 , n53285 );
and ( n22279 , C0 , RI1754c610_2);
or ( n53286 , n22278 , n22279 );
buf ( n53287 , n53286 );
not ( n53288 , n49053 );
and ( n53289 , n53288 , n43207 );
xor ( n53290 , n51113 , n53289 );
not ( n22280 , n29614 );
and ( n22281 , n22280 , RI1749fc90_957);
and ( n22282 , n53290 , n29614 );
or ( n53291 , n22281 , n22282 );
not ( n22283 , RI1754c610_2);
and ( n22284 , n22283 , n53291 );
and ( n22285 , C0 , RI1754c610_2);
or ( n53292 , n22284 , n22285 );
buf ( n53293 , n53292 );
not ( n53294 , n46856 );
xor ( n53295 , n36430 , n33935 );
xor ( n53296 , n53295 , n36287 );
and ( n53297 , n53294 , n53296 );
xor ( n53298 , n46853 , n53297 );
not ( n22286 , n29614 );
and ( n22287 , n22286 , RI17461080_1263);
and ( n22288 , n53298 , n29614 );
or ( n53299 , n22287 , n22288 );
not ( n22289 , RI1754c610_2);
and ( n22290 , n22289 , n53299 );
and ( n22291 , C0 , RI1754c610_2);
or ( n53300 , n22290 , n22291 );
buf ( n53301 , n53300 );
not ( n53302 , n38038 );
and ( n53303 , n53302 , n43324 );
xor ( n53304 , n37944 , n53303 );
not ( n22292 , n29614 );
and ( n22293 , n22292 , RI174a2dc8_942);
and ( n22294 , n53304 , n29614 );
or ( n53305 , n22293 , n22294 );
not ( n22295 , RI1754c610_2);
and ( n22296 , n22295 , n53305 );
and ( n22297 , C0 , RI1754c610_2);
or ( n53306 , n22296 , n22297 );
buf ( n53307 , n53306 );
not ( n53308 , n42520 );
and ( n53309 , n53308 , n42522 );
xor ( n53310 , n46648 , n53309 );
not ( n22298 , n29614 );
and ( n22299 , n22298 , RI173e2ca8_1650);
and ( n22300 , n53310 , n29614 );
or ( n53311 , n22299 , n22300 );
not ( n22301 , RI1754c610_2);
and ( n22302 , n22301 , n53311 );
and ( n22303 , C0 , RI1754c610_2);
or ( n53312 , n22302 , n22303 );
buf ( n53313 , n53312 );
not ( n53314 , n40217 );
and ( n53315 , n53314 , n48412 );
xor ( n53316 , n40211 , n53315 );
not ( n22304 , n29614 );
and ( n22305 , n22304 , RI1747c1a0_1131);
and ( n22306 , n53316 , n29614 );
or ( n53317 , n22305 , n22306 );
not ( n22307 , RI1754c610_2);
and ( n22308 , n22307 , n53317 );
and ( n22309 , C0 , RI1754c610_2);
or ( n53318 , n22308 , n22309 );
buf ( n53319 , n53318 );
buf ( n53320 , RI174ae240_887);
buf ( n53321 , RI174ce8b0_768);
not ( n53322 , n46971 );
and ( n53323 , n53322 , n50402 );
xor ( n53324 , n46968 , n53323 );
not ( n22310 , n29614 );
and ( n22311 , n22310 , RI173465e8_2098);
and ( n22312 , n53324 , n29614 );
or ( n53325 , n22311 , n22312 );
not ( n22313 , RI1754c610_2);
and ( n22314 , n22313 , n53325 );
and ( n22315 , C0 , RI1754c610_2);
or ( n53326 , n22314 , n22315 );
buf ( n53327 , n53326 );
buf ( n53328 , RI17490330_1033);
buf ( n53329 , RI174a4b50_933);
and ( n53330 , RI1754b170_46 , n34844 );
and ( n53331 , RI1754b170_46 , n34847 );
or ( n53332 , n53330 , n53331 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n22316 , n34859 );
and ( n22317 , n22316 , n53332 );
and ( n22318 , RI1754b170_46 , n34859 );
or ( n53333 , n22317 , n22318 );
not ( n22319 , RI19a22f70_2797);
and ( n22320 , n22319 , n53333 );
and ( n22321 , C0 , RI19a22f70_2797);
or ( n53334 , n22320 , n22321 );
not ( n22322 , n27683 );
and ( n22323 , n22322 , RI19ac0a40_2326);
and ( n22324 , n53334 , n27683 );
or ( n53335 , n22323 , n22324 );
not ( n22325 , RI1754c610_2);
and ( n22326 , n22325 , n53335 );
and ( n22327 , C0 , RI1754c610_2);
or ( n53336 , n22326 , n22327 );
buf ( n53337 , n53336 );
not ( n53338 , n45942 );
and ( n53339 , n53338 , n45944 );
xor ( n53340 , n51271 , n53339 );
not ( n22328 , n29614 );
and ( n22329 , n22328 , RI174a4b50_933);
and ( n22330 , n53340 , n29614 );
or ( n53341 , n22329 , n22330 );
not ( n22331 , RI1754c610_2);
and ( n22332 , n22331 , n53341 );
and ( n22333 , C0 , RI1754c610_2);
or ( n53342 , n22332 , n22333 );
buf ( n53343 , n53342 );
not ( n53344 , n49770 );
and ( n53345 , n53344 , n49772 );
xor ( n53346 , n48451 , n53345 );
not ( n22334 , n29614 );
and ( n22335 , n22334 , RI174118c8_1422);
and ( n22336 , n53346 , n29614 );
or ( n53347 , n22335 , n22336 );
not ( n22337 , RI1754c610_2);
and ( n22338 , n22337 , n53347 );
and ( n22339 , C0 , RI1754c610_2);
or ( n53348 , n22338 , n22339 );
buf ( n53349 , n53348 );
not ( n53350 , n45009 );
and ( n53351 , n53350 , n50018 );
xor ( n53352 , n45006 , n53351 );
not ( n22340 , n29614 );
and ( n22341 , n22340 , RI174a0668_954);
and ( n22342 , n53352 , n29614 );
or ( n53353 , n22341 , n22342 );
not ( n22343 , RI1754c610_2);
and ( n22344 , n22343 , n53353 );
and ( n22345 , C0 , RI1754c610_2);
or ( n53354 , n22344 , n22345 );
buf ( n53355 , n53354 );
not ( n53356 , n46738 );
and ( n53357 , n53356 , n50276 );
xor ( n53358 , n46735 , n53357 );
not ( n22346 , n29614 );
and ( n22347 , n22346 , RI17451090_1341);
and ( n22348 , n53358 , n29614 );
or ( n53359 , n22347 , n22348 );
not ( n22349 , RI1754c610_2);
and ( n22350 , n22349 , n53359 );
and ( n22351 , C0 , RI1754c610_2);
or ( n53360 , n22350 , n22351 );
buf ( n53361 , n53360 );
not ( n53362 , n41505 );
and ( n53363 , n53362 , n45331 );
xor ( n53364 , n41480 , n53363 );
not ( n22352 , n29614 );
and ( n22353 , n22352 , RI173e7190_1629);
and ( n22354 , n53364 , n29614 );
or ( n53365 , n22353 , n22354 );
not ( n22355 , RI1754c610_2);
and ( n22356 , n22355 , n53365 );
and ( n22357 , C0 , RI1754c610_2);
or ( n53366 , n22356 , n22357 );
buf ( n53367 , n53366 );
not ( n53368 , n43057 );
and ( n53369 , n53368 , n43059 );
xor ( n53370 , n45440 , n53369 );
not ( n22358 , n29614 );
and ( n22359 , n22358 , RI1747f620_1115);
and ( n22360 , n53370 , n29614 );
or ( n53371 , n22359 , n22360 );
not ( n22361 , RI1754c610_2);
and ( n22362 , n22361 , n53371 );
and ( n22363 , C0 , RI1754c610_2);
or ( n53372 , n22362 , n22363 );
buf ( n53373 , n53372 );
not ( n22364 , n34859 );
and ( n22365 , n22364 , C0 );
and ( n22366 , RI1754aae0_60 , n34859 );
or ( n53374 , n22365 , n22366 );
not ( n22367 , RI19a22f70_2797);
and ( n22368 , n22367 , n53374 );
and ( n22369 , C0 , RI19a22f70_2797);
or ( n53375 , n22368 , n22369 );
not ( n22370 , n27683 );
and ( n22371 , n22370 , RI19a86de0_2746);
and ( n22372 , n53375 , n27683 );
or ( n53376 , n22371 , n22372 );
not ( n22373 , RI1754c610_2);
and ( n22374 , n22373 , n53376 );
and ( n22375 , C0 , RI1754c610_2);
or ( n53377 , n22374 , n22375 );
buf ( n53378 , n53377 );
and ( n53379 , RI1754acc0_56 , n34844 );
buf ( n53380 , n53379 );
not ( n22376 , n34859 );
and ( n22377 , n22376 , n53380 );
and ( n22378 , RI1754acc0_56 , n34859 );
or ( n53381 , n22377 , n22378 );
not ( n22379 , RI19a22f70_2797);
and ( n22380 , n22379 , n53381 );
and ( n22381 , C0 , RI19a22f70_2797);
or ( n53382 , n22380 , n22381 );
not ( n22382 , n27683 );
and ( n22383 , n22382 , RI19a23c18_2790);
and ( n22384 , n53382 , n27683 );
or ( n53383 , n22383 , n22384 );
not ( n22385 , RI1754c610_2);
and ( n22386 , n22385 , n53383 );
and ( n22387 , C0 , RI1754c610_2);
or ( n53384 , n22386 , n22387 );
buf ( n53385 , n53384 );
buf ( n53386 , RI17465f40_1239);
buf ( n53387 , RI17475be8_1162);
not ( n53388 , n47816 );
and ( n53389 , n53388 , n47744 );
xor ( n53390 , n45113 , n53389 );
not ( n22388 , n29614 );
and ( n22389 , n22388 , RI174565e0_1315);
and ( n22390 , n53390 , n29614 );
or ( n53391 , n22389 , n22390 );
not ( n22391 , RI1754c610_2);
and ( n22392 , n22391 , n53391 );
and ( n22393 , C0 , RI1754c610_2);
or ( n53392 , n22392 , n22393 );
buf ( n53393 , n53392 );
not ( n22394 , n27683 );
and ( n22395 , n22394 , RI19a87b78_2740);
and ( n22396 , RI19ad0238_2210 , n27683 );
or ( n53394 , n22395 , n22396 );
not ( n22397 , RI1754c610_2);
and ( n22398 , n22397 , n53394 );
and ( n22399 , C0 , RI1754c610_2);
or ( n53395 , n22398 , n22399 );
buf ( n53396 , n53395 );
not ( n22400 , n27683 );
and ( n22401 , n22400 , RI19a82f88_2773);
and ( n22402 , RI19ab2508_2437 , n27683 );
or ( n53397 , n22401 , n22402 );
not ( n22403 , RI1754c610_2);
and ( n22404 , n22403 , n53397 );
and ( n22405 , C0 , RI1754c610_2);
or ( n53398 , n22404 , n22405 );
buf ( n53399 , n53398 );
not ( n53400 , n43584 );
and ( n53401 , n53400 , n43586 );
xor ( n53402 , n49080 , n53401 );
not ( n22406 , n29614 );
and ( n22407 , n22406 , RI173a39f0_1958);
and ( n22408 , n53402 , n29614 );
or ( n53403 , n22407 , n22408 );
not ( n22409 , RI1754c610_2);
and ( n22410 , n22409 , n53403 );
and ( n22411 , C0 , RI1754c610_2);
or ( n53404 , n22410 , n22411 );
buf ( n53405 , n53404 );
not ( n53406 , n45331 );
and ( n53407 , n53406 , n45333 );
xor ( n53408 , n41505 , n53407 );
not ( n22412 , n29614 );
and ( n22413 , n22412 , RI173f5740_1559);
and ( n22414 , n53408 , n29614 );
or ( n53409 , n22413 , n22414 );
not ( n22415 , RI1754c610_2);
and ( n22416 , n22415 , n53409 );
and ( n22417 , C0 , RI1754c610_2);
or ( n53410 , n22416 , n22417 );
buf ( n53411 , n53410 );
not ( n53412 , n47012 );
and ( n53413 , n53412 , n51271 );
xor ( n53414 , n45947 , n53413 );
not ( n22418 , n29614 );
and ( n22419 , n22418 , RI17487ca8_1074);
and ( n22420 , n53414 , n29614 );
or ( n53415 , n22419 , n22420 );
not ( n22421 , RI1754c610_2);
and ( n22422 , n22421 , n53415 );
and ( n22423 , C0 , RI1754c610_2);
or ( n53416 , n22422 , n22423 );
buf ( n53417 , n53416 );
not ( n22424 , n27683 );
and ( n22425 , n22424 , RI19ac1a30_2317);
and ( n22426 , RI19acaf40_2248 , n27683 );
or ( n53418 , n22425 , n22426 );
not ( n22427 , RI1754c610_2);
and ( n22428 , n22427 , n53418 );
and ( n22429 , C0 , RI1754c610_2);
or ( n53419 , n22428 , n22429 );
buf ( n53420 , n53419 );
not ( n22430 , n27683 );
and ( n22431 , n22430 , RI19a8faf8_2685);
and ( n22432 , RI19a99d28_2613 , n27683 );
or ( n53421 , n22431 , n22432 );
not ( n22433 , RI1754c610_2);
and ( n22434 , n22433 , n53421 );
and ( n22435 , C0 , RI1754c610_2);
or ( n53422 , n22434 , n22435 );
buf ( n53423 , n53422 );
buf ( n53424 , RI1749f600_959);
buf ( n53425 , RI174b3ad8_860);
not ( n53426 , n49454 );
and ( n53427 , n53426 , n49456 );
xor ( n53428 , n42350 , n53427 );
not ( n22436 , n29614 );
and ( n22437 , n22436 , RI173c5758_1793);
and ( n22438 , n53428 , n29614 );
or ( n53429 , n22437 , n22438 );
not ( n22439 , RI1754c610_2);
and ( n22440 , n22439 , n53429 );
and ( n22441 , C0 , RI1754c610_2);
or ( n53430 , n22440 , n22441 );
buf ( n53431 , n53430 );
buf ( n53432 , RI17502e70_751);
buf ( n53433 , RI17489058_1068);
not ( n53434 , n45624 );
and ( n53435 , n53434 , n45626 );
xor ( n53436 , n48830 , n53435 );
not ( n22442 , n29614 );
and ( n22443 , n22442 , RI17507628_743);
and ( n22444 , n53436 , n29614 );
or ( n53437 , n22443 , n22444 );
not ( n22445 , RI1754c610_2);
and ( n22446 , n22445 , n53437 );
and ( n22447 , C0 , RI1754c610_2);
or ( n53438 , n22446 , n22447 );
buf ( n53439 , n53438 );
not ( n53440 , n47181 );
and ( n53441 , n53440 , n41017 );
xor ( n53442 , n50365 , n53441 );
not ( n22448 , n29614 );
and ( n22449 , n22448 , RI174620e8_1258);
and ( n22450 , n53442 , n29614 );
or ( n53443 , n22449 , n22450 );
not ( n22451 , RI1754c610_2);
and ( n22452 , n22451 , n53443 );
and ( n22453 , C0 , RI1754c610_2);
or ( n53444 , n22452 , n22453 );
buf ( n53445 , n53444 );
not ( n22454 , n27683 );
and ( n22455 , n22454 , RI19ac2f48_2307);
and ( n22456 , RI19acbe40_2240 , n27683 );
or ( n53446 , n22455 , n22456 );
not ( n22457 , RI1754c610_2);
and ( n22458 , n22457 , n53446 );
and ( n22459 , C0 , RI1754c610_2);
or ( n53447 , n22458 , n22459 );
buf ( n53448 , n53447 );
not ( n22460 , n27683 );
and ( n22461 , n22460 , RI19ab4380_2422);
and ( n22462 , RI19abdbd8_2352 , n27683 );
or ( n53449 , n22461 , n22462 );
not ( n22463 , RI1754c610_2);
and ( n22464 , n22463 , n53449 );
and ( n22465 , C0 , RI1754c610_2);
or ( n53450 , n22464 , n22465 );
buf ( n53451 , n53450 );
not ( n53452 , n40978 );
and ( n53453 , n53452 , n40980 );
xor ( n53454 , n40383 , n53453 );
not ( n22466 , n29614 );
and ( n22467 , n22466 , RI174b6c10_845);
and ( n22468 , n53454 , n29614 );
or ( n53455 , n22467 , n22468 );
not ( n22469 , RI1754c610_2);
and ( n22470 , n22469 , n53455 );
and ( n22471 , C0 , RI1754c610_2);
or ( n53456 , n22470 , n22471 );
buf ( n53457 , n53456 );
not ( n53458 , n44665 );
and ( n53459 , n53458 , n40062 );
xor ( n53460 , n44662 , n53459 );
not ( n22472 , n29614 );
and ( n22473 , n22472 , RI17334bb8_2184);
and ( n22474 , n53460 , n29614 );
or ( n53461 , n22473 , n22474 );
not ( n22475 , RI1754c610_2);
and ( n22476 , n22475 , n53461 );
and ( n22477 , C0 , RI1754c610_2);
or ( n53462 , n22476 , n22477 );
buf ( n53463 , n53462 );
not ( n53464 , n30742 );
xor ( n53465 , n35350 , n41005 );
xor ( n53466 , n53465 , n40585 );
and ( n53467 , n53464 , n53466 );
xor ( n53468 , n30462 , n53467 );
not ( n22478 , n29614 );
and ( n22479 , n22478 , RI1738e7f8_2061);
and ( n22480 , n53468 , n29614 );
or ( n53469 , n22479 , n22480 );
not ( n22481 , RI1754c610_2);
and ( n22482 , n22481 , n53469 );
and ( n22483 , C0 , RI1754c610_2);
or ( n53470 , n22482 , n22483 );
buf ( n53471 , n53470 );
not ( n53472 , n44176 );
and ( n53473 , n53472 , n51282 );
xor ( n53474 , n44173 , n53473 );
not ( n22484 , n29614 );
and ( n22485 , n22484 , RI173d4a40_1719);
and ( n22486 , n53474 , n29614 );
or ( n53475 , n22485 , n22486 );
not ( n22487 , RI1754c610_2);
and ( n22488 , n22487 , n53475 );
and ( n22489 , C0 , RI1754c610_2);
or ( n53476 , n22488 , n22489 );
buf ( n53477 , n53476 );
not ( n22490 , RI1754c610_2);
and ( n22491 , n22490 , RI17536d88_596);
and ( n22492 , C0 , RI1754c610_2);
or ( n53478 , n22491 , n22492 );
buf ( n53479 , n53478 );
not ( n53480 , n51121 );
and ( n53481 , n53480 , n51123 );
xor ( n53482 , n46783 , n53481 );
not ( n22493 , n29614 );
and ( n22494 , n22493 , RI173ac3c0_1916);
and ( n22495 , n53482 , n29614 );
or ( n53483 , n22494 , n22495 );
not ( n22496 , RI1754c610_2);
and ( n22497 , n22496 , n53483 );
and ( n22498 , C0 , RI1754c610_2);
or ( n53484 , n22497 , n22498 );
buf ( n53485 , n53484 );
buf ( n53486 , RI174bd768_821);
buf ( n53487 , RI1750fc38_717);
buf ( n53488 , RI174820c8_1102);
buf ( n53489 , RI1749add0_981);
not ( n53490 , n48937 );
and ( n53491 , n53490 , n51152 );
xor ( n53492 , n48934 , n53491 );
not ( n22499 , n29614 );
and ( n22500 , n22499 , RI17405730_1481);
and ( n22501 , n53492 , n29614 );
or ( n53493 , n22500 , n22501 );
not ( n22502 , RI1754c610_2);
and ( n22503 , n22502 , n53493 );
and ( n22504 , C0 , RI1754c610_2);
or ( n53494 , n22503 , n22504 );
buf ( n53495 , n53494 );
not ( n22505 , n27683 );
and ( n22506 , n22505 , RI19aae110_2467);
and ( n22507 , RI19ab7da0_2396 , n27683 );
or ( n53496 , n22506 , n22507 );
not ( n22508 , RI1754c610_2);
and ( n22509 , n22508 , n53496 );
and ( n22510 , C0 , RI1754c610_2);
or ( n53497 , n22509 , n22510 );
buf ( n53498 , n53497 );
not ( n53499 , n48233 );
and ( n53500 , n53499 , n49973 );
xor ( n53501 , n40120 , n53500 );
not ( n22511 , n29614 );
and ( n22512 , n22511 , RI173a0570_1974);
and ( n22513 , n53501 , n29614 );
or ( n53502 , n22512 , n22513 );
not ( n22514 , RI1754c610_2);
and ( n22515 , n22514 , n53502 );
and ( n22516 , C0 , RI1754c610_2);
or ( n53503 , n22515 , n22516 );
buf ( n53504 , n53503 );
not ( n53505 , n52251 );
and ( n53506 , n53505 , n52253 );
xor ( n53507 , n46663 , n53506 );
not ( n22517 , n29614 );
and ( n22518 , n22517 , RI173bc3b0_1838);
and ( n22519 , n53507 , n29614 );
or ( n53508 , n22518 , n22519 );
not ( n22520 , RI1754c610_2);
and ( n22521 , n22520 , n53508 );
and ( n22522 , C0 , RI1754c610_2);
or ( n53509 , n22521 , n22522 );
buf ( n53510 , n53509 );
not ( n53511 , n45248 );
and ( n53512 , n53511 , n45250 );
xor ( n53513 , n37815 , n53512 );
not ( n22523 , n29614 );
and ( n22524 , n22523 , RI173fd0a8_1522);
and ( n22525 , n53513 , n29614 );
or ( n53514 , n22524 , n22525 );
not ( n22526 , RI1754c610_2);
and ( n22527 , n22526 , n53514 );
and ( n22528 , C0 , RI1754c610_2);
or ( n53515 , n22527 , n22528 );
buf ( n53516 , n53515 );
not ( n53517 , n43402 );
and ( n53518 , n53517 , n45752 );
xor ( n53519 , n43399 , n53518 );
not ( n22529 , n29614 );
and ( n22530 , n22529 , RI17338380_2167);
and ( n22531 , n53519 , n29614 );
or ( n53520 , n22530 , n22531 );
not ( n22532 , RI1754c610_2);
and ( n22533 , n22532 , n53520 );
and ( n22534 , C0 , RI1754c610_2);
or ( n53521 , n22533 , n22534 );
buf ( n53522 , n53521 );
buf ( n53523 , RI1746c840_1207);
not ( n22535 , n27683 );
and ( n22536 , n22535 , RI19aaaa38_2491);
and ( n22537 , RI19ab4740_2420 , n27683 );
or ( n53524 , n22536 , n22537 );
not ( n22538 , RI1754c610_2);
and ( n22539 , n22538 , n53524 );
and ( n22540 , C0 , RI1754c610_2);
or ( n53525 , n22539 , n22540 );
buf ( n53526 , n53525 );
not ( n53527 , n43850 );
and ( n53528 , n53527 , n43745 );
xor ( n53529 , n43847 , n53528 );
not ( n22541 , n29614 );
and ( n22542 , n22541 , RI174658b0_1241);
and ( n22543 , n53529 , n29614 );
or ( n53530 , n22542 , n22543 );
not ( n22544 , RI1754c610_2);
and ( n22545 , n22544 , n53530 );
and ( n22546 , C0 , RI1754c610_2);
or ( n53531 , n22545 , n22546 );
buf ( n53532 , n53531 );
not ( n53533 , n48549 );
and ( n53534 , n53533 , n47430 );
xor ( n53535 , n48546 , n53534 );
not ( n22547 , n29614 );
and ( n22548 , n22547 , RI173a7ed8_1937);
and ( n22549 , n53535 , n29614 );
or ( n53536 , n22548 , n22549 );
not ( n22550 , RI1754c610_2);
and ( n22551 , n22550 , n53536 );
and ( n22552 , C0 , RI1754c610_2);
or ( n53537 , n22551 , n22552 );
buf ( n53538 , n53537 );
not ( n53539 , n41745 );
and ( n53540 , n53539 , n49524 );
xor ( n53541 , n41742 , n53540 );
not ( n22553 , n29614 );
and ( n22554 , n22553 , RI1748f610_1037);
and ( n22555 , n53541 , n29614 );
or ( n53542 , n22554 , n22555 );
not ( n22556 , RI1754c610_2);
and ( n22557 , n22556 , n53542 );
and ( n22558 , C0 , RI1754c610_2);
or ( n53543 , n22557 , n22558 );
buf ( n53544 , n53543 );
not ( n53545 , n41462 );
and ( n53546 , n53545 , n41480 );
xor ( n53547 , n45333 , n53546 );
not ( n22559 , n29614 );
and ( n22560 , n22559 , RI173c9c40_1772);
and ( n22561 , n53547 , n29614 );
or ( n53548 , n22560 , n22561 );
not ( n22562 , RI1754c610_2);
and ( n22563 , n22562 , n53548 );
and ( n22564 , C0 , RI1754c610_2);
or ( n53549 , n22563 , n22564 );
buf ( n53550 , n53549 );
not ( n53551 , n49021 );
and ( n53552 , n53551 , n41431 );
xor ( n53553 , n47050 , n53552 );
not ( n22565 , n29614 );
and ( n22566 , n22565 , RI17392ce0_2040);
and ( n22567 , n53553 , n29614 );
or ( n53554 , n22566 , n22567 );
not ( n22568 , RI1754c610_2);
and ( n22569 , n22568 , n53554 );
and ( n22570 , C0 , RI1754c610_2);
or ( n53555 , n22569 , n22570 );
buf ( n53556 , n53555 );
not ( n53557 , n46903 );
and ( n53558 , n53557 , n51794 );
xor ( n53559 , n45546 , n53558 );
not ( n22571 , n29614 );
and ( n22572 , n22571 , RI173eeaf8_1592);
and ( n22573 , n53559 , n29614 );
or ( n53560 , n22572 , n22573 );
not ( n22574 , RI1754c610_2);
and ( n22575 , n22574 , n53560 );
and ( n22576 , C0 , RI1754c610_2);
or ( n53561 , n22575 , n22576 );
buf ( n53562 , n53561 );
not ( n22577 , n34859 );
and ( n22578 , n22577 , C0 );
and ( n22579 , RI1754a978_63 , n34859 );
or ( n53563 , n22578 , n22579 );
not ( n22580 , RI19a22f70_2797);
and ( n22581 , n22580 , n53563 );
and ( n22582 , C0 , RI19a22f70_2797);
or ( n53564 , n22581 , n22582 );
not ( n22583 , n27683 );
and ( n22584 , n22583 , RI19aa40c0_2537);
and ( n22585 , n53564 , n27683 );
or ( n53565 , n22584 , n22585 );
not ( n22586 , RI1754c610_2);
and ( n22587 , n22586 , n53565 );
and ( n22588 , C0 , RI1754c610_2);
or ( n53566 , n22587 , n22588 );
buf ( n53567 , n53566 );
not ( n22589 , n27683 );
and ( n22590 , n22589 , RI19ace618_2222);
and ( n22591 , RI19a981f8_2625 , n27683 );
or ( n53568 , n22590 , n22591 );
not ( n22592 , RI1754c610_2);
and ( n22593 , n22592 , n53568 );
and ( n22594 , C0 , RI1754c610_2);
or ( n53569 , n22593 , n22594 );
buf ( n53570 , n53569 );
not ( n22595 , RI1754c610_2);
and ( n22596 , n22595 , RI19ad1588_2202);
and ( n22597 , C0 , RI1754c610_2);
or ( n53571 , n22596 , n22597 );
buf ( n53572 , n53571 );
not ( n22598 , n27683 );
and ( n22599 , n22598 , RI19a8b250_2717);
and ( n22600 , RI19a954f8_2645 , n27683 );
or ( n53573 , n22599 , n22600 );
not ( n22601 , RI1754c610_2);
and ( n22602 , n22601 , n53573 );
and ( n22603 , C0 , RI1754c610_2);
or ( n53574 , n22602 , n22603 );
buf ( n53575 , n53574 );
not ( n53576 , n52095 );
and ( n53577 , n53576 , n46851 );
xor ( n53578 , n53296 , n53577 );
not ( n22604 , n29614 );
and ( n22605 , n22604 , RI1740d728_1442);
and ( n22606 , n53578 , n29614 );
or ( n53579 , n22605 , n22606 );
not ( n22607 , RI1754c610_2);
and ( n22608 , n22607 , n53579 );
and ( n22609 , C0 , RI1754c610_2);
or ( n53580 , n22608 , n22609 );
buf ( n53581 , n53580 );
not ( n53582 , n49070 );
and ( n53583 , n53582 , n52503 );
xor ( n53584 , n49067 , n53583 );
not ( n22610 , n29614 );
and ( n22611 , n22610 , RI173df828_1666);
and ( n22612 , n53584 , n29614 );
or ( n53585 , n22611 , n22612 );
not ( n22613 , RI1754c610_2);
and ( n22614 , n22613 , n53585 );
and ( n22615 , C0 , RI1754c610_2);
or ( n53586 , n22614 , n22615 );
buf ( n53587 , n53586 );
not ( n53588 , n45873 );
and ( n53589 , n53588 , n45875 );
xor ( n53590 , n52337 , n53589 );
not ( n22616 , n29614 );
and ( n22617 , n22616 , RI175236c0_656);
and ( n22618 , n53590 , n29614 );
or ( n53591 , n22617 , n22618 );
not ( n22619 , RI1754c610_2);
and ( n22620 , n22619 , n53591 );
and ( n22621 , C0 , RI1754c610_2);
or ( n53592 , n22620 , n22621 );
buf ( n53593 , n53592 );
not ( n53594 , n52515 );
and ( n53595 , n53594 , n43872 );
xor ( n53596 , n44051 , n53595 );
not ( n22622 , n29614 );
and ( n22623 , n22622 , RI1750dd48_723);
and ( n22624 , n53596 , n29614 );
or ( n53597 , n22623 , n22624 );
not ( n22625 , RI1754c610_2);
and ( n22626 , n22625 , n53597 );
and ( n22627 , C0 , RI1754c610_2);
or ( n53598 , n22626 , n22627 );
buf ( n53599 , n53598 );
not ( n22628 , n27683 );
and ( n22629 , n22628 , RI19ac96e0_2259);
and ( n22630 , RI19a84950_2762 , n27683 );
or ( n53600 , n22629 , n22630 );
not ( n22631 , RI1754c610_2);
and ( n22632 , n22631 , n53600 );
and ( n22633 , C0 , RI1754c610_2);
or ( n53601 , n22632 , n22633 );
buf ( n53602 , n53601 );
not ( n53603 , n52879 );
and ( n53604 , n53603 , n49217 );
xor ( n53605 , n48173 , n53604 );
not ( n22634 , n29614 );
and ( n22635 , n22634 , RI174b2098_868);
and ( n22636 , n53605 , n29614 );
or ( n53606 , n22635 , n22636 );
not ( n22637 , RI1754c610_2);
and ( n22638 , n22637 , n53606 );
and ( n22639 , C0 , RI1754c610_2);
or ( n53607 , n22638 , n22639 );
buf ( n53608 , n53607 );
buf ( n53609 , RI174c86b8_787);
buf ( n53610 , RI1746dbf0_1201);
buf ( n53611 , RI17490678_1032);
not ( n22640 , n27683 );
and ( n22641 , n22640 , RI19ac0d88_2324);
and ( n22642 , RI19aca040_2255 , n27683 );
or ( n53612 , n22641 , n22642 );
not ( n22643 , RI1754c610_2);
and ( n22644 , n22643 , n53612 );
and ( n22645 , C0 , RI1754c610_2);
or ( n53613 , n22644 , n22645 );
buf ( n53614 , n53613 );
not ( n53615 , n36160 );
and ( n53616 , n53615 , n48640 );
xor ( n53617 , n36154 , n53616 );
not ( n22646 , n29614 );
and ( n22647 , n22646 , RI174aef60_883);
and ( n22648 , n53617 , n29614 );
or ( n53618 , n22647 , n22648 );
not ( n22649 , RI1754c610_2);
and ( n22650 , n22649 , n53618 );
and ( n22651 , C0 , RI1754c610_2);
or ( n53619 , n22650 , n22651 );
buf ( n53620 , n53619 );
not ( n53621 , n36402 );
and ( n53622 , n53621 , n51409 );
xor ( n53623 , n36383 , n53622 );
not ( n22652 , n29614 );
and ( n22653 , n22652 , RI17495880_1007);
and ( n22654 , n53623 , n29614 );
or ( n53624 , n22653 , n22654 );
not ( n22655 , RI1754c610_2);
and ( n22656 , n22655 , n53624 );
and ( n22657 , C0 , RI1754c610_2);
or ( n53625 , n22656 , n22657 );
buf ( n53626 , n53625 );
not ( n53627 , n46461 );
and ( n53628 , n53627 , n52286 );
xor ( n53629 , n44690 , n53628 );
not ( n22658 , n29614 );
and ( n22659 , n22658 , RI1739bd40_1996);
and ( n22660 , n53629 , n29614 );
or ( n53630 , n22659 , n22660 );
not ( n22661 , RI1754c610_2);
and ( n22662 , n22661 , n53630 );
and ( n22663 , C0 , RI1754c610_2);
or ( n53631 , n22662 , n22663 );
buf ( n53632 , n53631 );
not ( n53633 , n46678 );
and ( n53634 , n53633 , n45082 );
xor ( n53635 , n49716 , n53634 );
not ( n22664 , n29614 );
and ( n22665 , n22664 , RI174b4168_858);
and ( n22666 , n53635 , n29614 );
or ( n53636 , n22665 , n22666 );
not ( n22667 , RI1754c610_2);
and ( n22668 , n22667 , n53636 );
and ( n22669 , C0 , RI1754c610_2);
or ( n53637 , n22668 , n22669 );
buf ( n53638 , n53637 );
not ( n53639 , n46892 );
and ( n53640 , n53639 , n49362 );
xor ( n53641 , n46889 , n53640 );
not ( n22670 , n29614 );
and ( n22671 , n22670 , RI17408ef8_1464);
and ( n22672 , n53641 , n29614 );
or ( n53642 , n22671 , n22672 );
not ( n22673 , RI1754c610_2);
and ( n22674 , n22673 , n53642 );
and ( n22675 , C0 , RI1754c610_2);
or ( n53643 , n22674 , n22675 );
buf ( n53644 , n53643 );
and ( n53645 , RI1754b620_36 , n34844 );
and ( n53646 , RI1754b620_36 , n34847 );
and ( n53647 , RI1754b620_36 , n34850 );
or ( n53648 , n53645 , n53646 , n53647 , C0 , C0 , C0 , C0 , C0 );
not ( n22676 , n34859 );
and ( n22677 , n22676 , n53648 );
and ( n22678 , RI1754b620_36 , n34859 );
or ( n53649 , n22677 , n22678 );
not ( n22679 , RI19a22f70_2797);
and ( n22680 , n22679 , n53649 );
and ( n22681 , C0 , RI19a22f70_2797);
or ( n53650 , n22680 , n22681 );
not ( n22682 , n27683 );
and ( n22683 , n22682 , RI19ab2508_2437);
and ( n22684 , n53650 , n27683 );
or ( n53651 , n22683 , n22684 );
not ( n22685 , RI1754c610_2);
and ( n22686 , n22685 , n53651 );
and ( n22687 , C0 , RI1754c610_2);
or ( n53652 , n22686 , n22687 );
buf ( n53653 , n53652 );
and ( n53654 , RI1754bd28_21 , n34844 );
and ( n53655 , RI1754bd28_21 , n34847 );
and ( n53656 , RI1754bd28_21 , n34850 );
and ( n53657 , RI1754bd28_21 , n34852 );
and ( n53658 , RI1754bd28_21 , n34854 );
or ( n53659 , n53654 , n53655 , n53656 , n53657 , n53658 , C0 , C0 , C0 );
not ( n22688 , n34859 );
and ( n22689 , n22688 , n53659 );
and ( n22690 , RI1754bd28_21 , n34859 );
or ( n53660 , n22689 , n22690 );
not ( n22691 , RI19a22f70_2797);
and ( n22692 , n22691 , n53660 );
and ( n22693 , C0 , RI19a22f70_2797);
or ( n53661 , n22692 , n22693 );
not ( n22694 , n27683 );
and ( n22695 , n22694 , RI19a9b420_2603);
and ( n22696 , n53661 , n27683 );
or ( n53662 , n22695 , n22696 );
not ( n22697 , RI1754c610_2);
and ( n22698 , n22697 , n53662 );
and ( n22699 , C0 , RI1754c610_2);
or ( n53663 , n22698 , n22699 );
buf ( n53664 , n53663 );
buf ( n53665 , RI17509a40_736);
buf ( n53666 , RI1746ae00_1215);
buf ( n53667 , RI17485f20_1083);
not ( n53668 , n46212 );
and ( n53669 , n53668 , n41216 );
xor ( n53670 , n39066 , n53669 );
not ( n22700 , n29614 );
and ( n22701 , n22700 , RI17485bd8_1084);
and ( n22702 , n53670 , n29614 );
or ( n53671 , n22701 , n22702 );
not ( n22703 , RI1754c610_2);
and ( n22704 , n22703 , n53671 );
and ( n22705 , C0 , RI1754c610_2);
or ( n53672 , n22704 , n22705 );
buf ( n53673 , n53672 );
not ( n53674 , n52411 );
and ( n53675 , n53674 , n36885 );
xor ( n53676 , n51970 , n53675 );
not ( n22706 , n29614 );
and ( n22707 , n22706 , RI17344518_2108);
and ( n22708 , n53676 , n29614 );
or ( n53677 , n22707 , n22708 );
not ( n22709 , RI1754c610_2);
and ( n22710 , n22709 , n53677 );
and ( n22711 , C0 , RI1754c610_2);
or ( n53678 , n22710 , n22711 );
buf ( n53679 , n53678 );
not ( n53680 , n44040 );
and ( n53681 , n53680 , n39688 );
xor ( n53682 , n44037 , n53681 );
not ( n22712 , n29614 );
and ( n22713 , n22712 , RI17494188_1014);
and ( n22714 , n53682 , n29614 );
or ( n53683 , n22713 , n22714 );
not ( n22715 , RI1754c610_2);
and ( n22716 , n22715 , n53683 );
and ( n22717 , C0 , RI1754c610_2);
or ( n53684 , n22716 , n22717 );
buf ( n53685 , n53684 );
not ( n53686 , n50692 );
and ( n53687 , n53686 , n36210 );
xor ( n53688 , n42692 , n53687 );
not ( n22718 , n29614 );
and ( n22719 , n22718 , RI173dfeb8_1664);
and ( n22720 , n53688 , n29614 );
or ( n53689 , n22719 , n22720 );
not ( n22721 , RI1754c610_2);
and ( n22722 , n22721 , n53689 );
and ( n22723 , C0 , RI1754c610_2);
or ( n53690 , n22722 , n22723 );
buf ( n53691 , n53690 );
buf ( n53692 , RI175066b0_746);
buf ( n53693 , RI17469d98_1220);
buf ( n53694 , RI17487ff0_1073);
not ( n53695 , n51997 );
and ( n53696 , n53695 , n45922 );
xor ( n53697 , n47888 , n53696 );
not ( n22724 , n29614 );
and ( n22725 , n22724 , RI1751fe08_667);
and ( n22726 , n53697 , n29614 );
or ( n53698 , n22725 , n22726 );
not ( n22727 , RI1754c610_2);
and ( n22728 , n22727 , n53698 );
and ( n22729 , C0 , RI1754c610_2);
or ( n53699 , n22728 , n22729 );
buf ( n53700 , n53699 );
not ( n53701 , n50580 );
and ( n53702 , n53701 , n49028 );
xor ( n53703 , n47783 , n53702 );
not ( n22730 , n29614 );
and ( n22731 , n22730 , RI17464500_1247);
and ( n22732 , n53703 , n29614 );
or ( n53704 , n22731 , n22732 );
not ( n22733 , RI1754c610_2);
and ( n22734 , n22733 , n53704 );
and ( n22735 , C0 , RI1754c610_2);
or ( n53705 , n22734 , n22735 );
buf ( n53706 , n53705 );
not ( n22736 , n27683 );
and ( n22737 , n22736 , RI19ab63d8_2407);
and ( n22738 , RI19abf870_2336 , n27683 );
or ( n53707 , n22737 , n22738 );
not ( n22739 , RI1754c610_2);
and ( n22740 , n22739 , n53707 );
and ( n22741 , C0 , RI1754c610_2);
or ( n53708 , n22740 , n22741 );
buf ( n53709 , n53708 );
not ( n53710 , n43292 );
and ( n53711 , n53710 , n43294 );
xor ( n53712 , n47445 , n53711 );
not ( n22742 , n29614 );
and ( n22743 , n22742 , RI1749a0b0_985);
and ( n22744 , n53712 , n29614 );
or ( n53713 , n22743 , n22744 );
not ( n22745 , RI1754c610_2);
and ( n22746 , n22745 , n53713 );
and ( n22747 , C0 , RI1754c610_2);
or ( n53714 , n22746 , n22747 );
buf ( n53715 , n53714 );
not ( n53716 , n38794 );
and ( n53717 , n53716 , n38818 );
xor ( n53718 , n43141 , n53717 );
not ( n22748 , n29614 );
and ( n22749 , n22748 , RI17516da8_695);
and ( n22750 , n53718 , n29614 );
or ( n53719 , n22749 , n22750 );
not ( n22751 , RI1754c610_2);
and ( n22752 , n22751 , n53719 );
and ( n22753 , C0 , RI1754c610_2);
or ( n53720 , n22752 , n22753 );
buf ( n53721 , n53720 );
not ( n22754 , n27683 );
and ( n22755 , n22754 , RI19ac34e8_2304);
and ( n22756 , RI19acc3e0_2237 , n27683 );
or ( n53722 , n22755 , n22756 );
not ( n22757 , RI1754c610_2);
and ( n22758 , n22757 , n53722 );
and ( n22759 , C0 , RI1754c610_2);
or ( n53723 , n22758 , n22759 );
buf ( n53724 , n53723 );
not ( n53725 , n47659 );
and ( n53726 , n53725 , n45017 );
xor ( n53727 , n41153 , n53726 );
not ( n22760 , n29614 );
and ( n22761 , n22760 , RI17392998_2041);
and ( n22762 , n53727 , n29614 );
or ( n53728 , n22761 , n22762 );
not ( n22763 , RI1754c610_2);
and ( n22764 , n22763 , n53728 );
and ( n22765 , C0 , RI1754c610_2);
or ( n53729 , n22764 , n22765 );
buf ( n53730 , n53729 );
not ( n53731 , n42409 );
and ( n53732 , n53731 , n42411 );
xor ( n53733 , n46010 , n53732 );
or ( n53734 , RI17539830_589 , RI17539218_590);
or ( n53735 , n53734 , RI17537fd0_593);
or ( n53736 , n53735 , RI175379b8_594);
xor ( n53737 , n53733 , n53736 );
not ( n22766 , n29614 );
and ( n22767 , n22766 , RI1746f630_1193);
and ( n22768 , n53737 , n29614 );
or ( n53738 , n22767 , n22768 );
not ( n22769 , RI1754c610_2);
and ( n22770 , n22769 , n53738 );
and ( n22771 , C0 , RI1754c610_2);
or ( n53739 , n22770 , n22771 );
buf ( n53740 , n53739 );
not ( n22772 , n27683 );
and ( n22773 , n22772 , RI19acaf40_2248);
and ( n22774 , RI19a864f8_2750 , n27683 );
or ( n53741 , n22773 , n22774 );
not ( n22775 , RI1754c610_2);
and ( n22776 , n22775 , n53741 );
and ( n22777 , C0 , RI1754c610_2);
or ( n53742 , n22776 , n22777 );
buf ( n53743 , n53742 );
not ( n22778 , n27683 );
and ( n22779 , n22778 , RI19ac8768_2266);
and ( n22780 , RI19a83690_2770 , n27683 );
or ( n53744 , n22779 , n22780 );
not ( n22781 , RI1754c610_2);
and ( n22782 , n22781 , n53744 );
and ( n22783 , C0 , RI1754c610_2);
or ( n53745 , n22782 , n22783 );
buf ( n53746 , n53745 );
not ( n22784 , n27683 );
and ( n22785 , n22784 , RI19aa7888_2513);
and ( n22786 , RI19ab16f8_2443 , n27683 );
or ( n53747 , n22785 , n22786 );
not ( n22787 , RI1754c610_2);
and ( n22788 , n22787 , n53747 );
and ( n22789 , C0 , RI1754c610_2);
or ( n53748 , n22788 , n22789 );
buf ( n53749 , n53748 );
not ( n53750 , n46432 );
and ( n53751 , n53750 , n49234 );
xor ( n53752 , n46429 , n53751 );
not ( n22790 , n29614 );
and ( n22791 , n22790 , RI17497950_997);
and ( n22792 , n53752 , n29614 );
or ( n53753 , n22791 , n22792 );
not ( n22793 , RI1754c610_2);
and ( n22794 , n22793 , n53753 );
and ( n22795 , C0 , RI1754c610_2);
or ( n53754 , n22794 , n22795 );
buf ( n53755 , n53754 );
not ( n53756 , n51246 );
and ( n53757 , n53756 , n50822 );
xor ( n53758 , n41626 , n53757 );
not ( n22796 , n29614 );
and ( n22797 , n22796 , RI1748bb00_1055);
and ( n22798 , n53758 , n29614 );
or ( n53759 , n22797 , n22798 );
not ( n22799 , RI1754c610_2);
and ( n22800 , n22799 , n53759 );
and ( n22801 , C0 , RI1754c610_2);
or ( n53760 , n22800 , n22801 );
buf ( n53761 , n53760 );
and ( n53762 , RI1754b9e0_28 , n34844 );
and ( n53763 , RI1754b9e0_28 , n34847 );
and ( n53764 , RI1754b9e0_28 , n34850 );
and ( n53765 , RI1754b9e0_28 , n34852 );
or ( n53766 , n53762 , n53763 , n53764 , n53765 , C0 , C0 , C0 , C0 );
not ( n22802 , n34859 );
and ( n22803 , n22802 , n53766 );
and ( n22804 , RI1754b9e0_28 , n34859 );
or ( n53767 , n22803 , n22804 );
not ( n22805 , RI19a22f70_2797);
and ( n22806 , n22805 , n53767 );
and ( n22807 , C0 , RI19a22f70_2797);
or ( n53768 , n22806 , n22807 );
not ( n22808 , n27683 );
and ( n22809 , n22808 , RI19aa5a88_2525);
and ( n22810 , n53768 , n27683 );
or ( n53769 , n22809 , n22810 );
not ( n22811 , RI1754c610_2);
and ( n22812 , n22811 , n53769 );
and ( n22813 , C0 , RI1754c610_2);
or ( n53770 , n22812 , n22813 );
buf ( n53771 , n53770 );
not ( n53772 , n42589 );
and ( n53773 , n53772 , n42620 );
xor ( n53774 , n43613 , n53773 );
not ( n22814 , n29614 );
and ( n22815 , n22814 , RI1740b310_1453);
and ( n22816 , n53774 , n29614 );
or ( n53775 , n22815 , n22816 );
not ( n22817 , RI1754c610_2);
and ( n22818 , n22817 , n53775 );
and ( n22819 , C0 , RI1754c610_2);
or ( n53776 , n22818 , n22819 );
buf ( n53777 , n53776 );
not ( n53778 , n41820 );
and ( n53779 , n53778 , n42399 );
xor ( n53780 , n41801 , n53779 );
not ( n22820 , n29614 );
and ( n22821 , n22820 , RI173e4058_1644);
and ( n22822 , n53780 , n29614 );
or ( n53781 , n22821 , n22822 );
not ( n22823 , RI1754c610_2);
and ( n22824 , n22823 , n53781 );
and ( n22825 , C0 , RI1754c610_2);
or ( n53782 , n22824 , n22825 );
buf ( n53783 , n53782 );
and ( n53784 , RI1754bb48_25 , n34844 );
and ( n53785 , RI1754bb48_25 , n34847 );
and ( n53786 , RI1754bb48_25 , n34850 );
and ( n53787 , RI1754bb48_25 , n34852 );
and ( n53788 , RI1754bb48_25 , n34854 );
or ( n53789 , n53784 , n53785 , n53786 , n53787 , n53788 , C0 , C0 , C0 );
not ( n22826 , n34859 );
and ( n22827 , n22826 , n53789 );
and ( n22828 , RI1754bb48_25 , n34859 );
or ( n53790 , n22827 , n22828 );
not ( n22829 , RI19a22f70_2797);
and ( n22830 , n22829 , n53790 );
and ( n22831 , C0 , RI19a22f70_2797);
or ( n53791 , n22830 , n22831 );
not ( n22832 , n27683 );
and ( n22833 , n22832 , RI19aa12d0_2559);
and ( n22834 , n53791 , n27683 );
or ( n53792 , n22833 , n22834 );
not ( n22835 , RI1754c610_2);
and ( n22836 , n22835 , n53792 );
and ( n22837 , C0 , RI1754c610_2);
or ( n53793 , n22836 , n22837 );
buf ( n53794 , n53793 );
not ( n53795 , n47694 );
and ( n53796 , n53795 , n46978 );
xor ( n53797 , n48296 , n53796 );
not ( n22838 , n29614 );
and ( n22839 , n22838 , RI174ab450_901);
and ( n22840 , n53797 , n29614 );
or ( n53798 , n22839 , n22840 );
not ( n22841 , RI1754c610_2);
and ( n22842 , n22841 , n53798 );
and ( n22843 , C0 , RI1754c610_2);
or ( n53799 , n22842 , n22843 );
buf ( n53800 , n53799 );
not ( n53801 , n46008 );
and ( n53802 , n53801 , n46010 );
xor ( n53803 , n42414 , n53802 );
not ( n22844 , n29614 );
and ( n22845 , n22844 , RI1749b118_980);
and ( n22846 , n53803 , n29614 );
or ( n53804 , n22845 , n22846 );
not ( n22847 , RI1754c610_2);
and ( n22848 , n22847 , n53804 );
and ( n22849 , C0 , RI1754c610_2);
or ( n53805 , n22848 , n22849 );
buf ( n53806 , n53805 );
buf ( n53807 , RI17512fc8_707);
buf ( n53808 , RI17480340_1111);
not ( n53809 , n50240 );
and ( n53810 , n53809 , n42468 );
xor ( n53811 , n49596 , n53810 );
not ( n22850 , n29614 );
and ( n22851 , n22850 , RI175134f0_706);
and ( n22852 , n53811 , n29614 );
or ( n53812 , n22851 , n22852 );
not ( n22853 , RI1754c610_2);
and ( n22854 , n22853 , n53812 );
and ( n22855 , C0 , RI1754c610_2);
or ( n53813 , n22854 , n22855 );
buf ( n53814 , n53813 );
not ( n53815 , n48612 );
and ( n53816 , n53815 , n46812 );
xor ( n53817 , n50812 , n53816 );
not ( n22856 , n29614 );
and ( n22857 , n22856 , RI173f53f8_1560);
and ( n22858 , n53817 , n29614 );
or ( n53818 , n22857 , n22858 );
not ( n22859 , RI1754c610_2);
and ( n22860 , n22859 , n53818 );
and ( n22861 , C0 , RI1754c610_2);
or ( n53819 , n22860 , n22861 );
buf ( n53820 , n53819 );
not ( n53821 , n43188 );
and ( n53822 , n53821 , n45679 );
xor ( n53823 , n40587 , n53822 );
not ( n22862 , n29614 );
and ( n22863 , n22862 , RI1747a418_1140);
and ( n22864 , n53823 , n29614 );
or ( n53824 , n22863 , n22864 );
not ( n22865 , RI1754c610_2);
and ( n22866 , n22865 , n53824 );
and ( n22867 , C0 , RI1754c610_2);
or ( n53825 , n22866 , n22867 );
buf ( n53826 , n53825 );
buf ( n53827 , RI19a240c8_2788);
not ( n22868 , n34859 );
and ( n22869 , n22868 , n53827 );
and ( n22870 , RI1754ab58_59 , n34859 );
or ( n53828 , n22869 , n22870 );
not ( n22871 , RI19a22f70_2797);
and ( n22872 , n22871 , n53828 );
and ( n22873 , RI19a240c8_2788 , RI19a22f70_2797);
or ( n53829 , n22872 , n22873 );
not ( n22874 , n27683 );
and ( n22875 , n22874 , RI19a85508_2757);
and ( n22876 , n53829 , n27683 );
or ( n53830 , n22875 , n22876 );
not ( n22877 , RI1754c610_2);
and ( n22878 , n22877 , n53830 );
and ( n22879 , C0 , RI1754c610_2);
or ( n53831 , n22878 , n22879 );
buf ( n53832 , n53831 );
not ( n53833 , n47515 );
and ( n53834 , n53833 , n41837 );
xor ( n53835 , n47512 , n53834 );
not ( n22880 , n29614 );
and ( n22881 , n22880 , RI174a1d60_947);
and ( n22882 , n53835 , n29614 );
or ( n53836 , n22881 , n22882 );
not ( n22883 , RI1754c610_2);
and ( n22884 , n22883 , n53836 );
and ( n22885 , C0 , RI1754c610_2);
or ( n53837 , n22884 , n22885 );
buf ( n53838 , n53837 );
not ( n53839 , n38726 );
and ( n53840 , n53839 , n50967 );
xor ( n53841 , n38683 , n53840 );
not ( n22886 , n29614 );
and ( n22887 , n22886 , RI174a9380_911);
and ( n22888 , n53841 , n29614 );
or ( n53842 , n22887 , n22888 );
not ( n22889 , RI1754c610_2);
and ( n22890 , n22889 , n53842 );
and ( n22891 , C0 , RI1754c610_2);
or ( n53843 , n22890 , n22891 );
buf ( n53844 , n53843 );
not ( n53845 , n40968 );
and ( n53846 , n53845 , n50163 );
xor ( n53847 , n40952 , n53846 );
not ( n22892 , n29614 );
and ( n22893 , n22892 , RI173a1c68_1967);
and ( n22894 , n53847 , n29614 );
or ( n53848 , n22893 , n22894 );
not ( n22895 , RI1754c610_2);
and ( n22896 , n22895 , n53848 );
and ( n22897 , C0 , RI1754c610_2);
or ( n53849 , n22896 , n22897 );
buf ( n53850 , n53849 );
not ( n53851 , n44408 );
and ( n53852 , n53851 , n44410 );
xor ( n53853 , n41171 , n53852 );
not ( n22898 , n29614 );
and ( n22899 , n22898 , RI173d7830_1705);
and ( n22900 , n53853 , n29614 );
or ( n53854 , n22899 , n22900 );
not ( n22901 , RI1754c610_2);
and ( n22902 , n22901 , n53854 );
and ( n22903 , C0 , RI1754c610_2);
or ( n53855 , n22902 , n22903 );
buf ( n53856 , n53855 );
not ( n53857 , n42468 );
and ( n53858 , n53857 , n42470 );
xor ( n53859 , n50240 , n53858 );
not ( n22904 , n29614 );
and ( n22905 , n22904 , RI17529de0_636);
and ( n22906 , n53859 , n29614 );
or ( n53860 , n22905 , n22906 );
not ( n22907 , RI1754c610_2);
and ( n22908 , n22907 , n53860 );
and ( n22909 , C0 , RI1754c610_2);
or ( n53861 , n22908 , n22909 );
buf ( n53862 , n53861 );
not ( n53863 , n49497 );
and ( n53864 , n53863 , n50135 );
xor ( n53865 , n49494 , n53864 );
not ( n22910 , n29614 );
and ( n22911 , n22910 , RI1739c088_1995);
and ( n22912 , n53865 , n29614 );
or ( n53866 , n22911 , n22912 );
not ( n22913 , RI1754c610_2);
and ( n22914 , n22913 , n53866 );
and ( n22915 , C0 , RI1754c610_2);
or ( n53867 , n22914 , n22915 );
buf ( n53868 , n53867 );
not ( n53869 , n47247 );
and ( n53870 , n53869 , n45789 );
xor ( n53871 , n50541 , n53870 );
not ( n22916 , n29614 );
and ( n22917 , n22916 , RI1738fba8_2055);
and ( n22918 , n53871 , n29614 );
or ( n53872 , n22917 , n22918 );
not ( n22919 , RI1754c610_2);
and ( n22920 , n22919 , n53872 );
and ( n22921 , C0 , RI1754c610_2);
or ( n53873 , n22920 , n22921 );
buf ( n53874 , n53873 );
not ( n53875 , n45699 );
and ( n53876 , n53875 , n36412 );
xor ( n53877 , n45095 , n53876 );
not ( n22922 , n29614 );
and ( n22923 , n22922 , RI174c5d78_795);
and ( n22924 , n53877 , n29614 );
or ( n53878 , n22923 , n22924 );
not ( n22925 , RI1754c610_2);
and ( n22926 , n22925 , n53878 );
and ( n22927 , C0 , RI1754c610_2);
or ( n53879 , n22926 , n22927 );
buf ( n53880 , n53879 );
not ( n53881 , n41400 );
and ( n53882 , n53881 , n41402 );
xor ( n53883 , n52596 , n53882 );
not ( n22928 , n29614 );
and ( n22929 , n22928 , RI17472420_1179);
and ( n22930 , n53883 , n29614 );
or ( n53884 , n22929 , n22930 );
not ( n22931 , RI1754c610_2);
and ( n22932 , n22931 , n53884 );
and ( n22933 , C0 , RI1754c610_2);
or ( n53885 , n22932 , n22933 );
buf ( n53886 , n53885 );
not ( n22934 , n27683 );
and ( n22935 , n22934 , RI19ac4910_2295);
and ( n22936 , RI19acd5b0_2229 , n27683 );
or ( n53887 , n22935 , n22936 );
not ( n22937 , RI1754c610_2);
and ( n22938 , n22937 , n53887 );
and ( n22939 , C0 , RI1754c610_2);
or ( n53888 , n22938 , n22939 );
buf ( n53889 , n53888 );
not ( n53890 , n45755 );
and ( n53891 , n53890 , n43397 );
xor ( n53892 , n45752 , n53891 );
not ( n22940 , n29614 );
and ( n22941 , n22940 , RI174ca5a8_781);
and ( n22942 , n53892 , n29614 );
or ( n53893 , n22941 , n22942 );
not ( n22943 , RI1754c610_2);
and ( n22944 , n22943 , n53893 );
and ( n22945 , C0 , RI1754c610_2);
or ( n53894 , n22944 , n22945 );
buf ( n53895 , n53894 );
not ( n22946 , n27683 );
and ( n22947 , n22946 , RI19ab4038_2423);
and ( n22948 , RI19abd9f8_2353 , n27683 );
or ( n53896 , n22947 , n22948 );
not ( n22949 , RI1754c610_2);
and ( n22950 , n22949 , n53896 );
and ( n22951 , C0 , RI1754c610_2);
or ( n53897 , n22950 , n22951 );
buf ( n53898 , n53897 );
not ( n53899 , n46877 );
and ( n53900 , n53899 , n44983 );
xor ( n53901 , n49340 , n53900 );
not ( n22952 , n29614 );
and ( n22953 , n22952 , RI1747e270_1121);
and ( n22954 , n53901 , n29614 );
or ( n53902 , n22953 , n22954 );
not ( n22955 , RI1754c610_2);
and ( n22956 , n22955 , n53902 );
and ( n22957 , C0 , RI1754c610_2);
or ( n53903 , n22956 , n22957 );
buf ( n53904 , n53903 );
not ( n53905 , n43219 );
and ( n53906 , n53905 , n38845 );
xor ( n53907 , n45982 , n53906 );
not ( n22958 , n29614 );
and ( n22959 , n22958 , RI173ceb00_1748);
and ( n22960 , n53907 , n29614 );
or ( n53908 , n22959 , n22960 );
not ( n22961 , RI1754c610_2);
and ( n22962 , n22961 , n53908 );
and ( n22963 , C0 , RI1754c610_2);
or ( n53909 , n22962 , n22963 );
buf ( n53910 , n53909 );
not ( n53911 , n42898 );
and ( n53912 , n53911 , n42900 );
xor ( n53913 , n46557 , n53912 );
not ( n22964 , n29614 );
and ( n22965 , n22964 , RI1733df60_2139);
and ( n22966 , n53913 , n29614 );
or ( n53914 , n22965 , n22966 );
not ( n22967 , RI1754c610_2);
and ( n22968 , n22967 , n53914 );
and ( n22969 , C0 , RI1754c610_2);
or ( n53915 , n22968 , n22969 );
buf ( n53916 , n53915 );
not ( n53917 , n50052 );
and ( n53918 , n53917 , n50054 );
xor ( n53919 , n50231 , n53918 );
not ( n22970 , n29614 );
and ( n22971 , n22970 , RI175038c0_749);
and ( n22972 , n53919 , n29614 );
or ( n53920 , n22971 , n22972 );
not ( n22973 , RI1754c610_2);
and ( n22974 , n22973 , n53920 );
and ( n22975 , C0 , RI1754c610_2);
or ( n53921 , n22974 , n22975 );
buf ( n53922 , n53921 );
not ( n53923 , n43297 );
and ( n53924 , n53923 , n47442 );
xor ( n53925 , n43294 , n53924 );
not ( n22976 , n29614 );
and ( n22977 , n22976 , RI1746e280_1199);
and ( n22978 , n53925 , n29614 );
or ( n53926 , n22977 , n22978 );
not ( n22979 , RI1754c610_2);
and ( n22980 , n22979 , n53926 );
and ( n22981 , C0 , RI1754c610_2);
or ( n53927 , n22980 , n22981 );
buf ( n53928 , n53927 );
not ( n22982 , n27683 );
and ( n22983 , n22982 , RI19a99f80_2612);
and ( n22984 , RI19aa3580_2542 , n27683 );
or ( n53929 , n22983 , n22984 );
not ( n22985 , RI1754c610_2);
and ( n22986 , n22985 , n53929 );
and ( n22987 , C0 , RI1754c610_2);
or ( n53930 , n22986 , n22987 );
buf ( n53931 , n53930 );
not ( n22988 , n27683 );
and ( n22989 , n22988 , RI19a93ba8_2656);
and ( n22990 , RI19a9de50_2585 , n27683 );
or ( n53932 , n22989 , n22990 );
not ( n22991 , RI1754c610_2);
and ( n22992 , n22991 , n53932 );
and ( n22993 , C0 , RI1754c610_2);
or ( n53933 , n22992 , n22993 );
buf ( n53934 , n53933 );
not ( n53935 , n45612 );
and ( n53936 , n53935 , n45614 );
xor ( n53937 , n48748 , n53936 );
not ( n22994 , n29614 );
and ( n22995 , n22994 , RI17474838_1168);
and ( n22996 , n53937 , n29614 );
or ( n53938 , n22995 , n22996 );
not ( n22997 , RI1754c610_2);
and ( n22998 , n22997 , n53938 );
and ( n22999 , C0 , RI1754c610_2);
or ( n53939 , n22998 , n22999 );
buf ( n53940 , n53939 );
not ( n23000 , n27683 );
and ( n23001 , n23000 , RI19aac040_2482);
and ( n23002 , RI19ab5d48_2410 , n27683 );
or ( n53941 , n23001 , n23002 );
not ( n23003 , RI1754c610_2);
and ( n23004 , n23003 , n53941 );
and ( n23005 , C0 , RI1754c610_2);
or ( n53942 , n23004 , n23005 );
buf ( n53943 , n53942 );
not ( n53944 , n44706 );
and ( n53945 , n53944 , n46093 );
xor ( n53946 , n42510 , n53945 );
not ( n23006 , n29614 );
and ( n23007 , n23006 , RI173da620_1691);
and ( n23008 , n53946 , n29614 );
or ( n53947 , n23007 , n23008 );
not ( n23009 , RI1754c610_2);
and ( n23010 , n23009 , n53947 );
and ( n23011 , C0 , RI1754c610_2);
or ( n53948 , n23010 , n23011 );
buf ( n53949 , n53948 );
not ( n53950 , n47076 );
and ( n53951 , n53950 , n52892 );
xor ( n53952 , n46632 , n53951 );
not ( n23012 , n29614 );
and ( n23013 , n23012 , RI17454ee8_1322);
and ( n23014 , n53952 , n29614 );
or ( n53953 , n23013 , n23014 );
not ( n23015 , RI1754c610_2);
and ( n23016 , n23015 , n53953 );
and ( n23017 , C0 , RI1754c610_2);
or ( n53954 , n23016 , n23017 );
buf ( n53955 , n53954 );
xor ( n53956 , n32335 , n41316 );
xor ( n53957 , n53956 , n35622 );
not ( n53958 , n53957 );
and ( n53959 , n53958 , n44115 );
xor ( n53960 , n42240 , n53959 );
not ( n23018 , n29614 );
and ( n23019 , n23018 , RI174a68d8_924);
and ( n23020 , n53960 , n29614 );
or ( n53961 , n23019 , n23020 );
not ( n23021 , RI1754c610_2);
and ( n23022 , n23021 , n53961 );
and ( n23023 , C0 , RI1754c610_2);
or ( n53962 , n23022 , n23023 );
buf ( n53963 , n53962 );
not ( n53964 , n48446 );
and ( n53965 , n53964 , n48448 );
xor ( n53966 , n49772 , n53965 );
not ( n23024 , n29614 );
and ( n23025 , n23024 , RI1745dc00_1279);
and ( n23026 , n53966 , n29614 );
or ( n53967 , n23025 , n23026 );
not ( n23027 , RI1754c610_2);
and ( n23028 , n23027 , n53967 );
and ( n23029 , C0 , RI1754c610_2);
or ( n53968 , n23028 , n23029 );
buf ( n53969 , n53968 );
not ( n53970 , n43957 );
and ( n53971 , n53970 , n43959 );
xor ( n53972 , n46104 , n53971 );
not ( n23030 , n29614 );
and ( n23031 , n23030 , RI174cd938_771);
and ( n23032 , n53972 , n29614 );
or ( n53973 , n23031 , n23032 );
not ( n23033 , RI1754c610_2);
and ( n23034 , n23033 , n53973 );
and ( n23035 , C0 , RI1754c610_2);
or ( n53974 , n23034 , n23035 );
buf ( n53975 , n53974 );
not ( n53976 , n52892 );
and ( n53977 , n53976 , n46627 );
xor ( n53978 , n47076 , n53977 );
not ( n23036 , n29614 );
and ( n23037 , n23036 , RI1747c4e8_1130);
and ( n23038 , n53978 , n29614 );
or ( n53979 , n23037 , n23038 );
not ( n23039 , RI1754c610_2);
and ( n23040 , n23039 , n53979 );
and ( n23041 , C0 , RI1754c610_2);
or ( n53980 , n23040 , n23041 );
buf ( n53981 , n53980 );
and ( n53982 , RI1754abd0_58 , n34844 );
buf ( n53983 , n34847 );
or ( n53984 , n53982 , n53983 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n23042 , n34859 );
and ( n23043 , n23042 , n53984 );
and ( n23044 , RI1754abd0_58 , n34859 );
or ( n53985 , n23043 , n23044 );
not ( n23045 , RI19a22f70_2797);
and ( n23046 , n23045 , n53985 );
and ( n23047 , C0 , RI19a22f70_2797);
or ( n53986 , n23046 , n23047 );
not ( n23048 , n27683 );
and ( n23049 , n23048 , RI19a83b40_2768);
and ( n23050 , n53986 , n27683 );
or ( n53987 , n23049 , n23050 );
not ( n23051 , RI1754c610_2);
and ( n23052 , n23051 , n53987 );
and ( n23053 , C0 , RI1754c610_2);
or ( n53988 , n23052 , n23053 );
buf ( n53989 , n53988 );
not ( n53990 , n44729 );
and ( n53991 , n53990 , n44731 );
xor ( n53992 , n42793 , n53991 );
not ( n23054 , n29614 );
and ( n23055 , n23054 , RI173c5de8_1791);
and ( n23056 , n53992 , n29614 );
or ( n53993 , n23055 , n23056 );
not ( n23057 , RI1754c610_2);
and ( n23058 , n23057 , n53993 );
and ( n23059 , C0 , RI1754c610_2);
or ( n53994 , n23058 , n23059 );
buf ( n53995 , n53994 );
not ( n53996 , n49890 );
and ( n53997 , n53996 , n40524 );
xor ( n53998 , n42310 , n53997 );
not ( n23060 , n29614 );
and ( n23061 , n23060 , RI17344ef0_2105);
and ( n23062 , n53998 , n29614 );
or ( n53999 , n23061 , n23062 );
not ( n23063 , RI1754c610_2);
and ( n23064 , n23063 , n53999 );
and ( n23065 , C0 , RI1754c610_2);
or ( n54000 , n23064 , n23065 );
buf ( n54001 , n54000 );
buf ( n54002 , RI1749f2b8_960);
buf ( n54003 , RI174b3e20_859);
not ( n54004 , n48799 );
and ( n54005 , n54004 , n48801 );
xor ( n54006 , n51582 , n54005 );
not ( n23066 , n29614 );
and ( n23067 , n23066 , RI173c95b0_1774);
and ( n23068 , n54006 , n29614 );
or ( n54007 , n23067 , n23068 );
not ( n23069 , RI1754c610_2);
and ( n23070 , n23069 , n54007 );
and ( n23071 , C0 , RI1754c610_2);
or ( n54008 , n23070 , n23071 );
buf ( n54009 , n54008 );
buf ( n54010 , RI174741a8_1170);
not ( n54011 , n49961 );
and ( n54012 , n54011 , n49963 );
xor ( n54013 , n50007 , n54012 );
not ( n23072 , n29614 );
and ( n23073 , n23072 , RI173eee40_1591);
and ( n23074 , n54013 , n29614 );
or ( n54014 , n23073 , n23074 );
not ( n23075 , RI1754c610_2);
and ( n23076 , n23075 , n54014 );
and ( n23077 , C0 , RI1754c610_2);
or ( n54015 , n23076 , n23077 );
buf ( n54016 , n54015 );
and ( n54017 , RI1754b2d8_43 , n34844 );
and ( n54018 , RI1754b2d8_43 , n34847 );
or ( n54019 , n54017 , n54018 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n23078 , n34859 );
and ( n23079 , n23078 , n54019 );
and ( n23080 , RI1754b2d8_43 , n34859 );
or ( n54020 , n23079 , n23080 );
not ( n23081 , RI19a22f70_2797);
and ( n23082 , n23081 , n54020 );
and ( n23083 , C0 , RI19a22f70_2797);
or ( n54021 , n23082 , n23083 );
not ( n23084 , n27683 );
and ( n23085 , n23084 , RI19abcfa8_2359);
and ( n23086 , n54021 , n27683 );
or ( n54022 , n23085 , n23086 );
not ( n23087 , RI1754c610_2);
and ( n23088 , n23087 , n54022 );
and ( n23089 , C0 , RI1754c610_2);
or ( n54023 , n23088 , n23089 );
buf ( n54024 , n54023 );
not ( n23090 , n27683 );
and ( n23091 , n23090 , RI19a9d1a8_2590);
and ( n23092 , RI19aa6988_2519 , n27683 );
or ( n54025 , n23091 , n23092 );
not ( n23093 , RI1754c610_2);
and ( n23094 , n23093 , n54025 );
and ( n23095 , C0 , RI1754c610_2);
or ( n54026 , n23094 , n23095 );
buf ( n54027 , n54026 );
not ( n23096 , n27683 );
and ( n23097 , n23096 , RI19abc8a0_2363);
and ( n23098 , RI19ac5108_2291 , n27683 );
or ( n54028 , n23097 , n23098 );
not ( n23099 , RI1754c610_2);
and ( n23100 , n23099 , n54028 );
and ( n23101 , C0 , RI1754c610_2);
or ( n54029 , n23100 , n23101 );
buf ( n54030 , n54029 );
not ( n54031 , n49427 );
and ( n54032 , n54031 , n51684 );
xor ( n54033 , n49424 , n54032 );
not ( n23102 , n29614 );
and ( n23103 , n23102 , RI174996d8_988);
and ( n23104 , n54033 , n29614 );
or ( n54034 , n23103 , n23104 );
not ( n23105 , RI1754c610_2);
and ( n23106 , n23105 , n54034 );
and ( n23107 , C0 , RI1754c610_2);
or ( n54035 , n23106 , n23107 );
buf ( n54036 , n54035 );
buf ( n54037 , RI174c00a8_813);
not ( n54038 , n46528 );
and ( n54039 , n54038 , n51636 );
xor ( n54040 , n46525 , n54039 );
not ( n23108 , n29614 );
and ( n23109 , n23108 , RI17450d48_1342);
and ( n23110 , n54040 , n29614 );
or ( n54041 , n23109 , n23110 );
not ( n23111 , RI1754c610_2);
and ( n23112 , n23111 , n54041 );
and ( n23113 , C0 , RI1754c610_2);
or ( n54042 , n23112 , n23113 );
buf ( n54043 , n54042 );
buf ( n54044 , RI17495f10_1005);
not ( n54045 , n47850 );
and ( n54046 , n54045 , n47852 );
xor ( n54047 , n52126 , n54046 );
not ( n23114 , n29614 );
and ( n23115 , n23114 , RI1739c3d0_1994);
and ( n23116 , n54047 , n29614 );
or ( n54048 , n23115 , n23116 );
not ( n23117 , RI1754c610_2);
and ( n23118 , n23117 , n54048 );
and ( n23119 , C0 , RI1754c610_2);
or ( n54049 , n23118 , n23119 );
buf ( n54050 , n54049 );
not ( n54051 , n46658 );
and ( n54052 , n54051 , n46660 );
xor ( n54053 , n52253 , n54052 );
not ( n23120 , n29614 );
and ( n23121 , n23120 , RI173908c8_2051);
and ( n23122 , n54053 , n29614 );
or ( n54054 , n23121 , n23122 );
not ( n23123 , RI1754c610_2);
and ( n23124 , n23123 , n54054 );
and ( n23125 , C0 , RI1754c610_2);
or ( n54055 , n23124 , n23125 );
buf ( n54056 , n54055 );
not ( n54057 , n48911 );
and ( n54058 , n54057 , n48913 );
xor ( n54059 , n51238 , n54058 );
not ( n23126 , n29614 );
and ( n23127 , n23126 , RI173eb330_1609);
and ( n23128 , n54059 , n29614 );
or ( n54060 , n23127 , n23128 );
not ( n23129 , RI1754c610_2);
and ( n23130 , n23129 , n54060 );
and ( n23131 , C0 , RI1754c610_2);
or ( n54061 , n23130 , n23131 );
buf ( n54062 , n54061 );
not ( n23132 , n27683 );
and ( n23133 , n23132 , RI19ab7a58_2397);
and ( n23134 , RI19ac0860_2327 , n27683 );
or ( n54063 , n23133 , n23134 );
not ( n23135 , RI1754c610_2);
and ( n23136 , n23135 , n54063 );
and ( n23137 , C0 , RI1754c610_2);
or ( n54064 , n23136 , n23137 );
buf ( n54065 , n54064 );
not ( n23138 , n27683 );
and ( n23139 , n23138 , RI19a92528_2666);
and ( n23140 , RI19a9c5f0_2595 , n27683 );
or ( n54066 , n23139 , n23140 );
not ( n23141 , RI1754c610_2);
and ( n23142 , n23141 , n54066 );
and ( n23143 , C0 , RI1754c610_2);
or ( n54067 , n23142 , n23143 );
buf ( n54068 , n54067 );
not ( n54069 , n39821 );
and ( n54070 , n54069 , n47959 );
xor ( n54071 , n39818 , n54070 );
not ( n23144 , n29614 );
and ( n23145 , n23144 , RI174025f8_1496);
and ( n23146 , n54071 , n29614 );
or ( n54072 , n23145 , n23146 );
not ( n23147 , RI1754c610_2);
and ( n23148 , n23147 , n54072 );
and ( n23149 , C0 , RI1754c610_2);
or ( n54073 , n23148 , n23149 );
buf ( n54074 , n54073 );
not ( n54075 , n41547 );
and ( n54076 , n54075 , n52112 );
xor ( n54077 , n41544 , n54076 );
not ( n23150 , n29614 );
and ( n23151 , n23150 , RI1745be78_1288);
and ( n23152 , n54077 , n29614 );
or ( n54078 , n23151 , n23152 );
not ( n23153 , RI1754c610_2);
and ( n23154 , n23153 , n54078 );
and ( n23155 , C0 , RI1754c610_2);
or ( n54079 , n23154 , n23155 );
buf ( n54080 , n54079 );
not ( n54081 , n46648 );
and ( n54082 , n54081 , n42520 );
xor ( n54083 , n46645 , n54082 );
not ( n23156 , n29614 );
and ( n23157 , n23156 , RI173d43b0_1721);
and ( n23158 , n54083 , n29614 );
or ( n54084 , n23157 , n23158 );
not ( n23159 , RI1754c610_2);
and ( n23160 , n23159 , n54084 );
and ( n23161 , C0 , RI1754c610_2);
or ( n54085 , n23160 , n23161 );
buf ( n54086 , n54085 );
not ( n54087 , n52568 );
and ( n54088 , n54087 , n48950 );
xor ( n54089 , n49447 , n54088 );
not ( n23162 , n29614 );
and ( n23163 , n23162 , RI1745efb0_1273);
and ( n23164 , n54089 , n29614 );
or ( n54090 , n23163 , n23164 );
not ( n23165 , RI1754c610_2);
and ( n23166 , n23165 , n54090 );
and ( n23167 , C0 , RI1754c610_2);
or ( n54091 , n23166 , n23167 );
buf ( n54092 , n54091 );
not ( n23168 , n27683 );
and ( n23169 , n23168 , RI19aa4ed0_2530);
and ( n23170 , RI19aaf268_2460 , n27683 );
or ( n54093 , n23169 , n23170 );
not ( n23171 , RI1754c610_2);
and ( n23172 , n23171 , n54093 );
and ( n23173 , C0 , RI1754c610_2);
or ( n54094 , n23172 , n23173 );
buf ( n54095 , n54094 );
not ( n54096 , n46566 );
and ( n54097 , n54096 , n50742 );
xor ( n54098 , n45534 , n54097 );
not ( n23174 , n29614 );
and ( n23175 , n23174 , RI173dc060_1683);
and ( n23176 , n54098 , n29614 );
or ( n54099 , n23175 , n23176 );
not ( n23177 , RI1754c610_2);
and ( n23178 , n23177 , n54099 );
and ( n23179 , C0 , RI1754c610_2);
or ( n54100 , n23178 , n23179 );
buf ( n54101 , n54100 );
xor ( n54102 , n38057 , n40091 );
xor ( n54103 , n54102 , n40111 );
not ( n54104 , n49561 );
and ( n54105 , n54104 , n49563 );
xor ( n54106 , n54103 , n54105 );
not ( n23180 , n29614 );
and ( n23181 , n23180 , RI174ac800_895);
and ( n23182 , n54106 , n29614 );
or ( n54107 , n23181 , n23182 );
not ( n23183 , RI1754c610_2);
and ( n23184 , n23183 , n54107 );
and ( n23185 , C0 , RI1754c610_2);
or ( n54108 , n23184 , n23185 );
buf ( n54109 , n54108 );
not ( n54110 , n40438 );
and ( n54111 , n54110 , n45141 );
xor ( n54112 , n40392 , n54111 );
not ( n23186 , n29614 );
and ( n23187 , n23186 , RI1751a138_685);
and ( n23188 , n54112 , n29614 );
or ( n54113 , n23187 , n23188 );
not ( n23189 , RI1754c610_2);
and ( n23190 , n23189 , n54113 );
and ( n23191 , C0 , RI1754c610_2);
or ( n54114 , n23190 , n23191 );
buf ( n54115 , n54114 );
not ( n54116 , n46542 );
and ( n54117 , n54116 , n46557 );
xor ( n54118 , n42903 , n54117 );
not ( n23192 , n29614 );
and ( n23193 , n23192 , RI173aa2f0_1926);
and ( n23194 , n54118 , n29614 );
or ( n54119 , n23193 , n23194 );
not ( n23195 , RI1754c610_2);
and ( n23196 , n23195 , n54119 );
and ( n23197 , C0 , RI1754c610_2);
or ( n54120 , n23196 , n23197 );
buf ( n54121 , n54120 );
and ( n54122 , RI1754c598_3 , n34844 );
and ( n54123 , RI1754c598_3 , n34847 );
and ( n54124 , RI1754c598_3 , n34850 );
and ( n54125 , RI1754c598_3 , n34852 );
and ( n54126 , RI1754c598_3 , n34854 );
and ( n54127 , RI1754c598_3 , n34856 );
and ( n54128 , RI1754c598_3 , n39233 );
or ( n54129 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , C0 );
not ( n23198 , n34859 );
and ( n23199 , n23198 , n54129 );
and ( n23200 , RI1754c598_3 , n34859 );
or ( n54130 , n23199 , n23200 );
not ( n23201 , RI19a22f70_2797);
and ( n23202 , n23201 , n54130 );
and ( n23203 , C0 , RI19a22f70_2797);
or ( n54131 , n23202 , n23203 );
not ( n23204 , n27683 );
and ( n23205 , n23204 , RI19a87dd0_2739);
and ( n23206 , n54131 , n27683 );
or ( n54132 , n23205 , n23206 );
not ( n23207 , RI1754c610_2);
and ( n23208 , n23207 , n54132 );
and ( n23209 , C0 , RI1754c610_2);
or ( n54133 , n23208 , n23209 );
buf ( n54134 , n54133 );
not ( n23210 , n27683 );
and ( n23211 , n23210 , RI19a98888_2622);
and ( n23212 , RI19aa2068_2552 , n27683 );
or ( n54135 , n23211 , n23212 );
not ( n23213 , RI1754c610_2);
and ( n23214 , n23213 , n54135 );
and ( n23215 , C0 , RI1754c610_2);
or ( n54136 , n23214 , n23215 );
buf ( n54137 , n54136 );
not ( n54138 , n44224 );
and ( n54139 , n54138 , n44226 );
xor ( n54140 , n50756 , n54139 );
not ( n23216 , n29614 );
and ( n23217 , n23216 , RI174a75f8_920);
and ( n23218 , n54140 , n29614 );
or ( n54141 , n23217 , n23218 );
not ( n23219 , RI1754c610_2);
and ( n23220 , n23219 , n54141 );
and ( n23221 , C0 , RI1754c610_2);
or ( n54142 , n23220 , n23221 );
buf ( n54143 , n54142 );
not ( n54144 , n48117 );
xor ( n54145 , n36543 , n37438 );
xor ( n54146 , n54145 , n30247 );
and ( n54147 , n54144 , n54146 );
xor ( n54148 , n48114 , n54147 );
not ( n23222 , n29614 );
and ( n23223 , n23222 , RI1740a5f0_1457);
and ( n23224 , n54148 , n29614 );
or ( n54149 , n23223 , n23224 );
not ( n23225 , RI1754c610_2);
and ( n23226 , n23225 , n54149 );
and ( n23227 , C0 , RI1754c610_2);
or ( n54150 , n23226 , n23227 );
buf ( n54151 , n54150 );
buf ( n54152 , RI1747aaa8_1138);
not ( n54153 , n43439 );
and ( n54154 , n54153 , n40267 );
xor ( n54155 , n50728 , n54154 );
not ( n23228 , n29614 );
and ( n23229 , n23228 , RI17493af8_1016);
and ( n23230 , n54155 , n29614 );
or ( n54156 , n23229 , n23230 );
not ( n23231 , RI1754c610_2);
and ( n23232 , n23231 , n54156 );
and ( n23233 , C0 , RI1754c610_2);
or ( n54157 , n23232 , n23233 );
buf ( n54158 , n54157 );
not ( n23234 , n27683 );
and ( n23235 , n23234 , RI19a84ba8_2761);
and ( n23236 , RI19ac1f58_2314 , n27683 );
or ( n54159 , n23235 , n23236 );
not ( n23237 , RI1754c610_2);
and ( n23238 , n23237 , n54159 );
and ( n23239 , C0 , RI1754c610_2);
or ( n54160 , n23238 , n23239 );
buf ( n54161 , n54160 );
not ( n23240 , n27683 );
and ( n23241 , n23240 , RI19aa8530_2507);
and ( n23242 , RI19ab2670_2436 , n27683 );
or ( n54162 , n23241 , n23242 );
not ( n23243 , RI1754c610_2);
and ( n23244 , n23243 , n54162 );
and ( n23245 , C0 , RI1754c610_2);
or ( n54163 , n23244 , n23245 );
buf ( n54164 , n54163 );
not ( n54165 , n46585 );
and ( n54166 , n54165 , n42189 );
xor ( n54167 , n50951 , n54166 );
not ( n23246 , n29614 );
and ( n23247 , n23246 , RI17497608_998);
and ( n23248 , n54167 , n29614 );
or ( n54168 , n23247 , n23248 );
not ( n23249 , RI1754c610_2);
and ( n23250 , n23249 , n54168 );
and ( n23251 , C0 , RI1754c610_2);
or ( n54169 , n23250 , n23251 );
buf ( n54170 , n54169 );
xor ( n54171 , n43459 , n40949 );
xor ( n54172 , n54171 , n34572 );
xor ( n54173 , n37370 , n33505 );
xor ( n54174 , n54173 , n39635 );
not ( n54175 , n54174 );
and ( n54176 , n54175 , n53211 );
xor ( n54177 , n54172 , n54176 );
not ( n23252 , n29614 );
and ( n23253 , n23252 , RI173afed0_1898);
and ( n23254 , n54177 , n29614 );
or ( n54178 , n23253 , n23254 );
not ( n23255 , RI1754c610_2);
and ( n23256 , n23255 , n54178 );
and ( n23257 , C0 , RI1754c610_2);
or ( n54179 , n23256 , n23257 );
buf ( n54180 , n54179 );
not ( n54181 , n49422 );
and ( n54182 , n54181 , n49424 );
xor ( n54183 , n51687 , n54182 );
not ( n23258 , n29614 );
and ( n23259 , n23258 , RI1747c830_1129);
and ( n23260 , n54183 , n29614 );
or ( n54184 , n23259 , n23260 );
not ( n23261 , RI1754c610_2);
and ( n23262 , n23261 , n54184 );
and ( n23263 , C0 , RI1754c610_2);
or ( n54185 , n23262 , n23263 );
buf ( n54186 , n54185 );
not ( n54187 , n44903 );
and ( n54188 , n54187 , n46802 );
xor ( n54189 , n44900 , n54188 );
not ( n23264 , n29614 );
and ( n23265 , n23264 , RI173a6e70_1942);
and ( n23266 , n54189 , n29614 );
or ( n54190 , n23265 , n23266 );
not ( n23267 , RI1754c610_2);
and ( n23268 , n23267 , n54190 );
and ( n23269 , C0 , RI1754c610_2);
or ( n54191 , n23268 , n23269 );
buf ( n54192 , n54191 );
not ( n54193 , n47702 );
and ( n54194 , n54193 , n34518 );
xor ( n54195 , n52072 , n54194 );
not ( n23270 , n29614 );
and ( n23271 , n23270 , RI173a36a8_1959);
and ( n23272 , n54195 , n29614 );
or ( n54196 , n23271 , n23272 );
not ( n23273 , RI1754c610_2);
and ( n23274 , n23273 , n54196 );
and ( n23275 , C0 , RI1754c610_2);
or ( n54197 , n23274 , n23275 );
buf ( n54198 , n54197 );
not ( n54199 , n49517 );
and ( n54200 , n54199 , n49585 );
xor ( n54201 , n49514 , n54200 );
not ( n23276 , n29614 );
and ( n23277 , n23276 , RI173f8bc0_1543);
and ( n23278 , n54201 , n29614 );
or ( n54202 , n23277 , n23278 );
not ( n23279 , RI1754c610_2);
and ( n23280 , n23279 , n54202 );
and ( n23281 , C0 , RI1754c610_2);
or ( n54203 , n23280 , n23281 );
buf ( n54204 , n54203 );
not ( n23282 , RI1754a720_68);
and ( n23283 , n23282 , RI19a822e0_2779);
and ( n23284 , C1 , RI1754a720_68);
or ( n54205 , n23283 , n23284 );
not ( n54206 , RI1754c610_2);
and ( n54207 , n54205 , n54206 );
buf ( n54208 , n54207 );
not ( n54209 , n50215 );
and ( n54210 , n54209 , n43148 );
xor ( n54211 , n51401 , n54210 );
not ( n23285 , n29614 );
and ( n23286 , n23285 , RI173b15c8_1891);
and ( n23287 , n54211 , n29614 );
or ( n54212 , n23286 , n23287 );
not ( n23288 , RI1754c610_2);
and ( n23289 , n23288 , n54212 );
and ( n23290 , C0 , RI1754c610_2);
or ( n54213 , n23289 , n23290 );
buf ( n54214 , n54213 );
not ( n23291 , n27683 );
and ( n23292 , n23291 , RI19aa0f10_2561);
and ( n23293 , RI19aaad80_2489 , n27683 );
or ( n54215 , n23292 , n23293 );
not ( n23294 , RI1754c610_2);
and ( n23295 , n23294 , n54215 );
and ( n23296 , C0 , RI1754c610_2);
or ( n54216 , n23295 , n23296 );
buf ( n54217 , n54216 );
xor ( n54218 , n39901 , n33397 );
xor ( n54219 , n54218 , n35710 );
not ( n54220 , n54219 );
and ( n54221 , n54220 , n48592 );
xor ( n54222 , n47068 , n54221 );
not ( n23297 , n29614 );
and ( n23298 , n23297 , RI174b6f58_844);
and ( n23299 , n54222 , n29614 );
or ( n54223 , n23298 , n23299 );
not ( n23300 , RI1754c610_2);
and ( n23301 , n23300 , n54223 );
and ( n23302 , C0 , RI1754c610_2);
or ( n54224 , n23301 , n23302 );
buf ( n54225 , n54224 );
not ( n54226 , n40891 );
and ( n54227 , n54226 , n44183 );
xor ( n54228 , n40869 , n54227 );
not ( n23303 , n29614 );
and ( n23304 , n23303 , RI17464848_1246);
and ( n23305 , n54228 , n29614 );
or ( n54229 , n23304 , n23305 );
not ( n23306 , RI1754c610_2);
and ( n23307 , n23306 , n54229 );
and ( n23308 , C0 , RI1754c610_2);
or ( n54230 , n23307 , n23308 );
buf ( n54231 , n54230 );
not ( n54232 , n43409 );
and ( n54233 , n54232 , n43411 );
xor ( n54234 , n46746 , n54233 );
not ( n23309 , n29614 );
and ( n23310 , n23309 , RI17403660_1491);
and ( n23311 , n54234 , n29614 );
or ( n54235 , n23310 , n23311 );
not ( n23312 , RI1754c610_2);
and ( n23313 , n23312 , n54235 );
and ( n23314 , C0 , RI1754c610_2);
or ( n54236 , n23313 , n23314 );
buf ( n54237 , n54236 );
not ( n54238 , n52072 );
and ( n54239 , n54238 , n47702 );
xor ( n54240 , n34645 , n54239 );
not ( n23315 , n29614 );
and ( n23316 , n23315 , RI17394a68_2031);
and ( n23317 , n54240 , n29614 );
or ( n54241 , n23316 , n23317 );
not ( n23318 , RI1754c610_2);
and ( n23319 , n23318 , n54241 );
and ( n23320 , C0 , RI1754c610_2);
or ( n54242 , n23319 , n23320 );
buf ( n54243 , n54242 );
not ( n54244 , n45438 );
and ( n54245 , n54244 , n45440 );
xor ( n54246 , n43062 , n54245 );
not ( n23321 , n29614 );
and ( n23322 , n23321 , RI17462430_1257);
and ( n23323 , n54246 , n29614 );
or ( n54247 , n23322 , n23323 );
not ( n23324 , RI1754c610_2);
and ( n23325 , n23324 , n54247 );
and ( n23326 , C0 , RI1754c610_2);
or ( n54248 , n23325 , n23326 );
buf ( n54249 , n54248 );
not ( n23327 , n27683 );
and ( n23328 , n23327 , RI19abd9f8_2353);
and ( n23329 , RI19ac6620_2282 , n27683 );
or ( n54250 , n23328 , n23329 );
not ( n23330 , RI1754c610_2);
and ( n23331 , n23330 , n54250 );
and ( n23332 , C0 , RI1754c610_2);
or ( n54251 , n23331 , n23332 );
buf ( n54252 , n54251 );
not ( n23333 , RI1754c610_2);
and ( n23334 , n23333 , RI19ad1858_2201);
and ( n23335 , C0 , RI1754c610_2);
or ( n54253 , n23334 , n23335 );
buf ( n54254 , n54253 );
buf ( n54255 , RI174a3458_940);
not ( n54256 , n43750 );
and ( n54257 , n54256 , n43847 );
xor ( n54258 , n43747 , n54257 );
not ( n23336 , n29614 );
and ( n23337 , n23336 , RI17415720_1403);
and ( n23338 , n54258 , n29614 );
or ( n54259 , n23337 , n23338 );
not ( n23339 , RI1754c610_2);
and ( n23340 , n23339 , n54259 );
and ( n23341 , C0 , RI1754c610_2);
or ( n54260 , n23340 , n23341 );
buf ( n54261 , n54260 );
buf ( n54262 , RI174afc80_879);
buf ( n54263 , RI17501ef8_754);
not ( n54264 , n48876 );
and ( n54265 , n54264 , n51582 );
xor ( n54266 , n48804 , n54265 );
not ( n23342 , n29614 );
and ( n23343 , n23342 , RI173f50b0_1561);
and ( n23344 , n54266 , n29614 );
or ( n54267 , n23343 , n23344 );
not ( n23345 , RI1754c610_2);
and ( n23346 , n23345 , n54267 );
and ( n23347 , C0 , RI1754c610_2);
or ( n54268 , n23346 , n23347 );
buf ( n54269 , n54268 );
buf ( n54270 , RI174896e8_1066);
not ( n54271 , n45063 );
and ( n54272 , n54271 , n42960 );
xor ( n54273 , n35598 , n54272 );
not ( n23348 , n29614 );
and ( n23349 , n23348 , RI17406450_1477);
and ( n23350 , n54273 , n29614 );
or ( n54274 , n23349 , n23350 );
not ( n23351 , RI1754c610_2);
and ( n23352 , n23351 , n54274 );
and ( n23353 , C0 , RI1754c610_2);
or ( n54275 , n23352 , n23353 );
buf ( n54276 , n54275 );
not ( n54277 , n45367 );
and ( n54278 , n54277 , n45369 );
xor ( n54279 , n46174 , n54278 );
not ( n23354 , n29614 );
and ( n23355 , n23354 , RI1739c718_1993);
and ( n23356 , n54279 , n29614 );
or ( n54280 , n23355 , n23356 );
not ( n23357 , RI1754c610_2);
and ( n23358 , n23357 , n54280 );
and ( n23359 , C0 , RI1754c610_2);
or ( n54281 , n23358 , n23359 );
buf ( n54282 , n54281 );
not ( n54283 , n35855 );
and ( n54284 , n54283 , n31622 );
xor ( n54285 , n42715 , n54284 );
not ( n23360 , n29614 );
and ( n23361 , n23360 , RI17343168_2114);
and ( n23362 , n54285 , n29614 );
or ( n54286 , n23361 , n23362 );
not ( n23363 , RI1754c610_2);
and ( n23364 , n23363 , n54286 );
and ( n23365 , C0 , RI1754c610_2);
or ( n54287 , n23364 , n23365 );
buf ( n54288 , n54287 );
not ( n54289 , n45291 );
and ( n54290 , n54289 , n43071 );
xor ( n54291 , n42849 , n54290 );
not ( n23366 , n29614 );
and ( n23367 , n23366 , RI174b0658_876);
and ( n23368 , n54291 , n29614 );
or ( n54292 , n23367 , n23368 );
not ( n23369 , RI1754c610_2);
and ( n23370 , n23369 , n54292 );
and ( n23371 , C0 , RI1754c610_2);
or ( n54293 , n23370 , n23371 );
buf ( n54294 , n54293 );
not ( n54295 , n37697 );
and ( n54296 , n54295 , n37745 );
xor ( n54297 , n45250 , n54296 );
not ( n23372 , n29614 );
and ( n23373 , n23372 , RI173d15c0_1735);
and ( n23374 , n54297 , n29614 );
or ( n54298 , n23373 , n23374 );
not ( n23375 , RI1754c610_2);
and ( n23376 , n23375 , n54298 );
and ( n23377 , C0 , RI1754c610_2);
or ( n54299 , n23376 , n23377 );
buf ( n54300 , n54299 );
not ( n54301 , n46959 );
and ( n54302 , n54301 , n52596 );
xor ( n54303 , n41405 , n54302 );
not ( n23378 , n29614 );
and ( n23379 , n23378 , RI1749df08_966);
and ( n23380 , n54303 , n29614 );
or ( n54304 , n23379 , n23380 );
not ( n23381 , RI1754c610_2);
and ( n23382 , n23381 , n54304 );
and ( n23383 , C0 , RI1754c610_2);
or ( n54305 , n23382 , n23383 );
buf ( n54306 , n54305 );
not ( n54307 , n49473 );
and ( n54308 , n54307 , n51230 );
xor ( n54309 , n49150 , n54308 );
not ( n23384 , n29614 );
and ( n23385 , n23384 , RI1751cfa0_676);
and ( n23386 , n54309 , n29614 );
or ( n54310 , n23385 , n23386 );
not ( n23387 , RI1754c610_2);
and ( n23388 , n23387 , n54310 );
and ( n23389 , C0 , RI1754c610_2);
or ( n54311 , n23388 , n23389 );
buf ( n54312 , n54311 );
not ( n54313 , n49292 );
and ( n54314 , n54313 , n49294 );
xor ( n54315 , n51312 , n54314 );
not ( n23390 , n29614 );
and ( n23391 , n23390 , RI17395e18_2025);
and ( n23392 , n54315 , n29614 );
or ( n54316 , n23391 , n23392 );
not ( n23393 , RI1754c610_2);
and ( n23394 , n23393 , n54316 );
and ( n23395 , C0 , RI1754c610_2);
or ( n54317 , n23394 , n23395 );
buf ( n54318 , n54317 );
not ( n54319 , n44910 );
and ( n54320 , n54319 , n44912 );
xor ( n54321 , n52807 , n54320 );
not ( n23396 , n29614 );
and ( n23397 , n23396 , RI17470d28_1186);
and ( n23398 , n54321 , n29614 );
or ( n54322 , n23397 , n23398 );
not ( n23399 , RI1754c610_2);
and ( n23400 , n23399 , n54322 );
and ( n23401 , C0 , RI1754c610_2);
or ( n54323 , n23400 , n23401 );
buf ( n54324 , n54323 );
not ( n54325 , n46093 );
and ( n54326 , n54325 , n42505 );
xor ( n54327 , n44706 , n54326 );
not ( n23402 , n29614 );
and ( n23403 , n23402 , RI173e8f18_1620);
and ( n23404 , n54327 , n29614 );
or ( n54328 , n23403 , n23404 );
not ( n23405 , RI1754c610_2);
and ( n23406 , n23405 , n54328 );
and ( n23407 , C0 , RI1754c610_2);
or ( n54329 , n23406 , n23407 );
buf ( n54330 , n54329 );
not ( n54331 , n45129 );
and ( n54332 , n54331 , n45131 );
xor ( n54333 , n52348 , n54332 );
not ( n23408 , n29614 );
and ( n23409 , n23408 , RI1748fca0_1035);
and ( n23410 , n54333 , n29614 );
or ( n54334 , n23409 , n23410 );
not ( n23411 , RI1754c610_2);
and ( n23412 , n23411 , n54334 );
and ( n23413 , C0 , RI1754c610_2);
or ( n54335 , n23412 , n23413 );
buf ( n54336 , n54335 );
not ( n54337 , n41626 );
and ( n54338 , n54337 , n51246 );
xor ( n54339 , n41623 , n54338 );
not ( n23414 , n29614 );
and ( n23415 , n23414 , RI1747d550_1125);
and ( n23416 , n54339 , n29614 );
or ( n54340 , n23415 , n23416 );
not ( n23417 , RI1754c610_2);
and ( n23418 , n23417 , n54340 );
and ( n23419 , C0 , RI1754c610_2);
or ( n54341 , n23418 , n23419 );
buf ( n54342 , n54341 );
and ( n54343 , RI1754b4b8_39 , n34844 );
and ( n54344 , RI1754b4b8_39 , n34847 );
and ( n54345 , RI1754b4b8_39 , n34850 );
or ( n54346 , n54343 , n54344 , n54345 , C0 , C0 , C0 , C0 , C0 );
not ( n23420 , n34859 );
and ( n23421 , n23420 , n54346 );
and ( n23422 , RI1754b4b8_39 , n34859 );
or ( n54347 , n23421 , n23422 );
not ( n23423 , RI19a22f70_2797);
and ( n23424 , n23423 , n54347 );
and ( n23425 , C0 , RI19a22f70_2797);
or ( n54348 , n23424 , n23425 );
not ( n23426 , n27683 );
and ( n23427 , n23426 , RI19ab6cc0_2403);
and ( n23428 , n54348 , n27683 );
or ( n54349 , n23427 , n23428 );
not ( n23429 , RI1754c610_2);
and ( n23430 , n23429 , n54349 );
and ( n23431 , C0 , RI1754c610_2);
or ( n54350 , n23430 , n23431 );
buf ( n54351 , n54350 );
not ( n23432 , n27683 );
and ( n23433 , n23432 , RI19aae458_2466);
and ( n23434 , RI19ab7f80_2395 , n27683 );
or ( n54352 , n23433 , n23434 );
not ( n23435 , RI1754c610_2);
and ( n23436 , n23435 , n54352 );
and ( n23437 , C0 , RI1754c610_2);
or ( n54353 , n23436 , n23437 );
buf ( n54354 , n54353 );
not ( n54355 , n48489 );
and ( n54356 , n54355 , n47984 );
xor ( n54357 , n52051 , n54356 );
not ( n23438 , n29614 );
and ( n23439 , n23438 , RI17481d80_1103);
and ( n23440 , n54357 , n29614 );
or ( n54358 , n23439 , n23440 );
not ( n23441 , RI1754c610_2);
and ( n23442 , n23441 , n54358 );
and ( n23443 , C0 , RI1754c610_2);
or ( n54359 , n23442 , n23443 );
buf ( n54360 , n54359 );
not ( n23444 , n27683 );
and ( n23445 , n23444 , RI19ace168_2224);
and ( n23446 , RI19a95048_2647 , n27683 );
or ( n54361 , n23445 , n23446 );
not ( n23447 , RI1754c610_2);
and ( n23448 , n23447 , n54361 );
and ( n23449 , C0 , RI1754c610_2);
or ( n54362 , n23448 , n23449 );
buf ( n54363 , n54362 );
not ( n54364 , n43626 );
and ( n54365 , n54364 , n48962 );
xor ( n54366 , n43623 , n54365 );
not ( n23450 , n29614 );
and ( n23451 , n23450 , RI173a95d0_1930);
and ( n23452 , n54366 , n29614 );
or ( n54367 , n23451 , n23452 );
not ( n23453 , RI1754c610_2);
and ( n23454 , n23453 , n54367 );
and ( n23455 , C0 , RI1754c610_2);
or ( n54368 , n23454 , n23455 );
buf ( n54369 , n54368 );
not ( n54370 , n45809 );
and ( n54371 , n54370 , n51802 );
xor ( n54372 , n45806 , n54371 );
not ( n23456 , n29614 );
and ( n23457 , n23456 , RI1744fce0_1347);
and ( n23458 , n54372 , n29614 );
or ( n54373 , n23457 , n23458 );
not ( n23459 , RI1754c610_2);
and ( n23460 , n23459 , n54373 );
and ( n23461 , C0 , RI1754c610_2);
or ( n54374 , n23460 , n23461 );
buf ( n54375 , n54374 );
not ( n54376 , n50982 );
and ( n54377 , n54376 , n45896 );
xor ( n54378 , n43826 , n54377 );
not ( n23462 , n29614 );
and ( n23463 , n23462 , RI173c43a8_1799);
and ( n23464 , n54378 , n29614 );
or ( n54379 , n23463 , n23464 );
not ( n23465 , RI1754c610_2);
and ( n23466 , n23465 , n54379 );
and ( n23467 , C0 , RI1754c610_2);
or ( n54380 , n23466 , n23467 );
buf ( n54381 , n54380 );
not ( n54382 , n44352 );
and ( n54383 , n54382 , n47573 );
xor ( n54384 , n44349 , n54383 );
not ( n23468 , n29614 );
and ( n23469 , n23468 , RI17397510_2018);
and ( n23470 , n54384 , n29614 );
or ( n54385 , n23469 , n23470 );
not ( n23471 , RI1754c610_2);
and ( n23472 , n23471 , n54385 );
and ( n23473 , C0 , RI1754c610_2);
or ( n54386 , n23472 , n23473 );
buf ( n54387 , n54386 );
not ( n23474 , n27683 );
and ( n23475 , n23474 , RI19ac4280_2298);
and ( n23476 , RI19accea8_2232 , n27683 );
or ( n54388 , n23475 , n23476 );
not ( n23477 , RI1754c610_2);
and ( n23478 , n23477 , n54388 );
and ( n23479 , C0 , RI1754c610_2);
or ( n54389 , n23478 , n23479 );
buf ( n54390 , n54389 );
not ( n23480 , n27683 );
and ( n23481 , n23480 , RI19ab3de0_2424);
and ( n23482 , RI19abd890_2354 , n27683 );
or ( n54391 , n23481 , n23482 );
not ( n23483 , RI1754c610_2);
and ( n23484 , n23483 , n54391 );
and ( n23485 , C0 , RI1754c610_2);
or ( n54392 , n23484 , n23485 );
buf ( n54393 , n54392 );
not ( n23486 , n27683 );
and ( n23487 , n23486 , RI19aac6d0_2480);
and ( n23488 , RI19ab5f28_2409 , n27683 );
or ( n54394 , n23487 , n23488 );
not ( n23489 , RI1754c610_2);
and ( n23490 , n23489 , n54394 );
and ( n23491 , C0 , RI1754c610_2);
or ( n54395 , n23490 , n23491 );
buf ( n54396 , n54395 );
not ( n54397 , n42485 );
and ( n54398 , n54397 , n52768 );
xor ( n54399 , n42482 , n54398 );
not ( n23492 , n29614 );
and ( n23493 , n23492 , RI17401248_1502);
and ( n23494 , n54399 , n29614 );
or ( n54400 , n23493 , n23494 );
not ( n23495 , RI1754c610_2);
and ( n23496 , n23495 , n54400 );
and ( n23497 , C0 , RI1754c610_2);
or ( n54401 , n23496 , n23497 );
buf ( n54402 , n54401 );
not ( n54403 , n47068 );
and ( n54404 , n54403 , n54219 );
xor ( n54405 , n47065 , n54404 );
not ( n23498 , n29614 );
and ( n23499 , n23498 , RI1733a108_2158);
and ( n23500 , n54405 , n29614 );
or ( n54406 , n23499 , n23500 );
not ( n23501 , RI1754c610_2);
and ( n23502 , n23501 , n54406 );
and ( n23503 , C0 , RI1754c610_2);
or ( n54407 , n23502 , n23503 );
buf ( n54408 , n54407 );
not ( n54409 , n50951 );
and ( n54410 , n54409 , n46585 );
xor ( n54411 , n42194 , n54410 );
not ( n23504 , n29614 );
and ( n23505 , n23504 , RI17488d10_1069);
and ( n23506 , n54411 , n29614 );
or ( n54412 , n23505 , n23506 );
not ( n23507 , RI1754c610_2);
and ( n23508 , n23507 , n54412 );
and ( n23509 , C0 , RI1754c610_2);
or ( n54413 , n23508 , n23509 );
buf ( n54414 , n54413 );
not ( n54415 , n50714 );
and ( n54416 , n54415 , n50480 );
xor ( n54417 , n52430 , n54416 );
not ( n23510 , n29614 );
and ( n23511 , n23510 , RI174a1388_950);
and ( n23512 , n54417 , n29614 );
or ( n54418 , n23511 , n23512 );
not ( n23513 , RI1754c610_2);
and ( n23514 , n23513 , n54418 );
and ( n23515 , C0 , RI1754c610_2);
or ( n54419 , n23514 , n23515 );
buf ( n54420 , n54419 );
not ( n54421 , n47019 );
and ( n54422 , n54421 , n47021 );
xor ( n54423 , n47908 , n54422 );
not ( n23516 , n29614 );
and ( n23517 , n23516 , RI174cfd50_764);
and ( n23518 , n54423 , n29614 );
or ( n54424 , n23517 , n23518 );
not ( n23519 , RI1754c610_2);
and ( n23520 , n23519 , n54424 );
and ( n23521 , C0 , RI1754c610_2);
or ( n54425 , n23520 , n23521 );
buf ( n54426 , n54425 );
not ( n54427 , n46516 );
and ( n54428 , n54427 , n49394 );
xor ( n54429 , n44760 , n54428 );
not ( n23522 , n29614 );
and ( n23523 , n23522 , RI173fafd8_1532);
and ( n23524 , n54429 , n29614 );
or ( n54430 , n23523 , n23524 );
not ( n23525 , RI1754c610_2);
and ( n23526 , n23525 , n54430 );
and ( n23527 , C0 , RI1754c610_2);
or ( n54431 , n23526 , n23527 );
buf ( n54432 , n54431 );
not ( n54433 , n49588 );
and ( n54434 , n54433 , n49512 );
xor ( n54435 , n49585 , n54434 );
not ( n23528 , n29614 );
and ( n23529 , n23528 , RI173cd0c0_1756);
and ( n23530 , n54435 , n29614 );
or ( n54436 , n23529 , n23530 );
not ( n23531 , RI1754c610_2);
and ( n23532 , n23531 , n54436 );
and ( n23533 , C0 , RI1754c610_2);
or ( n54437 , n23532 , n23533 );
buf ( n54438 , n54437 );
not ( n54439 , n54172 );
and ( n54440 , n54439 , n54174 );
xor ( n54441 , n53216 , n54440 );
not ( n23534 , n29614 );
and ( n23535 , n23534 , RI173a1920_1968);
and ( n23536 , n54441 , n29614 );
or ( n54442 , n23535 , n23536 );
not ( n23537 , RI1754c610_2);
and ( n23538 , n23537 , n54442 );
and ( n23539 , C0 , RI1754c610_2);
or ( n54443 , n23538 , n23539 );
buf ( n54444 , n54443 );
not ( n54445 , n48284 );
and ( n54446 , n54445 , n48286 );
xor ( n54447 , n52582 , n54446 );
not ( n23540 , n29614 );
and ( n23541 , n23540 , RI17515908_699);
and ( n23542 , n54447 , n29614 );
or ( n54448 , n23541 , n23542 );
not ( n23543 , RI1754c610_2);
and ( n23544 , n23543 , n54448 );
and ( n23545 , C0 , RI1754c610_2);
or ( n54449 , n23544 , n23545 );
buf ( n54450 , n54449 );
not ( n54451 , n41947 );
and ( n54452 , n54451 , n41949 );
xor ( n54453 , n51052 , n54452 );
not ( n23546 , n29614 );
and ( n23547 , n23546 , RI1739ca60_1992);
and ( n23548 , n54453 , n29614 );
or ( n54454 , n23547 , n23548 );
not ( n23549 , RI1754c610_2);
and ( n23550 , n23549 , n54454 );
and ( n23551 , C0 , RI1754c610_2);
or ( n54455 , n23550 , n23551 );
buf ( n54456 , n54455 );
not ( n54457 , n40898 );
and ( n54458 , n54457 , n40903 );
xor ( n54459 , n47554 , n54458 );
not ( n23552 , n29614 );
and ( n23553 , n23552 , RI173895f0_2086);
and ( n23554 , n54459 , n29614 );
or ( n54460 , n23553 , n23554 );
not ( n23555 , RI1754c610_2);
and ( n23556 , n23555 , n54460 );
and ( n23557 , C0 , RI1754c610_2);
or ( n54461 , n23556 , n23557 );
buf ( n54462 , n54461 );
not ( n23558 , n27683 );
and ( n23559 , n23558 , RI19abd188_2358);
and ( n23560 , RI19ac5978_2287 , n27683 );
or ( n54463 , n23559 , n23560 );
not ( n23561 , RI1754c610_2);
and ( n23562 , n23561 , n54463 );
and ( n23563 , C0 , RI1754c610_2);
or ( n54464 , n23562 , n23563 );
buf ( n54465 , n54464 );
not ( n23564 , n27683 );
and ( n23565 , n23564 , RI19aa1f00_2553);
and ( n23566 , RI19aac040_2482 , n27683 );
or ( n54466 , n23565 , n23566 );
not ( n23567 , RI1754c610_2);
and ( n23568 , n23567 , n54466 );
and ( n23569 , C0 , RI1754c610_2);
or ( n54467 , n23568 , n23569 );
buf ( n54468 , n54467 );
not ( n54469 , n39302 );
and ( n54470 , n54469 , n39304 );
xor ( n54471 , n44802 , n54470 );
not ( n23570 , n29614 );
and ( n23571 , n23570 , RI17391fc0_2044);
and ( n23572 , n54471 , n29614 );
or ( n54472 , n23571 , n23572 );
not ( n23573 , RI1754c610_2);
and ( n23574 , n23573 , n54472 );
and ( n23575 , C0 , RI1754c610_2);
or ( n54473 , n23574 , n23575 );
buf ( n54474 , n54473 );
not ( n54475 , n42777 );
and ( n54476 , n54475 , n41252 );
xor ( n54477 , n49696 , n54476 );
not ( n23576 , n29614 );
and ( n23577 , n23576 , RI17456fb8_1312);
and ( n23578 , n54477 , n29614 );
or ( n54478 , n23577 , n23578 );
not ( n23579 , RI1754c610_2);
and ( n23580 , n23579 , n54478 );
and ( n23581 , C0 , RI1754c610_2);
or ( n54479 , n23580 , n23581 );
buf ( n54480 , n54479 );
not ( n23582 , n27683 );
and ( n23583 , n23582 , RI19abe9e8_2344);
and ( n23584 , RI19ac7958_2273 , n27683 );
or ( n54481 , n23583 , n23584 );
not ( n23585 , RI1754c610_2);
and ( n23586 , n23585 , n54481 );
and ( n23587 , C0 , RI1754c610_2);
or ( n54482 , n23586 , n23587 );
buf ( n54483 , n54482 );
not ( n54484 , n48131 );
and ( n54485 , n54484 , n47544 );
xor ( n54486 , n44850 , n54485 );
not ( n23588 , n29614 );
and ( n23589 , n23588 , RI173dcd80_1679);
and ( n23590 , n54486 , n29614 );
or ( n54487 , n23589 , n23590 );
not ( n23591 , RI1754c610_2);
and ( n23592 , n23591 , n54487 );
and ( n23593 , C0 , RI1754c610_2);
or ( n54488 , n23592 , n23593 );
buf ( n54489 , n54488 );
not ( n54490 , n43962 );
and ( n54491 , n54490 , n46101 );
xor ( n54492 , n43959 , n54491 );
not ( n23594 , n29614 );
and ( n23595 , n23594 , RI1752c1f8_629);
and ( n23596 , n54492 , n29614 );
or ( n54493 , n23595 , n23596 );
not ( n23597 , RI1754c610_2);
and ( n23598 , n23597 , n54493 );
and ( n23599 , C0 , RI1754c610_2);
or ( n54494 , n23598 , n23599 );
buf ( n54495 , n54494 );
not ( n54496 , n50782 );
and ( n54497 , n54496 , n54103 );
xor ( n54498 , n49566 , n54497 );
not ( n23600 , n29614 );
and ( n23601 , n23600 , RI1751b0b0_682);
and ( n23602 , n54498 , n29614 );
or ( n54499 , n23601 , n23602 );
not ( n23603 , RI1754c610_2);
and ( n23604 , n23603 , n54499 );
and ( n23605 , C0 , RI1754c610_2);
or ( n54500 , n23604 , n23605 );
buf ( n54501 , n54500 );
not ( n54502 , n46174 );
and ( n54503 , n54502 , n45367 );
xor ( n54504 , n46171 , n54503 );
not ( n23606 , n29614 );
and ( n23607 , n23606 , RI1738de20_2064);
and ( n23608 , n54504 , n29614 );
or ( n54505 , n23607 , n23608 );
not ( n23609 , RI1754c610_2);
and ( n23610 , n23609 , n54505 );
and ( n23611 , C0 , RI1754c610_2);
or ( n54506 , n23610 , n23611 );
buf ( n54507 , n54506 );
not ( n54508 , n45498 );
and ( n54509 , n54508 , n45500 );
xor ( n54510 , n38190 , n54509 );
not ( n23612 , n29614 );
and ( n23613 , n23612 , RI173c4a38_1797);
and ( n23614 , n54510 , n29614 );
or ( n54511 , n23613 , n23614 );
not ( n23615 , RI1754c610_2);
and ( n23616 , n23615 , n54511 );
and ( n23617 , C0 , RI1754c610_2);
or ( n54512 , n23616 , n23617 );
buf ( n54513 , n54512 );
not ( n54514 , n46764 );
and ( n54515 , n54514 , n46615 );
xor ( n54516 , n36655 , n54515 );
not ( n23618 , n29614 );
and ( n23619 , n23618 , RI173ef188_1590);
and ( n23620 , n54516 , n29614 );
or ( n54517 , n23619 , n23620 );
not ( n23621 , RI1754c610_2);
and ( n23622 , n23621 , n54517 );
and ( n23623 , C0 , RI1754c610_2);
or ( n54518 , n23622 , n23623 );
buf ( n54519 , n54518 );
not ( n23624 , n27683 );
and ( n23625 , n23624 , RI19acb300_2246);
and ( n23626 , RI19a869a8_2748 , n27683 );
or ( n54520 , n23625 , n23626 );
not ( n23627 , RI1754c610_2);
and ( n23628 , n23627 , n54520 );
and ( n23629 , C0 , RI1754c610_2);
or ( n54521 , n23628 , n23629 );
buf ( n54522 , n54521 );
not ( n23630 , n27683 );
and ( n23631 , n23630 , RI19ac0680_2328);
and ( n23632 , RI19ac9938_2258 , n27683 );
or ( n54523 , n23631 , n23632 );
not ( n23633 , RI1754c610_2);
and ( n23634 , n23633 , n54523 );
and ( n23635 , C0 , RI1754c610_2);
or ( n54524 , n23634 , n23635 );
buf ( n54525 , n54524 );
not ( n54526 , n49237 );
and ( n54527 , n54526 , n46427 );
xor ( n54528 , n49234 , n54527 );
not ( n23636 , n29614 );
and ( n23637 , n23636 , RI173a0228_1975);
and ( n23638 , n54528 , n29614 );
or ( n54529 , n23637 , n23638 );
not ( n23639 , RI1754c610_2);
and ( n23640 , n23639 , n54529 );
and ( n23641 , C0 , RI1754c610_2);
or ( n54530 , n23640 , n23641 );
buf ( n54531 , n54530 );
not ( n23642 , n27683 );
and ( n23643 , n23642 , RI19a93fe0_2654);
and ( n23644 , RI19a9e288_2583 , n27683 );
or ( n54532 , n23643 , n23644 );
not ( n23645 , RI1754c610_2);
and ( n23646 , n23645 , n54532 );
and ( n23647 , C0 , RI1754c610_2);
or ( n54533 , n23646 , n23647 );
buf ( n54534 , n54533 );
not ( n54535 , n45721 );
and ( n54536 , n54535 , n51076 );
xor ( n54537 , n45718 , n54536 );
not ( n23648 , n29614 );
and ( n23649 , n23648 , RI174d0278_763);
and ( n23650 , n54537 , n29614 );
or ( n54538 , n23649 , n23650 );
not ( n23651 , RI1754c610_2);
and ( n23652 , n23651 , n54538 );
and ( n23653 , C0 , RI1754c610_2);
or ( n54539 , n23652 , n23653 );
buf ( n54540 , n54539 );
not ( n54541 , n52807 );
and ( n54542 , n54541 , n44910 );
xor ( n54543 , n47355 , n54542 );
not ( n23654 , n29614 );
and ( n23655 , n23654 , RI17453e80_1327);
and ( n23656 , n54543 , n29614 );
or ( n54544 , n23655 , n23656 );
not ( n23657 , RI1754c610_2);
and ( n23658 , n23657 , n54544 );
and ( n23659 , C0 , RI1754c610_2);
or ( n54545 , n23658 , n23659 );
buf ( n54546 , n54545 );
not ( n54547 , n49217 );
and ( n54548 , n54547 , n48168 );
xor ( n54549 , n52879 , n54548 );
not ( n23660 , n29614 );
and ( n23661 , n23660 , RI174c5850_796);
and ( n23662 , n54549 , n29614 );
or ( n54550 , n23661 , n23662 );
not ( n23663 , RI1754c610_2);
and ( n23664 , n23663 , n54550 );
and ( n23665 , C0 , RI1754c610_2);
or ( n54551 , n23664 , n23665 );
buf ( n54552 , n54551 );
and ( n54553 , RI1754b0f8_47 , n34844 );
and ( n54554 , RI1754b0f8_47 , n34847 );
or ( n54555 , n54553 , n54554 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n23666 , n34859 );
and ( n23667 , n23666 , n54555 );
and ( n23668 , RI1754b0f8_47 , n34859 );
or ( n54556 , n23667 , n23668 );
not ( n23669 , RI19a22f70_2797);
and ( n23670 , n23669 , n54556 );
and ( n23671 , C0 , RI19a22f70_2797);
or ( n54557 , n23670 , n23671 );
not ( n23672 , n27683 );
and ( n23673 , n23672 , RI19ac1f58_2314);
and ( n23674 , n54557 , n27683 );
or ( n54558 , n23673 , n23674 );
not ( n23675 , RI1754c610_2);
and ( n23676 , n23675 , n54558 );
and ( n23677 , C0 , RI1754c610_2);
or ( n54559 , n23676 , n23677 );
buf ( n54560 , n54559 );
not ( n54561 , n45229 );
and ( n54562 , n54561 , n46497 );
xor ( n54563 , n45226 , n54562 );
not ( n23678 , n29614 );
and ( n23679 , n23678 , RI17412c78_1416);
and ( n23680 , n54563 , n29614 );
or ( n54564 , n23679 , n23680 );
not ( n23681 , RI1754c610_2);
and ( n23682 , n23681 , n54564 );
and ( n23683 , C0 , RI1754c610_2);
or ( n54565 , n23682 , n23683 );
buf ( n54566 , n54565 );
not ( n54567 , n40770 );
and ( n54568 , n54567 , n40772 );
xor ( n54569 , n43015 , n54568 );
not ( n23684 , n29614 );
and ( n23685 , n23684 , RI173c6478_1789);
and ( n23686 , n54569 , n29614 );
or ( n54570 , n23685 , n23686 );
not ( n23687 , RI1754c610_2);
and ( n23688 , n23687 , n54570 );
and ( n23689 , C0 , RI1754c610_2);
or ( n54571 , n23688 , n23689 );
buf ( n54572 , n54571 );
not ( n54573 , n44030 );
and ( n54574 , n54573 , n42456 );
xor ( n54575 , n43790 , n54574 );
not ( n23690 , n29614 );
and ( n23691 , n23690 , RI173b7b80_1860);
and ( n23692 , n54575 , n29614 );
or ( n54576 , n23691 , n23692 );
not ( n23693 , RI1754c610_2);
and ( n23694 , n23693 , n54576 );
and ( n23695 , C0 , RI1754c610_2);
or ( n54577 , n23694 , n23695 );
buf ( n54578 , n54577 );
not ( n54579 , n43945 );
and ( n54580 , n54579 , n43947 );
xor ( n54581 , n50065 , n54580 );
not ( n23696 , n29614 );
and ( n23697 , n23696 , RI1751c028_679);
and ( n23698 , n54581 , n29614 );
or ( n54582 , n23697 , n23698 );
not ( n23699 , RI1754c610_2);
and ( n23700 , n23699 , n54582 );
and ( n23701 , C0 , RI1754c610_2);
or ( n54583 , n23700 , n23701 );
buf ( n54584 , n54583 );
not ( n54585 , n45886 );
and ( n54586 , n54585 , n49665 );
xor ( n54587 , n45420 , n54586 );
not ( n23702 , n29614 );
and ( n23703 , n23702 , RI17493468_1018);
and ( n23704 , n54587 , n29614 );
or ( n54588 , n23703 , n23704 );
not ( n23705 , RI1754c610_2);
and ( n23706 , n23705 , n54588 );
and ( n23707 , C0 , RI1754c610_2);
or ( n54589 , n23706 , n23707 );
buf ( n54590 , n54589 );
not ( n23708 , n27683 );
and ( n23709 , n23708 , RI19ac3b00_2301);
and ( n23710 , RI19acc818_2235 , n27683 );
or ( n54591 , n23709 , n23710 );
not ( n23711 , RI1754c610_2);
and ( n23712 , n23711 , n54591 );
and ( n23713 , C0 , RI1754c610_2);
or ( n54592 , n23712 , n23713 );
buf ( n54593 , n54592 );
buf ( n54594 , RI17497fe0_995);
buf ( n54595 , RI174bc7f0_824);
buf ( n54596 , RI17479d88_1142);
and ( n54597 , RI1754c0e8_13 , n34844 );
and ( n54598 , RI1754c0e8_13 , n34847 );
and ( n54599 , RI1754c0e8_13 , n34850 );
and ( n54600 , RI1754c0e8_13 , n34852 );
and ( n54601 , RI1754c0e8_13 , n34854 );
and ( n54602 , RI1754c0e8_13 , n34856 );
or ( n54603 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , C0 , C0 );
not ( n23714 , n34859 );
and ( n23715 , n23714 , n54603 );
and ( n23716 , RI1754c0e8_13 , n34859 );
or ( n54604 , n23715 , n23716 );
not ( n23717 , RI19a22f70_2797);
and ( n23718 , n23717 , n54604 );
and ( n23719 , C0 , RI19a22f70_2797);
or ( n54605 , n23718 , n23719 );
not ( n23720 , n27683 );
and ( n23721 , n23720 , RI19a8eb08_2692);
and ( n23722 , n54605 , n27683 );
or ( n54606 , n23721 , n23722 );
not ( n23723 , RI1754c610_2);
and ( n23724 , n23723 , n54606 );
and ( n23725 , C0 , RI1754c610_2);
or ( n54607 , n23724 , n23725 );
buf ( n54608 , n54607 );
not ( n54609 , n53466 );
and ( n54610 , n54609 , n51460 );
xor ( n54611 , n30742 , n54610 );
not ( n23726 , n29614 );
and ( n23727 , n23726 , RI1739cda8_1991);
and ( n23728 , n54611 , n29614 );
or ( n54612 , n23727 , n23728 );
not ( n23729 , RI1754c610_2);
and ( n23730 , n23729 , n54612 );
and ( n23731 , C0 , RI1754c610_2);
or ( n54613 , n23730 , n23731 );
buf ( n54614 , n54613 );
not ( n54615 , n42240 );
and ( n54616 , n54615 , n53957 );
xor ( n54617 , n42237 , n54616 );
not ( n23732 , n29614 );
and ( n23733 , n23732 , RI17497fe0_995);
and ( n23734 , n54617 , n29614 );
or ( n54618 , n23733 , n23734 );
not ( n23735 , RI1754c610_2);
and ( n23736 , n23735 , n54618 );
and ( n23737 , C0 , RI1754c610_2);
or ( n54619 , n23736 , n23737 );
buf ( n54620 , n54619 );
not ( n54621 , n33618 );
and ( n54622 , n54621 , n33698 );
xor ( n54623 , n44627 , n54622 );
not ( n23738 , n29614 );
and ( n23739 , n23738 , RI173e5a98_1636);
and ( n23740 , n54623 , n29614 );
or ( n54624 , n23739 , n23740 );
not ( n23741 , RI1754c610_2);
and ( n23742 , n23741 , n54624 );
and ( n23743 , C0 , RI1754c610_2);
or ( n54625 , n23742 , n23743 );
buf ( n54626 , n54625 );
not ( n54627 , n45025 );
and ( n54628 , n54627 , n37422 );
xor ( n54629 , n44237 , n54628 );
not ( n23744 , n29614 );
and ( n23745 , n23744 , RI17446c80_1391);
and ( n23746 , n54629 , n29614 );
or ( n54630 , n23745 , n23746 );
not ( n23747 , RI1754c610_2);
and ( n23748 , n23747 , n54630 );
and ( n23749 , C0 , RI1754c610_2);
or ( n54631 , n23748 , n23749 );
buf ( n54632 , n54631 );
not ( n54633 , n54146 );
and ( n54634 , n54633 , n49464 );
xor ( n54635 , n48117 , n54634 );
not ( n23750 , n29614 );
and ( n23751 , n23750 , RI173d0540_1740);
and ( n23752 , n54635 , n29614 );
or ( n54636 , n23751 , n23752 );
not ( n23753 , RI1754c610_2);
and ( n23754 , n23753 , n54636 );
and ( n23755 , C0 , RI1754c610_2);
or ( n54637 , n23754 , n23755 );
buf ( n54638 , n54637 );
not ( n54639 , n48180 );
and ( n54640 , n54639 , n48182 );
xor ( n54641 , n47311 , n54640 );
not ( n23756 , n29614 );
and ( n23757 , n23756 , RI17410ef0_1425);
and ( n23758 , n54641 , n29614 );
or ( n54642 , n23757 , n23758 );
not ( n23759 , RI1754c610_2);
and ( n23760 , n23759 , n54642 );
and ( n23761 , C0 , RI1754c610_2);
or ( n54643 , n23760 , n23761 );
buf ( n54644 , n54643 );
not ( n54645 , n50430 );
and ( n54646 , n54645 , n50464 );
xor ( n54647 , n50427 , n54646 );
not ( n23762 , n29614 );
and ( n23763 , n23762 , RI1748ceb0_1049);
and ( n23764 , n54647 , n29614 );
or ( n54648 , n23763 , n23764 );
not ( n23765 , RI1754c610_2);
and ( n23766 , n23765 , n54648 );
and ( n23767 , C0 , RI1754c610_2);
or ( n54649 , n23766 , n23767 );
buf ( n54650 , n54649 );
not ( n23768 , n27683 );
and ( n23769 , n23768 , RI19a8dfc8_2697);
and ( n23770 , RI19a98018_2626 , n27683 );
or ( n54651 , n23769 , n23770 );
not ( n23771 , RI1754c610_2);
and ( n23772 , n23771 , n54651 );
and ( n23773 , C0 , RI1754c610_2);
or ( n54652 , n23772 , n23773 );
buf ( n54653 , n54652 );
not ( n54654 , n38245 );
and ( n54655 , n54654 , n38250 );
xor ( n54656 , n43737 , n54655 );
not ( n23774 , n29614 );
and ( n23775 , n23774 , RI1738b378_2077);
and ( n23776 , n54656 , n29614 );
or ( n54657 , n23775 , n23776 );
not ( n23777 , RI1754c610_2);
and ( n23778 , n23777 , n54657 );
and ( n23779 , C0 , RI1754c610_2);
or ( n54658 , n23778 , n23779 );
buf ( n54659 , n54658 );
buf ( n54660 , RI1746d8a8_1202);
buf ( n54661 , RI17465220_1243);
not ( n54662 , n46802 );
and ( n54663 , n54662 , n46804 );
xor ( n54664 , n44903 , n54663 );
not ( n23780 , n29614 );
and ( n23781 , n23780 , RI173b5768_1871);
and ( n23782 , n54664 , n29614 );
or ( n54665 , n23781 , n23782 );
not ( n23783 , RI1754c610_2);
and ( n23784 , n23783 , n54665 );
and ( n23785 , C0 , RI1754c610_2);
or ( n54666 , n23784 , n23785 );
buf ( n54667 , n54666 );
not ( n54668 , n43337 );
and ( n54669 , n54668 , n43339 );
xor ( n54670 , n47288 , n54669 );
not ( n23786 , n29614 );
and ( n23787 , n23786 , RI1739d0f0_1990);
and ( n23788 , n54670 , n29614 );
or ( n54671 , n23787 , n23788 );
not ( n23789 , RI1754c610_2);
and ( n23790 , n23789 , n54671 );
and ( n23791 , C0 , RI1754c610_2);
or ( n54672 , n23790 , n23791 );
buf ( n54673 , n54672 );
not ( n23792 , n27683 );
and ( n23793 , n23792 , RI19ab6090_2408);
and ( n23794 , RI19abf4b0_2338 , n27683 );
or ( n54674 , n23793 , n23794 );
not ( n23795 , RI1754c610_2);
and ( n23796 , n23795 , n54674 );
and ( n23797 , C0 , RI1754c610_2);
or ( n54675 , n23796 , n23797 );
buf ( n54676 , n54675 );
not ( n54677 , n46746 );
and ( n54678 , n54677 , n43409 );
xor ( n54679 , n43556 , n54678 );
not ( n23798 , n29614 );
and ( n23799 , n23798 , RI173f4d68_1562);
and ( n23800 , n54679 , n29614 );
or ( n54680 , n23799 , n23800 );
not ( n23801 , RI1754c610_2);
and ( n23802 , n23801 , n54680 );
and ( n23803 , C0 , RI1754c610_2);
or ( n54681 , n23802 , n23803 );
buf ( n54682 , n54681 );
not ( n23804 , n27683 );
and ( n23805 , n23804 , RI19acfb30_2213);
and ( n23806 , RI19aa5a88_2525 , n27683 );
or ( n54683 , n23805 , n23806 );
not ( n23807 , RI1754c610_2);
and ( n23808 , n23807 , n54683 );
and ( n23809 , C0 , RI1754c610_2);
or ( n54684 , n23808 , n23809 );
buf ( n54685 , n54684 );
not ( n23810 , n27683 );
and ( n23811 , n23810 , RI19ac7d90_2271);
and ( n23812 , RI19a82b50_2775 , n27683 );
or ( n54686 , n23811 , n23812 );
not ( n23813 , RI1754c610_2);
and ( n23814 , n23813 , n54686 );
and ( n23815 , C0 , RI1754c610_2);
or ( n54687 , n23814 , n23815 );
buf ( n54688 , n54687 );
buf ( n54689 , RI17494b60_1011);
buf ( n54690 , RI174a4808_934);
buf ( n54691 , RI174ae8d0_885);
buf ( n54692 , RI174c1f98_807);
not ( n23816 , n27683 );
and ( n23817 , n23816 , RI19a85760_2756);
and ( n23818 , RI19a23330_2795 , n27683 );
or ( n54693 , n23817 , n23818 );
not ( n23819 , RI1754c610_2);
and ( n23820 , n23819 , n54693 );
and ( n23821 , C0 , RI1754c610_2);
or ( n54694 , n23820 , n23821 );
buf ( n54695 , n54694 );
buf ( n54696 , RI1749ef70_961);
not ( n54697 , n45651 );
and ( n54698 , n54697 , n51018 );
xor ( n54699 , n41964 , n54698 );
not ( n23822 , n29614 );
and ( n23823 , n23822 , RI174a8660_915);
and ( n23824 , n54699 , n29614 );
or ( n54700 , n23823 , n23824 );
not ( n23825 , RI1754c610_2);
and ( n23826 , n23825 , n54700 );
and ( n23827 , C0 , RI1754c610_2);
or ( n54701 , n23826 , n23827 );
buf ( n54702 , n54701 );
buf ( n54703 , RI174b4168_858);
not ( n54704 , n43695 );
xor ( n54705 , n34394 , n39989 );
xor ( n54706 , n54705 , n40009 );
and ( n54707 , n54704 , n54706 );
xor ( n54708 , n43692 , n54707 );
not ( n23828 , n29614 );
and ( n23829 , n23828 , RI1739d438_1989);
and ( n23830 , n54708 , n29614 );
or ( n54709 , n23829 , n23830 );
not ( n23831 , RI1754c610_2);
and ( n23832 , n23831 , n54709 );
and ( n23833 , C0 , RI1754c610_2);
or ( n54710 , n23832 , n23833 );
buf ( n54711 , n54710 );
not ( n54712 , n44935 );
and ( n54713 , n54712 , n48630 );
xor ( n54714 , n44932 , n54713 );
not ( n23834 , n29614 );
and ( n23835 , n23834 , RI1745fcd0_1269);
and ( n23836 , n54714 , n29614 );
or ( n54715 , n23835 , n23836 );
not ( n23837 , RI1754c610_2);
and ( n23838 , n23837 , n54715 );
and ( n23839 , C0 , RI1754c610_2);
or ( n54716 , n23838 , n23839 );
buf ( n54717 , n54716 );
not ( n54718 , n49183 );
and ( n54719 , n54718 , n47948 );
xor ( n54720 , n45488 , n54719 );
not ( n23840 , n29614 );
and ( n23841 , n23840 , RI17346fc0_2095);
and ( n23842 , n54720 , n29614 );
or ( n54721 , n23841 , n23842 );
not ( n23843 , RI1754c610_2);
and ( n23844 , n23843 , n54721 );
and ( n23845 , C0 , RI1754c610_2);
or ( n54722 , n23844 , n23845 );
buf ( n54723 , n54722 );
not ( n54724 , n47614 );
and ( n54725 , n54724 , n46573 );
xor ( n54726 , n47453 , n54725 );
not ( n23846 , n29614 );
and ( n23847 , n23846 , RI173fe7a0_1515);
and ( n23848 , n54726 , n29614 );
or ( n54727 , n23847 , n23848 );
not ( n23849 , RI1754c610_2);
and ( n23850 , n23849 , n54727 );
and ( n23851 , C0 , RI1754c610_2);
or ( n54728 , n23850 , n23851 );
buf ( n54729 , n54728 );
buf ( n54730 , RI174672f0_1233);
buf ( n54731 , RI17478d20_1147);
not ( n54732 , n48903 );
and ( n54733 , n54732 , n49908 );
xor ( n54734 , n48310 , n54733 );
not ( n23852 , n29614 );
and ( n23853 , n23852 , RI175014a8_756);
and ( n23854 , n54734 , n29614 );
or ( n54735 , n23853 , n23854 );
not ( n23855 , RI1754c610_2);
and ( n23856 , n23855 , n54735 );
and ( n23857 , C0 , RI1754c610_2);
or ( n54736 , n23856 , n23857 );
buf ( n54737 , n54736 );
not ( n54738 , n47989 );
and ( n54739 , n54738 , n52051 );
xor ( n54740 , n47986 , n54739 );
not ( n23858 , n29614 );
and ( n23859 , n23858 , RI17464b90_1245);
and ( n23860 , n54740 , n29614 );
or ( n54741 , n23859 , n23860 );
not ( n23861 , RI1754c610_2);
and ( n23862 , n23861 , n54741 );
and ( n23863 , C0 , RI1754c610_2);
or ( n54742 , n23862 , n23863 );
buf ( n54743 , n54742 );
and ( n54744 , RI1754bff8_15 , n34844 );
and ( n54745 , RI1754bff8_15 , n34847 );
and ( n54746 , RI1754bff8_15 , n34850 );
and ( n54747 , RI1754bff8_15 , n34852 );
and ( n54748 , RI1754bff8_15 , n34854 );
and ( n54749 , RI1754bff8_15 , n34856 );
or ( n54750 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , C0 , C0 );
not ( n23864 , n34859 );
and ( n23865 , n23864 , n54750 );
and ( n23866 , RI1754bff8_15 , n34859 );
or ( n54751 , n23865 , n23866 );
not ( n23867 , RI19a22f70_2797);
and ( n23868 , n23867 , n54751 );
and ( n23869 , C0 , RI19a22f70_2797);
or ( n54752 , n23868 , n23869 );
not ( n23870 , n27683 );
and ( n23871 , n23870 , RI19a91c40_2670);
and ( n23872 , n54752 , n27683 );
or ( n54753 , n23871 , n23872 );
not ( n23873 , RI1754c610_2);
and ( n23874 , n23873 , n54753 );
and ( n23875 , C0 , RI1754c610_2);
or ( n54754 , n23874 , n23875 );
buf ( n54755 , n54754 );
not ( n23876 , n27683 );
and ( n23877 , n23876 , RI19ab8d90_2389);
and ( n23878 , RI19ac1670_2319 , n27683 );
or ( n54756 , n23877 , n23878 );
not ( n23879 , RI1754c610_2);
and ( n23880 , n23879 , n54756 );
and ( n23881 , C0 , RI1754c610_2);
or ( n54757 , n23880 , n23881 );
buf ( n54758 , n54757 );
not ( n23882 , n27683 );
and ( n23883 , n23882 , RI19aa9868_2499);
and ( n23884 , RI19ab34f8_2429 , n27683 );
or ( n54759 , n23883 , n23884 );
not ( n23885 , RI1754c610_2);
and ( n23886 , n23885 , n54759 );
and ( n23887 , C0 , RI1754c610_2);
or ( n54760 , n23886 , n23887 );
buf ( n54761 , n54760 );
not ( n23888 , n27683 );
and ( n23889 , n23888 , RI19a90818_2679);
and ( n23890 , RI19a9a868_2608 , n27683 );
or ( n54762 , n23889 , n23890 );
not ( n23891 , RI1754c610_2);
and ( n23892 , n23891 , n54762 );
and ( n23893 , C0 , RI1754c610_2);
or ( n54763 , n23892 , n23893 );
buf ( n54764 , n54763 );
buf ( n54765 , n43086 );
not ( n23894 , n43088 );
and ( n23895 , n23894 , RI19a250b8_2781);
and ( n23896 , n54765 , n43088 );
or ( n54766 , n23895 , n23896 );
not ( n23897 , RI1754c610_2);
and ( n23898 , n23897 , n54766 );
and ( n23899 , C0 , RI1754c610_2);
or ( n54767 , n23898 , n23899 );
buf ( n54768 , n54767 );
buf ( n54769 , RI17495bc8_1006);
buf ( n54770 , RI1748d888_1046);
buf ( n54771 , RI174ccee8_773);
buf ( n54772 , RI174c62a0_794);
not ( n54773 , n50365 );
and ( n54774 , n54773 , n47181 );
xor ( n54775 , n41022 , n54774 );
not ( n23900 , n29614 );
and ( n23901 , n23900 , RI1749c4c8_974);
and ( n23902 , n54775 , n29614 );
or ( n54776 , n23901 , n23902 );
not ( n23903 , RI1754c610_2);
and ( n23904 , n23903 , n54776 );
and ( n23905 , C0 , RI1754c610_2);
or ( n54777 , n23904 , n23905 );
buf ( n54778 , n54777 );
not ( n54779 , n36149 );
and ( n54780 , n54779 , n36154 );
xor ( n54781 , n48643 , n54780 );
not ( n23906 , n29614 );
and ( n23907 , n23906 , RI1751ee90_670);
and ( n23908 , n54781 , n29614 );
or ( n54782 , n23907 , n23908 );
not ( n23909 , RI1754c610_2);
and ( n23910 , n23909 , n54782 );
and ( n23911 , C0 , RI1754c610_2);
or ( n54783 , n23910 , n23911 );
buf ( n54784 , n54783 );
not ( n54785 , n46783 );
and ( n54786 , n54785 , n51121 );
xor ( n54787 , n46780 , n54786 );
not ( n23912 , n29614 );
and ( n23913 , n23912 , RI1739d780_1988);
and ( n23914 , n54787 , n29614 );
or ( n54788 , n23913 , n23914 );
not ( n23915 , RI1754c610_2);
and ( n23916 , n23915 , n54788 );
and ( n23917 , C0 , RI1754c610_2);
or ( n54789 , n23916 , n23917 );
buf ( n54790 , n54789 );
not ( n54791 , n49409 );
and ( n54792 , n54791 , n45962 );
xor ( n54793 , n36875 , n54792 );
not ( n23918 , n29614 );
and ( n23919 , n23918 , RI1739dac8_1987);
and ( n23920 , n54793 , n29614 );
or ( n54794 , n23919 , n23920 );
not ( n23921 , RI1754c610_2);
and ( n23922 , n23921 , n54794 );
and ( n23923 , C0 , RI1754c610_2);
or ( n54795 , n23922 , n23923 );
buf ( n54796 , n54795 );
not ( n23924 , n27683 );
and ( n23925 , n23924 , RI19a998f0_2615);
and ( n23926 , RI19aa3238_2544 , n27683 );
or ( n54797 , n23925 , n23926 );
not ( n23927 , RI1754c610_2);
and ( n23928 , n23927 , n54797 );
and ( n23929 , C0 , RI1754c610_2);
or ( n54798 , n23928 , n23929 );
buf ( n54799 , n54798 );
not ( n23930 , n27683 );
and ( n23931 , n23930 , RI19a8cfd8_2704);
and ( n23932 , RI19a97208_2632 , n27683 );
or ( n54800 , n23931 , n23932 );
not ( n23933 , RI1754c610_2);
and ( n23934 , n23933 , n54800 );
and ( n23935 , C0 , RI1754c610_2);
or ( n54801 , n23934 , n23935 );
buf ( n54802 , n54801 );
not ( n54803 , n48345 );
and ( n54804 , n54803 , n47602 );
xor ( n54805 , n48342 , n54804 );
not ( n23936 , n29614 );
and ( n23937 , n23936 , RI173cfb68_1743);
and ( n23938 , n54805 , n29614 );
or ( n54806 , n23937 , n23938 );
not ( n23939 , RI1754c610_2);
and ( n23940 , n23939 , n54806 );
and ( n23941 , C0 , RI1754c610_2);
or ( n54807 , n23940 , n23941 );
buf ( n54808 , n54807 );
not ( n54809 , n44333 );
and ( n54810 , n54809 , n44335 );
xor ( n54811 , n50561 , n54810 );
not ( n23942 , n29614 );
and ( n23943 , n23942 , RI173b22e8_1887);
and ( n23944 , n54811 , n29614 );
or ( n54812 , n23943 , n23944 );
not ( n23945 , RI1754c610_2);
and ( n23946 , n23945 , n54812 );
and ( n23947 , C0 , RI1754c610_2);
or ( n54813 , n23946 , n23947 );
buf ( n54814 , n54813 );
not ( n54815 , n43901 );
and ( n54816 , n54815 , n43903 );
xor ( n54817 , n43802 , n54816 );
not ( n23948 , n29614 );
and ( n23949 , n23948 , RI173ad428_1911);
and ( n23950 , n54817 , n29614 );
or ( n54818 , n23949 , n23950 );
not ( n23951 , RI1754c610_2);
and ( n23952 , n23951 , n54818 );
and ( n23953 , C0 , RI1754c610_2);
or ( n54819 , n23952 , n23953 );
buf ( n54820 , n54819 );
not ( n23954 , n27683 );
and ( n23955 , n23954 , RI19a9aac0_2607);
and ( n23956 , RI19aa44f8_2535 , n27683 );
or ( n54821 , n23955 , n23956 );
not ( n23957 , RI1754c610_2);
and ( n23958 , n23957 , n54821 );
and ( n23959 , C0 , RI1754c610_2);
or ( n54822 , n23958 , n23959 );
buf ( n54823 , n54822 );
not ( n54824 , n43611 );
and ( n54825 , n54824 , n43613 );
xor ( n54826 , n42636 , n54825 );
not ( n23960 , n29614 );
and ( n23961 , n23960 , RI174609f0_1265);
and ( n23962 , n54826 , n29614 );
or ( n54827 , n23961 , n23962 );
not ( n23963 , RI1754c610_2);
and ( n23964 , n23963 , n54827 );
and ( n23965 , C0 , RI1754c610_2);
or ( n54828 , n23964 , n23965 );
buf ( n54829 , n54828 );
not ( n54830 , n51086 );
and ( n54831 , n54830 , n47634 );
xor ( n54832 , n49095 , n54831 );
not ( n23966 , n29614 );
and ( n23967 , n23966 , RI1752fab0_618);
and ( n23968 , n54832 , n29614 );
or ( n54833 , n23967 , n23968 );
not ( n23969 , RI1754c610_2);
and ( n23970 , n23969 , n54833 );
and ( n23971 , C0 , RI1754c610_2);
or ( n54834 , n23970 , n23971 );
buf ( n54835 , n54834 );
not ( n54836 , n51282 );
and ( n54837 , n54836 , n51284 );
xor ( n54838 , n44176 , n54837 );
not ( n23972 , n29614 );
and ( n23973 , n23972 , RI1740f168_1434);
and ( n23974 , n54838 , n29614 );
or ( n54839 , n23973 , n23974 );
not ( n23975 , RI1754c610_2);
and ( n23976 , n23975 , n54839 );
and ( n23977 , C0 , RI1754c610_2);
or ( n54840 , n23976 , n23977 );
buf ( n54841 , n54840 );
not ( n54842 , n40320 );
and ( n54843 , n54842 , n50728 );
xor ( n54844 , n40285 , n54843 );
not ( n23978 , n29614 );
and ( n23979 , n23978 , RI174765c0_1159);
and ( n23980 , n54844 , n29614 );
or ( n54845 , n23979 , n23980 );
not ( n23981 , RI1754c610_2);
and ( n23982 , n23981 , n54845 );
and ( n23983 , C0 , RI1754c610_2);
or ( n54846 , n23982 , n23983 );
buf ( n54847 , n54846 );
not ( n54848 , n40860 );
and ( n54849 , n54848 , n44645 );
xor ( n54850 , n40857 , n54849 );
or ( n54851 , n27689 , RI175385e8_592);
or ( n54852 , n54851 , RI17537fd0_593);
or ( n54853 , n54852 , RI175379b8_594);
or ( n54854 , n54853 , RI17536d88_596);
xor ( n54855 , n54850 , n54854 );
not ( n23984 , n29614 );
and ( n23985 , n23984 , RI1746f2e8_1194);
and ( n23986 , n54855 , n29614 );
or ( n54856 , n23985 , n23986 );
not ( n23987 , RI1754c610_2);
and ( n23988 , n23987 , n54856 );
and ( n23989 , C0 , RI1754c610_2);
or ( n54857 , n23988 , n23989 );
buf ( n54858 , n54857 );
not ( n54859 , n51018 );
and ( n54860 , n54859 , n41959 );
xor ( n54861 , n45651 , n54860 );
not ( n23990 , n29614 );
and ( n23991 , n23990 , RI1746df38_1200);
and ( n23992 , n54861 , n29614 );
or ( n54862 , n23991 , n23992 );
not ( n23993 , RI1754c610_2);
and ( n23994 , n23993 , n54862 );
and ( n23995 , C0 , RI1754c610_2);
or ( n54863 , n23994 , n23995 );
buf ( n54864 , n54863 );
not ( n23996 , n27683 );
and ( n23997 , n23996 , RI19ac7250_2276);
and ( n23998 , RI19acfd88_2212 , n27683 );
or ( n54865 , n23997 , n23998 );
not ( n23999 , RI1754c610_2);
and ( n24000 , n23999 , n54865 );
and ( n24001 , C0 , RI1754c610_2);
or ( n54866 , n24000 , n24001 );
buf ( n54867 , n54866 );
buf ( n54868 , RI174a68d8_924);
not ( n54869 , n38952 );
and ( n54870 , n54869 , n44004 );
xor ( n54871 , n38949 , n54870 );
not ( n24002 , n29614 );
and ( n24003 , n24002 , RI174b44b0_857);
and ( n24004 , n54871 , n29614 );
or ( n54872 , n24003 , n24004 );
not ( n24005 , RI1754c610_2);
and ( n24006 , n24005 , n54872 );
and ( n24007 , C0 , RI1754c610_2);
or ( n54873 , n24006 , n24007 );
buf ( n54874 , n54873 );
not ( n54875 , n49464 );
and ( n54876 , n54875 , n48112 );
xor ( n54877 , n54146 , n54876 );
not ( n24008 , n29614 );
and ( n24009 , n24008 , RI173deb08_1670);
and ( n24010 , n54877 , n29614 );
or ( n54878 , n24009 , n24010 );
not ( n24011 , RI1754c610_2);
and ( n24012 , n24011 , n54878 );
and ( n24013 , C0 , RI1754c610_2);
or ( n54879 , n24012 , n24013 );
buf ( n54880 , n54879 );
buf ( n54881 , RI174acb48_894);
not ( n24014 , n27683 );
and ( n24015 , n24014 , RI19aa5dd0_2524);
and ( n24016 , RI19ab0000_2454 , n27683 );
or ( n54882 , n24015 , n24016 );
not ( n24017 , RI1754c610_2);
and ( n24018 , n24017 , n54882 );
and ( n24019 , C0 , RI1754c610_2);
or ( n54883 , n24018 , n24019 );
buf ( n54884 , n54883 );
not ( n54885 , n41717 );
and ( n54886 , n54885 , n45385 );
xor ( n54887 , n41714 , n54886 );
not ( n24020 , n29614 );
and ( n24021 , n24020 , RI173aee68_1903);
and ( n24022 , n54887 , n29614 );
or ( n54888 , n24021 , n24022 );
not ( n24023 , RI1754c610_2);
and ( n24024 , n24023 , n54888 );
and ( n24025 , C0 , RI1754c610_2);
or ( n54889 , n24024 , n24025 );
buf ( n54890 , n54889 );
not ( n54891 , n48412 );
and ( n54892 , n54891 , n48266 );
xor ( n54893 , n40217 , n54892 );
not ( n24026 , n29614 );
and ( n24027 , n24026 , RI1748aa98_1060);
and ( n24028 , n54893 , n29614 );
or ( n54894 , n24027 , n24028 );
not ( n24029 , RI1754c610_2);
and ( n24030 , n24029 , n54894 );
and ( n24031 , C0 , RI1754c610_2);
or ( n54895 , n24030 , n24031 );
buf ( n54896 , n54895 );
not ( n24032 , n27683 );
and ( n24033 , n24032 , RI19ac6080_2284);
and ( n24034 , RI19aced20_2219 , n27683 );
or ( n54897 , n24033 , n24034 );
not ( n24035 , RI1754c610_2);
and ( n24036 , n24035 , n54897 );
and ( n24037 , C0 , RI1754c610_2);
or ( n54898 , n24036 , n24037 );
buf ( n54899 , n54898 );
not ( n54900 , n42636 );
and ( n54901 , n54900 , n43611 );
xor ( n54902 , n42620 , n54901 );
not ( n24038 , n29614 );
and ( n24039 , n24038 , RI174520f8_1336);
and ( n24040 , n54902 , n29614 );
or ( n54903 , n24039 , n24040 );
not ( n24041 , RI1754c610_2);
and ( n24042 , n24041 , n54903 );
and ( n24043 , C0 , RI1754c610_2);
or ( n54904 , n24042 , n24043 );
buf ( n54905 , n54904 );
not ( n54906 , n49505 );
and ( n54907 , n54906 , n51312 );
xor ( n54908 , n49297 , n54907 );
not ( n24044 , n29614 );
and ( n24045 , n24044 , RI173c1900_1812);
and ( n24046 , n54908 , n29614 );
or ( n54909 , n24045 , n24046 );
not ( n24047 , RI1754c610_2);
and ( n24048 , n24047 , n54909 );
and ( n24049 , C0 , RI1754c610_2);
or ( n54910 , n24048 , n24049 );
buf ( n54911 , n54910 );
not ( n54912 , n47888 );
and ( n54913 , n54912 , n51997 );
xor ( n54914 , n45927 , n54913 );
not ( n24050 , n29614 );
and ( n24051 , n24050 , RI17508ff0_738);
and ( n24052 , n54914 , n29614 );
or ( n54915 , n24051 , n24052 );
not ( n24053 , RI1754c610_2);
and ( n24054 , n24053 , n54915 );
and ( n24055 , C0 , RI1754c610_2);
or ( n54916 , n24054 , n24055 );
buf ( n54917 , n54916 );
not ( n54918 , n44432 );
and ( n54919 , n54918 , n44434 );
xor ( n54920 , n46442 , n54919 );
not ( n24056 , n29614 );
and ( n24057 , n24056 , RI17487618_1076);
and ( n24058 , n54920 , n29614 );
or ( n54921 , n24057 , n24058 );
not ( n24059 , RI1754c610_2);
and ( n24060 , n24059 , n54921 );
and ( n24061 , C0 , RI1754c610_2);
or ( n54922 , n24060 , n24061 );
buf ( n54923 , n54922 );
and ( n54924 , RI1754b698_35 , n34844 );
and ( n54925 , RI1754b698_35 , n34847 );
and ( n54926 , RI1754b698_35 , n34850 );
or ( n54927 , n54924 , n54925 , n54926 , C0 , C0 , C0 , C0 , C0 );
not ( n24062 , n34859 );
and ( n24063 , n24062 , n54927 );
and ( n24064 , RI1754b698_35 , n34859 );
or ( n54928 , n24063 , n24064 );
not ( n24065 , RI19a22f70_2797);
and ( n24066 , n24065 , n54928 );
and ( n24067 , C0 , RI19a22f70_2797);
or ( n54929 , n24066 , n24067 );
not ( n24068 , n27683 );
and ( n24069 , n24068 , RI19ab0c30_2448);
and ( n24070 , n54929 , n27683 );
or ( n54930 , n24069 , n24070 );
not ( n24071 , RI1754c610_2);
and ( n24072 , n24071 , n54930 );
and ( n24073 , C0 , RI1754c610_2);
or ( n54931 , n24072 , n24073 );
buf ( n54932 , n54931 );
not ( n24074 , n27683 );
and ( n24075 , n24074 , RI19abbc70_2369);
and ( n24076 , RI19ac4280_2298 , n27683 );
or ( n54933 , n24075 , n24076 );
not ( n24077 , RI1754c610_2);
and ( n24078 , n24077 , n54933 );
and ( n24079 , C0 , RI1754c610_2);
or ( n54934 , n24078 , n24079 );
buf ( n54935 , n54934 );
not ( n24080 , n27683 );
and ( n24081 , n24080 , RI19aa6988_2519);
and ( n24082 , RI19ab0a50_2449 , n27683 );
or ( n54936 , n24081 , n24082 );
not ( n24083 , RI1754c610_2);
and ( n24084 , n24083 , n54936 );
and ( n24085 , C0 , RI1754c610_2);
or ( n54937 , n24084 , n24085 );
buf ( n54938 , n54937 );
not ( n54939 , n42125 );
and ( n54940 , n54939 , n41571 );
xor ( n54941 , n45239 , n54940 );
not ( n24086 , n29614 );
and ( n24087 , n24086 , RI173892a8_2087);
and ( n24088 , n54941 , n29614 );
or ( n54942 , n24087 , n24088 );
not ( n24089 , RI1754c610_2);
and ( n24090 , n24089 , n54942 );
and ( n24091 , C0 , RI1754c610_2);
or ( n54943 , n24090 , n24091 );
buf ( n54944 , n54943 );
buf ( n54945 , RI17475210_1165);
not ( n24092 , n27683 );
and ( n24093 , n24092 , RI19a91808_2672);
and ( n24094 , RI19a9bb28_2600 , n27683 );
or ( n54946 , n24093 , n24094 );
not ( n24095 , RI1754c610_2);
and ( n24096 , n24095 , n54946 );
and ( n24097 , C0 , RI1754c610_2);
or ( n54947 , n24096 , n24097 );
buf ( n54948 , n54947 );
not ( n54949 , n44483 );
and ( n54950 , n54949 , n34671 );
xor ( n54951 , n47866 , n54950 );
not ( n24098 , n29614 );
and ( n24099 , n24098 , RI173ef4d0_1589);
and ( n24100 , n54951 , n29614 );
or ( n54952 , n24099 , n24100 );
not ( n24101 , RI1754c610_2);
and ( n24102 , n24101 , n54952 );
and ( n24103 , C0 , RI1754c610_2);
or ( n54953 , n24102 , n24103 );
buf ( n54954 , n54953 );
not ( n54955 , n47595 );
and ( n54956 , n54955 , n37170 );
xor ( n54957 , n46020 , n54956 );
not ( n24104 , n29614 );
and ( n24105 , n24104 , RI173e74d8_1628);
and ( n24106 , n54957 , n29614 );
or ( n54958 , n24105 , n24106 );
not ( n24107 , RI1754c610_2);
and ( n24108 , n24107 , n54958 );
and ( n24109 , C0 , RI1754c610_2);
or ( n54959 , n24108 , n24109 );
buf ( n54960 , n54959 );
not ( n54961 , n44722 );
and ( n54962 , n54961 , n44058 );
xor ( n54963 , n38373 , n54962 );
not ( n24110 , n29614 );
and ( n24111 , n24110 , RI1750a9b8_733);
and ( n24112 , n54963 , n29614 );
or ( n54964 , n24111 , n24112 );
not ( n24113 , RI1754c610_2);
and ( n24114 , n24113 , n54964 );
and ( n24115 , C0 , RI1754c610_2);
or ( n54965 , n24114 , n24115 );
buf ( n54966 , n54965 );
not ( n24116 , n27683 );
and ( n24117 , n24116 , RI19a9c398_2596);
and ( n24118 , RI19aa5dd0_2524 , n27683 );
or ( n54967 , n24117 , n24118 );
not ( n24119 , RI1754c610_2);
and ( n24120 , n24119 , n54967 );
and ( n24121 , C0 , RI1754c610_2);
or ( n54968 , n24120 , n24121 );
buf ( n54969 , n54968 );
not ( n54970 , n52768 );
and ( n54971 , n54970 , n51561 );
xor ( n54972 , n42485 , n54971 );
not ( n24122 , n29614 );
and ( n24123 , n24122 , RI173c6b08_1787);
and ( n24124 , n54972 , n29614 );
or ( n54973 , n24123 , n24124 );
not ( n24125 , RI1754c610_2);
and ( n24126 , n24125 , n54973 );
and ( n24127 , C0 , RI1754c610_2);
or ( n54974 , n24126 , n24127 );
buf ( n54975 , n54974 );
not ( n54976 , n38821 );
and ( n54977 , n54976 , n43138 );
xor ( n54978 , n38818 , n54977 );
not ( n24128 , n29614 );
and ( n24129 , n24128 , RI1733b170_2153);
and ( n24130 , n54978 , n29614 );
or ( n54979 , n24129 , n24130 );
not ( n24131 , RI1754c610_2);
and ( n24132 , n24131 , n54979 );
and ( n24133 , C0 , RI1754c610_2);
or ( n54980 , n24132 , n24133 );
buf ( n54981 , n54980 );
not ( n54982 , n46111 );
and ( n54983 , n54982 , n46113 );
xor ( n54984 , n48894 , n54983 );
not ( n24134 , n29614 );
and ( n24135 , n24134 , RI1738cdb8_2069);
and ( n24136 , n54984 , n29614 );
or ( n54985 , n24135 , n24136 );
not ( n24137 , RI1754c610_2);
and ( n24138 , n24137 , n54985 );
and ( n24139 , C0 , RI1754c610_2);
or ( n54986 , n24138 , n24139 );
buf ( n54987 , n54986 );
not ( n24140 , RI1754c610_2);
and ( n24141 , n24140 , RI19ad1c18_2200);
and ( n24142 , C0 , RI1754c610_2);
or ( n54988 , n24141 , n24142 );
buf ( n54989 , n54988 );
xor ( n54990 , n39608 , n35272 );
xor ( n54991 , n54990 , n35009 );
not ( n54992 , n54991 );
and ( n54993 , n54992 , n52181 );
xor ( n54994 , n52989 , n54993 );
not ( n24143 , n29614 );
and ( n24144 , n24143 , RI175361d0_598);
and ( n24145 , n54994 , n29614 );
or ( n54995 , n24144 , n24145 );
not ( n24146 , RI1754c610_2);
and ( n24147 , n24146 , n54995 );
and ( n24148 , C0 , RI1754c610_2);
or ( n54996 , n24147 , n24148 );
buf ( n54997 , n54996 );
not ( n54998 , n40867 );
and ( n54999 , n54998 , n40869 );
xor ( n55000 , n44185 , n54999 );
not ( n24149 , n29614 );
and ( n24150 , n24149 , RI17490330_1033);
and ( n24151 , n55000 , n29614 );
or ( n55001 , n24150 , n24151 );
not ( n24152 , RI1754c610_2);
and ( n24153 , n24152 , n55001 );
and ( n24154 , C0 , RI1754c610_2);
or ( n55002 , n24153 , n24154 );
buf ( n55003 , n55002 );
and ( n55004 , RI1754c520_4 , n34844 );
and ( n55005 , RI1754c520_4 , n34847 );
and ( n55006 , RI1754c520_4 , n34850 );
and ( n55007 , RI1754c520_4 , n34852 );
and ( n55008 , RI1754c520_4 , n34854 );
and ( n55009 , RI1754c520_4 , n34856 );
and ( n55010 , RI1754c520_4 , n39233 );
or ( n55011 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , C0 );
not ( n24155 , n34859 );
and ( n24156 , n24155 , n55011 );
and ( n24157 , RI1754c520_4 , n34859 );
or ( n55012 , n24156 , n24157 );
not ( n24158 , RI19a22f70_2797);
and ( n24159 , n24158 , n55012 );
and ( n24160 , C0 , RI19a22f70_2797);
or ( n55013 , n24159 , n24160 );
not ( n24161 , n27683 );
and ( n24162 , n24161 , RI19a88028_2738);
and ( n24163 , n55013 , n27683 );
or ( n55014 , n24162 , n24163 );
not ( n24164 , RI1754c610_2);
and ( n24165 , n24164 , n55014 );
and ( n24166 , C0 , RI1754c610_2);
or ( n55015 , n24165 , n24166 );
buf ( n55016 , n55015 );
not ( n24167 , n27683 );
and ( n24168 , n24167 , RI19abad70_2375);
and ( n24169 , RI19ac34e8_2304 , n27683 );
or ( n55017 , n24168 , n24169 );
not ( n24170 , RI1754c610_2);
and ( n24171 , n24170 , n55017 );
and ( n24172 , C0 , RI1754c610_2);
or ( n55018 , n24171 , n24172 );
buf ( n55019 , n55018 );
not ( n55020 , n44476 );
and ( n55021 , n55020 , n44942 );
xor ( n55022 , n44473 , n55021 );
not ( n24173 , n29614 );
and ( n24174 , n24173 , RI174ca080_782);
and ( n24175 , n55022 , n29614 );
or ( n55023 , n24174 , n24175 );
not ( n24176 , RI1754c610_2);
and ( n24177 , n24176 , n55023 );
and ( n24178 , C0 , RI1754c610_2);
or ( n55024 , n24177 , n24178 );
buf ( n55025 , n55024 );
not ( n55026 , n46372 );
and ( n55027 , n55026 , n45279 );
xor ( n55028 , n47761 , n55027 );
not ( n24179 , n29614 );
and ( n24180 , n24179 , RI1744c1d0_1365);
and ( n24181 , n55028 , n29614 );
or ( n55029 , n24180 , n24181 );
not ( n24182 , RI1754c610_2);
and ( n24183 , n24182 , n55029 );
and ( n24184 , C0 , RI1754c610_2);
or ( n55030 , n24183 , n24184 );
buf ( n55031 , n55030 );
not ( n55032 , n51460 );
and ( n55033 , n55032 , n29982 );
xor ( n55034 , n53466 , n55033 );
not ( n24185 , n29614 );
and ( n24186 , n24185 , RI173ab6a0_1920);
and ( n24187 , n55034 , n29614 );
or ( n55035 , n24186 , n24187 );
not ( n24188 , RI1754c610_2);
and ( n24189 , n24188 , n55035 );
and ( n24190 , C0 , RI1754c610_2);
or ( n55036 , n24189 , n24190 );
buf ( n55037 , n55036 );
not ( n55038 , n51076 );
and ( n55039 , n55038 , n51078 );
xor ( n55040 , n45721 , n55039 );
not ( n24191 , n29614 );
and ( n24192 , n24191 , RI17517d20_692);
and ( n24193 , n55040 , n29614 );
or ( n55041 , n24192 , n24193 );
not ( n24194 , RI1754c610_2);
and ( n24195 , n24194 , n55041 );
and ( n24196 , C0 , RI1754c610_2);
or ( n55042 , n24195 , n24196 );
buf ( n55043 , n55042 );
and ( n55044 , RI1754b968_29 , n34844 );
and ( n55045 , RI1754b968_29 , n34847 );
and ( n55046 , RI1754b968_29 , n34850 );
and ( n55047 , RI1754b968_29 , n34852 );
or ( n55048 , n55044 , n55045 , n55046 , n55047 , C0 , C0 , C0 , C0 );
not ( n24197 , n34859 );
and ( n24198 , n24197 , n55048 );
and ( n24199 , RI1754b968_29 , n34859 );
or ( n55049 , n24198 , n24199 );
not ( n24200 , RI19a22f70_2797);
and ( n24201 , n24200 , n55049 );
and ( n24202 , C0 , RI19a22f70_2797);
or ( n55050 , n24201 , n24202 );
not ( n24203 , n27683 );
and ( n24204 , n24203 , RI19aa7540_2514);
and ( n24205 , n55050 , n27683 );
or ( n55051 , n24204 , n24205 );
not ( n24206 , RI1754c610_2);
and ( n24207 , n24206 , n55051 );
and ( n24208 , C0 , RI1754c610_2);
or ( n55052 , n24207 , n24208 );
buf ( n55053 , n55052 );
not ( n24209 , n27683 );
and ( n24210 , n24209 , RI19acdcb8_2226);
and ( n24211 , RI19a91c40_2670 , n27683 );
or ( n55054 , n24210 , n24211 );
not ( n24212 , RI1754c610_2);
and ( n24213 , n24212 , n55054 );
and ( n24214 , C0 , RI1754c610_2);
or ( n55055 , n24213 , n24214 );
buf ( n55056 , n55055 );
not ( n24215 , n27683 );
and ( n24216 , n24215 , RI19a94490_2652);
and ( n24217 , RI19a9e8a0_2580 , n27683 );
or ( n55057 , n24216 , n24217 );
not ( n24218 , RI1754c610_2);
and ( n24219 , n24218 , n55057 );
and ( n24220 , C0 , RI1754c610_2);
or ( n55058 , n24219 , n24220 );
buf ( n55059 , n55058 );
buf ( n55060 , RI17483478_1096);
not ( n55061 , n36885 );
and ( n55062 , n55061 , n36892 );
xor ( n55063 , n52411 , n55062 );
not ( n24221 , n29614 );
and ( n24222 , n24221 , RI174458d0_1397);
and ( n24223 , n55063 , n29614 );
or ( n55064 , n24222 , n24223 );
not ( n24224 , RI1754c610_2);
and ( n24225 , n24224 , n55064 );
and ( n24226 , C0 , RI1754c610_2);
or ( n55065 , n24225 , n24226 );
buf ( n55066 , n55065 );
buf ( n55067 , RI17513f40_704);
buf ( n55068 , RI17461a58_1260);
not ( n55069 , n41431 );
and ( n55070 , n55069 , n41433 );
xor ( n55071 , n49021 , n55070 );
not ( n24227 , n29614 );
and ( n24228 , n24227 , RI173a15d8_1969);
and ( n24229 , n55071 , n29614 );
or ( n55072 , n24228 , n24229 );
not ( n24230 , RI1754c610_2);
and ( n24231 , n24230 , n55072 );
and ( n24232 , C0 , RI1754c610_2);
or ( n55073 , n24231 , n24232 );
buf ( n55074 , n55073 );
not ( n55075 , n46104 );
and ( n55076 , n55075 , n43957 );
xor ( n55077 , n46101 , n55076 );
not ( n24233 , n29614 );
and ( n24234 , n24233 , RI174b72a0_843);
and ( n24235 , n55077 , n29614 );
or ( n55078 , n24234 , n24235 );
not ( n24236 , RI1754c610_2);
and ( n24237 , n24236 , n55078 );
and ( n24238 , C0 , RI1754c610_2);
or ( n55079 , n24237 , n24238 );
buf ( n55080 , n55079 );
not ( n55081 , n52755 );
and ( n55082 , n55081 , n47255 );
xor ( n55083 , n38595 , n55082 );
not ( n24239 , n29614 );
and ( n24240 , n24239 , RI1740ddb8_1440);
and ( n24241 , n55083 , n29614 );
or ( n55084 , n24240 , n24241 );
not ( n24242 , RI1754c610_2);
and ( n24243 , n24242 , n55084 );
and ( n24244 , C0 , RI1754c610_2);
or ( n55085 , n24243 , n24244 );
buf ( n55086 , n55085 );
not ( n55087 , n39093 );
and ( n55088 , n55087 , n39095 );
xor ( n55089 , n45217 , n55088 );
not ( n24245 , n29614 );
and ( n24246 , n24245 , RI173a7b90_1938);
and ( n24247 , n55089 , n29614 );
or ( n55090 , n24246 , n24247 );
not ( n24248 , RI1754c610_2);
and ( n24249 , n24248 , n55090 );
and ( n24250 , C0 , RI1754c610_2);
or ( n55091 , n24249 , n24250 );
buf ( n55092 , n55091 );
not ( n55093 , n42388 );
and ( n55094 , n55093 , n32974 );
xor ( n55095 , n48986 , n55094 );
not ( n24251 , n29614 );
and ( n24252 , n24251 , RI17337cf0_2169);
and ( n24253 , n55095 , n29614 );
or ( n55096 , n24252 , n24253 );
not ( n24254 , RI1754c610_2);
and ( n24255 , n24254 , n55096 );
and ( n24256 , C0 , RI1754c610_2);
or ( n55097 , n24255 , n24256 );
buf ( n55098 , n55097 );
not ( n55099 , n38602 );
and ( n55100 , n55099 , n38604 );
xor ( n55101 , n44811 , n55100 );
not ( n24257 , n29614 );
and ( n24258 , n24257 , RI17479a40_1143);
and ( n24259 , n55101 , n29614 );
or ( n55102 , n24258 , n24259 );
not ( n24260 , RI1754c610_2);
and ( n24261 , n24260 , n55102 );
and ( n24262 , C0 , RI1754c610_2);
or ( n55103 , n24261 , n24262 );
buf ( n55104 , n55103 );
buf ( n55105 , RI1748ef80_1039);
not ( n55106 , n37923 );
and ( n55107 , n55106 , n37944 );
xor ( n55108 , n43327 , n55107 );
not ( n24263 , n29614 );
and ( n24264 , n24263 , RI1744a790_1373);
and ( n24265 , n55108 , n29614 );
or ( n55109 , n24264 , n24265 );
not ( n24266 , RI1754c610_2);
and ( n24267 , n24266 , n55109 );
and ( n24268 , C0 , RI1754c610_2);
or ( n55110 , n24267 , n24268 );
buf ( n55111 , n55110 );
not ( n55112 , n44930 );
and ( n55113 , n55112 , n44932 );
xor ( n55114 , n48633 , n55113 );
not ( n24269 , n29614 );
and ( n24270 , n24269 , RI17413ce0_1411);
and ( n24271 , n55114 , n29614 );
or ( n55115 , n24270 , n24271 );
not ( n24272 , RI1754c610_2);
and ( n24273 , n24272 , n55115 );
and ( n24274 , C0 , RI1754c610_2);
or ( n55116 , n24273 , n24274 );
buf ( n55117 , n55116 );
buf ( n55118 , RI174caff8_779);
not ( n55119 , n51199 );
and ( n55120 , n55119 , n48209 );
xor ( n55121 , n48029 , n55120 );
not ( n24275 , n29614 );
and ( n24276 , n24275 , RI173a3360_1960);
and ( n24277 , n55121 , n29614 );
or ( n55122 , n24276 , n24277 );
not ( n24278 , RI1754c610_2);
and ( n24279 , n24278 , n55122 );
and ( n24280 , C0 , RI1754c610_2);
or ( n55123 , n24279 , n24280 );
buf ( n55124 , n55123 );
buf ( n55125 , RI17473b18_1172);
not ( n24281 , n27683 );
and ( n24282 , n24281 , RI19ac9b90_2257);
and ( n24283 , RI19a84e00_2760 , n27683 );
or ( n55126 , n24282 , n24283 );
not ( n24284 , RI1754c610_2);
and ( n24285 , n24284 , n55126 );
and ( n24286 , C0 , RI1754c610_2);
or ( n55127 , n24285 , n24286 );
buf ( n55128 , n55127 );
not ( n55129 , n40070 );
and ( n55130 , n55129 , n44662 );
xor ( n55131 , n40064 , n55130 );
not ( n24287 , n29614 );
and ( n24288 , n24287 , RI1750c380_728);
and ( n24289 , n55131 , n29614 );
or ( n55132 , n24288 , n24289 );
not ( n24290 , RI1754c610_2);
and ( n24291 , n24290 , n55132 );
and ( n24292 , C0 , RI1754c610_2);
or ( n55133 , n24291 , n24292 );
buf ( n55134 , n55133 );
not ( n55135 , n48375 );
and ( n55136 , n55135 , n48377 );
xor ( n55137 , n51422 , n55136 );
not ( n24293 , n29614 );
and ( n24294 , n24293 , RI1740e790_1437);
and ( n24295 , n55137 , n29614 );
or ( n55138 , n24294 , n24295 );
not ( n24296 , RI1754c610_2);
and ( n24297 , n24296 , n55138 );
and ( n24298 , C0 , RI1754c610_2);
or ( n55139 , n24297 , n24298 );
buf ( n55140 , n55139 );
not ( n55141 , n35274 );
and ( n55142 , n55141 , n46235 );
xor ( n55143 , n35217 , n55142 );
not ( n24299 , n29614 );
and ( n24300 , n24299 , RI17359008_2091);
and ( n24301 , n55143 , n29614 );
or ( n55144 , n24300 , n24301 );
not ( n24302 , RI1754c610_2);
and ( n24303 , n24302 , n55144 );
and ( n24304 , C0 , RI1754c610_2);
or ( n55145 , n24303 , n24304 );
buf ( n55146 , n55145 );
not ( n55147 , n41160 );
and ( n55148 , n55147 , n41165 );
xor ( n55149 , n44410 , n55148 );
not ( n24305 , n29614 );
and ( n24306 , n24305 , RI173f4a20_1563);
and ( n24307 , n55149 , n29614 );
xor ( n55150 , n24306 , n24307 );
not ( n24308 , RI1754c610_2);
nand ( n24309 , n24308 , n55150 );
nand ( n24310 , C0 , RI1754c610_2);
nor ( n55151 , n24309 , n24310 );
buf ( n55152 , n55151 );
not ( n24311 , n27683 );
nand ( n24312 , n24311 , RI19aaac18_2490);
nand ( n24313 , RI19ab48a8_2419 , n27683 );
nor ( n55153 , n24312 , n24313 );
not ( n24314 , RI1754c610_2);
nand ( n24315 , n24314 , n55153 );
nand ( n24316 , C0 , RI1754c610_2);
xor ( n55154 , n24315 , n24316 );
buf ( n55155 , n55154 );
not ( n55156 , RI174a89a8_914);
buf ( n55157 , RI174aaa78_904);
not ( n55158 , n49916 );
and ( n55159 , n55158 , n49065 );
xor ( n55160 , n52503 , n55159 );
not ( n24317 , n29614 );
and ( n24318 , n24317 , RI173fcd60_1523);
and ( n24319 , n55160 , n29614 );
or ( n55161 , n24318 , n24319 );
not ( n24320 , RI1754c610_2);
and ( n24321 , n24320 , n55161 );
and ( n24322 , C0 , RI1754c610_2);
or ( n55162 , n24321 , n24322 );
buf ( n55163 , n55162 );
buf ( n55164 , RI17464848_1246);
not ( n55165 , n49749 );
and ( n55166 , n55165 , n49573 );
xor ( n55167 , n51619 , n55166 );
not ( n24323 , n29614 );
and ( n24324 , n24323 , RI17462778_1256);
and ( n24325 , n55167 , n29614 );
or ( n55168 , n24324 , n24325 );
not ( n24326 , RI1754c610_2);
and ( n24327 , n24326 , n55168 );
and ( n24328 , C0 , RI1754c610_2);
or ( n55169 , n24327 , n24328 );
buf ( n55170 , n55169 );
not ( n55171 , n45541 );
and ( n55172 , n55171 , n45543 );
xor ( n55173 , n51794 , n55172 );
not ( n24329 , n29614 );
and ( n24330 , n24329 , RI1740bce8_1450);
and ( n24331 , n55173 , n29614 );
or ( n55174 , n24330 , n24331 );
not ( n24332 , RI1754c610_2);
and ( n24333 , n24332 , n55174 );
and ( n24334 , C0 , RI1754c610_2);
or ( n55175 , n24333 , n24334 );
buf ( n55176 , n55175 );
not ( n55177 , n47370 );
and ( n55178 , n55177 , n47372 );
xor ( n55179 , n47337 , n55178 );
not ( n24335 , n29614 );
and ( n24336 , n24335 , RI173bb348_1843);
and ( n24337 , n55179 , n29614 );
or ( n55180 , n24336 , n24337 );
not ( n24338 , RI1754c610_2);
and ( n24339 , n24338 , n55180 );
and ( n24340 , C0 , RI1754c610_2);
or ( n55181 , n24339 , n24340 );
buf ( n55182 , n55181 );
not ( n55183 , n44550 );
and ( n55184 , n55183 , n42910 );
xor ( n55185 , n44547 , n55184 );
not ( n24341 , n29614 );
and ( n24342 , n24341 , RI1733c868_2146);
and ( n24343 , n55185 , n29614 );
or ( n55186 , n24342 , n24343 );
not ( n24344 , RI1754c610_2);
and ( n24345 , n24344 , n55186 );
and ( n24346 , C0 , RI1754c610_2);
or ( n55187 , n24345 , n24346 );
buf ( n55188 , n55187 );
not ( n55189 , n50789 );
and ( n55190 , n55189 , n44831 );
xor ( n55191 , n42837 , n55190 );
not ( n24347 , n29614 );
and ( n24348 , n24347 , RI17342790_2117);
and ( n24349 , n55191 , n29614 );
or ( n55192 , n24348 , n24349 );
not ( n24350 , RI1754c610_2);
and ( n24351 , n24350 , n55192 );
and ( n24352 , C0 , RI1754c610_2);
or ( n55193 , n24351 , n24352 );
buf ( n55194 , n55193 );
not ( n24353 , n27683 );
and ( n24354 , n24353 , RI19aae7a0_2465);
and ( n24355 , RI19ab82c8_2394 , n27683 );
or ( n55195 , n24354 , n24355 );
not ( n24356 , RI1754c610_2);
and ( n24357 , n24356 , n55195 );
and ( n24358 , C0 , RI1754c610_2);
or ( n55196 , n24357 , n24358 );
buf ( n55197 , n55196 );
not ( n55198 , n45095 );
and ( n55199 , n55198 , n45699 );
xor ( n55200 , n36465 , n55199 );
not ( n24359 , n29614 );
and ( n24360 , n24359 , RI174b23e0_867);
and ( n24361 , n55200 , n29614 );
or ( n55201 , n24360 , n24361 );
not ( n24362 , RI1754c610_2);
and ( n24363 , n24362 , n55201 );
and ( n24364 , C0 , RI1754c610_2);
or ( n55202 , n24363 , n24364 );
buf ( n55203 , n55202 );
not ( n55204 , n51453 );
and ( n55205 , n55204 , n52126 );
xor ( n55206 , n47855 , n55205 );
not ( n24365 , n29614 );
and ( n24366 , n24365 , RI1733e938_2136);
and ( n24367 , n55206 , n29614 );
or ( n55207 , n24366 , n24367 );
not ( n24368 , RI1754c610_2);
and ( n24369 , n24368 , n55207 );
and ( n24370 , C0 , RI1754c610_2);
or ( n55208 , n24369 , n24370 );
buf ( n55209 , n55208 );
not ( n24371 , n27683 );
and ( n24372 , n24371 , RI19acb648_2244);
and ( n24373 , RI19a86fc0_2745 , n27683 );
or ( n55210 , n24372 , n24373 );
not ( n24374 , RI1754c610_2);
and ( n24375 , n24374 , n55210 );
and ( n24376 , C0 , RI1754c610_2);
or ( n55211 , n24375 , n24376 );
buf ( n55212 , n55211 );
not ( n55213 , n43709 );
and ( n55214 , n55213 , n43711 );
xor ( n55215 , n50854 , n55214 );
not ( n24377 , n29614 );
and ( n24378 , n24377 , RI17448378_1384);
and ( n24379 , n55215 , n29614 );
or ( n55216 , n24378 , n24379 );
not ( n24380 , RI1754c610_2);
and ( n24381 , n24380 , n55216 );
and ( n24382 , C0 , RI1754c610_2);
or ( n55217 , n24381 , n24382 );
buf ( n55218 , n55217 );
not ( n55219 , n53216 );
and ( n55220 , n55219 , n54172 );
xor ( n55221 , n53213 , n55220 );
not ( n24383 , n29614 );
and ( n24384 , n24383 , RI17393028_2039);
and ( n24385 , n55221 , n29614 );
or ( n55222 , n24384 , n24385 );
not ( n24386 , RI1754c610_2);
and ( n24387 , n24386 , n55222 );
and ( n24388 , C0 , RI1754c610_2);
or ( n55223 , n24387 , n24388 );
buf ( n55224 , n55223 );
not ( n55225 , n44171 );
and ( n55226 , n55225 , n44173 );
xor ( n55227 , n51284 , n55226 );
not ( n24389 , n29614 );
and ( n24390 , n24389 , RI1745b4a0_1291);
and ( n24391 , n55227 , n29614 );
or ( n55228 , n24390 , n24391 );
not ( n24392 , RI1754c610_2);
and ( n24393 , n24392 , n55228 );
and ( n24394 , C0 , RI1754c610_2);
or ( n55229 , n24393 , n24394 );
buf ( n55230 , n55229 );
not ( n55231 , n44237 );
and ( n55232 , n55231 , n45025 );
xor ( n55233 , n37491 , n55232 );
not ( n24395 , n29614 );
and ( n24396 , n24395 , RI1745a0f0_1297);
and ( n24397 , n55233 , n29614 );
or ( n55234 , n24396 , n24397 );
not ( n24398 , RI1754c610_2);
and ( n24399 , n24398 , n55234 );
and ( n24400 , C0 , RI1754c610_2);
or ( n55235 , n24399 , n24400 );
buf ( n55236 , n55235 );
not ( n24401 , n27683 );
and ( n24402 , n24401 , RI19a9d9a0_2587);
and ( n24403 , RI19aa7090_2516 , n27683 );
or ( n55237 , n24402 , n24403 );
not ( n24404 , RI1754c610_2);
and ( n24405 , n24404 , n55237 );
and ( n24406 , C0 , RI1754c610_2);
or ( n55238 , n24405 , n24406 );
buf ( n55239 , n55238 );
buf ( n55240 , RI17483e50_1093);
buf ( n55241 , RI17497608_998);
not ( n55242 , n45831 );
xor ( n55243 , n36115 , n39131 );
xor ( n55244 , n55243 , n39151 );
and ( n55245 , n55242 , n55244 );
xor ( n55246 , n45828 , n55245 );
not ( n24407 , n29614 );
and ( n24408 , n24407 , RI174a4178_936);
and ( n24409 , n55246 , n29614 );
or ( n55247 , n24408 , n24409 );
not ( n24410 , RI1754c610_2);
and ( n24411 , n24410 , n55247 );
and ( n24412 , C0 , RI1754c610_2);
or ( n55248 , n24411 , n24412 );
buf ( n55249 , n55248 );
not ( n55250 , n37527 );
and ( n55251 , n55250 , n37580 );
xor ( n55252 , n44603 , n55251 );
not ( n24413 , n29614 );
and ( n24414 , n24413 , RI17530500_616);
and ( n24415 , n55252 , n29614 );
or ( n55253 , n24414 , n24415 );
not ( n24416 , RI1754c610_2);
and ( n24417 , n24416 , n55253 );
and ( n24418 , C0 , RI1754c610_2);
or ( n55254 , n24417 , n24418 );
buf ( n55255 , n55254 );
not ( n55256 , n41868 );
and ( n55257 , n55256 , n41870 );
xor ( n55258 , n46595 , n55257 );
not ( n24419 , n29614 );
and ( n24420 , n24419 , RI1739de10_1986);
and ( n24421 , n55258 , n29614 );
or ( n55259 , n24420 , n24421 );
not ( n24422 , RI1754c610_2);
and ( n24423 , n24422 , n55259 );
and ( n24424 , C0 , RI1754c610_2);
or ( n55260 , n24423 , n24424 );
buf ( n55261 , n55260 );
not ( n55262 , n43280 );
and ( n55263 , n55262 , n43282 );
xor ( n55264 , n47771 , n55263 );
not ( n24425 , n29614 );
and ( n24426 , n24425 , RI17526a50_646);
and ( n24427 , n55264 , n29614 );
or ( n55265 , n24426 , n24427 );
not ( n24428 , RI1754c610_2);
xor ( n24429 , n24428 , n55265 );
and ( n24430 , C0 , RI1754c610_2);
nor ( n55266 , n24429 , n24430 );
buf ( n55267 , n55266 );
not ( n55268 , RI174c3438_803);
buf ( n55269 , RI1750cdd0_726);
not ( n55270 , n41858 );
or ( n55271 , n55270 , n47512 );
or ( n55272 , n41855 , n55271 );
not ( n24431 , n29614 );
and ( n24432 , n24431 , RI17484b70_1089);
and ( n24433 , n55272 , n29614 );
or ( n55273 , n24432 , n24433 );
not ( n24434 , RI1754c610_2);
and ( n24435 , n24434 , n55273 );
and ( n24436 , C0 , RI1754c610_2);
or ( n55274 , n24435 , n24436 );
buf ( n55275 , n55274 );
not ( n55276 , n45004 );
and ( n55277 , n55276 , n45006 );
xor ( n55278 , n50021 , n55277 );
not ( n24437 , n29614 );
and ( n24438 , n24437 , RI174837c0_1095);
and ( n24439 , n55278 , n29614 );
or ( n55279 , n24438 , n24439 );
not ( n24440 , RI1754c610_2);
and ( n24441 , n24440 , n55279 );
and ( n24442 , C0 , RI1754c610_2);
or ( n55280 , n24441 , n24442 );
buf ( n55281 , n55280 );
not ( n24443 , n27683 );
and ( n24444 , n24443 , RI19a831e0_2772);
and ( n24445 , RI19ab3c00_2425 , n27683 );
or ( n55282 , n24444 , n24445 );
not ( n24446 , RI1754c610_2);
and ( n24447 , n24446 , n55282 );
and ( n24448 , C0 , RI1754c610_2);
or ( n55283 , n24447 , n24448 );
buf ( n55284 , n55283 );
not ( n24449 , n27683 );
and ( n24450 , n24449 , RI19abf0f0_2340);
and ( n24451 , RI19ac81c8_2269 , n27683 );
or ( n55285 , n24450 , n24451 );
not ( n24452 , RI1754c610_2);
and ( n24453 , n24452 , n55285 );
and ( n24454 , C0 , RI1754c610_2);
or ( n55286 , n24453 , n24454 );
buf ( n55287 , n55286 );
not ( n55288 , n45690 );
and ( n55289 , n55288 , n44524 );
xor ( n55290 , n45687 , n55289 );
not ( n24455 , n29614 );
and ( n24456 , n24455 , RI1744bb40_1367);
and ( n24457 , n55290 , n29614 );
or ( n55291 , n24456 , n24457 );
not ( n24458 , RI1754c610_2);
and ( n24459 , n24458 , n55291 );
and ( n24460 , C0 , RI1754c610_2);
or ( n55292 , n24459 , n24460 );
buf ( n55293 , n55292 );
not ( n55294 , n48056 );
and ( n55295 , n55294 , n48467 );
xor ( n55296 , n46831 , n55295 );
not ( n24461 , n29614 );
and ( n24462 , n24461 , RI173f8878_1544);
and ( n24463 , n55296 , n29614 );
or ( n55297 , n24462 , n24463 );
not ( n24464 , RI1754c610_2);
and ( n24465 , n24464 , n55297 );
and ( n24466 , C0 , RI1754c610_2);
or ( n55298 , n24465 , n24466 );
buf ( n55299 , n55298 );
buf ( n55300 , RI17462430_1257);
buf ( n55301 , RI174772e0_1155);
not ( n55302 , n44557 );
and ( n55303 , n55302 , n44559 );
xor ( n55304 , n29611 , n55303 );
not ( n24467 , n29614 );
and ( n24468 , n24467 , RI17482758_1100);
and ( n24469 , n55304 , n29614 );
or ( n55305 , n24468 , n24469 );
not ( n24470 , RI1754c610_2);
and ( n24471 , n24470 , n55305 );
and ( n24472 , C0 , RI1754c610_2);
or ( n55306 , n24471 , n24472 );
buf ( n55307 , n55306 );
not ( n55308 , n50123 );
and ( n55309 , n55308 , n50125 );
xor ( n55310 , n52935 , n55309 );
not ( n24473 , n29614 );
and ( n24474 , n24473 , RI17464ed8_1244);
and ( n24475 , n55310 , n29614 );
or ( n55311 , n24474 , n24475 );
not ( n24476 , RI1754c610_2);
and ( n24477 , n24476 , n55311 );
and ( n24478 , C0 , RI1754c610_2);
or ( n55312 , n24477 , n24478 );
buf ( n55313 , n55312 );
not ( n55314 , n52181 );
and ( n55315 , n55314 , n52183 );
xor ( n55316 , n54991 , n55315 );
not ( n24479 , n29614 );
and ( n24480 , n24479 , RI1744ae20_1371);
and ( n24481 , n55316 , n29614 );
or ( n55317 , n24480 , n24481 );
not ( n24482 , RI1754c610_2);
and ( n24483 , n24482 , n55317 );
and ( n24484 , C0 , RI1754c610_2);
or ( n55318 , n24483 , n24484 );
buf ( n55319 , n55318 );
not ( n55320 , n53296 );
and ( n55321 , n55320 , n52095 );
xor ( n55322 , n46856 , n55321 );
not ( n24485 , n29614 );
and ( n24486 , n24485 , RI1733b4b8_2152);
and ( n24487 , n55322 , n29614 );
or ( n55323 , n24486 , n24487 );
not ( n24488 , RI1754c610_2);
and ( n24489 , n24488 , n55323 );
and ( n24490 , C0 , RI1754c610_2);
or ( n55324 , n24489 , n24490 );
buf ( n55325 , n55324 );
not ( n55326 , n51510 );
and ( n55327 , n55326 , n45826 );
xor ( n55328 , n55244 , n55327 );
not ( n24491 , n29614 );
and ( n24492 , n24491 , RI174789d8_1148);
and ( n24493 , n55328 , n29614 );
or ( n55329 , n24492 , n24493 );
not ( n24494 , RI1754c610_2);
and ( n24495 , n24494 , n55329 );
and ( n24496 , C0 , RI1754c610_2);
or ( n55330 , n24495 , n24496 );
buf ( n55331 , n55330 );
not ( n55332 , n47576 );
and ( n55333 , n55332 , n44347 );
xor ( n55334 , n47573 , n55333 );
not ( n24497 , n29614 );
and ( n24498 , n24497 , RI173b43b8_1877);
and ( n24499 , n55334 , n29614 );
or ( n55335 , n24498 , n24499 );
not ( n24500 , RI1754c610_2);
and ( n24501 , n24500 , n55335 );
and ( n24502 , C0 , RI1754c610_2);
or ( n55336 , n24501 , n24502 );
buf ( n55337 , n55336 );
not ( n55338 , n52112 );
and ( n55339 , n55338 , n52040 );
xor ( n55340 , n41547 , n55339 );
not ( n24503 , n29614 );
and ( n24504 , n24503 , RI174c5328_797);
and ( n24505 , n55340 , n29614 );
or ( n55341 , n24504 , n24505 );
not ( n24506 , RI1754c610_2);
and ( n24507 , n24506 , n55341 );
and ( n24508 , C0 , RI1754c610_2);
or ( n55342 , n24507 , n24508 );
buf ( n55343 , n55342 );
not ( n55344 , n46507 );
and ( n55345 , n55344 , n35640 );
xor ( n55346 , n35070 , n55345 );
not ( n24509 , n29614 );
and ( n24510 , n24509 , RI173db340_1687);
and ( n24511 , n55346 , n29614 );
or ( n55347 , n24510 , n24511 );
not ( n24512 , RI1754c610_2);
and ( n24513 , n24512 , n55347 );
and ( n24514 , C0 , RI1754c610_2);
or ( n55348 , n24513 , n24514 );
buf ( n55349 , n55348 );
not ( n55350 , n43981 );
and ( n55351 , n55350 , n43996 );
xor ( n55352 , n39887 , n55351 );
not ( n24515 , n29614 );
and ( n24516 , n24515 , RI173d2970_1729);
and ( n24517 , n55352 , n29614 );
or ( n55353 , n24516 , n24517 );
not ( n24518 , RI1754c610_2);
and ( n24519 , n24518 , n55353 );
and ( n24520 , C0 , RI1754c610_2);
or ( n55354 , n24519 , n24520 );
buf ( n55355 , n55354 );
not ( n55356 , n47255 );
and ( n55357 , n55356 , n38533 );
xor ( n55358 , n52755 , n55357 );
not ( n24521 , n29614 );
and ( n24522 , n24521 , RI1744b4b0_1369);
and ( n24523 , n55358 , n29614 );
or ( n55359 , n24522 , n24523 );
not ( n24524 , RI1754c610_2);
and ( n24525 , n24524 , n55359 );
and ( n24526 , C0 , RI1754c610_2);
or ( n55360 , n24525 , n24526 );
buf ( n55361 , n55360 );
not ( n55362 , n49145 );
and ( n55363 , n55362 , n49147 );
xor ( n55364 , n51230 , n55363 );
not ( n24527 , n29614 );
and ( n24528 , n24527 , RI174adbb0_889);
and ( n24529 , n55364 , n29614 );
or ( n55365 , n24528 , n24529 );
not ( n24530 , RI1754c610_2);
and ( n24531 , n24530 , n55365 );
and ( n24532 , C0 , RI1754c610_2);
or ( n55366 , n24531 , n24532 );
buf ( n55367 , n55366 );
not ( n55368 , n44514 );
and ( n55369 , n55368 , n44516 );
xor ( n55370 , n40747 , n55369 );
not ( n24533 , n29614 );
and ( n24534 , n24533 , RI1747fff8_1112);
and ( n24535 , n55370 , n29614 );
or ( n55371 , n24534 , n24535 );
not ( n24536 , RI1754c610_2);
and ( n24537 , n24536 , n55371 );
and ( n24538 , C0 , RI1754c610_2);
or ( n55372 , n24537 , n24538 );
buf ( n55373 , n55372 );
not ( n55374 , n45982 );
nand ( n55375 , n55374 , n43219 );
or ( n55376 , n38890 , n55375 );
not ( n24539 , n29614 );
nand ( n24540 , n24539 , RI17408bb0_1465);
nand ( n24541 , n55376 , n29614 );
xor ( n55377 , n24540 , n24541 );
not ( n24542 , RI1754c610_2);
and ( n24543 , n24542 , n55377 );
and ( n24544 , C0 , RI1754c610_2);
xor ( n55378 , n24543 , n24544 );
buf ( n55379 , n55378 );
not ( n55380 , n45912 );
and ( n55381 , n55380 , n45914 );
xor ( n55382 , n43099 , n55381 );
not ( n24545 , n29614 );
and ( n24546 , n24545 , RI17397858_2017);
and ( n24547 , n55382 , n29614 );
or ( n55383 , n24546 , n24547 );
not ( n24548 , RI1754c610_2);
and ( n24549 , n24548 , n55383 );
and ( n24550 , C0 , RI1754c610_2);
or ( n55384 , n24549 , n24550 );
buf ( n55385 , n55384 );
not ( n55386 , n47139 );
and ( n55387 , n55386 , n46670 );
xor ( n55388 , n42434 , n55387 );
not ( n24551 , n29614 );
and ( n24552 , n24551 , RI1747b138_1136);
and ( n24553 , n55388 , n29614 );
or ( n55389 , n24552 , n24553 );
not ( n24554 , RI1754c610_2);
and ( n24555 , n24554 , n55389 );
and ( n24556 , C0 , RI1754c610_2);
or ( n55390 , n24555 , n24556 );
buf ( n55391 , n55390 );
not ( n55392 , n55244 );
and ( n55393 , n55392 , n51510 );
xor ( n55394 , n45831 , n55393 );
not ( n24557 , n29614 );
and ( n24558 , n24557 , RI17469d98_1220);
and ( n24559 , n55394 , n29614 );
or ( n55395 , n24558 , n24559 );
not ( n24560 , RI1754c610_2);
and ( n24561 , n24560 , n55395 );
and ( n24562 , C0 , RI1754c610_2);
or ( n55396 , n24561 , n24562 );
buf ( n55397 , n55396 );
not ( n24563 , n27683 );
and ( n24564 , n24563 , RI19abff78_2332);
and ( n24565 , RI19ac90c8_2262 , n27683 );
or ( n55398 , n24564 , n24565 );
not ( n24566 , RI1754c610_2);
and ( n24567 , n24566 , n55398 );
and ( n24568 , C0 , RI1754c610_2);
or ( n55399 , n24567 , n24568 );
buf ( n55400 , n55399 );
not ( n55401 , n46040 );
and ( n55402 , n55401 , n51062 );
xor ( n55403 , n46037 , n55402 );
not ( n24569 , n29614 );
and ( n24570 , n24569 , RI1752a830_634);
and ( n24571 , n55403 , n29614 );
or ( n55404 , n24570 , n24571 );
not ( n24572 , RI1754c610_2);
and ( n24573 , n24572 , n55404 );
and ( n24574 , C0 , RI1754c610_2);
or ( n55405 , n24573 , n24574 );
buf ( n55406 , n55405 );
buf ( n55407 , RI1748a0c0_1063);
buf ( n55408 , RI17488680_1071);
buf ( n55409 , RI17492dd8_1020);
buf ( n55410 , RI174916e0_1027);
buf ( n55411 , RI174c7218_791);
buf ( n55412 , RI174c48d8_799);
not ( n55413 , n47552 );
and ( n55414 , n55413 , n47554 );
xor ( n55415 , n40916 , n55414 );
not ( n24575 , n29614 );
and ( n24576 , n24575 , RI17495538_1008);
and ( n24577 , n55415 , n29614 );
or ( n55416 , n24576 , n24577 );
not ( n24578 , RI1754c610_2);
and ( n24579 , n24578 , n55416 );
and ( n24580 , C0 , RI1754c610_2);
or ( n55417 , n24579 , n24580 );
buf ( n55418 , n55417 );
buf ( n55419 , RI17503de8_748);
buf ( n55420 , RI175014a8_756);
not ( n55421 , n50485 );
and ( n55422 , n55421 , n52430 );
xor ( n55423 , n50482 , n55422 );
not ( n24581 , n29614 );
and ( n24582 , n24581 , RI17484198_1092);
and ( n24583 , n55423 , n29614 );
or ( n55424 , n24582 , n24583 );
not ( n24584 , RI1754c610_2);
and ( n24585 , n24584 , n55424 );
and ( n24586 , C0 , RI1754c610_2);
or ( n55425 , n24585 , n24586 );
buf ( n55426 , n55425 );
not ( n24587 , n27683 );
and ( n24588 , n24587 , RI19a94940_2650);
and ( n24589 , RI19a9ed50_2578 , n27683 );
or ( n55427 , n24588 , n24589 );
not ( n24590 , RI1754c610_2);
and ( n24591 , n24590 , n55427 );
and ( n24592 , C0 , RI1754c610_2);
or ( n55428 , n24591 , n24592 );
buf ( n55429 , n55428 );
not ( n24593 , n27683 );
and ( n24594 , n24593 , RI19a92960_2664);
and ( n24595 , RI19a9ca28_2593 , n27683 );
or ( n55430 , n24594 , n24595 );
not ( n24596 , RI1754c610_2);
and ( n24597 , n24596 , n55430 );
and ( n24598 , C0 , RI1754c610_2);
or ( n55431 , n24597 , n24598 );
buf ( n55432 , n55431 );
not ( n55433 , n39831 );
and ( n55434 , n55433 , n39833 );
xor ( n55435 , n43996 , n55434 );
not ( n24599 , n29614 );
and ( n24600 , n24599 , RI173ef818_1588);
and ( n24601 , n55435 , n29614 );
or ( n55436 , n24600 , n24601 );
not ( n24602 , RI1754c610_2);
and ( n24603 , n24602 , n55436 );
and ( n24604 , C0 , RI1754c610_2);
or ( n55437 , n24603 , n24604 );
buf ( n55438 , n55437 );
not ( n55439 , n53211 );
and ( n55440 , n55439 , n53213 );
xor ( n55441 , n54174 , n55440 );
not ( n24605 , n29614 );
and ( n24606 , n24605 , RI173beb10_1826);
and ( n24607 , n55441 , n29614 );
or ( n55442 , n24606 , n24607 );
not ( n24608 , RI1754c610_2);
and ( n24609 , n24608 , n55442 );
and ( n24610 , C0 , RI1754c610_2);
or ( n55443 , n24609 , n24610 );
buf ( n55444 , n55443 );
not ( n24611 , n27683 );
and ( n24612 , n24611 , RI19aa46d8_2534);
and ( n24613 , RI19aae980_2464 , n27683 );
or ( n55445 , n24612 , n24613 );
not ( n24614 , RI1754c610_2);
and ( n24615 , n24614 , n55445 );
and ( n24616 , C0 , RI1754c610_2);
or ( n55446 , n24615 , n24616 );
buf ( n55447 , n55446 );
not ( n55448 , n48592 );
and ( n55449 , n55448 , n47063 );
xor ( n55450 , n54219 , n55449 );
not ( n24617 , n29614 );
and ( n24618 , n24617 , RI174cd410_772);
and ( n24619 , n55450 , n29614 );
or ( n55451 , n24618 , n24619 );
not ( n24620 , RI1754c610_2);
and ( n24621 , n24620 , n55451 );
and ( n24622 , C0 , RI1754c610_2);
or ( n55452 , n24621 , n24622 );
buf ( n55453 , n55452 );
not ( n55454 , n43571 );
and ( n55455 , n55454 , n48659 );
xor ( n55456 , n43568 , n55455 );
not ( n24623 , n29614 );
and ( n24624 , n24623 , RI173b8558_1857);
and ( n24625 , n55456 , n29614 );
or ( n55457 , n24624 , n24625 );
not ( n24626 , RI1754c610_2);
and ( n24627 , n24626 , n55457 );
and ( n24628 , C0 , RI1754c610_2);
or ( n55458 , n24627 , n24628 );
buf ( n55459 , n55458 );
not ( n55460 , n49883 );
and ( n55461 , n55460 , n50044 );
xor ( n55462 , n49554 , n55461 );
not ( n24629 , n29614 );
and ( n24630 , n24629 , RI1750f1e8_719);
and ( n24631 , n55462 , n29614 );
or ( n55463 , n24630 , n24631 );
not ( n24632 , RI1754c610_2);
and ( n24633 , n24632 , n55463 );
and ( n24634 , C0 , RI1754c610_2);
or ( n55464 , n24633 , n24634 );
buf ( n55465 , n55464 );
not ( n55466 , n48305 );
and ( n55467 , n55466 , n48307 );
xor ( n55468 , n49908 , n55467 );
not ( n24635 , n29614 );
and ( n24636 , n24635 , RI17530f50_614);
and ( n24637 , n55468 , n29614 );
or ( n55469 , n24636 , n24637 );
not ( n24638 , RI1754c610_2);
and ( n24639 , n24638 , n55469 );
and ( n24640 , C0 , RI1754c610_2);
or ( n55470 , n24639 , n24640 );
buf ( n55471 , n55470 );
not ( n24641 , n27683 );
and ( n24642 , n24641 , RI19ab7878_2398);
and ( n24643 , RI19ac0680_2328 , n27683 );
or ( n55472 , n24642 , n24643 );
not ( n24644 , RI1754c610_2);
and ( n24645 , n24644 , n55472 );
and ( n24646 , C0 , RI1754c610_2);
or ( n55473 , n24645 , n24646 );
buf ( n55474 , n55473 );
not ( n55475 , n45591 );
and ( n55476 , n55475 , n43160 );
xor ( n55477 , n45588 , n55476 );
not ( n24647 , n29614 );
and ( n24648 , n24647 , RI1744e2a0_1355);
and ( n24649 , n55477 , n29614 );
or ( n55478 , n24648 , n24649 );
not ( n24650 , RI1754c610_2);
and ( n24651 , n24650 , n55478 );
and ( n24652 , C0 , RI1754c610_2);
or ( n55479 , n24651 , n24652 );
buf ( n55480 , n55479 );
not ( n55481 , n41724 );
and ( n55482 , n55481 , n41742 );
xor ( n55483 , n49527 , n55482 );
not ( n24653 , n29614 );
and ( n24654 , n24653 , RI174720d8_1180);
and ( n24655 , n55483 , n29614 );
or ( n55484 , n24654 , n24655 );
not ( n24656 , RI1754c610_2);
and ( n24657 , n24656 , n55484 );
and ( n24658 , C0 , RI1754c610_2);
or ( n55485 , n24657 , n24658 );
buf ( n55486 , n55485 );
not ( n55487 , n44997 );
and ( n55488 , n55487 , n45204 );
xor ( n55489 , n43928 , n55488 );
not ( n24659 , n29614 );
and ( n24660 , n24659 , RI175323f0_610);
and ( n24661 , n55489 , n29614 );
or ( n55490 , n24660 , n24661 );
not ( n24662 , RI1754c610_2);
and ( n24663 , n24662 , n55490 );
and ( n24664 , C0 , RI1754c610_2);
or ( n55491 , n24663 , n24664 );
buf ( n55492 , n55491 );
buf ( n55493 , RI17484eb8_1088);
buf ( n55494 , RI174a3110_941);
buf ( n55495 , RI174affc8_878);
buf ( n55496 , RI17510bb0_714);
not ( n24665 , n27683 );
and ( n24666 , n24665 , RI19a97dc0_2627);
and ( n24667 , RI19aa17f8_2556 , n27683 );
or ( n55497 , n24666 , n24667 );
not ( n24668 , RI1754c610_2);
and ( n24669 , n24668 , n55497 );
and ( n24670 , C0 , RI1754c610_2);
or ( n55498 , n24669 , n24670 );
buf ( n55499 , n55498 );
not ( n55500 , n47544 );
and ( n55501 , n55500 , n44845 );
xor ( n55502 , n48131 , n55501 );
not ( n24671 , n29614 );
and ( n24672 , n24671 , RI173eb9c0_1607);
and ( n24673 , n55502 , n29614 );
or ( n55503 , n24672 , n24673 );
not ( n24674 , RI1754c610_2);
and ( n24675 , n24674 , n55503 );
and ( n24676 , C0 , RI1754c610_2);
or ( n55504 , n24675 , n24676 );
buf ( n55505 , n55504 );
not ( n55506 , n40255 );
and ( n55507 , n55506 , n40257 );
xor ( n55508 , n44585 , n55507 );
not ( n24677 , n29614 );
and ( n24678 , n24677 , RI173e1c40_1655);
and ( n24679 , n55508 , n29614 );
or ( n55509 , n24678 , n24679 );
not ( n24680 , RI1754c610_2);
and ( n24681 , n24680 , n55509 );
and ( n24682 , C0 , RI1754c610_2);
or ( n55510 , n24681 , n24682 );
buf ( n55511 , n55510 );
not ( n55512 , n47948 );
and ( n55513 , n55512 , n45483 );
xor ( n55514 , n49183 , n55513 );
not ( n24683 , n29614 );
and ( n24684 , n24683 , RI17396160_2024);
and ( n24685 , n55514 , n29614 );
or ( n55515 , n24684 , n24685 );
not ( n24686 , RI1754c610_2);
and ( n24687 , n24686 , n55515 );
and ( n24688 , C0 , RI1754c610_2);
or ( n55516 , n24687 , n24688 );
buf ( n55517 , n55516 );
not ( n55518 , n54103 );
and ( n55519 , n55518 , n49561 );
xor ( n55520 , n50782 , n55519 );
not ( n24689 , n29614 );
and ( n24690 , n24689 , RI175319a0_612);
and ( n24691 , n55520 , n29614 );
or ( n55521 , n24690 , n24691 );
not ( n24692 , RI1754c610_2);
and ( n24693 , n24692 , n55521 );
and ( n24694 , C0 , RI1754c610_2);
or ( n55522 , n24693 , n24694 );
buf ( n55523 , n55522 );
not ( n55524 , n43397 );
and ( n55525 , n55524 , n43399 );
xor ( n55526 , n45755 , n55525 );
not ( n24695 , n29614 );
and ( n24696 , n24695 , RI17511b28_711);
and ( n24697 , n55526 , n29614 );
or ( n55527 , n24696 , n24697 );
not ( n24698 , RI1754c610_2);
and ( n24699 , n24698 , n55527 );
and ( n24700 , C0 , RI1754c610_2);
or ( n55528 , n24699 , n24700 );
buf ( n55529 , n55528 );
buf ( n55530 , RI174a23f0_945);
buf ( n55531 , RI174b44b0_857);
not ( n55532 , n41898 );
and ( n55533 , n55532 , n47362 );
xor ( n55534 , n41895 , n55533 );
not ( n24701 , n29614 );
and ( n24702 , n24701 , RI17457990_1309);
and ( n24703 , n55534 , n29614 );
or ( n55535 , n24702 , n24703 );
not ( n24704 , RI1754c610_2);
and ( n24705 , n24704 , n55535 );
and ( n24706 , C0 , RI1754c610_2);
or ( n55536 , n24705 , n24706 );
buf ( n55537 , n55536 );
buf ( n55538 , RI17463e70_1249);
not ( n24707 , n27683 );
and ( n24708 , n24707 , RI19ac12b0_2321);
and ( n24709 , RI19aca748_2252 , n27683 );
or ( n55539 , n24708 , n24709 );
not ( n24710 , RI1754c610_2);
and ( n24711 , n24710 , n55539 );
and ( n24712 , C0 , RI1754c610_2);
or ( n55540 , n24711 , n24712 );
buf ( n55541 , n55540 );
not ( n55542 , n47866 );
and ( n55543 , n55542 , n44483 );
xor ( n55544 , n34838 , n55543 );
not ( n24713 , n29614 );
and ( n24714 , n24713 , RI173e0bd8_1660);
and ( n24715 , n55544 , n29614 );
or ( n55545 , n24714 , n24715 );
not ( n24716 , RI1754c610_2);
and ( n24717 , n24716 , n55545 );
and ( n24718 , C0 , RI1754c610_2);
or ( n55546 , n24717 , n24718 );
buf ( n55547 , n55546 );
not ( n55548 , n50259 );
and ( n55549 , n55548 , n52935 );
xor ( n55550 , n50128 , n55549 );
not ( n24719 , n29614 );
and ( n24720 , n24719 , RI174909c0_1031);
and ( n24721 , n55550 , n29614 );
or ( n55551 , n24720 , n24721 );
not ( n24722 , RI1754c610_2);
and ( n24723 , n24722 , n55551 );
and ( n24724 , C0 , RI1754c610_2);
or ( n55552 , n24723 , n24724 );
buf ( n55553 , n55552 );
not ( n24725 , n27683 );
and ( n24726 , n24725 , RI19aa27e8_2549);
and ( n24727 , RI19aacbf8_2477 , n27683 );
or ( n55554 , n24726 , n24727 );
not ( n24728 , RI1754c610_2);
and ( n24729 , n24728 , n55554 );
and ( n24730 , C0 , RI1754c610_2);
or ( n55555 , n24729 , n24730 );
buf ( n55556 , n55555 );
not ( n24731 , n27683 );
and ( n24732 , n24731 , RI19a983d8_2624);
and ( n24733 , RI19aa1d20_2554 , n27683 );
or ( n55557 , n24732 , n24733 );
not ( n24734 , RI1754c610_2);
and ( n24735 , n24734 , n55557 );
and ( n24736 , C0 , RI1754c610_2);
or ( n55558 , n24735 , n24736 );
buf ( n55559 , n55558 );
not ( n55560 , n42788 );
and ( n55561 , n55560 , n42790 );
xor ( n55562 , n44731 , n55561 );
not ( n24737 , n29614 );
and ( n24738 , n24737 , RI173e2ff0_1649);
and ( n24739 , n55562 , n29614 );
or ( n55563 , n24738 , n24739 );
not ( n24740 , RI1754c610_2);
and ( n24741 , n24740 , n55563 );
and ( n24742 , C0 , RI1754c610_2);
or ( n55564 , n24741 , n24742 );
buf ( n55565 , n55564 );
not ( n55566 , n42702 );
and ( n55567 , n55566 , n37049 );
xor ( n55568 , n50655 , n55567 );
not ( n24743 , n29614 );
and ( n24744 , n24743 , RI1752cc48_627);
and ( n24745 , n55568 , n29614 );
or ( n55569 , n24744 , n24745 );
not ( n24746 , RI1754c610_2);
and ( n24747 , n24746 , n55569 );
and ( n24748 , C0 , RI1754c610_2);
or ( n55570 , n24747 , n24748 );
buf ( n55571 , n55570 );
not ( n55572 , n42310 );
and ( n55573 , n55572 , n49890 );
xor ( n55574 , n40529 , n55573 );
not ( n24749 , n29614 );
and ( n24750 , n24749 , RI173bfb78_1821);
and ( n24751 , n55574 , n29614 );
or ( n55575 , n24750 , n24751 );
not ( n24752 , RI1754c610_2);
and ( n24753 , n24752 , n55575 );
and ( n24754 , C0 , RI1754c610_2);
or ( n55576 , n24753 , n24754 );
buf ( n55577 , n55576 );
not ( n55578 , n42837 );
and ( n55579 , n55578 , n50789 );
xor ( n55580 , n42834 , n55579 );
not ( n24755 , n29614 );
and ( n24756 , n24755 , RI173bd418_1833);
and ( n24757 , n55580 , n29614 );
or ( n55581 , n24756 , n24757 );
not ( n24758 , RI1754c610_2);
and ( n24759 , n24758 , n55581 );
and ( n24760 , C0 , RI1754c610_2);
or ( n55582 , n24759 , n24760 );
buf ( n55583 , n55582 );
not ( n24761 , n27683 );
and ( n24762 , n24761 , RI19acd808_2228);
and ( n24763 , RI19a8eb08_2692 , n27683 );
or ( n55584 , n24762 , n24763 );
not ( n24764 , RI1754c610_2);
and ( n24765 , n24764 , n55584 );
and ( n24766 , C0 , RI1754c610_2);
or ( n55585 , n24765 , n24766 );
buf ( n55586 , n55585 );
not ( n24767 , n27683 );
and ( n24768 , n24767 , RI19aa0970_2564);
and ( n24769 , RI19aaa510_2493 , n27683 );
or ( n55587 , n24768 , n24769 );
not ( n24770 , RI1754c610_2);
and ( n24771 , n24770 , n55587 );
and ( n24772 , C0 , RI1754c610_2);
or ( n55588 , n24771 , n24772 );
buf ( n55589 , n55588 );
not ( n55590 , n45804 );
and ( n55591 , n55590 , n45806 );
xor ( n55592 , n51805 , n55591 );
not ( n24773 , n29614 );
and ( n24774 , n24773 , RI173f46d8_1564);
and ( n24775 , n55592 , n29614 );
or ( n55593 , n24774 , n24775 );
not ( n24776 , RI1754c610_2);
and ( n24777 , n24776 , n55593 );
and ( n24778 , C0 , RI1754c610_2);
or ( n55594 , n24777 , n24778 );
buf ( n55595 , n55594 );
not ( n55596 , n43655 );
and ( n55597 , n55596 , n46069 );
xor ( n55598 , n43652 , n55597 );
not ( n24779 , n29614 );
and ( n24780 , n24779 , RI1751df18_673);
and ( n24781 , n55598 , n29614 );
or ( n55599 , n24780 , n24781 );
not ( n24782 , RI1754c610_2);
and ( n24783 , n24782 , n55599 );
and ( n24784 , C0 , RI1754c610_2);
or ( n55600 , n24783 , n24784 );
buf ( n55601 , n55600 );
not ( n55602 , n43638 );
and ( n55603 , n55602 , n46082 );
xor ( n55604 , n43635 , n55603 );
not ( n24785 , n29614 );
and ( n24786 , n24785 , RI173a1290_1970);
and ( n24787 , n55604 , n29614 );
or ( n55605 , n24786 , n24787 );
not ( n24788 , RI1754c610_2);
and ( n24789 , n24788 , n55605 );
and ( n24790 , C0 , RI1754c610_2);
or ( n55606 , n24789 , n24790 );
buf ( n55607 , n55606 );
not ( n24791 , n27683 );
and ( n24792 , n24791 , RI19a8c948_2707);
and ( n24793 , RI19a96bf0_2635 , n27683 );
or ( n55608 , n24792 , n24793 );
not ( n24794 , RI1754c610_2);
and ( n24795 , n24794 , n55608 );
and ( n24796 , C0 , RI1754c610_2);
or ( n55609 , n24795 , n24796 );
buf ( n55610 , n55609 );
not ( n55611 , n43249 );
and ( n55612 , n55611 , n36378 );
xor ( n55613 , n51409 , n55612 );
not ( n24797 , n29614 );
and ( n24798 , n24797 , RI17469a50_1221);
and ( n24799 , n55613 , n29614 );
or ( n55614 , n24798 , n24799 );
not ( n24800 , RI1754c610_2);
and ( n24801 , n24800 , n55614 );
and ( n24802 , C0 , RI1754c610_2);
or ( n55615 , n24801 , n24802 );
buf ( n55616 , n55615 );
not ( n24803 , n27683 );
and ( n24804 , n24803 , RI19abf870_2336);
and ( n24805 , RI19ac8768_2266 , n27683 );
or ( n55617 , n24804 , n24805 );
not ( n24806 , RI1754c610_2);
and ( n24807 , n24806 , n55617 );
and ( n24808 , C0 , RI1754c610_2);
or ( n55618 , n24807 , n24808 );
buf ( n55619 , n55618 );
buf ( n55620 , RI1748ffe8_1034);
not ( n55621 , n52227 );
and ( n55622 , n55621 , n52582 );
xor ( n55623 , n48289 , n55622 );
not ( n24809 , n29614 );
and ( n24810 , n24809 , RI174b7930_841);
and ( n24811 , n55623 , n29614 );
or ( n55624 , n24810 , n24811 );
not ( n24812 , RI1754c610_2);
and ( n24813 , n24812 , n55624 );
and ( n24814 , C0 , RI1754c610_2);
or ( n55625 , n24813 , n24814 );
buf ( n55626 , n55625 );
buf ( n55627 , RI174cedd8_767);
not ( n55628 , n43667 );
and ( n55629 , n55628 , n44323 );
xor ( n55630 , n43664 , n55629 );
not ( n24815 , n29614 );
and ( n24816 , n24815 , RI173a6b28_1943);
and ( n24817 , n55630 , n29614 );
or ( n55631 , n24816 , n24817 );
not ( n24818 , RI1754c610_2);
and ( n24819 , n24818 , n55631 );
and ( n24820 , C0 , RI1754c610_2);
or ( n55632 , n24819 , n24820 );
buf ( n55633 , n55632 );
not ( n55634 , n49078 );
and ( n55635 , n55634 , n49080 );
xor ( n55636 , n43589 , n55635 );
not ( n24821 , n29614 );
and ( n24822 , n24821 , RI17345c10_2101);
and ( n24823 , n55636 , n29614 );
or ( n55637 , n24822 , n24823 );
not ( n24824 , RI1754c610_2);
and ( n24825 , n24824 , n55637 );
and ( n24826 , C0 , RI1754c610_2);
or ( n55638 , n24825 , n24826 );
buf ( n55639 , n55638 );
not ( n55640 , n52316 );
and ( n55641 , n55640 , n43690 );
xor ( n55642 , n54706 , n55641 );
not ( n24827 , n29614 );
and ( n24828 , n24827 , RI173ba970_1846);
and ( n24829 , n55642 , n29614 );
or ( n55643 , n24828 , n24829 );
not ( n24830 , RI1754c610_2);
and ( n24831 , n24830 , n55643 );
and ( n24832 , C0 , RI1754c610_2);
or ( n55644 , n24831 , n24832 );
buf ( n55645 , n55644 );
not ( n55646 , n42076 );
and ( n55647 , n55646 , n45453 );
xor ( n55648 , n42073 , n55647 );
not ( n24833 , n29614 );
and ( n24834 , n24833 , RI173ddde8_1674);
and ( n24835 , n55648 , n29614 );
or ( n55649 , n24834 , n24835 );
not ( n24836 , RI1754c610_2);
and ( n24837 , n24836 , n55649 );
and ( n24838 , C0 , RI1754c610_2);
or ( n55650 , n24837 , n24838 );
buf ( n55651 , n55650 );
not ( n55652 , n48429 );
and ( n55653 , n55652 , n46197 );
xor ( n55654 , n49201 , n55653 );
not ( n24839 , n29614 );
and ( n24840 , n24839 , RI174af2a8_882);
and ( n24841 , n55654 , n29614 );
or ( n55655 , n24840 , n24841 );
not ( n24842 , RI1754c610_2);
and ( n24843 , n24842 , n55655 );
and ( n24844 , C0 , RI1754c610_2);
or ( n55656 , n24843 , n24844 );
buf ( n55657 , n55656 );
not ( n55658 , n54706 );
and ( n55659 , n55658 , n52316 );
xor ( n55660 , n43695 , n55659 );
not ( n24845 , n29614 );
and ( n24846 , n24845 , RI173ac078_1917);
and ( n24847 , n55660 , n29614 );
or ( n55661 , n24846 , n24847 );
not ( n24848 , RI1754c610_2);
and ( n24849 , n24848 , n55661 );
and ( n24850 , C0 , RI1754c610_2);
or ( n55662 , n24849 , n24850 );
buf ( n55663 , n55662 );
not ( n55664 , n39103 );
and ( n55665 , n55664 , n45214 );
xor ( n55666 , n39095 , n55665 );
not ( n24851 , n29614 );
and ( n24852 , n24851 , RI1733b800_2151);
and ( n24853 , n55666 , n29614 );
or ( n55667 , n24852 , n24853 );
not ( n24854 , RI1754c610_2);
and ( n24855 , n24854 , n55667 );
and ( n24856 , C0 , RI1754c610_2);
or ( n55668 , n24855 , n24856 );
buf ( n55669 , n55668 );
not ( n24857 , n27683 );
and ( n24858 , n24857 , RI19ab5f28_2409);
and ( n24859 , RI19abf2d0_2339 , n27683 );
or ( n55670 , n24858 , n24859 );
not ( n24860 , RI1754c610_2);
and ( n24861 , n24860 , n55670 );
and ( n24862 , C0 , RI1754c610_2);
or ( n55671 , n24861 , n24862 );
buf ( n55672 , n55671 );
not ( n24863 , n27683 );
and ( n24864 , n24863 , RI19aac838_2479);
and ( n24865 , RI19ab6090_2408 , n27683 );
or ( n55673 , n24864 , n24865 );
not ( n24866 , RI1754c610_2);
and ( n24867 , n24866 , n55673 );
and ( n24868 , C0 , RI1754c610_2);
or ( n55674 , n24867 , n24868 );
buf ( n55675 , n55674 );
not ( n24869 , RI1754c610_2);
and ( n24870 , n24869 , RI19ad1ee8_2199);
and ( n24871 , C0 , RI1754c610_2);
or ( n55676 , n24870 , n24871 );
buf ( n55677 , n55676 );
not ( n24872 , n27683 );
and ( n24873 , n24872 , RI19acba08_2242);
and ( n24874 , RI19a87470_2743 , n27683 );
or ( n55678 , n24873 , n24874 );
not ( n24875 , RI1754c610_2);
and ( n24876 , n24875 , n55678 );
and ( n24877 , C0 , RI1754c610_2);
or ( n55679 , n24876 , n24877 );
buf ( n55680 , n55679 );
not ( n55681 , n42449 );
and ( n55682 , n55681 , n45473 );
xor ( n55683 , n42446 , n55682 );
not ( n24878 , n29614 );
and ( n24879 , n24878 , RI17465220_1243);
and ( n24880 , n55683 , n29614 );
or ( n55684 , n24879 , n24880 );
not ( n24881 , RI1754c610_2);
and ( n24882 , n24881 , n55684 );
and ( n24883 , C0 , RI1754c610_2);
or ( n55685 , n24882 , n24883 );
buf ( n55686 , n55685 );
not ( n55687 , n43035 );
and ( n55688 , n55687 , n43037 );
xor ( n55689 , n47160 , n55688 );
not ( n24884 , n29614 );
and ( n24885 , n24884 , RI1744f650_1349);
and ( n24886 , n55689 , n29614 );
or ( n55690 , n24885 , n24886 );
not ( n24887 , RI1754c610_2);
and ( n24888 , n24887 , n55690 );
and ( n24889 , C0 , RI1754c610_2);
or ( n55691 , n24888 , n24889 );
buf ( n55692 , n55691 );
not ( n55693 , n43524 );
and ( n55694 , n55693 , n43526 );
xor ( n55695 , n43180 , n55694 );
not ( n24890 , n29614 );
and ( n24891 , n24890 , RI17522748_659);
and ( n24892 , n55695 , n29614 );
or ( n55696 , n24891 , n24892 );
not ( n24893 , RI1754c610_2);
and ( n24894 , n24893 , n55696 );
and ( n24895 , C0 , RI1754c610_2);
or ( n55697 , n24894 , n24895 );
buf ( n55698 , n55697 );
not ( n55699 , n48977 );
and ( n55700 , n55699 , n41296 );
xor ( n55701 , n48974 , n55700 );
not ( n24896 , n29614 );
and ( n24897 , n24896 , RI17507100_744);
and ( n24898 , n55701 , n29614 );
or ( n55702 , n24897 , n24898 );
not ( n24899 , RI1754c610_2);
and ( n24900 , n24899 , n55702 );
and ( n24901 , C0 , RI1754c610_2);
or ( n55703 , n24900 , n24901 );
buf ( n55704 , n55703 );
not ( n24902 , n27683 );
and ( n24903 , n24902 , RI19a84e00_2760);
and ( n24904 , RI19ac36c8_2303 , n27683 );
or ( n55705 , n24903 , n24904 );
not ( n24905 , RI1754c610_2);
and ( n24906 , n24905 , n55705 );
and ( n24907 , C0 , RI1754c610_2);
or ( n55706 , n24906 , n24907 );
buf ( n55707 , n55706 );
not ( n24908 , n27683 );
and ( n24909 , n24908 , RI19ac8c18_2264);
and ( n24910 , RI19a83d20_2767 , n27683 );
or ( n55708 , n24909 , n24910 );
not ( n24911 , RI1754c610_2);
and ( n24912 , n24911 , n55708 );
and ( n24913 , C0 , RI1754c610_2);
or ( n55709 , n24912 , n24913 );
buf ( n55710 , n55709 );
buf ( n55711 , RI1747c830_1129);
not ( n55712 , n42421 );
and ( n55713 , n55712 , n38934 );
xor ( n55714 , n44004 , n55713 );
not ( n24914 , n29614 );
and ( n24915 , n24914 , RI17510688_715);
and ( n24916 , n55714 , n29614 );
or ( n55715 , n24915 , n24916 );
not ( n24917 , RI1754c610_2);
and ( n24918 , n24917 , n55715 );
and ( n24919 , C0 , RI1754c610_2);
or ( n55716 , n24918 , n24919 );
buf ( n55717 , n55716 );
buf ( n55718 , RI1746f2e8_1194);
not ( n55719 , n51445 );
and ( n55720 , n55719 , n44147 );
xor ( n55721 , n51442 , n55720 );
not ( n24920 , n29614 );
and ( n24921 , n24920 , RI17496f78_1000);
and ( n24922 , n55721 , n29614 );
or ( n55722 , n24921 , n24922 );
not ( n24923 , RI1754c610_2);
and ( n24924 , n24923 , n55722 );
and ( n24925 , C0 , RI1754c610_2);
or ( n55723 , n24924 , n24925 );
buf ( n55724 , n55723 );
not ( n55725 , n47288 );
and ( n55726 , n55725 , n43337 );
xor ( n55727 , n46450 , n55726 );
not ( n24926 , n29614 );
and ( n24927 , n24926 , RI1738eb40_2060);
and ( n24928 , n55727 , n29614 );
or ( n55728 , n24927 , n24928 );
not ( n24929 , RI1754c610_2);
and ( n24930 , n24929 , n55728 );
and ( n24931 , C0 , RI1754c610_2);
or ( n55729 , n24930 , n24931 );
buf ( n55730 , n55729 );
not ( n55731 , n47453 );
and ( n55732 , n55731 , n47614 );
xor ( n55733 , n46578 , n55732 );
not ( n24932 , n29614 );
and ( n24933 , n24932 , RI173efb60_1587);
and ( n24934 , n55733 , n29614 );
or ( n55734 , n24933 , n24934 );
not ( n24935 , RI1754c610_2);
and ( n24936 , n24935 , n55734 );
and ( n24937 , C0 , RI1754c610_2);
or ( n55735 , n24936 , n24937 );
buf ( n55736 , n55735 );
not ( n55737 , n44095 );
and ( n55738 , n55737 , n44097 );
xor ( n55739 , n45184 , n55738 );
not ( n24938 , n29614 );
and ( n24939 , n24938 , RI173d8f28_1698);
and ( n24940 , n55739 , n29614 );
or ( n55740 , n24939 , n24940 );
not ( n24941 , RI1754c610_2);
and ( n24942 , n24941 , n55740 );
and ( n24943 , C0 , RI1754c610_2);
or ( n55741 , n24942 , n24943 );
buf ( n55742 , n55741 );
not ( n55743 , n36210 );
and ( n55744 , n55743 , n36228 );
xor ( n55745 , n50692 , n55744 );
not ( n24944 , n29614 );
and ( n24945 , n24944 , RI17410518_1428);
and ( n24946 , n55745 , n29614 );
or ( n55746 , n24945 , n24946 );
not ( n24947 , RI1754c610_2);
and ( n24948 , n24947 , n55746 );
and ( n24949 , C0 , RI1754c610_2);
or ( n55747 , n24948 , n24949 );
buf ( n55748 , n55747 );
and ( n55749 , RI1754b008_49 , n34844 );
and ( n55750 , RI1754b008_49 , n34847 );
or ( n55751 , n55749 , n55750 , C0 , C0 , C0 , C0 , C0 , C0 );
not ( n24950 , n34859 );
and ( n24951 , n24950 , n55751 );
and ( n24952 , RI1754b008_49 , n34859 );
or ( n55752 , n24951 , n24952 );
not ( n24953 , RI19a22f70_2797);
and ( n24954 , n24953 , n55752 );
and ( n24955 , C0 , RI19a22f70_2797);
or ( n55753 , n24954 , n24955 );
not ( n24956 , n27683 );
and ( n24957 , n24956 , RI19ac4f28_2292);
and ( n24958 , n55753 , n27683 );
or ( n55754 , n24957 , n24958 );
not ( n24959 , RI1754c610_2);
and ( n24960 , n24959 , n55754 );
and ( n24961 , C0 , RI1754c610_2);
or ( n55755 , n24960 , n24961 );
buf ( n55756 , n55755 );
not ( n24962 , n27683 );
and ( n24963 , n24962 , RI19a8ffa8_2683);
and ( n24964 , RI19a9a160_2611 , n27683 );
or ( n55757 , n24963 , n24964 );
not ( n24965 , RI1754c610_2);
and ( n24966 , n24965 , n55757 );
and ( n24967 , C0 , RI1754c610_2);
or ( n55758 , n24966 , n24967 );
buf ( n55759 , n55758 );
buf ( n55760 , RI1747b480_1135);
buf ( n55761 , RI174865b0_1081);
buf ( n55762 , RI17508ff0_738);
not ( n55763 , n51687 );
and ( n55764 , n55763 , n49422 );
xor ( n55765 , n51684 , n55764 );
or ( n55766 , n27689 , RI17538c00_591);
or ( n55767 , n55766 , RI17537fd0_593);
or ( n55768 , n55767 , RI175373a0_595);
or ( n55769 , n55768 , RI17536770_597);
xor ( n55770 , n55765 , n55769 );
not ( n24968 , n29614 );
and ( n24969 , n24968 , RI1746dbf0_1201);
and ( n24970 , n55770 , n29614 );
or ( n55771 , n24969 , n24970 );
not ( n24971 , RI1754c610_2);
and ( n24972 , n24971 , n55771 );
and ( n24973 , C0 , RI1754c610_2);
or ( n55772 , n24972 , n24973 );
buf ( n55773 , n55772 );
not ( n55774 , n39221 );
and ( n55775 , n55774 , n43935 );
xor ( n55776 , n39215 , n55775 );
not ( n24974 , n29614 );
and ( n24975 , n24974 , RI173f4390_1565);
and ( n24976 , n55776 , n29614 );
or ( n55777 , n24975 , n24976 );
not ( n24977 , RI1754c610_2);
and ( n24978 , n24977 , n55777 );
and ( n24979 , C0 , RI1754c610_2);
or ( n55778 , n24978 , n24979 );
buf ( n55779 , n55778 );
and ( n55780 , RI1754c4a8_5 , n34844 );
and ( n55781 , RI1754c4a8_5 , n34847 );
and ( n55782 , RI1754c4a8_5 , n34850 );
and ( n55783 , RI1754c4a8_5 , n34852 );
and ( n55784 , RI1754c4a8_5 , n34854 );
and ( n55785 , RI1754c4a8_5 , n34856 );
and ( n55786 , RI1754c4a8_5 , n39233 );
or ( n55787 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , C0 );
not ( n24980 , n34859 );
and ( n24981 , n24980 , n55787 );
and ( n24982 , RI1754c4a8_5 , n34859 );
or ( n55788 , n24981 , n24982 );
not ( n24983 , RI19a22f70_2797);
and ( n24984 , n24983 , n55788 );
and ( n24985 , C0 , RI19a22f70_2797);
or ( n55789 , n24984 , n24985 );
not ( n24986 , n27683 );
and ( n24987 , n24986 , RI19a88208_2737);
and ( n24988 , n55789 , n27683 );
or ( n55790 , n24987 , n24988 );
not ( n24989 , RI1754c610_2);
and ( n24990 , n24989 , n55790 );
and ( n24991 , C0 , RI1754c610_2);
or ( n55791 , n24990 , n24991 );
buf ( n55792 , n55791 );
not ( n55793 , n51884 );
and ( n55794 , n55793 , n48685 );
xor ( n55795 , n51881 , n55794 );
not ( n24992 , n29614 );
and ( n24993 , n24992 , RI17399928_2007);
and ( n24994 , n55795 , n29614 );
or ( n55796 , n24993 , n24994 );
not ( n24995 , RI1754c610_2);
and ( n24996 , n24995 , n55796 );
and ( n24997 , C0 , RI1754c610_2);
or ( n55797 , n24996 , n24997 );
buf ( n55798 , n55797 );
not ( n55799 , n42350 );
and ( n55800 , n55799 , n49454 );
xor ( n55801 , n42347 , n55800 );
not ( n24998 , n29614 );
and ( n24999 , n24998 , RI173ffb50_1509);
and ( n25000 , n55801 , n29614 );
or ( n55802 , n24999 , n25000 );
not ( n25001 , RI1754c610_2);
and ( n25002 , n25001 , n55802 );
and ( n25003 , C0 , RI1754c610_2);
or ( n55803 , n25002 , n25003 );
buf ( n55804 , n55803 );
not ( n55805 , n45456 );
and ( n55806 , n55805 , n42071 );
xor ( n55807 , n45453 , n55806 );
not ( n25004 , n29614 );
and ( n25005 , n25004 , RI173fac90_1533);
and ( n25006 , n55807 , n29614 );
or ( n55808 , n25005 , n25006 );
not ( n25007 , RI1754c610_2);
and ( n25008 , n25007 , n55808 );
and ( n25009 , C0 , RI1754c610_2);
or ( n55809 , n25008 , n25009 );
buf ( n55810 , n55809 );
not ( n25010 , n27683 );
and ( n25011 , n25010 , RI19a9b8d0_2601);
and ( n25012 , RI19aa4ed0_2530 , n27683 );
or ( n55811 , n25011 , n25012 );
not ( n25013 , RI1754c610_2);
and ( n25014 , n25013 , n55811 );
and ( n25015 , C0 , RI1754c610_2);
or ( n55812 , n25014 , n25015 );
buf ( n55813 , n55812 );
not ( n55814 , n40719 );
and ( n55815 , n55814 , n42083 );
xor ( n55816 , n40700 , n55815 );
not ( n25016 , n29614 );
and ( n25017 , n25016 , RI1740afc8_1454);
and ( n25018 , n55816 , n29614 );
or ( n55817 , n25017 , n25018 );
not ( n25019 , RI1754c610_2);
and ( n25020 , n25019 , n55817 );
and ( n25021 , C0 , RI1754c610_2);
or ( n55818 , n25020 , n25021 );
buf ( n55819 , n55818 );
not ( n55820 , n49853 );
and ( n55821 , n55820 , n48932 );
xor ( n55822 , n51152 , n55821 );
not ( n25022 , n29614 );
and ( n25023 , n25022 , RI173d9c48_1694);
and ( n25024 , n55822 , n29614 );
or ( n55823 , n25023 , n25024 );
not ( n25025 , RI1754c610_2);
and ( n25026 , n25025 , n55823 );
and ( n25027 , C0 , RI1754c610_2);
or ( n55824 , n25026 , n25027 );
buf ( n55825 , n55824 );
not ( n55826 , n41952 );
and ( n55827 , n55826 , n51050 );
xor ( n55828 , n41949 , n55827 );
not ( n25028 , n29614 );
and ( n25029 , n25028 , RI173b9f98_1849);
and ( n25030 , n55828 , n29614 );
or ( n55829 , n25029 , n25030 );
not ( n25031 , RI1754c610_2);
and ( n25032 , n25031 , n55829 );
and ( n25033 , C0 , RI1754c610_2);
or ( n55830 , n25032 , n25033 );
buf ( n55831 , n55830 );
and ( n55832 , RI1754b710_34 , n34844 );
and ( n55833 , RI1754b710_34 , n34847 );
and ( n55834 , RI1754b710_34 , n34850 );
and ( n55835 , RI1754b710_34 , n34852 );
buf ( n55836 , n34854 );
or ( n55837 , n55832 , n55833 , n55834 , n55835 , n55836 , C0 , C0 , C0 );
not ( n25034 , n34859 );
and ( n25035 , n25034 , n55837 );
and ( n25036 , RI1754b710_34 , n34859 );
or ( n55838 , n25035 , n25036 );
not ( n25037 , RI19a22f70_2797);
and ( n25038 , n25037 , n55838 );
and ( n25039 , C0 , RI19a22f70_2797);
or ( n55839 , n25038 , n25039 );
not ( n25040 , n27683 );
and ( n25041 , n25040 , RI19aaf448_2459);
and ( n25042 , n55839 , n27683 );
or ( n55840 , n25041 , n25042 );
not ( n25043 , RI1754c610_2);
and ( n25044 , n25043 , n55840 );
and ( n25045 , C0 , RI1754c610_2);
or ( n55841 , n25044 , n25045 );
buf ( n55842 , n55841 );
not ( n55843 , n43872 );
and ( n55844 , n55843 , n43874 );
xor ( n55845 , n52515 , n55844 );
not ( n25046 , n29614 );
and ( n25047 , n25046 , RI17525088_651);
and ( n25048 , n55845 , n29614 );
or ( n55846 , n25047 , n25048 );
not ( n25049 , RI1754c610_2);
and ( n25050 , n25049 , n55846 );
and ( n25051 , C0 , RI1754c610_2);
or ( n55847 , n25050 , n25051 );
buf ( n55848 , n55847 );
not ( n55849 , n42071 );
and ( n55850 , n55849 , n42073 );
xor ( n55851 , n45456 , n55850 );
not ( n25052 , n29614 );
and ( n25053 , n25052 , RI174098d0_1461);
and ( n25054 , n55851 , n29614 );
or ( n55852 , n25053 , n25054 );
not ( n25055 , RI1754c610_2);
and ( n25056 , n25055 , n55852 );
and ( n25057 , C0 , RI1754c610_2);
or ( n55853 , n25056 , n25057 );
buf ( n55854 , n55853 );
not ( n55855 , n47306 );
and ( n55856 , n55855 , n47308 );
xor ( n55857 , n48182 , n55856 );
not ( n25058 , n29614 );
and ( n25059 , n25058 , RI1745d228_1282);
and ( n25060 , n55857 , n29614 );
or ( n55858 , n25059 , n25060 );
not ( n25061 , RI1754c610_2);
and ( n25062 , n25061 , n55858 );
and ( n25063 , C0 , RI1754c610_2);
or ( n55859 , n25062 , n25063 );
buf ( n55860 , n55859 );
not ( n55861 , n46350 );
and ( n55862 , n55861 , n44857 );
xor ( n55863 , n42997 , n55862 );
not ( n25064 , n29614 );
and ( n25065 , n25064 , RI174744f0_1169);
and ( n25066 , n55863 , n29614 );
or ( n55864 , n25065 , n25066 );
not ( n25067 , RI1754c610_2);
and ( n25068 , n25067 , n55864 );
and ( n25069 , C0 , RI1754c610_2);
or ( n55865 , n25068 , n25069 );
buf ( n55866 , n55865 );
not ( n55867 , n46838 );
and ( n55868 , n55867 , n46840 );
xor ( n55869 , n44206 , n55868 );
not ( n25070 , n29614 );
and ( n25071 , n25070 , RI17469708_1222);
and ( n25072 , n55869 , n29614 );
or ( n55870 , n25071 , n25072 );
not ( n25073 , RI1754c610_2);
and ( n25074 , n25073 , n55870 );
and ( n25075 , C0 , RI1754c610_2);
or ( n55871 , n25074 , n25075 );
buf ( n55872 , n55871 );
not ( n25076 , n34859 );
and ( n25077 , n25076 , C0 );
and ( n25078 , RI1754a9f0_62 , n34859 );
or ( n55873 , n25077 , n25078 );
not ( n25079 , RI19a22f70_2797);
and ( n25080 , n25079 , n55873 );
and ( n25081 , C0 , RI19a22f70_2797);
or ( n55874 , n25080 , n25081 );
not ( n25082 , n27683 );
and ( n25083 , n25082 , RI19a94df0_2648);
and ( n25084 , n55874 , n27683 );
or ( n55875 , n25083 , n25084 );
not ( n25085 , RI1754c610_2);
and ( n25086 , n25085 , n55875 );
and ( n25087 , C0 , RI1754c610_2);
or ( n55876 , n25086 , n25087 );
buf ( n55877 , n55876 );
and ( n55878 , RI19a247d0_2785 , n43086 );
not ( n25088 , n43088 );
and ( n25089 , n25088 , RI19a24578_2786);
and ( n25090 , n55878 , n43088 );
or ( n55879 , n25089 , n25090 );
not ( n25091 , RI1754c610_2);
and ( n25092 , n25091 , n55879 );
and ( n25093 , C0 , RI1754c610_2);
or ( n55880 , n25092 , n25093 );
buf ( n55881 , n55880 );
not ( n55882 , n42158 );
and ( n55883 , n55882 , n42160 );
xor ( n55884 , n44072 , n55883 );
not ( n25094 , n29614 );
and ( n25095 , n25094 , RI173e43a0_1643);
and ( n25096 , n55884 , n29614 );
or ( n55885 , n25095 , n25096 );
not ( n25097 , RI1754c610_2);
and ( n25098 , n25097 , n55885 );
and ( n25099 , C0 , RI1754c610_2);
or ( n55886 , n25098 , n25099 );
buf ( n55887 , n55886 );
not ( n55888 , n51401 );
and ( n55889 , n55888 , n50215 );
xor ( n55890 , n43153 , n55889 );
not ( n25100 , n29614 );
and ( n25101 , n25100 , RI173a3018_1961);
and ( n25102 , n55890 , n29614 );
or ( n55891 , n25101 , n25102 );
not ( n25103 , RI1754c610_2);
and ( n25104 , n25103 , n55891 );
and ( n25105 , C0 , RI1754c610_2);
or ( n55892 , n25104 , n25105 );
buf ( n55893 , n55892 );
and ( n55894 , RI1754b8f0_30 , n34844 );
and ( n55895 , RI1754b8f0_30 , n34847 );
and ( n55896 , RI1754b8f0_30 , n34850 );
and ( n55897 , RI1754b8f0_30 , n34852 );
or ( n55898 , n55894 , n55895 , n55896 , n55897 , C0 , C0 , C0 , C0 );
not ( n25106 , n34859 );
and ( n25107 , n25106 , n55898 );
and ( n25108 , RI1754b8f0_30 , n34859 );
or ( n55899 , n25107 , n25108 );
not ( n25109 , RI19a22f70_2797);
and ( n25110 , n25109 , n55899 );
and ( n25111 , C0 , RI19a22f70_2797);
or ( n55900 , n25110 , n25111 );
not ( n25112 , n27683 );
and ( n25113 , n25112 , RI19aa8f80_2503);
and ( n25114 , n55900 , n27683 );
or ( n55901 , n25113 , n25114 );
not ( n25115 , RI1754c610_2);
and ( n25116 , n25115 , n55901 );
and ( n25117 , C0 , RI1754c610_2);
or ( n55902 , n25116 , n25117 );
buf ( n55903 , n55902 );
not ( n25118 , n27683 );
and ( n25119 , n25118 , RI19ab9c18_2382);
and ( n25120 , RI19ac2840_2310 , n27683 );
or ( n55904 , n25119 , n25120 );
not ( n25121 , RI1754c610_2);
and ( n25122 , n25121 , n55904 );
and ( n25123 , C0 , RI1754c610_2);
or ( n55905 , n25122 , n25123 );
buf ( n55906 , n55905 );
not ( n25124 , n27683 );
and ( n25125 , n25124 , RI19a8f3f0_2688);
and ( n25126 , RI19a99440_2617 , n27683 );
or ( n55907 , n25125 , n25126 );
not ( n25127 , RI1754c610_2);
and ( n25128 , n25127 , n55907 );
and ( n25129 , C0 , RI1754c610_2);
or ( n55908 , n25128 , n25129 );
buf ( n55909 , n55908 );
not ( n55910 , n48380 );
and ( n55911 , n55910 , n51420 );
xor ( n55912 , n48377 , n55911 );
not ( n25130 , n29614 );
nand ( n25131 , n25130 , RI1745aac8_1294);
nand ( n25132 , n55912 , n29614 );
xor ( n55913 , n25131 , n25132 );
not ( n25133 , RI1754c610_2);
and ( n25134 , n25133 , n55913 );
and ( n25135 , C0 , RI1754c610_2);
or ( n55914 , n25134 , n25135 );
buf ( n55915 , n55914 );
not ( n55916 , n49037 );
and ( n55917 , n55916 , n51238 );
xor ( n55918 , n48916 , n55917 );
not ( n25136 , n29614 );
and ( n25137 , n25136 , RI173ce470_1750);
and ( n25138 , n55918 , n29614 );
or ( n55919 , n25137 , n25138 );
not ( n25139 , RI1754c610_2);
and ( n25140 , n25139 , n55919 );
and ( n25141 , C0 , RI1754c610_2);
or ( n55920 , n25140 , n25141 );
buf ( n55921 , n55920 );
not ( n25142 , RI1754c610_2);
and ( n25143 , n25142 , RI17538c00_591);
and ( n25144 , C0 , RI1754c610_2);
or ( n55922 , n25143 , n25144 );
buf ( n55923 , n55922 );
not ( n25145 , n27683 );
and ( n25146 , n25145 , RI19aae980_2464);
and ( n25147 , RI19ab8430_2393 , n27683 );
or ( n55924 , n25146 , n25147 );
not ( n25148 , RI1754c610_2);
and ( n25149 , n25148 , n55924 );
and ( n25150 , C0 , RI1754c610_2);
or ( n55925 , n25149 , n25150 );
buf ( n55926 , n55925 );
not ( n55927 , n41886 );
and ( n55928 , n55927 , n46593 );
xor ( n55929 , n41870 , n55928 );
not ( n25151 , n29614 );
and ( n25152 , n25151 , RI17447310_1389);
and ( n25153 , n55929 , n29614 );
or ( n55930 , n25152 , n25153 );
not ( n25154 , RI1754c610_2);
and ( n25155 , n25154 , n55930 );
and ( n25156 , C0 , RI1754c610_2);
or ( n55931 , n25155 , n25156 );
buf ( n55932 , n55931 );
not ( n55933 , n45716 );
and ( n55934 , n55933 , n45718 );
xor ( n55935 , n51078 , n55934 );
not ( n25157 , n29614 );
and ( n25158 , n25157 , RI174aa730_905);
and ( n25159 , n55935 , n29614 );
or ( n55936 , n25158 , n25159 );
not ( n25160 , RI1754c610_2);
and ( n25161 , n25160 , n55936 );
and ( n25162 , C0 , RI1754c610_2);
or ( n55937 , n25161 , n25162 );
buf ( n55938 , n55937 );
not ( n55939 , n44685 );
and ( n55940 , n55939 , n44687 );
xor ( n55941 , n52286 , n55940 );
not ( n25163 , n29614 );
and ( n25164 , n25163 , RI173b8f30_1854);
and ( n25165 , n55941 , n29614 );
or ( n55942 , n25164 , n25165 );
not ( n25166 , RI1754c610_2);
and ( n25167 , n25166 , n55942 );
and ( n25168 , C0 , RI1754c610_2);
or ( n55943 , n25167 , n25168 );
buf ( n55944 , n55943 );
not ( n55945 , n40829 );
and ( n55946 , n55945 , n40831 );
xor ( n55947 , n39953 , n55946 );
not ( n25169 , n29614 );
and ( n25170 , n25169 , RI173b3698_1881);
and ( n25171 , n55947 , n29614 );
or ( n55948 , n25170 , n25171 );
not ( n25172 , RI1754c610_2);
and ( n25173 , n25172 , n55948 );
and ( n25174 , C0 , RI1754c610_2);
or ( n55949 , n25173 , n25174 );
buf ( n55950 , n55949 );
not ( n55951 , n50967 );
and ( n55952 , n55951 , n47839 );
xor ( n55953 , n38726 , n55952 );
not ( n25175 , n29614 );
and ( n25176 , n25175 , RI1746efa0_1195);
and ( n25177 , n55953 , n29614 );
or ( n55954 , n25176 , n25177 );
not ( n25178 , RI1754c610_2);
and ( n25179 , n25178 , n55954 );
and ( n25180 , C0 , RI1754c610_2);
or ( n55955 , n25179 , n25180 );
buf ( n55956 , n55955 );
not ( n55957 , n44115 );
and ( n55958 , n55957 , n42235 );
xor ( n55959 , n53957 , n55958 );
not ( n25181 , n29614 );
and ( n25182 , n25181 , RI1746c1b0_1209);
and ( n25183 , n55959 , n29614 );
or ( n55960 , n25182 , n25183 );
not ( n25184 , RI1754c610_2);
and ( n25185 , n25184 , n55960 );
and ( n25186 , C0 , RI1754c610_2);
or ( n55961 , n25185 , n25186 );
buf ( n55962 , n55961 );
not ( n55963 , n38838 );
and ( n55964 , n55963 , n45164 );
xor ( n55965 , n38835 , n55964 );
not ( n25187 , n29614 );
and ( n25188 , n25187 , RI17462ac0_1255);
and ( n25189 , n55965 , n29614 );
or ( n55966 , n25188 , n25189 );
not ( n25190 , RI1754c610_2);
and ( n25191 , n25190 , n55966 );
and ( n25192 , C0 , RI1754c610_2);
or ( n55967 , n25191 , n25192 );
buf ( n55968 , n55967 );
not ( n25193 , n27683 );
and ( n25194 , n25193 , RI19acd358_2230);
and ( n25195 , RI19a8b958_2714 , n27683 );
or ( n55969 , n25194 , n25195 );
not ( n25196 , RI1754c610_2);
and ( n25197 , n25196 , n55969 );
and ( n25198 , C0 , RI1754c610_2);
or ( n55970 , n25197 , n25198 );
buf ( n55971 , n55970 );
not ( n55972 , n52989 );
and ( n55973 , n55972 , n54991 );
xor ( n55974 , n52186 , n55973 );
not ( n25199 , n29614 );
and ( n25200 , n25199 , RI173c2620_1808);
and ( n25201 , n55974 , n29614 );
or ( n55975 , n25200 , n25201 );
not ( n25202 , RI1754c610_2);
and ( n25203 , n25202 , n55975 );
and ( n25204 , C0 , RI1754c610_2);
or ( n55976 , n25203 , n25204 );
buf ( n55977 , n55976 );
not ( n55978 , n39291 );
and ( n55979 , n55978 , n42225 );
xor ( n55980 , n39285 , n55979 );
not ( n25205 , n29614 );
and ( n25206 , n25205 , RI1738fef0_2054);
and ( n25207 , n55980 , n29614 );
or ( n55981 , n25206 , n25207 );
not ( n25208 , RI1754c610_2);
and ( n25209 , n25208 , n55981 );
and ( n25210 , C0 , RI1754c610_2);
or ( n55982 , n25209 , n25210 );
buf ( n55983 , n55982 );
not ( n25211 , RI1754c610_2);
and ( n25212 , n25211 , RI19ad0958_2207);
and ( n25213 , C0 , RI1754c610_2);
or ( n55984 , n25212 , n25213 );
buf ( n55985 , n55984 );
not ( n55986 , n35070 );
and ( n55987 , n55986 , n46507 );
xor ( n55988 , n35011 , n55987 );
not ( n25214 , n29614 );
and ( n25215 , n25214 , RI173cca30_1758);
and ( n25216 , n55988 , n29614 );
or ( n55989 , n25215 , n25216 );
not ( n25217 , RI1754c610_2);
and ( n25218 , n25217 , n55989 );
and ( n25219 , C0 , RI1754c610_2);
or ( n55990 , n25218 , n25219 );
buf ( n55991 , n55990 );
not ( n55992 , n51357 );
and ( n55993 , n55992 , n42873 );
xor ( n55994 , n51354 , n55993 );
not ( n25220 , n29614 );
and ( n25221 , n25220 , RI17407e90_1469);
and ( n25222 , n55994 , n29614 );
or ( n55995 , n25221 , n25222 );
not ( n25223 , RI1754c610_2);
and ( n25224 , n25223 , n55995 );
and ( n25225 , C0 , RI1754c610_2);
or ( n55996 , n25224 , n25225 );
buf ( n55997 , n55996 );
not ( n55998 , n50163 );
and ( n55999 , n55998 , n41692 );
xor ( n56000 , n40968 , n55999 );
not ( n25226 , n29614 );
and ( n25227 , n25226 , RI173b0560_1896);
and ( n25228 , n56000 , n29614 );
or ( n56001 , n25227 , n25228 );
not ( n25229 , RI1754c610_2);
and ( n25230 , n25229 , n56001 );
and ( n25231 , C0 , RI1754c610_2);
or ( n56002 , n25230 , n25231 );
buf ( n56003 , n56002 );
not ( n56004 , n49095 );
and ( n56005 , n56004 , n51086 );
xor ( n56006 , n47639 , n56005 );
not ( n25232 , n29614 );
and ( n25233 , n25232 , RI17518c98_689);
and ( n25234 , n56006 , n29614 );
or ( n56007 , n25233 , n25234 );
not ( n25235 , RI1754c610_2);
and ( n25236 , n25235 , n56007 );
and ( n25237 , C0 , RI1754c610_2);
or ( n56008 , n25236 , n25237 );
buf ( n56009 , n56008 );
buf ( n56010 , RI1746df38_1200);
buf ( n56011 , RI174989b8_992);
not ( n56012 , n48737 );
and ( n56013 , n56012 , n50028 );
xor ( n56014 , n48734 , n56013 );
not ( n25238 , n29614 );
and ( n25239 , n25238 , RI1749baf0_977);
and ( n25240 , n56014 , n29614 );
or ( n56015 , n25239 , n25240 );
not ( n25241 , RI1754c610_2);
and ( n25242 , n25241 , n56015 );
and ( n25243 , C0 , RI1754c610_2);
or ( n56016 , n25242 , n25243 );
buf ( n56017 , n56016 );
buf ( n56018 , RI174bb878_827);
not ( n56019 , n48451 );
and ( n56020 , n56019 , n49770 );
xor ( n56021 , n48448 , n56020 );
not ( n25244 , n29614 );
and ( n25245 , n25244 , RI173eda90_1597);
and ( n25246 , n56021 , n29614 );
or ( n56022 , n25245 , n25246 );
not ( n25247 , RI1754c610_2);
and ( n25248 , n25247 , n56022 );
and ( n25249 , C0 , RI1754c610_2);
or ( n56023 , n25248 , n25249 );
buf ( n56024 , n56023 );
not ( n25250 , n27683 );
and ( n25251 , n25250 , RI19a9e030_2584);
and ( n25252 , RI19aa7a68_2512 , n27683 );
or ( n56025 , n25251 , n25252 );
not ( n25253 , RI1754c610_2);
and ( n25254 , n25253 , n56025 );
and ( n25255 , C0 , RI1754c610_2);
or ( n56026 , n25254 , n25255 );
buf ( n56027 , n56026 );
not ( n56028 , n50065 );
and ( n56029 , n56028 , n43945 );
xor ( n56030 , n48048 , n56029 );
not ( n25256 , n29614 );
and ( n25257 , n25256 , RI17503398_750);
and ( n25258 , n56030 , n29614 );
or ( n56031 , n25257 , n25258 );
not ( n25259 , RI1754c610_2);
and ( n25260 , n25259 , n56031 );
and ( n25261 , C0 , RI1754c610_2);
or ( n56032 , n25260 , n25261 );
buf ( n56033 , n56032 );
not ( n56034 , n52027 );
and ( n56035 , n56034 , n52337 );
xor ( n56036 , n45878 , n56035 );
not ( n25262 , n29614 );
and ( n25263 , n25262 , RI174c4e00_798);
and ( n25264 , n56036 , n29614 );
or ( n56037 , n25263 , n25264 );
not ( n25265 , RI1754c610_2);
and ( n25266 , n25265 , n56037 );
and ( n25267 , C0 , RI1754c610_2);
or ( n56038 , n25266 , n25267 );
buf ( n56039 , n56038 );
not ( n56040 , n49696 );
and ( n56041 , n56040 , n42777 );
xor ( n56042 , n41257 , n56041 );
not ( n25268 , n29614 );
and ( n25269 , n25268 , RI17448a08_1382);
and ( n25270 , n56042 , n29614 );
or ( n56043 , n25269 , n25270 );
not ( n25271 , RI1754c610_2);
and ( n25272 , n25271 , n56043 );
and ( n25273 , C0 , RI1754c610_2);
or ( n56044 , n25272 , n25273 );
buf ( n56045 , n56044 );
not ( n56046 , n46934 );
and ( n56047 , n56046 , n39314 );
xor ( n56048 , n46791 , n56047 );
not ( n25274 , n29614 );
and ( n25275 , n25274 , RI1738a658_2081);
and ( n25276 , n56048 , n29614 );
or ( n56049 , n25275 , n25276 );
not ( n25277 , RI1754c610_2);
and ( n25278 , n25277 , n56049 );
and ( n25279 , C0 , RI1754c610_2);
or ( n56050 , n25278 , n25279 );
buf ( n56051 , n56050 );
not ( n25280 , n27683 );
and ( n25281 , n25280 , RI19acbe40_2240);
and ( n25282 , RI19a87920_2741 , n27683 );
or ( n56052 , n25281 , n25282 );
not ( n25283 , RI1754c610_2);
and ( n25284 , n25283 , n56052 );
and ( n25285 , C0 , RI1754c610_2);
or ( n56053 , n25284 , n25285 );
buf ( n56054 , n56053 );
not ( n25286 , n27683 );
and ( n25287 , n25286 , RI19aa7a68_2512);
and ( n25288 , RI19ab1860_2442 , n27683 );
or ( n56055 , n25287 , n25288 );
not ( n25289 , RI1754c610_2);
and ( n25290 , n25289 , n56055 );
and ( n25291 , C0 , RI1754c610_2);
or ( n56056 , n25290 , n25291 );
buf ( n56057 , n56056 );
not ( n56058 , n46116 );
and ( n56059 , n56058 , n48892 );
xor ( n56060 , n46113 , n56059 );
not ( n25292 , n29614 );
and ( n25293 , n25292 , RI173a9fa8_1927);
and ( n25294 , n56060 , n29614 );
or ( n56061 , n25293 , n25294 );
not ( n25295 , RI1754c610_2);
and ( n25296 , n25295 , n56061 );
and ( n25297 , C0 , RI1754c610_2);
or ( n56062 , n25296 , n25297 );
buf ( n56063 , n56062 );
not ( n56064 , n41069 );
and ( n56065 , n56064 , n49705 );
xor ( n56066 , n41050 , n56065 );
not ( n25298 , n29614 );
and ( n25299 , n25298 , RI174693c0_1223);
and ( n25300 , n56066 , n29614 );
or ( n56067 , n25299 , n25300 );
not ( n25301 , RI1754c610_2);
and ( n25302 , n25301 , n56067 );
and ( n25303 , C0 , RI1754c610_2);
or ( n56068 , n25302 , n25303 );
buf ( n56069 , n56068 );
not ( n56070 , n48986 );
and ( n56071 , n56070 , n42388 );
xor ( n56072 , n33176 , n56071 );
not ( n25304 , n29614 );
and ( n25305 , n25304 , RI17528418_641);
and ( n25306 , n56072 , n29614 );
or ( n56073 , n25305 , n25306 );
not ( n25307 , RI1754c610_2);
and ( n25308 , n25307 , n56073 );
and ( n25309 , C0 , RI1754c610_2);
or ( n56074 , n25308 , n25309 );
buf ( n56075 , n56074 );
not ( n25310 , n27683 );
and ( n25311 , n25310 , RI19a8c240_2710);
and ( n25312 , RI19a96290_2639 , n27683 );
or ( n56076 , n25311 , n25312 );
not ( n25313 , RI1754c610_2);
and ( n25314 , n25313 , n56076 );
and ( n25315 , C0 , RI1754c610_2);
or ( n56077 , n25314 , n25315 );
buf ( n56078 , n56077 );
and ( C0 , n27688 , RI1753aa78_586 );
or ( C1 , n27688 , RI1753aa78_586 );
endmodule

