//NOTE: no-implementation module stub

module GtCLK_NOT (
    output Z,
    input A
);

endmodule
