// IWLS benchmark module "z4ml" printed on Wed May 29 17:30:39 2002
module z4ml(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \24 , \25 , \26 , \27 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ;
output
  \24 ,
  \25 ,
  \26 ,
  \27 ;
wire
  \[2] ,
  \[12] ,
  \[3] ,
  \[8] ,
  \[4] ,
  \[9] ,
  \[10] ,
  \[1] ;
assign
  \[2]  = (\[8]  & (~\[3]  & (\5  & \2 ))) | ((\6  & (\5  & (\3  & \2 ))) | ((\[8]  & (~\[3]  & ~\[1] )) | ((~\[1]  & (\6  & \3 )) | (\[10]  & ~\[1] )))),
  \[12]  = (~\4  & ~\1 ) | (\4  & \1 ),
  \[3]  = (~\[9]  & ~\[8] ) | (\[9]  & \[8] ),
  \[8]  = (~\[4]  & \1 ) | (\7  & \4 ),
  \[4]  = (~\[12]  & ~\7 ) | (\[12]  & \7 ),
  \[9]  = (~\6  & ~\3 ) | (\6  & \3 ),
  \24  = \[1] ,
  \25  = \[2] ,
  \26  = \[3] ,
  \27  = \[4] ,
  \[10]  = \5  | \2 ,
  \[1]  = (\[10]  & (\[8]  & \6 )) | ((\[10]  & (~\[3]  & \3 )) | (\5  & \2 ));
endmodule

