module add_2_6_8(a, b, c);
  input [1:0] a;
  input [5:0] b;
  output [7:0] c;
  assign c = a + b;
endmodule
