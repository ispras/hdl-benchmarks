//NOTE: no-implementation module stub

module EMC (
    input `ifdef FD_EVB PERICLK, `else DSPCLK, `endif
    input GRST,
    input PPclr_h,
    input [15:0] DMDin,
    input T_selECM,
    input PM_bdry_sel,
    input GO_Fx,
    input GO_Ex,
    input GO_EC,
    input ECYC,
    input BGn,
    input [7:0] PMOVL_dsp,
    input [3:0] DMOVL_dsp,
    input Dummy_E,
    input [10:0] IOaddr,
    input Double_E,
    input accCM_E,
    input rdCM_E,
    input [13:0] DMA,
    input [13:0] PMA,
    input WSCR_we,
    input WSCR_ext_we,
    input EXTC_Eg,
    input Pread_Ei,
    input Pwrite_Ei,
    input Dread_Ei,
    input Dwrite_Ei,
    input IOcmd_Ei,
    input IOread_Ei,
    input IOwrite_Ei,
    input MMR_web,
    input [13:0] CMAin,
    input [1:0] ECMAWAIT,
    input [23:0] IDR,
    input [7:0] T_EA,
    input [15:0] T_ED,
    input [15:0] PMDin,
    input [23:0] CM_rd,
    input BDMAmode,
    input [7:0] BMpage,
    input BDIR,
    input [7:0] BWdataBUF,
    input BWRn,
    input [13:0] BEAD,
    input BSreq,
    input BSack,
    input BWend,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input EA_oe,
    input [14:0] EA_do,
    input ED_oe,
    input [15:0] ED_do,
    input PMSn,
    input DMSn,
    input IOSn,
    input BMSn,
    input CMSn,
    input RDn,
    input WRn,
    input ECMSn,
    input ECMA_EN,
    input eRDY,
    input [14:0] WSCR,
    input [7:0] WSCR_ext,
    input emcDMD_oe,
    input [15:0] emcDMD_do,
    input emcPMD_oe,
    input [15:0] emcPMD_do,
    input [23:0] CM_rdata,
    input ENS12,
    input ECS12,
    input ENS13,
    input ECS13,
    input ENS14,
    input ECS14,
    input ENS0,
    input BMcs
);

endmodule
