module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 ;
output g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 ;
wire t_0 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( n199 , g198 );
buf ( n200 , g199 );
buf ( n201 , g200 );
buf ( n202 , g201 );
buf ( n203 , g202 );
buf ( n204 , g203 );
buf ( n205 , g204 );
buf ( n206 , g205 );
buf ( n207 , g206 );
buf ( n208 , g207 );
buf ( n209 , g208 );
buf ( n210 , g209 );
buf ( n211 , g210 );
buf ( n212 , g211 );
buf ( n213 , g212 );
buf ( n214 , g213 );
buf ( n215 , g214 );
buf ( n216 , g215 );
buf ( n217 , g216 );
buf ( n218 , g217 );
buf ( n219 , g218 );
buf ( n220 , g219 );
buf ( n221 , g220 );
buf ( n222 , g221 );
buf ( n223 , g222 );
buf ( n224 , g223 );
buf ( n225 , g224 );
buf ( n226 , g225 );
buf ( n227 , g226 );
buf ( n228 , g227 );
buf ( n229 , g228 );
buf ( n230 , g229 );
buf ( n231 , g230 );
buf ( n232 , g231 );
buf ( n233 , g232 );
buf ( n234 , g233 );
buf ( n235 , g234 );
buf ( n236 , g235 );
buf ( n237 , g236 );
buf ( n238 , g237 );
buf ( n239 , g238 );
buf ( n240 , g239 );
buf ( n241 , g240 );
buf ( n242 , g241 );
buf ( n243 , g242 );
buf ( n244 , g243 );
buf ( n245 , g244 );
buf ( g245 , n246 );
buf ( g246 , n247 );
buf ( g247 , n248 );
buf ( g248 , n249 );
buf ( g249 , n250 );
buf ( g250 , n251 );
buf ( g251 , n252 );
buf ( g252 , n253 );
buf ( g253 , n254 );
buf ( g254 , n255 );
buf ( g255 , n256 );
buf ( g256 , n257 );
buf ( g257 , n258 );
buf ( g258 , n259 );
buf ( g259 , n260 );
buf ( g260 , n261 );
buf ( g261 , n262 );
buf ( g262 , n263 );
buf ( g263 , n264 );
buf ( g264 , n265 );
buf ( g265 , n266 );
buf ( g266 , n267 );
buf ( g267 , n268 );
buf ( g268 , n269 );
buf ( g269 , n270 );
buf ( g270 , n271 );
buf ( g271 , n272 );
buf ( g272 , n273 );
buf ( g273 , n274 );
buf ( g274 , n275 );
buf ( g275 , n276 );
buf ( g276 , n277 );
buf ( g277 , n278 );
buf ( g278 , n279 );
buf ( g279 , n280 );
buf ( g280 , n281 );
buf ( g281 , n282 );
buf ( g282 , n283 );
buf ( g283 , n284 );
buf ( g284 , n285 );
buf ( g285 , n286 );
buf ( g286 , n287 );
buf ( g287 , n288 );
buf ( g288 , n289 );
buf ( g289 , n290 );
buf ( g290 , n291 );
buf ( g291 , n292 );
buf ( g292 , n293 );
buf ( g293 , n294 );
buf ( g294 , n295 );
buf ( g295 , n296 );
buf ( g296 , n297 );
buf ( g297 , n298 );
buf ( g298 , n299 );
buf ( g299 , n300 );
buf ( g300 , n301 );
buf ( g301 , n302 );
buf ( g302 , n303 );
buf ( g303 , n304 );
buf ( g304 , n305 );
buf ( g305 , n306 );
buf ( g306 , n307 );
buf ( g307 , n308 );
buf ( g308 , n309 );
buf ( g309 , n310 );
buf ( g310 , n311 );
buf ( g311 , n312 );
buf ( g312 , n313 );
buf ( g313 , n314 );
buf ( g314 , n315 );
buf ( g315 , n316 );
buf ( g316 , n317 );
buf ( g317 , n318 );
buf ( g318 , n319 );
buf ( g319 , n320 );
buf ( g320 , n321 );
buf ( g321 , n322 );
buf ( g322 , n323 );
buf ( g323 , n324 );
buf ( g324 , n325 );
buf ( g325 , n326 );
buf ( g326 , n327 );
buf ( g327 , n328 );
buf ( g328 , n329 );
buf ( g329 , n330 );
buf ( g330 , n331 );
buf ( g331 , n332 );
buf ( g332 , n333 );
buf ( g333 , n334 );
buf ( g334 , n335 );
buf ( g335 , n336 );
buf ( g336 , n337 );
buf ( g337 , n338 );
buf ( g338 , n339 );
buf ( g339 , n340 );
buf ( g340 , n341 );
buf ( g341 , n342 );
buf ( g342 , n343 );
buf ( g343 , n344 );
buf ( g344 , n345 );
buf ( n246 , n3244 );
buf ( n247 , n3292 );
buf ( n248 , n3389 );
buf ( n249 , n3453 );
buf ( n250 , n3635 );
buf ( n251 , n3582 );
buf ( n252 , n3758 );
buf ( n253 , n3861 );
buf ( n254 , n3510 );
buf ( n255 , n3549 );
buf ( n256 , n3820 );
buf ( n257 , n3519 );
buf ( n258 , n3825 );
buf ( n259 , n3649 );
buf ( n260 , n3671 );
buf ( n261 , n3867 );
buf ( n262 , n3737 );
buf ( n263 , n3747 );
buf ( n264 , n3836 );
buf ( n265 , n3345 );
buf ( n266 , n3715 );
buf ( n267 , n3801 );
buf ( n268 , n3726 );
buf ( n269 , n3768 );
buf ( n270 , n3847 );
buf ( n271 , n4665 );
buf ( n272 , n3918 );
buf ( n273 , n3879 );
buf ( n274 , n3888 );
buf ( n275 , n3924 );
buf ( n276 , n3893 );
buf ( n277 , n3912 );
buf ( n278 , n3929 );
buf ( n279 , n3964 );
buf ( n280 , n3954 );
buf ( n281 , n2906 );
buf ( n282 , n3968 );
buf ( n283 , n3973 );
buf ( n284 , n4675 );
buf ( n285 , n3898 );
buf ( n286 , n3903 );
buf ( n287 , n3978 );
buf ( n288 , n3982 );
buf ( n289 , n3997 );
buf ( n290 , n3934 );
buf ( n291 , n3939 );
buf ( n292 , n3959 );
buf ( n293 , n3944 );
buf ( n294 , n3988 );
buf ( n295 , n3993 );
buf ( n296 , n4630 );
buf ( n297 , n4635 );
buf ( n298 , n3949 );
buf ( n299 , n4639 );
buf ( n300 , n4661 );
buf ( n301 , n4259 );
buf ( n302 , n4284 );
buf ( n303 , n4310 );
buf ( n304 , n4328 );
buf ( n305 , n4363 );
buf ( n306 , n4382 );
buf ( n307 , n4402 );
buf ( n308 , n4417 );
buf ( n309 , n4438 );
buf ( n310 , n4453 );
buf ( n311 , n4471 );
buf ( n312 , n4486 );
buf ( n313 , n4507 );
buf ( n314 , n4524 );
buf ( n315 , n4543 );
buf ( n316 , n4568 );
buf ( n317 , n4585 );
buf ( n318 , n4603 );
buf ( n319 , n4613 );
buf ( n320 , n4626 );
buf ( n321 , n3883 );
buf ( n322 , n4670 );
buf ( n323 , n4643 );
buf ( n324 , n4647 );
buf ( n325 , n4651 );
buf ( n326 , n4654 );
buf ( n327 , n4657 );
buf ( n328 , n4744 );
buf ( n329 , n4716 );
buf ( n330 , n4749 );
buf ( n331 , n4721 );
buf ( n332 , n4741 );
buf ( n333 , n4731 );
buf ( n334 , n4752 );
buf ( n335 , n4761 );
buf ( n336 , n4681 );
buf ( n337 , n4701 );
buf ( n338 , n4706 );
buf ( n339 , n4696 );
buf ( n340 , n4691 );
buf ( n341 , n4726 );
buf ( n342 , n4711 );
buf ( n343 , n4736 );
buf ( n344 , n4686 );
buf ( n345 , n4757 );
not ( n348 , n1 );
and ( n349 , n348 , n31 );
not ( n350 , n348 );
not ( n351 , n31 );
nor ( n352 , n6 , n7 );
nor ( n353 , n4 , n12 );
nor ( n354 , n5 , n13 );
nand ( n355 , n352 , n353 , n354 );
not ( n356 , n355 );
nor ( n357 , n8 , n14 );
nor ( n358 , n15 , n17 );
nor ( n359 , n2 , n11 );
nor ( n360 , n9 , n16 );
nand ( n361 , n358 , n359 , n360 );
not ( n362 , n3 );
not ( n363 , n10 );
nand ( n364 , n362 , n363 );
nor ( n365 , n361 , n364 );
nand ( n366 , n356 , n357 , n365 );
not ( n367 , n366 );
nor ( n368 , n28 , n32 );
not ( n369 , n368 );
not ( n370 , n29 );
not ( n371 , n20 );
nor ( n372 , n18 , n19 );
nand ( n373 , n370 , n371 , n372 );
nor ( n374 , n369 , n373 );
nand ( n375 , n367 , n374 );
nor ( n376 , n30 , n375 );
not ( n377 , n376 );
or ( n378 , n351 , n377 );
or ( n379 , n376 , n31 );
nand ( n380 , n378 , n379 );
and ( n381 , n350 , n380 );
nor ( n382 , n349 , n381 );
not ( n383 , n382 );
not ( n384 , n383 );
not ( n385 , n27 );
not ( n386 , n25 );
not ( n387 , n26 );
not ( n388 , n24 );
not ( n389 , n23 );
nor ( n390 , n21 , n22 );
nand ( n391 , n388 , n389 , n390 );
not ( n392 , n391 );
not ( n393 , n392 );
not ( n394 , n393 );
nand ( n395 , n360 , n359 , n358 );
not ( n396 , n395 );
nor ( n397 , n8 , n14 );
nor ( n398 , n3 , n10 );
nand ( n399 , n396 , n356 , n397 , n398 );
buf ( n400 , n399 );
not ( n401 , n400 );
not ( n402 , n29 );
not ( n403 , n20 );
nor ( n404 , n18 , n19 );
nand ( n405 , n402 , n403 , n404 );
not ( n406 , n405 );
not ( n407 , n30 );
not ( n408 , n31 );
nand ( n409 , n406 , n368 , n407 , n408 );
not ( n410 , n409 );
nand ( n411 , n401 , n410 );
not ( n412 , n411 );
and ( n413 , n386 , n387 , n394 , n412 );
nand ( n414 , n385 , n1 , n413 );
not ( n415 , n414 );
buf ( n416 , n415 );
not ( n417 , n416 );
not ( n418 , n1 );
and ( n419 , n418 , n32 );
not ( n420 , n418 );
not ( n421 , n373 );
not ( n422 , n366 );
and ( n423 , n421 , n422 );
and ( n424 , n423 , n32 );
not ( n425 , n423 );
not ( n426 , n32 );
and ( n427 , n425 , n426 );
nor ( n428 , n424 , n427 );
not ( n429 , n428 );
and ( n430 , n420 , n429 );
nor ( n431 , n419 , n430 );
not ( n432 , n1 );
and ( n433 , n432 , n30 );
not ( n434 , n432 );
not ( n435 , n30 );
and ( n436 , n375 , n435 );
not ( n437 , n375 );
and ( n438 , n437 , n30 );
nor ( n439 , n436 , n438 );
not ( n440 , n439 );
and ( n441 , n434 , n440 );
nor ( n442 , n433 , n441 );
and ( n443 , n431 , n442 );
not ( n444 , n1 );
nand ( n445 , n29 , n444 );
not ( n446 , n29 );
not ( n447 , n20 );
not ( n448 , n400 );
and ( n449 , n446 , n447 , n372 , n448 );
not ( n450 , n449 );
not ( n451 , n20 );
not ( n452 , n451 );
not ( n453 , n399 );
and ( n454 , n372 , n453 );
not ( n455 , n454 );
or ( n456 , n452 , n455 );
nand ( n457 , n456 , n29 );
nand ( n458 , n450 , n457 , n1 );
and ( n459 , n445 , n458 );
not ( n460 , n1 );
and ( n461 , n460 , n28 );
not ( n462 , n460 );
not ( n463 , n32 );
not ( n464 , n400 );
nand ( n465 , n463 , n421 , n464 );
not ( n466 , n28 );
and ( n467 , n465 , n466 );
not ( n468 , n465 );
and ( n469 , n468 , n28 );
nor ( n470 , n467 , n469 );
not ( n471 , n470 );
and ( n472 , n462 , n471 );
nor ( n473 , n461 , n472 );
and ( n474 , n443 , n459 , n473 );
nor ( n475 , n417 , n474 );
not ( n476 , n1 );
not ( n477 , n7 );
not ( n478 , n6 );
not ( n479 , n8 );
not ( n480 , n9 );
nand ( n481 , n477 , n478 , n479 , n480 );
not ( n482 , n481 );
nor ( n483 , n4 , n5 );
nor ( n484 , n2 , n3 );
nand ( n485 , n482 , n483 , n484 );
not ( n486 , n485 );
nor ( n487 , n12 , n13 );
nor ( n488 , n10 , n11 );
nand ( n489 , n486 , n487 , n488 );
not ( n490 , n14 );
and ( n491 , n489 , n490 );
not ( n492 , n489 );
and ( n493 , n492 , n14 );
nor ( n494 , n491 , n493 );
not ( n495 , n494 );
not ( n496 , n495 );
or ( n497 , n476 , n496 );
not ( n498 , n1 );
nand ( n499 , n14 , n498 );
nand ( n500 , n497 , n499 );
not ( n501 , n8 );
buf ( n502 , n352 );
nand ( n503 , n501 , n502 );
and ( n504 , n503 , n1 );
xor ( n505 , n504 , n9 );
not ( n506 , n505 );
not ( n507 , n506 );
not ( n508 , n5 );
buf ( n509 , n477 );
not ( n510 , n6 );
not ( n511 , n8 );
not ( n512 , n9 );
nand ( n513 , n510 , n511 , n512 );
not ( n514 , n513 );
nand ( n515 , n508 , n484 , n509 , n514 );
not ( n516 , n515 );
not ( n517 , n484 );
nand ( n518 , n509 , n514 );
nor ( n519 , n517 , n518 );
nor ( n520 , n519 , n508 );
nor ( n521 , n516 , n520 );
and ( n522 , n1 , n521 );
not ( n523 , n1 );
and ( n524 , n523 , n5 );
or ( n525 , n522 , n524 );
nor ( n526 , n507 , n525 );
not ( n527 , n1 );
nand ( n528 , n527 , n11 );
nor ( n529 , n485 , n11 );
not ( n530 , n529 );
nand ( n531 , n11 , n485 );
nand ( n532 , n530 , n531 , n1 );
and ( n533 , n528 , n532 );
not ( n534 , n1 );
and ( n535 , n534 , n13 );
not ( n536 , n534 );
not ( n537 , n13 );
not ( n538 , n10 );
not ( n539 , n11 );
nand ( n540 , n538 , n539 );
not ( n541 , n7 );
not ( n542 , n6 );
not ( n543 , n8 );
not ( n544 , n9 );
nand ( n545 , n541 , n542 , n543 , n544 );
not ( n546 , n545 );
nor ( n547 , n2 , n3 );
nand ( n548 , n546 , n483 , n547 );
nor ( n549 , n540 , n548 );
not ( n550 , n549 );
or ( n551 , n537 , n550 );
nor ( n552 , n540 , n485 );
or ( n553 , n552 , n13 );
nand ( n554 , n551 , n553 );
and ( n555 , n536 , n554 );
nor ( n556 , n535 , n555 );
nand ( n557 , n526 , n533 , n556 );
not ( n558 , n8 );
not ( n559 , n1 );
not ( n560 , n559 );
or ( n561 , n558 , n560 );
not ( n562 , n8 );
nor ( n563 , n562 , n502 );
not ( n564 , n563 );
nand ( n565 , n564 , n1 , n503 );
nand ( n566 , n561 , n565 );
buf ( n567 , n566 );
not ( n568 , n1 );
not ( n569 , n18 );
not ( n570 , n569 );
not ( n571 , n19 );
nand ( n572 , n571 , n448 );
not ( n573 , n572 );
or ( n574 , n570 , n573 );
nor ( n575 , n3 , n10 );
nand ( n576 , n575 , n357 , n353 , n354 );
not ( n577 , n576 );
nor ( n578 , n15 , n17 );
nor ( n579 , n2 , n11 );
nor ( n580 , n9 , n16 );
nand ( n581 , n578 , n579 , n580 );
nor ( n582 , n569 , n581 );
nand ( n583 , n577 , n582 , n571 , n502 );
nand ( n584 , n574 , n583 );
not ( n585 , n584 );
or ( n586 , n568 , n585 );
or ( n587 , n569 , n1 );
nand ( n588 , n586 , n587 );
nor ( n589 , n567 , n588 );
not ( n590 , n1 );
and ( n591 , n590 , n10 );
not ( n592 , n590 );
not ( n593 , n10 );
not ( n594 , n529 );
or ( n595 , n593 , n594 );
or ( n596 , n10 , n529 );
nand ( n597 , n595 , n596 );
and ( n598 , n592 , n597 );
nor ( n599 , n591 , n598 );
not ( n600 , n1 );
and ( n601 , n600 , n20 );
not ( n602 , n600 );
and ( n603 , n454 , n20 );
not ( n604 , n454 );
not ( n605 , n20 );
and ( n606 , n604 , n605 );
nor ( n607 , n603 , n606 );
not ( n608 , n607 );
and ( n609 , n602 , n608 );
nor ( n610 , n601 , n609 );
nand ( n611 , n589 , n599 , n610 );
nor ( n612 , n500 , n557 , n611 );
not ( n613 , n612 );
not ( n614 , n6 );
not ( n615 , n515 );
not ( n616 , n4 );
nor ( n617 , n615 , n616 );
not ( n618 , n616 );
not ( n619 , n515 );
not ( n620 , n619 );
or ( n621 , n618 , n620 );
nand ( n622 , n621 , n1 );
or ( n623 , n617 , n622 );
not ( n624 , n1 );
nand ( n625 , n4 , n624 );
nand ( n626 , n623 , n625 );
not ( n627 , n626 );
nand ( n628 , n614 , n627 );
not ( n629 , n1 );
not ( n630 , n481 );
nor ( n631 , n629 , n630 );
not ( n632 , n2 );
xor ( n633 , n631 , n632 );
or ( n634 , n518 , n2 );
nand ( n635 , n634 , n1 );
xnor ( n636 , n635 , n3 );
not ( n637 , n636 );
and ( n638 , n633 , n637 );
not ( n639 , n509 );
not ( n640 , n639 );
not ( n641 , n1 );
not ( n642 , n641 );
or ( n643 , n640 , n642 );
not ( n644 , n509 );
nor ( n645 , n6 , n644 );
not ( n646 , n645 );
not ( n647 , n509 );
nand ( n648 , n6 , n647 );
nand ( n649 , n646 , n648 , n1 );
nand ( n650 , n643 , n649 );
not ( n651 , n650 );
not ( n652 , n1 );
nand ( n653 , n19 , n652 );
and ( n654 , n400 , n19 );
not ( n655 , n654 );
nand ( n656 , n655 , n1 , n572 );
and ( n657 , n653 , n656 );
nand ( n658 , n638 , n651 , n657 );
nor ( n659 , n628 , n658 );
not ( n660 , n12 );
not ( n661 , n13 );
nand ( n662 , n661 , n549 );
xnor ( n663 , n660 , n662 );
and ( n664 , n1 , n663 );
not ( n665 , n1 );
and ( n666 , n665 , n12 );
or ( n667 , n664 , n666 );
not ( n668 , n548 );
nand ( n669 , n668 , n487 , n488 );
not ( n670 , n669 );
nor ( n671 , n14 , n16 );
nand ( n672 , n670 , n671 );
not ( n673 , n17 );
and ( n674 , n672 , n673 );
not ( n675 , n672 );
and ( n676 , n675 , n17 );
nor ( n677 , n674 , n676 );
and ( n678 , n1 , n677 );
not ( n679 , n1 );
and ( n680 , n679 , n673 );
nor ( n681 , n678 , n680 );
nor ( n682 , n667 , n681 );
not ( n683 , n1 );
and ( n684 , n683 , n16 );
not ( n685 , n683 );
not ( n686 , n489 );
nand ( n687 , n686 , n490 );
not ( n688 , n16 );
and ( n689 , n687 , n688 );
not ( n690 , n687 );
and ( n691 , n690 , n16 );
nor ( n692 , n689 , n691 );
not ( n693 , n692 );
and ( n694 , n685 , n693 );
nor ( n695 , n684 , n694 );
not ( n696 , n669 );
nand ( n697 , n696 , n673 , n671 );
not ( n698 , n15 );
and ( n699 , n697 , n698 );
not ( n700 , n697 );
and ( n701 , n700 , n15 );
nor ( n702 , n699 , n701 );
not ( n703 , n702 );
and ( n704 , n1 , n703 );
not ( n705 , n1 );
and ( n706 , n705 , n15 );
nor ( n707 , n704 , n706 );
and ( n708 , n659 , n682 , n695 , n707 );
not ( n709 , n708 );
or ( n710 , n613 , n709 );
nand ( n711 , n710 , n416 );
not ( n712 , n711 );
nor ( n713 , n475 , n712 );
xor ( n714 , n384 , n713 );
not ( n715 , n714 );
not ( n716 , n473 );
not ( n717 , n716 );
not ( n718 , n717 );
not ( n719 , n431 );
not ( n720 , n719 );
not ( n721 , n459 );
nand ( n722 , n721 , n712 );
nor ( n723 , n720 , n722 );
not ( n724 , n723 );
and ( n725 , n718 , n724 );
and ( n726 , n717 , n723 );
nor ( n727 , n725 , n726 );
not ( n728 , n727 );
not ( n729 , n716 );
not ( n730 , n729 );
nand ( n731 , n730 , n723 );
and ( n732 , n731 , n442 );
not ( n733 , n731 );
not ( n734 , n442 );
and ( n735 , n733 , n734 );
nor ( n736 , n732 , n735 );
nand ( n737 , n728 , n736 );
not ( n738 , n737 );
not ( n739 , n738 );
not ( n740 , n739 );
not ( n741 , n740 );
nor ( n742 , n715 , n741 );
nor ( n743 , n736 , n727 , n715 );
or ( n744 , n742 , n743 );
not ( n745 , n744 );
nand ( n746 , n532 , n702 );
not ( n747 , n746 );
nor ( n748 , n597 , n663 );
nand ( n749 , n747 , n458 , n748 );
not ( n750 , n6 );
nand ( n751 , n750 , n428 );
nor ( n752 , n751 , n380 );
nand ( n753 , n410 , n453 );
not ( n754 , n753 );
not ( n755 , n754 );
not ( n756 , n22 );
and ( n757 , n755 , n756 );
not ( n758 , n411 );
and ( n759 , n758 , n22 );
nor ( n760 , n757 , n759 );
nand ( n761 , n633 , n607 , n760 );
not ( n762 , n761 );
not ( n763 , n753 );
not ( n764 , n22 );
nand ( n765 , n763 , n764 );
not ( n766 , n21 );
and ( n767 , n765 , n766 );
not ( n768 , n765 );
and ( n769 , n768 , n21 );
nor ( n770 , n767 , n769 );
nand ( n771 , n752 , n762 , n470 , n770 );
nor ( n772 , n749 , n771 );
not ( n773 , n772 );
nor ( n774 , n505 , n650 );
nand ( n775 , n677 , n774 , n656 );
not ( n776 , n775 );
nor ( n777 , n566 , n584 );
nand ( n778 , n776 , n777 , n692 , n439 );
not ( n779 , n1 );
and ( n780 , n779 , n387 );
not ( n781 , n779 );
nand ( n782 , n453 , n392 , n410 );
and ( n783 , n782 , n387 );
not ( n784 , n782 );
and ( n785 , n784 , n26 );
nor ( n786 , n783 , n785 );
and ( n787 , n781 , n786 );
nor ( n788 , n780 , n787 );
not ( n789 , n788 );
not ( n790 , n24 );
nor ( n791 , n21 , n22 );
not ( n792 , n23 );
nand ( n793 , n791 , n792 , n410 );
not ( n794 , n464 );
nor ( n795 , n793 , n794 );
not ( n796 , n795 );
not ( n797 , n796 );
or ( n798 , n790 , n797 );
nand ( n799 , n791 , n792 , n410 );
not ( n800 , n799 );
not ( n801 , n24 );
and ( n802 , n800 , n801 , n464 );
not ( n803 , n1 );
nor ( n804 , n802 , n803 );
nand ( n805 , n798 , n804 );
nor ( n806 , n525 , n626 );
nor ( n807 , n636 , n554 );
nand ( n808 , n422 , n791 , n410 );
and ( n809 , n808 , n792 );
not ( n810 , n808 );
not ( n811 , n792 );
and ( n812 , n810 , n811 );
nor ( n813 , n809 , n812 );
nand ( n814 , n807 , n494 , n813 );
not ( n815 , n814 );
nand ( n816 , n789 , n805 , n806 , n815 );
nor ( n817 , n778 , n816 );
not ( n818 , n817 );
or ( n819 , n773 , n818 );
nand ( n820 , n819 , n415 );
not ( n821 , n25 );
not ( n822 , n1 );
not ( n823 , n822 );
or ( n824 , n821 , n823 );
not ( n825 , n412 );
nor ( n826 , n825 , n25 , n26 , n393 );
not ( n827 , n826 );
nand ( n828 , n387 , n394 , n412 );
nand ( n829 , n25 , n828 );
nand ( n830 , n827 , n829 , n1 );
nand ( n831 , n824 , n830 );
not ( n832 , n831 );
and ( n833 , n820 , n832 );
not ( n834 , n820 );
not ( n835 , n832 );
and ( n836 , n834 , n835 );
nor ( n837 , n833 , n836 );
not ( n838 , n831 );
not ( n839 , n838 );
nand ( n840 , n772 , n817 );
nand ( n841 , n839 , n840 , n415 );
not ( n842 , n841 );
not ( n843 , n27 );
not ( n844 , n1 );
not ( n845 , n844 );
or ( n846 , n843 , n845 );
not ( n847 , n27 );
nor ( n848 , n847 , n826 );
not ( n849 , n848 );
not ( n850 , n27 );
nand ( n851 , n850 , n413 );
nand ( n852 , n849 , n1 , n851 );
nand ( n853 , n846 , n852 );
and ( n854 , n842 , n853 );
not ( n855 , n842 );
not ( n856 , n853 );
and ( n857 , n855 , n856 );
nor ( n858 , n854 , n857 );
nand ( n859 , n837 , n858 );
not ( n860 , n859 );
not ( n861 , n860 );
not ( n862 , n861 );
nand ( n863 , n47 , n862 );
not ( n864 , n841 );
not ( n865 , n856 );
or ( n866 , n864 , n865 );
or ( n867 , n856 , n841 );
nand ( n868 , n866 , n867 );
nand ( n869 , n868 , n837 );
buf ( n870 , n869 );
not ( n871 , n870 );
nand ( n872 , n46 , n871 );
not ( n873 , n837 );
nand ( n874 , n873 , n868 );
buf ( n875 , n874 );
not ( n876 , n875 );
nand ( n877 , n45 , n876 );
nand ( n878 , n873 , n858 );
buf ( n879 , n878 );
not ( n880 , n879 );
nand ( n881 , n48 , n880 );
nand ( n882 , n863 , n872 , n877 , n881 );
buf ( n883 , n859 );
not ( n884 , n883 );
nand ( n885 , n884 , n51 );
not ( n886 , n870 );
nand ( n887 , n886 , n50 );
not ( n888 , n875 );
nand ( n889 , n888 , n52 );
not ( n890 , n878 );
not ( n891 , n890 );
not ( n892 , n891 );
nand ( n893 , n892 , n49 );
nand ( n894 , n885 , n887 , n889 , n893 );
nand ( n895 , n882 , n894 );
not ( n896 , n41 );
nand ( n897 , n868 , n837 );
not ( n898 , n897 );
not ( n899 , n898 );
or ( n900 , n896 , n899 );
nand ( n901 , n873 , n868 );
not ( n902 , n901 );
nand ( n903 , n44 , n902 );
nand ( n904 , n900 , n903 );
not ( n905 , n42 );
not ( n906 , n890 );
or ( n907 , n905 , n906 );
nand ( n908 , n837 , n858 );
not ( n909 , n908 );
nand ( n910 , n43 , n909 );
nand ( n911 , n907 , n910 );
nor ( n912 , n904 , n911 );
not ( n913 , n34 );
not ( n914 , n869 );
not ( n915 , n914 );
or ( n916 , n913 , n915 );
nand ( n917 , n35 , n860 );
nand ( n918 , n916 , n917 );
not ( n919 , n36 );
not ( n920 , n901 );
not ( n921 , n920 );
or ( n922 , n919 , n921 );
not ( n923 , n837 );
nand ( n924 , n923 , n858 );
not ( n925 , n924 );
nand ( n926 , n33 , n925 );
nand ( n927 , n922 , n926 );
nor ( n928 , n918 , n927 );
nor ( n929 , n912 , n928 );
not ( n930 , n883 );
not ( n931 , n930 );
not ( n932 , n931 );
not ( n933 , n861 );
nand ( n934 , n39 , n933 );
not ( n935 , n38 );
buf ( n936 , n869 );
nor ( n937 , n935 , n936 );
not ( n938 , n937 );
not ( n939 , n40 );
nor ( n940 , n939 , n875 );
not ( n941 , n940 );
not ( n942 , n37 );
nor ( n943 , n942 , n879 );
not ( n944 , n943 );
nand ( n945 , n934 , n938 , n941 , n944 );
nand ( n946 , n929 , n932 , n945 );
nor ( n947 , n895 , n946 );
not ( n948 , n947 );
not ( n949 , n948 );
not ( n950 , n949 );
nand ( n951 , n57 , n880 );
not ( n952 , n860 );
not ( n953 , n952 );
nand ( n954 , n59 , n953 );
nand ( n955 , n60 , n876 );
not ( n956 , n936 );
nand ( n957 , n956 , n58 );
nand ( n958 , n951 , n954 , n955 , n957 );
not ( n959 , n958 );
not ( n960 , n959 );
buf ( n961 , n960 );
and ( n962 , n950 , n961 );
not ( n963 , n950 );
not ( n964 , n961 );
and ( n965 , n963 , n964 );
nor ( n966 , n962 , n965 );
not ( n967 , n533 );
not ( n968 , n967 );
not ( n969 , n1 );
nand ( n970 , n24 , n969 );
and ( n971 , n970 , n805 );
not ( n972 , n789 );
nor ( n973 , n971 , n972 );
not ( n974 , n973 );
not ( n975 , n971 );
not ( n976 , n1 );
and ( n977 , n976 , n21 );
not ( n978 , n976 );
not ( n979 , n770 );
and ( n980 , n978 , n979 );
nor ( n981 , n977 , n980 );
not ( n982 , n1 );
and ( n983 , n982 , n811 );
not ( n984 , n982 );
not ( n985 , n813 );
and ( n986 , n984 , n985 );
nor ( n987 , n983 , n986 );
nand ( n988 , n981 , n987 );
and ( n989 , n1 , n760 );
not ( n990 , n1 );
and ( n991 , n990 , n764 );
or ( n992 , n989 , n991 );
nand ( n993 , n382 , n992 , n474 );
or ( n994 , n988 , n993 );
nand ( n995 , n994 , n416 );
nand ( n996 , n995 , n711 );
nor ( n997 , n975 , n996 );
not ( n998 , n997 );
not ( n999 , n971 );
nand ( n1000 , n999 , n996 );
nand ( n1001 , n998 , n1000 );
nand ( n1002 , n971 , n972 );
nand ( n1003 , n974 , n1001 , n1002 );
buf ( n1004 , n1003 );
not ( n1005 , n1004 );
not ( n1006 , n1005 );
or ( n1007 , n968 , n1006 );
nand ( n1008 , n164 , n1004 );
nand ( n1009 , n1007 , n1008 );
nor ( n1010 , n966 , n1009 );
not ( n1011 , n1010 );
not ( n1012 , n1004 );
and ( n1013 , n1012 , n599 );
not ( n1014 , n1012 );
not ( n1015 , n163 );
and ( n1016 , n1014 , n1015 );
or ( n1017 , n1013 , n1016 );
not ( n1018 , n1017 );
not ( n1019 , n891 );
nand ( n1020 , n53 , n1019 );
not ( n1021 , n883 );
nand ( n1022 , n55 , n1021 );
not ( n1023 , n875 );
nand ( n1024 , n1023 , n56 );
nand ( n1025 , n54 , n956 );
nand ( n1026 , n1020 , n1022 , n1024 , n1025 );
not ( n1027 , n1026 );
not ( n1028 , n1027 );
nand ( n1029 , n960 , n949 );
not ( n1030 , n1029 );
and ( n1031 , n1028 , n1030 );
not ( n1032 , n1028 );
and ( n1033 , n1032 , n1029 );
or ( n1034 , n1031 , n1033 );
nor ( n1035 , n1018 , n1034 );
not ( n1036 , n1035 );
nand ( n1037 , n1011 , n1036 );
not ( n1038 , n1037 );
buf ( n1039 , n875 );
not ( n1040 , n1039 );
nand ( n1041 , n1040 , n68 );
nand ( n1042 , n67 , n930 );
nand ( n1043 , n66 , n956 );
not ( n1044 , n891 );
nand ( n1045 , n65 , n1044 );
nand ( n1046 , n1041 , n1042 , n1043 , n1045 );
not ( n1047 , n62 );
not ( n1048 , n879 );
not ( n1049 , n1048 );
or ( n1050 , n1047 , n1049 );
not ( n1051 , n883 );
nand ( n1052 , n61 , n1051 );
nand ( n1053 , n1050 , n1052 );
not ( n1054 , n1053 );
not ( n1055 , n63 );
not ( n1056 , n914 );
nor ( n1057 , n1055 , n1056 );
not ( n1058 , n64 );
nor ( n1059 , n1058 , n1039 );
nor ( n1060 , n1057 , n1059 );
nand ( n1061 , n1054 , n1060 );
nand ( n1062 , n1046 , n1061 );
not ( n1063 , n1062 );
nor ( n1064 , n959 , n1027 );
nand ( n1065 , n947 , n1063 , n1064 );
not ( n1066 , n1065 );
buf ( n1067 , n1066 );
not ( n1068 , n72 );
not ( n1069 , n875 );
not ( n1070 , n1069 );
or ( n1071 , n1068 , n1070 );
nand ( n1072 , n70 , n898 );
nand ( n1073 , n1071 , n1072 );
not ( n1074 , n69 );
not ( n1075 , n890 );
or ( n1076 , n1074 , n1075 );
not ( n1077 , n908 );
nand ( n1078 , n1077 , n71 );
nand ( n1079 , n1076 , n1078 );
nor ( n1080 , n1073 , n1079 );
not ( n1081 , n76 );
not ( n1082 , n920 );
or ( n1083 , n1081 , n1082 );
nand ( n1084 , n74 , n898 );
nand ( n1085 , n1083 , n1084 );
not ( n1086 , n73 );
not ( n1087 , n925 );
or ( n1088 , n1086 , n1087 );
not ( n1089 , n908 );
nand ( n1090 , n1089 , n75 );
nand ( n1091 , n1088 , n1090 );
nor ( n1092 , n1085 , n1091 );
nor ( n1093 , n1080 , n1092 );
buf ( n1094 , n1093 );
nand ( n1095 , n1067 , n1094 );
not ( n1096 , n1056 );
nand ( n1097 , n82 , n1096 );
nand ( n1098 , n83 , n930 );
nand ( n1099 , n84 , n1023 );
nand ( n1100 , n81 , n1044 );
nand ( n1101 , n1097 , n1098 , n1099 , n1100 );
buf ( n1102 , n1101 );
not ( n1103 , n1102 );
buf ( n1104 , n1103 );
and ( n1105 , n1095 , n1104 );
not ( n1106 , n1095 );
not ( n1107 , n1104 );
and ( n1108 , n1106 , n1107 );
nor ( n1109 , n1105 , n1108 );
not ( n1110 , n1109 );
not ( n1111 , n681 );
not ( n1112 , n1111 );
not ( n1113 , n1112 );
not ( n1114 , n1113 );
buf ( n1115 , n1004 );
not ( n1116 , n1115 );
and ( n1117 , n1114 , n1116 );
not ( n1118 , n1005 );
and ( n1119 , n183 , n1118 );
nor ( n1120 , n1117 , n1119 );
not ( n1121 , n1120 );
not ( n1122 , n1121 );
not ( n1123 , n1122 );
nor ( n1124 , n1110 , n1123 );
not ( n1125 , n707 );
not ( n1126 , n1125 );
not ( n1127 , n1126 );
not ( n1128 , n1127 );
not ( n1129 , n1128 );
buf ( n1130 , n1003 );
not ( n1131 , n1130 );
not ( n1132 , n1131 );
not ( n1133 , n1132 );
not ( n1134 , n1133 );
or ( n1135 , n1129 , n1134 );
not ( n1136 , n182 );
nand ( n1137 , n1136 , n1115 );
nand ( n1138 , n1135 , n1137 );
not ( n1139 , n1138 );
nand ( n1140 , n1101 , n1093 );
not ( n1141 , n1140 );
nand ( n1142 , n1067 , n1141 );
not ( n1143 , n80 );
buf ( n1144 , n876 );
not ( n1145 , n1144 );
or ( n1146 , n1143 , n1145 );
not ( n1147 , n883 );
not ( n1148 , n1147 );
not ( n1149 , n1148 );
nand ( n1150 , n77 , n1149 );
nand ( n1151 , n1146 , n1150 );
not ( n1152 , n1151 );
not ( n1153 , n79 );
buf ( n1154 , n870 );
not ( n1155 , n1154 );
not ( n1156 , n1155 );
or ( n1157 , n1153 , n1156 );
not ( n1158 , n1048 );
not ( n1159 , n1158 );
nand ( n1160 , n78 , n1159 );
nand ( n1161 , n1157 , n1160 );
not ( n1162 , n1161 );
and ( n1163 , n1152 , n1162 );
and ( n1164 , n1142 , n1163 );
not ( n1165 , n1142 );
not ( n1166 , n1163 );
and ( n1167 , n1165 , n1166 );
nor ( n1168 , n1164 , n1167 );
not ( n1169 , n1168 );
nor ( n1170 , n1139 , n1169 );
nor ( n1171 , n1124 , n1170 );
not ( n1172 , n1067 );
nor ( n1173 , n1085 , n1091 );
not ( n1174 , n1173 );
not ( n1175 , n1174 );
not ( n1176 , n1175 );
and ( n1177 , n1172 , n1176 );
not ( n1178 , n1172 );
and ( n1179 , n1178 , n1175 );
nor ( n1180 , n1177 , n1179 );
not ( n1181 , n1180 );
not ( n1182 , n185 );
not ( n1183 , n1182 );
not ( n1184 , n1131 );
not ( n1185 , n1184 );
or ( n1186 , n1183 , n1185 );
or ( n1187 , n500 , n1132 );
nand ( n1188 , n1186 , n1187 );
not ( n1189 , n1188 );
not ( n1190 , n1189 );
nand ( n1191 , n1181 , n1190 );
not ( n1192 , n695 );
not ( n1193 , n1192 );
not ( n1194 , n1193 );
not ( n1195 , n1005 );
not ( n1196 , n1195 );
not ( n1197 , n1196 );
or ( n1198 , n1194 , n1197 );
not ( n1199 , n184 );
nand ( n1200 , n1199 , n1115 );
nand ( n1201 , n1198 , n1200 );
not ( n1202 , n1201 );
nor ( n1203 , n1073 , n1079 );
not ( n1204 , n1203 );
not ( n1205 , n1204 );
not ( n1206 , n1066 );
not ( n1207 , n1206 );
nand ( n1208 , n1207 , n1174 );
xnor ( n1209 , n1205 , n1208 );
nor ( n1210 , n1202 , n1209 );
not ( n1211 , n1210 );
nand ( n1212 , n1171 , n1191 , n1211 );
not ( n1213 , n1212 );
not ( n1214 , n556 );
not ( n1215 , n1214 );
not ( n1216 , n1215 );
buf ( n1217 , n1130 );
not ( n1218 , n1217 );
not ( n1219 , n1218 );
or ( n1220 , n1216 , n1219 );
not ( n1221 , n162 );
not ( n1222 , n1004 );
not ( n1223 , n1222 );
nand ( n1224 , n1221 , n1223 );
nand ( n1225 , n1220 , n1224 );
not ( n1226 , n1225 );
not ( n1227 , n1226 );
not ( n1228 , n1227 );
not ( n1229 , n1228 );
not ( n1230 , n948 );
buf ( n1231 , n1064 );
and ( n1232 , n1230 , n1231 );
not ( n1233 , n1232 );
not ( n1234 , n1053 );
nand ( n1235 , n1060 , n1234 );
not ( n1236 , n1235 );
and ( n1237 , n1233 , n1236 );
not ( n1238 , n1233 );
and ( n1239 , n1238 , n1235 );
nor ( n1240 , n1237 , n1239 );
nand ( n1241 , n1229 , n1240 );
nand ( n1242 , n1232 , n1235 );
not ( n1243 , n1242 );
and ( n1244 , n1041 , n1042 );
and ( n1245 , n1043 , n1045 );
nand ( n1246 , n1244 , n1245 );
not ( n1247 , n1246 );
not ( n1248 , n1247 );
not ( n1249 , n1248 );
and ( n1250 , n1243 , n1249 );
not ( n1251 , n1247 );
and ( n1252 , n1242 , n1251 );
nor ( n1253 , n1250 , n1252 );
not ( n1254 , n1253 );
not ( n1255 , n667 );
not ( n1256 , n1255 );
not ( n1257 , n1256 );
not ( n1258 , n1257 );
not ( n1259 , n1133 );
or ( n1260 , n1258 , n1259 );
not ( n1261 , n186 );
nand ( n1262 , n1261 , n1115 );
nand ( n1263 , n1260 , n1262 );
not ( n1264 , n1263 );
not ( n1265 , n1264 );
nand ( n1266 , n1254 , n1265 );
nand ( n1267 , n1241 , n1266 );
not ( n1268 , n1267 );
not ( n1269 , n525 );
not ( n1270 , n1269 );
or ( n1271 , n1270 , n1217 );
not ( n1272 , n166 );
nand ( n1273 , n1272 , n1132 );
nand ( n1274 , n1271 , n1273 );
not ( n1275 , n1274 );
not ( n1276 , n1275 );
not ( n1277 , n931 );
not ( n1278 , n952 );
not ( n1279 , n39 );
not ( n1280 , n1279 );
and ( n1281 , n1278 , n1280 );
nor ( n1282 , n1281 , n937 );
nor ( n1283 , n943 , n940 );
nand ( n1284 , n1282 , n1283 );
nand ( n1285 , n1277 , n1284 );
not ( n1286 , n1285 );
not ( n1287 , n1286 );
nor ( n1288 , n1287 , n895 );
not ( n1289 , n918 );
not ( n1290 , n927 );
and ( n1291 , n1289 , n1290 );
buf ( n1292 , n1291 );
not ( n1293 , n1292 );
and ( n1294 , n1288 , n1293 );
not ( n1295 , n1288 );
and ( n1296 , n1295 , n1292 );
nor ( n1297 , n1294 , n1296 );
nand ( n1298 , n1276 , n1297 );
not ( n1299 , n627 );
not ( n1300 , n1299 );
not ( n1301 , n1131 );
or ( n1302 , n1300 , n1301 );
not ( n1303 , n1222 );
nand ( n1304 , n165 , n1303 );
nand ( n1305 , n1302 , n1304 );
not ( n1306 , n1305 );
not ( n1307 , n1306 );
not ( n1308 , n1307 );
not ( n1309 , n1291 );
nor ( n1310 , n1285 , n895 );
nand ( n1311 , n1309 , n1310 );
not ( n1312 , n904 );
not ( n1313 , n911 );
and ( n1314 , n1312 , n1313 );
xor ( n1315 , n1311 , n1314 );
nand ( n1316 , n1308 , n1315 );
and ( n1317 , n1298 , n1316 );
not ( n1318 , n637 );
not ( n1319 , n1318 );
or ( n1320 , n1319 , n1217 );
nand ( n1321 , n167 , n1130 );
nand ( n1322 , n1320 , n1321 );
not ( n1323 , n1322 );
not ( n1324 , n1323 );
not ( n1325 , n882 );
not ( n1326 , n1325 );
not ( n1327 , n1285 );
and ( n1328 , n1326 , n1327 );
nand ( n1329 , n887 , n885 , n889 , n893 );
buf ( n1330 , n1329 );
xnor ( n1331 , n1328 , n1330 );
nand ( n1332 , n1324 , n1331 );
not ( n1333 , n633 );
buf ( n1334 , n1333 );
or ( n1335 , n1334 , n1115 );
not ( n1336 , n168 );
not ( n1337 , n1131 );
nand ( n1338 , n1336 , n1337 );
nand ( n1339 , n1335 , n1338 );
not ( n1340 , n1339 );
not ( n1341 , n1340 );
not ( n1342 , n1286 );
not ( n1343 , n1325 );
not ( n1344 , n1343 );
and ( n1345 , n1342 , n1344 );
not ( n1346 , n1342 );
and ( n1347 , n1346 , n1343 );
nor ( n1348 , n1345 , n1347 );
buf ( n1349 , n1348 );
nor ( n1350 , n1341 , n1349 );
not ( n1351 , n1324 );
not ( n1352 , n1331 );
nand ( n1353 , n1351 , n1352 );
nand ( n1354 , n1350 , n1353 );
nand ( n1355 , n1332 , n1354 );
and ( n1356 , n1317 , n1355 );
not ( n1357 , n1307 );
nor ( n1358 , n1357 , n1315 );
not ( n1359 , n1358 );
not ( n1360 , n1359 );
nor ( n1361 , n1356 , n1360 );
not ( n1362 , n1340 );
nand ( n1363 , n1362 , n1348 );
and ( n1364 , n1363 , n1353 );
not ( n1365 , n567 );
not ( n1366 , n973 );
nand ( n1367 , n1366 , n1002 , n1001 );
not ( n1368 , n1367 );
and ( n1369 , n1365 , n1368 );
not ( n1370 , n170 );
and ( n1371 , n1370 , n1003 );
nor ( n1372 , n1369 , n1371 );
not ( n1373 , n154 );
not ( n1374 , n1021 );
or ( n1375 , n1373 , n1374 );
nand ( n1376 , n157 , n871 );
nand ( n1377 , n1375 , n1376 );
not ( n1378 , n155 );
not ( n1379 , n1019 );
or ( n1380 , n1378 , n1379 );
nand ( n1381 , n156 , n876 );
nand ( n1382 , n1380 , n1381 );
nor ( n1383 , n1377 , n1382 );
not ( n1384 , n1383 );
not ( n1385 , n1384 );
nand ( n1386 , n1372 , n1385 );
not ( n1387 , n1386 );
not ( n1388 , n507 );
not ( n1389 , n1388 );
not ( n1390 , n1004 );
and ( n1391 , n1389 , n1390 );
and ( n1392 , n169 , n1130 );
nor ( n1393 , n1391 , n1392 );
not ( n1394 , n1393 );
not ( n1395 , n1394 );
not ( n1396 , n1395 );
not ( n1397 , n1277 );
not ( n1398 , n1397 );
not ( n1399 , n1398 );
not ( n1400 , n1284 );
nand ( n1401 , n1399 , n1400 );
not ( n1402 , n1401 );
nor ( n1403 , n1402 , n1327 );
not ( n1404 , n1403 );
nor ( n1405 , n1396 , n1404 );
not ( n1406 , n1405 );
nand ( n1407 , n1387 , n1406 );
nand ( n1408 , n1396 , n1404 );
not ( n1409 , n1367 );
and ( n1410 , n1409 , n651 );
not ( n1411 , n1409 );
not ( n1412 , n171 );
and ( n1413 , n1411 , n1412 );
nor ( n1414 , n1410 , n1413 );
not ( n1415 , n1414 );
not ( n1416 , n1415 );
not ( n1417 , n150 );
not ( n1418 , n930 );
or ( n1419 , n1417 , n1418 );
nand ( n1420 , n152 , n956 );
nand ( n1421 , n1419 , n1420 );
not ( n1422 , n153 );
not ( n1423 , n1044 );
or ( n1424 , n1422 , n1423 );
nand ( n1425 , n151 , n1023 );
nand ( n1426 , n1424 , n1425 );
nor ( n1427 , n1421 , n1426 );
not ( n1428 , n1427 );
not ( n1429 , n1428 );
nand ( n1430 , n1416 , n1429 );
not ( n1431 , n6 );
and ( n1432 , n1222 , n1431 );
not ( n1433 , n1222 );
not ( n1434 , n172 );
and ( n1435 , n1433 , n1434 );
nor ( n1436 , n1432 , n1435 );
not ( n1437 , n1436 );
not ( n1438 , n146 );
not ( n1439 , n1438 );
not ( n1440 , n931 );
and ( n1441 , n1439 , n1440 );
not ( n1442 , n1144 );
not ( n1443 , n1442 );
and ( n1444 , n149 , n1443 );
nor ( n1445 , n1441 , n1444 );
not ( n1446 , n147 );
not ( n1447 , n1446 );
not ( n1448 , n1159 );
not ( n1449 , n1448 );
and ( n1450 , n1447 , n1449 );
not ( n1451 , n1155 );
not ( n1452 , n1451 );
and ( n1453 , n148 , n1452 );
nor ( n1454 , n1450 , n1453 );
nand ( n1455 , n1445 , n1454 );
nand ( n1456 , n1437 , n1455 );
nand ( n1457 , n1415 , n1428 );
not ( n1458 , n1457 );
not ( n1459 , n1458 );
not ( n1460 , n1459 );
not ( n1461 , n1460 );
nand ( n1462 , n1456 , n1461 );
nand ( n1463 , n1430 , n1462 );
not ( n1464 , n1372 );
not ( n1465 , n1464 );
not ( n1466 , n1384 );
nor ( n1467 , n1465 , n1466 );
not ( n1468 , n1467 );
not ( n1469 , n1468 );
not ( n1470 , n1469 );
nand ( n1471 , n1463 , n1470 , n1406 );
nand ( n1472 , n1407 , n1408 , n1471 );
nand ( n1473 , n1364 , n1472 , n1317 );
nor ( n1474 , n1276 , n1297 );
nand ( n1475 , n1474 , n1316 );
nand ( n1476 , n1361 , n1473 , n1475 );
nand ( n1477 , n1038 , n1213 , n1268 , n1476 );
not ( n1478 , n966 );
not ( n1479 , n1009 );
nor ( n1480 , n1478 , n1479 );
and ( n1481 , n1480 , n1036 );
nand ( n1482 , n1034 , n1018 );
not ( n1483 , n1482 );
nor ( n1484 , n1481 , n1483 );
or ( n1485 , n1267 , n1484 );
nor ( n1486 , n1240 , n1227 );
and ( n1487 , n1486 , n1266 );
not ( n1488 , n1263 );
nand ( n1489 , n1488 , n1253 );
not ( n1490 , n1489 );
nor ( n1491 , n1487 , n1490 );
nand ( n1492 , n1485 , n1491 );
and ( n1493 , n1492 , n1213 );
not ( n1494 , n1189 );
not ( n1495 , n1494 );
nand ( n1496 , n1495 , n1180 );
or ( n1497 , n1496 , n1210 );
nand ( n1498 , n1202 , n1209 );
nand ( n1499 , n1497 , n1498 );
and ( n1500 , n1499 , n1171 );
nor ( n1501 , n1493 , n1500 );
nor ( n1502 , n1122 , n1109 );
not ( n1503 , n1170 );
and ( n1504 , n1502 , n1503 );
nor ( n1505 , n1168 , n1138 );
not ( n1506 , n1505 );
not ( n1507 , n1506 );
nor ( n1508 , n1504 , n1507 );
nand ( n1509 , n1477 , n1501 , n1508 );
not ( n1510 , n1196 );
nand ( n1511 , n193 , n1510 );
not ( n1512 , n1511 );
nand ( n1513 , n115 , n933 );
nand ( n1514 , n112 , n880 );
not ( n1515 , n870 );
nand ( n1516 , n113 , n1515 );
nand ( n1517 , n876 , n114 );
nand ( n1518 , n1513 , n1514 , n1516 , n1517 );
nand ( n1519 , n888 , n108 );
nand ( n1520 , n110 , n871 );
nand ( n1521 , n1147 , n111 );
nand ( n1522 , n1048 , n109 );
nand ( n1523 , n1519 , n1520 , n1521 , n1522 );
nand ( n1524 , n1518 , n1523 );
not ( n1525 , n119 );
not ( n1526 , n1525 );
not ( n1527 , n883 );
and ( n1528 , n1526 , n1527 );
not ( n1529 , n875 );
and ( n1530 , n116 , n1529 );
nor ( n1531 , n1528 , n1530 );
not ( n1532 , n925 );
not ( n1533 , n118 );
nor ( n1534 , n1532 , n1533 );
not ( n1535 , n898 );
not ( n1536 , n117 );
nor ( n1537 , n1535 , n1536 );
nor ( n1538 , n1534 , n1537 );
nand ( n1539 , n1531 , n1538 );
not ( n1540 , n122 );
nor ( n1541 , n1540 , n870 );
not ( n1542 , n120 );
not ( n1543 , n920 );
nor ( n1544 , n1542 , n1543 );
nor ( n1545 , n1541 , n1544 );
not ( n1546 , n924 );
not ( n1547 , n1546 );
not ( n1548 , n121 );
nor ( n1549 , n1547 , n1548 );
not ( n1550 , n909 );
not ( n1551 , n123 );
nor ( n1552 , n1550 , n1551 );
nor ( n1553 , n1549 , n1552 );
nand ( n1554 , n1545 , n1553 );
nand ( n1555 , n1539 , n1554 );
nor ( n1556 , n1524 , n1555 );
not ( n1557 , n135 );
not ( n1558 , n876 );
or ( n1559 , n1557 , n1558 );
nand ( n1560 , n132 , n1048 );
nand ( n1561 , n1559 , n1560 );
not ( n1562 , n133 );
not ( n1563 , n871 );
or ( n1564 , n1562 , n1563 );
nand ( n1565 , n134 , n1147 );
nand ( n1566 , n1564 , n1565 );
nor ( n1567 , n1561 , n1566 );
not ( n1568 , n131 );
not ( n1569 , n1023 );
or ( n1570 , n1568 , n1569 );
nand ( n1571 , n128 , n1021 );
nand ( n1572 , n1570 , n1571 );
not ( n1573 , n129 );
not ( n1574 , n956 );
or ( n1575 , n1573 , n1574 );
nand ( n1576 , n130 , n1019 );
nand ( n1577 , n1575 , n1576 );
nor ( n1578 , n1572 , n1577 );
nor ( n1579 , n1567 , n1578 );
nand ( n1580 , n1556 , n1579 );
not ( n1581 , n1580 );
not ( n1582 , n105 );
not ( n1583 , n956 );
or ( n1584 , n1582 , n1583 );
nand ( n1585 , n107 , n1023 );
nand ( n1586 , n1584 , n1585 );
not ( n1587 , n106 );
not ( n1588 , n1044 );
or ( n1589 , n1587 , n1588 );
nand ( n1590 , n104 , n953 );
nand ( n1591 , n1589 , n1590 );
nor ( n1592 , n1586 , n1591 );
not ( n1593 , n101 );
not ( n1594 , n1096 );
or ( n1595 , n1593 , n1594 );
not ( n1596 , n1039 );
nand ( n1597 , n102 , n1596 );
nand ( n1598 , n1595 , n1597 );
not ( n1599 , n100 );
not ( n1600 , n1044 );
or ( n1601 , n1599 , n1600 );
nand ( n1602 , n103 , n930 );
nand ( n1603 , n1601 , n1602 );
nor ( n1604 , n1598 , n1603 );
nor ( n1605 , n1592 , n1604 );
nand ( n1606 , n1581 , n1605 );
nor ( n1607 , n1062 , n1140 );
nor ( n1608 , n1151 , n1161 );
nor ( n1609 , n1608 , n1325 );
nand ( n1610 , n929 , n932 , n1284 );
nand ( n1611 , n1329 , n1026 , n958 );
nor ( n1612 , n1610 , n1611 );
nand ( n1613 , n1607 , n1609 , n1612 );
nor ( n1614 , n1606 , n1613 );
not ( n1615 , n1614 );
not ( n1616 , n1615 );
not ( n1617 , n141 );
not ( n1618 , n1144 );
or ( n1619 , n1617 , n1618 );
not ( n1620 , n1148 );
nand ( n1621 , n142 , n1620 );
nand ( n1622 , n1619 , n1621 );
not ( n1623 , n139 );
not ( n1624 , n1155 );
or ( n1625 , n1623 , n1624 );
not ( n1626 , n1158 );
nand ( n1627 , n140 , n1626 );
nand ( n1628 , n1625 , n1627 );
nor ( n1629 , n1622 , n1628 );
buf ( n1630 , n1629 );
not ( n1631 , n1630 );
not ( n1632 , n1631 );
xor ( n1633 , n1616 , n1632 );
not ( n1634 , n1633 );
not ( n1635 , n1634 );
or ( n1636 , n1512 , n1635 );
not ( n1637 , n1222 );
nand ( n1638 , n194 , n1637 );
not ( n1639 , n1638 );
not ( n1640 , n1639 );
nand ( n1641 , n126 , n1144 );
nand ( n1642 , n125 , n1155 );
nand ( n1643 , n127 , n1149 );
nand ( n1644 , n124 , n1626 );
nand ( n1645 , n1641 , n1642 , n1643 , n1644 );
buf ( n1646 , n1645 );
nand ( n1647 , n1631 , n1616 );
xor ( n1648 , n1646 , n1647 );
not ( n1649 , n1648 );
nand ( n1650 , n1640 , n1649 );
nand ( n1651 , n1636 , n1650 );
not ( n1652 , n1651 );
not ( n1653 , n85 );
not ( n1654 , n1096 );
or ( n1655 , n1653 , n1654 );
nand ( n1656 , n88 , n1596 );
nand ( n1657 , n1655 , n1656 );
not ( n1658 , n87 );
not ( n1659 , n930 );
or ( n1660 , n1658 , n1659 );
nand ( n1661 , n86 , n1044 );
nand ( n1662 , n1660 , n1661 );
nor ( n1663 , n1657 , n1662 );
not ( n1664 , n1663 );
not ( n1665 , n1664 );
not ( n1666 , n1665 );
not ( n1667 , n1645 );
nor ( n1668 , n1667 , n1629 );
buf ( n1669 , n1668 );
nand ( n1670 , n1666 , n1616 , n1669 );
not ( n1671 , n90 );
not ( n1672 , n1096 );
or ( n1673 , n1671 , n1672 );
nand ( n1674 , n91 , n1023 );
nand ( n1675 , n1673 , n1674 );
not ( n1676 , n89 );
not ( n1677 , n1044 );
or ( n1678 , n1676 , n1677 );
nand ( n1679 , n92 , n953 );
nand ( n1680 , n1678 , n1679 );
nor ( n1681 , n1675 , n1680 );
not ( n1682 , n1681 );
not ( n1683 , n1682 );
and ( n1684 , n1670 , n1683 );
not ( n1685 , n1670 );
not ( n1686 , n1683 );
and ( n1687 , n1685 , n1686 );
nor ( n1688 , n1684 , n1687 );
not ( n1689 , n1688 );
buf ( n1690 , n1337 );
nand ( n1691 , n191 , n1690 );
not ( n1692 , n1691 );
nor ( n1693 , n1689 , n1692 );
nand ( n1694 , n192 , n1303 );
not ( n1695 , n1694 );
not ( n1696 , n1606 );
and ( n1697 , n1609 , n1607 , n1612 );
buf ( n1698 , n1697 );
nand ( n1699 , n1696 , n1698 , n1669 );
and ( n1700 , n1699 , n1665 );
not ( n1701 , n1699 );
not ( n1702 , n1665 );
and ( n1703 , n1701 , n1702 );
nor ( n1704 , n1700 , n1703 );
not ( n1705 , n1704 );
nor ( n1706 , n1695 , n1705 );
nor ( n1707 , n1693 , n1706 );
nand ( n1708 , n1652 , n1707 );
not ( n1709 , n94 );
not ( n1710 , n956 );
or ( n1711 , n1709 , n1710 );
nand ( n1712 , n96 , n1040 );
nand ( n1713 , n1711 , n1712 );
not ( n1714 , n95 );
not ( n1715 , n1021 );
or ( n1716 , n1714 , n1715 );
nand ( n1717 , n93 , n1044 );
nand ( n1718 , n1716 , n1717 );
nor ( n1719 , n1713 , n1718 );
not ( n1720 , n1719 );
not ( n1721 , n1720 );
not ( n1722 , n1721 );
nor ( n1723 , n1663 , n1681 );
nand ( n1724 , n1668 , n1723 );
nor ( n1725 , n1615 , n1724 );
nand ( n1726 , n1722 , n1725 );
not ( n1727 , n98 );
nor ( n1728 , n1727 , n1154 );
not ( n1729 , n97 );
not ( n1730 , n876 );
or ( n1731 , n1729 , n1730 );
nand ( n1732 , n99 , n1048 );
nand ( n1733 , n1731 , n1732 );
nor ( n1734 , n1728 , n1733 );
not ( n1735 , n1734 );
xor ( n1736 , n1726 , n1735 );
not ( n1737 , n1736 );
nand ( n1738 , n187 , n1303 );
buf ( n1739 , n1738 );
buf ( n1740 , n1739 );
buf ( n1741 , n1740 );
nand ( n1742 , n1737 , n1741 );
nand ( n1743 , n188 , n1118 );
not ( n1744 , n1743 );
not ( n1745 , n1744 );
not ( n1746 , n1725 );
not ( n1747 , n1722 );
xnor ( n1748 , n1746 , n1747 );
not ( n1749 , n1748 );
nand ( n1750 , n1745 , n1749 );
nand ( n1751 , n189 , n1637 );
not ( n1752 , n1751 );
not ( n1753 , n1724 );
nor ( n1754 , n1734 , n1719 );
nand ( n1755 , n1753 , n1614 , n1754 );
not ( n1756 , n1448 );
nand ( n1757 , n137 , n1756 );
not ( n1758 , n1451 );
nand ( n1759 , n136 , n1758 );
not ( n1760 , n1442 );
nand ( n1761 , n1760 , n138 );
nand ( n1762 , n1757 , n1759 , n1761 );
buf ( n1763 , n1762 );
not ( n1764 , n1763 );
and ( n1765 , n1755 , n1764 );
not ( n1766 , n1755 );
and ( n1767 , n1766 , n1763 );
nor ( n1768 , n1765 , n1767 );
not ( n1769 , n1768 );
nor ( n1770 , n1752 , n1769 );
nand ( n1771 , n190 , n1223 );
not ( n1772 , n1613 );
nor ( n1773 , n1572 , n1577 );
not ( n1774 , n1773 );
not ( n1775 , n1524 );
nand ( n1776 , n1762 , n1774 , n1645 , n1775 );
nor ( n1777 , n1622 , n1628 );
not ( n1778 , n1555 );
not ( n1779 , n1778 );
nor ( n1780 , n1777 , n1779 );
nand ( n1781 , n1780 , n1754 , n1723 , n1605 );
nor ( n1782 , n1776 , n1781 );
not ( n1783 , n1567 );
nand ( n1784 , n1772 , n1782 , n1783 );
nand ( n1785 , n145 , n1756 );
nand ( n1786 , n143 , n1452 );
nand ( n1787 , n144 , n1443 );
nand ( n1788 , n1785 , n1786 , n1787 );
and ( n1789 , n1784 , n1788 );
not ( n1790 , n1784 );
not ( n1791 , n1788 );
and ( n1792 , n1790 , n1791 );
nor ( n1793 , n1789 , n1792 );
not ( n1794 , n1793 );
nor ( n1795 , n1771 , n1794 );
nor ( n1796 , n1770 , n1795 );
nand ( n1797 , n1742 , n1750 , n1796 );
nor ( n1798 , n1708 , n1797 );
not ( n1799 , n1580 );
nand ( n1800 , n1697 , n1799 );
not ( n1801 , n1592 );
not ( n1802 , n1801 );
buf ( n1803 , n1802 );
xor ( n1804 , n1800 , n1803 );
not ( n1805 , n1804 );
nand ( n1806 , n196 , n1115 );
not ( n1807 , n1806 );
nor ( n1808 , n1805 , n1807 );
not ( n1809 , n1808 );
nand ( n1810 , n195 , n1301 );
not ( n1811 , n1800 );
nand ( n1812 , n1811 , n1801 );
not ( n1813 , n1604 );
not ( n1814 , n1813 );
and ( n1815 , n1812 , n1814 );
not ( n1816 , n1812 );
not ( n1817 , n1814 );
and ( n1818 , n1816 , n1817 );
nor ( n1819 , n1815 , n1818 );
nand ( n1820 , n1810 , n1819 );
nand ( n1821 , n1809 , n1820 );
nand ( n1822 , n198 , n1118 );
not ( n1823 , n1556 );
not ( n1824 , n1823 );
nand ( n1825 , n1698 , n1824 );
not ( n1826 , n1774 );
not ( n1827 , n1826 );
buf ( n1828 , n1827 );
not ( n1829 , n1828 );
and ( n1830 , n1825 , n1829 );
not ( n1831 , n1825 );
and ( n1832 , n1831 , n1828 );
nor ( n1833 , n1830 , n1832 );
nand ( n1834 , n1822 , n1833 );
not ( n1835 , n1823 );
not ( n1836 , n1826 );
nand ( n1837 , n1835 , n1836 );
not ( n1838 , n1837 );
nand ( n1839 , n1838 , n1698 );
not ( n1840 , n1783 );
not ( n1841 , n1840 );
and ( n1842 , n1839 , n1841 );
not ( n1843 , n1839 );
not ( n1844 , n1841 );
and ( n1845 , n1843 , n1844 );
nor ( n1846 , n1842 , n1845 );
not ( n1847 , n1846 );
not ( n1848 , n1218 );
nand ( n1849 , n197 , n1848 );
nand ( n1850 , n1847 , n1849 );
nand ( n1851 , n1834 , n1850 );
nor ( n1852 , n1821 , n1851 );
not ( n1853 , n1852 );
not ( n1854 , n1778 );
not ( n1855 , n1854 );
nand ( n1856 , n1698 , n1855 );
not ( n1857 , n1518 );
not ( n1858 , n1857 );
and ( n1859 , n1856 , n1858 );
not ( n1860 , n1856 );
not ( n1861 , n1858 );
and ( n1862 , n1860 , n1861 );
nor ( n1863 , n1859 , n1862 );
not ( n1864 , n1863 );
not ( n1865 , n610 );
not ( n1866 , n1865 );
or ( n1867 , n1866 , n1690 );
nand ( n1868 , n201 , n1223 );
nand ( n1869 , n1867 , n1868 );
not ( n1870 , n1869 );
nand ( n1871 , n1864 , n1870 );
nor ( n1872 , n1857 , n1854 );
nand ( n1873 , n1698 , n1872 );
and ( n1874 , n1520 , n1519 );
and ( n1875 , n1521 , n1522 );
nand ( n1876 , n1874 , n1875 );
and ( n1877 , n1873 , n1876 );
not ( n1878 , n1873 );
not ( n1879 , n1876 );
and ( n1880 , n1878 , n1879 );
nor ( n1881 , n1877 , n1880 );
not ( n1882 , n1881 );
not ( n1883 , n721 );
not ( n1884 , n1883 );
or ( n1885 , n1884 , n1690 );
not ( n1886 , n202 );
nand ( n1887 , n1886 , n1132 );
nand ( n1888 , n1885 , n1887 );
nand ( n1889 , n1882 , n1888 );
and ( n1890 , n1871 , n1889 );
not ( n1891 , n1890 );
nor ( n1892 , n1853 , n1891 );
not ( n1893 , n657 );
not ( n1894 , n1893 );
not ( n1895 , n1894 );
not ( n1896 , n1895 );
or ( n1897 , n1690 , n1896 );
nand ( n1898 , n199 , n1195 );
nand ( n1899 , n1897 , n1898 );
not ( n1900 , n1899 );
not ( n1901 , n1900 );
nand ( n1902 , n1545 , n1553 );
not ( n1903 , n1902 );
not ( n1904 , n1903 );
not ( n1905 , n1698 );
or ( n1906 , n1904 , n1905 );
not ( n1907 , n1903 );
not ( n1908 , n1907 );
or ( n1909 , n1908 , n1698 );
nand ( n1910 , n1906 , n1909 );
not ( n1911 , n1910 );
or ( n1912 , n1901 , n1911 );
nand ( n1913 , n1698 , n1902 );
nand ( n1914 , n1531 , n1538 );
and ( n1915 , n1913 , n1914 );
not ( n1916 , n1913 );
not ( n1917 , n1914 );
and ( n1918 , n1916 , n1917 );
nor ( n1919 , n1915 , n1918 );
not ( n1920 , n1919 );
not ( n1921 , n588 );
not ( n1922 , n1921 );
not ( n1923 , n1922 );
not ( n1924 , n1923 );
not ( n1925 , n1924 );
or ( n1926 , n1925 , n1637 );
nand ( n1927 , n200 , n1217 );
nand ( n1928 , n1926 , n1927 );
not ( n1929 , n1928 );
nand ( n1930 , n1920 , n1929 );
nand ( n1931 , n1912 , n1930 );
not ( n1932 , n1931 );
nand ( n1933 , n1509 , n1798 , n1892 , n1932 );
not ( n1934 , n1511 );
nand ( n1935 , n1934 , n1633 );
nand ( n1936 , n1639 , n1648 );
and ( n1937 , n1935 , n1936 );
not ( n1938 , n1937 );
nand ( n1939 , n1707 , n1650 , n1938 );
nor ( n1940 , n1704 , n1694 );
buf ( n1941 , n1940 );
not ( n1942 , n1693 );
and ( n1943 , n1941 , n1942 );
and ( n1944 , n1692 , n1689 );
nor ( n1945 , n1943 , n1944 );
nand ( n1946 , n1939 , n1945 );
not ( n1947 , n1797 );
nand ( n1948 , n1946 , n1947 );
not ( n1949 , n1793 );
nand ( n1950 , n1949 , n1771 );
nand ( n1951 , n1948 , n1950 );
nand ( n1952 , n1769 , n1752 );
nor ( n1953 , n1795 , n1952 );
nor ( n1954 , n1951 , n1953 );
not ( n1955 , n1833 );
not ( n1956 , n1822 );
nand ( n1957 , n1955 , n1956 );
not ( n1958 , n1957 );
and ( n1959 , n1958 , n1850 );
not ( n1960 , n1846 );
nor ( n1961 , n1960 , n1849 );
not ( n1962 , n1961 );
not ( n1963 , n1962 );
nor ( n1964 , n1959 , n1963 );
or ( n1965 , n1964 , n1821 );
nor ( n1966 , n1810 , n1819 );
not ( n1967 , n1966 );
nand ( n1968 , n1965 , n1967 );
not ( n1969 , n1968 );
not ( n1970 , n1899 );
not ( n1971 , n1910 );
not ( n1972 , n1971 );
or ( n1973 , n1970 , n1972 );
not ( n1974 , n1919 );
nor ( n1975 , n1974 , n1929 );
not ( n1976 , n1975 );
nand ( n1977 , n1973 , n1976 );
nand ( n1978 , n1977 , n1930 , n1890 );
not ( n1979 , n1978 );
nand ( n1980 , n1869 , n1863 );
not ( n1981 , n1980 );
and ( n1982 , n1981 , n1889 );
not ( n1983 , n1888 );
nand ( n1984 , n1983 , n1881 );
not ( n1985 , n1984 );
nor ( n1986 , n1982 , n1985 );
not ( n1987 , n1986 );
or ( n1988 , n1979 , n1987 );
nand ( n1989 , n1988 , n1852 );
nor ( n1990 , n1804 , n1806 );
nand ( n1991 , n1990 , n1820 );
nand ( n1992 , n1969 , n1989 , n1991 );
and ( n1993 , n1992 , n1798 );
not ( n1994 , n1740 );
nand ( n1995 , n1736 , n1994 );
not ( n1996 , n1995 );
not ( n1997 , n1996 );
nand ( n1998 , n1744 , n1748 );
not ( n1999 , n1998 );
nand ( n2000 , n1999 , n1742 );
and ( n2001 , n1997 , n2000 );
not ( n2002 , n1796 );
nor ( n2003 , n2001 , n2002 );
nor ( n2004 , n1993 , n2003 );
nand ( n2005 , n1933 , n1954 , n2004 );
not ( n2006 , n2005 );
not ( n2007 , n2006 );
or ( n2008 , n745 , n2007 );
nand ( n2009 , n158 , n742 );
nand ( n2010 , n2008 , n2009 );
and ( n2011 , n712 , n1883 );
not ( n2012 , n712 );
and ( n2013 , n2012 , n721 );
nor ( n2014 , n2011 , n2013 );
not ( n2015 , n719 );
xor ( n2016 , n722 , n2015 );
nor ( n2017 , n2014 , n2016 );
nand ( n2018 , n161 , n2017 );
not ( n2019 , n2018 );
nand ( n2020 , n2010 , n2019 );
not ( n2021 , n2014 );
nor ( n2022 , n2021 , n2016 );
and ( n2023 , n161 , n2022 );
and ( n2024 , n2023 , n743 );
not ( n2025 , n2024 );
not ( n2026 , n2005 );
or ( n2027 , n2025 , n2026 );
and ( n2028 , n2021 , n161 , n2016 );
and ( n2029 , n736 , n727 , n714 );
not ( n2030 , n2029 );
and ( n2031 , n1738 , n1735 );
not ( n2032 , n1751 );
not ( n2033 , n1763 );
and ( n2034 , n2032 , n2033 );
and ( n2035 , n1751 , n1763 );
nor ( n2036 , n2034 , n2035 );
or ( n2037 , n2031 , n2036 );
nand ( n2038 , n2031 , n2036 );
nand ( n2039 , n1691 , n1682 );
not ( n2040 , n1743 );
not ( n2041 , n2040 );
not ( n2042 , n1721 );
or ( n2043 , n2041 , n2042 );
nand ( n2044 , n1743 , n1720 );
nand ( n2045 , n2043 , n2044 );
xor ( n2046 , n2039 , n2045 );
nand ( n2047 , n2037 , n2038 , n2046 );
nand ( n2048 , n1638 , n1645 );
not ( n2049 , n1695 );
not ( n2050 , n1665 );
or ( n2051 , n2049 , n2050 );
nand ( n2052 , n1694 , n1664 );
nand ( n2053 , n2051 , n2052 );
nand ( n2054 , n2048 , n2053 );
or ( n2055 , n2048 , n2053 );
not ( n2056 , n1202 );
not ( n2057 , n1205 );
or ( n2058 , n2056 , n2057 );
nand ( n2059 , n1201 , n1204 );
nand ( n2060 , n2058 , n2059 );
nand ( n2061 , n1188 , n1174 );
and ( n2062 , n2060 , n2061 );
not ( n2063 , n2060 );
not ( n2064 , n2061 );
and ( n2065 , n2063 , n2064 );
nor ( n2066 , n2062 , n2065 );
nand ( n2067 , n2054 , n2055 , n2066 );
nor ( n2068 , n2047 , n2067 );
not ( n2069 , n1771 );
and ( n2070 , n2069 , n1791 );
and ( n2071 , n1771 , n1788 );
nor ( n2072 , n2070 , n2071 );
or ( n2073 , n2035 , n2072 );
not ( n2074 , n1840 );
nand ( n2075 , n1849 , n2074 );
not ( n2076 , n1807 );
not ( n2077 , n1802 );
or ( n2078 , n2076 , n2077 );
nand ( n2079 , n1806 , n1801 );
nand ( n2080 , n2078 , n2079 );
xor ( n2081 , n2075 , n2080 );
nand ( n2082 , n2035 , n2072 );
nand ( n2083 , n2073 , n2081 , n2082 );
nand ( n2084 , n1888 , n1876 );
or ( n2085 , n1822 , n1827 );
nand ( n2086 , n1822 , n1827 );
nand ( n2087 , n2085 , n2086 );
or ( n2088 , n2084 , n2087 );
not ( n2089 , n1139 );
not ( n2090 , n1163 );
or ( n2091 , n2089 , n2090 );
not ( n2092 , n1163 );
nand ( n2093 , n1138 , n2092 );
nand ( n2094 , n2091 , n2093 );
nand ( n2095 , n1120 , n1102 );
and ( n2096 , n2094 , n2095 );
not ( n2097 , n2094 );
not ( n2098 , n2095 );
and ( n2099 , n2097 , n2098 );
nor ( n2100 , n2096 , n2099 );
nand ( n2101 , n2084 , n2087 );
nand ( n2102 , n2088 , n2100 , n2101 );
nor ( n2103 , n2083 , n2102 );
nor ( n2104 , n1849 , n1783 );
not ( n2105 , n2104 );
nand ( n2106 , n2105 , n2075 );
nand ( n2107 , n2086 , n2106 );
or ( n2108 , n2086 , n2106 );
nand ( n2109 , n1263 , n1246 );
or ( n2110 , n1263 , n1246 );
nand ( n2111 , n2109 , n2110 );
nand ( n2112 , n1225 , n1235 );
and ( n2113 , n2111 , n2112 );
not ( n2114 , n2111 );
not ( n2115 , n2112 );
and ( n2116 , n2114 , n2115 );
nor ( n2117 , n2113 , n2116 );
nand ( n2118 , n2107 , n2108 , n2117 );
not ( n2119 , n1630 );
nand ( n2120 , n1511 , n2119 );
or ( n2121 , n1638 , n1646 );
nand ( n2122 , n2121 , n2048 );
or ( n2123 , n2120 , n2122 );
nand ( n2124 , n2120 , n2122 );
not ( n2125 , n2109 );
not ( n2126 , n2125 );
nor ( n2127 , n1188 , n1174 );
not ( n2128 , n2127 );
nand ( n2129 , n2128 , n2061 );
not ( n2130 , n2129 );
or ( n2131 , n2126 , n2130 );
or ( n2132 , n2125 , n2129 );
nand ( n2133 , n2131 , n2132 );
nand ( n2134 , n2123 , n2124 , n2133 );
nor ( n2135 , n2118 , n2134 );
or ( n2136 , n1810 , n1813 );
nand ( n2137 , n1810 , n1813 );
nand ( n2138 , n2136 , n2137 );
or ( n2139 , n2079 , n2138 );
nand ( n2140 , n2079 , n2138 );
not ( n2141 , n1121 );
not ( n2142 , n1103 );
or ( n2143 , n2141 , n2142 );
nand ( n2144 , n2143 , n2095 );
and ( n2145 , n2144 , n2059 );
not ( n2146 , n2144 );
not ( n2147 , n2059 );
and ( n2148 , n2146 , n2147 );
nor ( n2149 , n2145 , n2148 );
nand ( n2150 , n2139 , n2140 , n2149 );
or ( n2151 , n1869 , n1857 );
or ( n2152 , n1888 , n1876 );
nand ( n2153 , n2152 , n2084 );
or ( n2154 , n2151 , n2153 );
nand ( n2155 , n2151 , n2153 );
nand ( n2156 , n1929 , n1914 );
not ( n2157 , n1869 );
not ( n2158 , n1858 );
not ( n2159 , n2158 );
or ( n2160 , n2157 , n2159 );
nand ( n2161 , n2160 , n2151 );
nand ( n2162 , n2156 , n2161 );
nand ( n2163 , n2154 , n2155 , n2162 );
nor ( n2164 , n2150 , n2163 );
and ( n2165 , n2068 , n2103 , n2135 , n2164 );
nand ( n2166 , n1017 , n1028 );
not ( n2167 , n1226 );
not ( n2168 , n1235 );
not ( n2169 , n2168 );
or ( n2170 , n2167 , n2169 );
nand ( n2171 , n2170 , n2112 );
and ( n2172 , n2166 , n2171 );
or ( n2173 , n2166 , n2171 );
not ( n2174 , n1394 );
not ( n2175 , n2174 );
buf ( n2176 , n1400 );
and ( n2177 , n2176 , n1398 );
not ( n2178 , n2176 );
and ( n2179 , n2178 , n1397 );
nor ( n2180 , n2177 , n2179 );
not ( n2181 , n2180 );
not ( n2182 , n2181 );
and ( n2183 , n2175 , n2182 );
and ( n2184 , n1395 , n2181 );
nor ( n2185 , n2183 , n2184 );
nand ( n2186 , n2173 , n2185 );
nor ( n2187 , n2172 , n2186 );
nand ( n2188 , n1900 , n1902 );
or ( n2189 , n1929 , n1914 );
nand ( n2190 , n2189 , n2156 );
and ( n2191 , n2188 , n2190 );
or ( n2192 , n2156 , n2161 );
or ( n2193 , n2188 , n2190 );
nand ( n2194 , n2192 , n2193 );
nor ( n2195 , n2191 , n2194 );
not ( n2196 , n1344 );
nand ( n2197 , n1339 , n2196 );
not ( n2198 , n1324 );
not ( n2199 , n1330 );
not ( n2200 , n2199 );
or ( n2201 , n2198 , n2200 );
nand ( n2202 , n1323 , n1330 );
nand ( n2203 , n2201 , n2202 );
and ( n2204 , n2197 , n2203 );
nand ( n2205 , n149 , n1443 );
nand ( n2206 , n146 , n1277 );
nand ( n2207 , n148 , n1452 );
nand ( n2208 , n147 , n1756 );
and ( n2209 , n2205 , n2206 , n2207 , n2208 );
nand ( n2210 , n1436 , n2209 );
nand ( n2211 , n1456 , n2210 );
nor ( n2212 , n2204 , n2211 );
buf ( n2213 , n2093 );
not ( n2214 , n1899 );
not ( n2215 , n1903 );
or ( n2216 , n2214 , n2215 );
nand ( n2217 , n2216 , n2188 );
and ( n2218 , n2213 , n2217 );
or ( n2219 , n2217 , n2213 );
or ( n2220 , n2197 , n2203 );
nand ( n2221 , n2219 , n2220 );
nor ( n2222 , n2218 , n2221 );
and ( n2223 , n2187 , n2195 , n2212 , n2222 );
or ( n2224 , n1691 , n1682 );
nand ( n2225 , n2224 , n2039 );
and ( n2226 , n2052 , n2225 );
or ( n2227 , n2052 , n2225 );
not ( n2228 , n1275 );
not ( n2229 , n1292 );
not ( n2230 , n2229 );
not ( n2231 , n2230 );
or ( n2232 , n2228 , n2231 );
not ( n2233 , n1274 );
not ( n2234 , n2233 );
nand ( n2235 , n2234 , n2229 );
nand ( n2236 , n2232 , n2235 );
not ( n2237 , n2202 );
not ( n2238 , n2237 );
and ( n2239 , n2236 , n2238 );
not ( n2240 , n2236 );
and ( n2241 , n2240 , n2237 );
nor ( n2242 , n2239 , n2241 );
nand ( n2243 , n2227 , n2242 );
nor ( n2244 , n2226 , n2243 );
or ( n2245 , n1511 , n1631 );
nand ( n2246 , n2245 , n2120 );
and ( n2247 , n2137 , n2246 );
or ( n2248 , n2137 , n2246 );
not ( n2249 , n1009 );
not ( n2250 , n961 );
not ( n2251 , n2250 );
or ( n2252 , n2249 , n2251 );
nand ( n2253 , n960 , n1479 );
nand ( n2254 , n2252 , n2253 );
not ( n2255 , n1314 );
nand ( n2256 , n1306 , n2255 );
and ( n2257 , n2254 , n2256 );
not ( n2258 , n2254 );
not ( n2259 , n2256 );
and ( n2260 , n2258 , n2259 );
nor ( n2261 , n2257 , n2260 );
nand ( n2262 , n2248 , n2261 );
nor ( n2263 , n2247 , n2262 );
and ( n2264 , n2244 , n2263 );
not ( n2265 , n1340 );
not ( n2266 , n2196 );
not ( n2267 , n2266 );
or ( n2268 , n2265 , n2267 );
nand ( n2269 , n2268 , n2197 );
not ( n2270 , n2253 );
not ( n2271 , n2270 );
not ( n2272 , n1018 );
not ( n2273 , n1028 );
not ( n2274 , n2273 );
or ( n2275 , n2272 , n2274 );
nand ( n2276 , n2275 , n2166 );
not ( n2277 , n2276 );
not ( n2278 , n1314 );
nor ( n2279 , n1306 , n2278 );
not ( n2280 , n2279 );
nand ( n2281 , n2280 , n2256 );
nor ( n2282 , n1414 , n1428 );
not ( n2283 , n2282 );
not ( n2284 , n1427 );
nand ( n2285 , n2284 , n1414 );
nand ( n2286 , n2283 , n2285 );
nor ( n2287 , n1372 , n1384 );
not ( n2288 , n2287 );
not ( n2289 , n1383 );
nand ( n2290 , n2289 , n1372 );
nand ( n2291 , n2288 , n2290 );
nand ( n2292 , n2165 , n2223 , n2264 , t_0 );
not ( n2293 , n2292 );
or ( n2294 , n2030 , n2293 );
nand ( n2295 , n158 , n2029 );
nand ( n2296 , n2294 , n2295 );
nand ( n2297 , n2028 , n2296 );
nand ( n2298 , n2027 , n2297 );
not ( n2299 , n2021 );
nand ( n2300 , n2299 , n161 , n2016 );
not ( n2301 , n2023 );
and ( n2302 , n2300 , n2018 , n2301 );
nor ( n2303 , n2302 , n2295 );
not ( n2304 , n2303 );
not ( n2305 , n736 );
nand ( n2306 , n727 , n2305 );
nor ( n2307 , n715 , n2306 );
nand ( n2308 , n2028 , n2307 , n2292 );
nand ( n2309 , n2304 , n2308 );
nor ( n2310 , n2298 , n2309 );
nand ( n2311 , n2020 , n2310 );
nand ( n2312 , n742 , n2005 );
and ( n2313 , n2009 , n2312 );
nor ( n2314 , n2313 , n2301 );
nor ( n2315 , n2311 , n2314 );
nand ( n2316 , n1980 , n1984 );
nor ( n2317 , n2316 , n1975 );
and ( n2318 , n2317 , n1931 );
or ( n2319 , n1871 , n1985 );
nand ( n2320 , n2319 , n1889 );
nor ( n2321 , n2318 , n2320 );
nor ( n2322 , n1966 , n1990 );
nand ( n2323 , n1962 , n1957 , n2322 );
or ( n2324 , n2321 , n2323 );
nand ( n2325 , n1808 , n1967 );
nand ( n2326 , n2324 , n2325 );
not ( n2327 , n2322 );
or ( n2328 , n1834 , n1961 );
nand ( n2329 , n2328 , n1850 );
not ( n2330 , n2329 );
or ( n2331 , n2327 , n2330 );
nand ( n2332 , n2331 , n1820 );
or ( n2333 , n2326 , n2332 );
nor ( n2334 , n1688 , n1691 );
nor ( n2335 , n2334 , n1940 );
nand ( n2336 , n2335 , n1937 );
and ( n2337 , n1952 , n1950 );
nand ( n2338 , n2337 , n1998 , n1995 );
nor ( n2339 , n2336 , n2338 );
nand ( n2340 , n2333 , n2339 );
nand ( n2341 , n1950 , n1770 );
or ( n2342 , n1996 , n1750 );
nand ( n2343 , n2342 , n1742 );
nand ( n2344 , n2337 , n2343 );
nand ( n2345 , n2340 , n2341 , n2344 );
not ( n2346 , n2345 );
not ( n2347 , n2323 );
and ( n2348 , n2339 , n2347 );
not ( n2349 , n1977 );
not ( n2350 , n1386 );
nand ( n2351 , n2210 , n1430 );
nand ( n2352 , n1459 , n2351 );
not ( n2353 , n2352 );
or ( n2354 , n2350 , n2353 );
nand ( n2355 , n2354 , n1468 );
and ( n2356 , n2355 , n1408 );
nor ( n2357 , n2356 , n1405 );
nor ( n2358 , n1350 , n2357 );
nor ( n2359 , n1474 , n1358 );
nand ( n2360 , n2358 , n1332 , n2359 );
not ( n2361 , n1353 );
not ( n2362 , n1363 );
nand ( n2363 , n2362 , n1332 );
not ( n2364 , n2363 );
or ( n2365 , n2361 , n2364 );
nand ( n2366 , n2365 , n2359 );
not ( n2367 , n1298 );
nand ( n2368 , n2367 , n1359 );
nand ( n2369 , n2360 , n2366 , n1316 , n2368 );
nor ( n2370 , n1502 , n1505 );
and ( n2371 , n2370 , n1496 , n1498 );
not ( n2372 , n1486 );
nand ( n2373 , n2372 , n1489 );
nor ( n2374 , n2373 , n1480 );
not ( n2375 , n1483 );
nand ( n2376 , n2369 , n2371 , n2374 , n2375 );
not ( n2377 , n1498 );
or ( n2378 , n1191 , n2377 );
nand ( n2379 , n2378 , n1211 );
nand ( n2380 , n2379 , n2370 );
and ( n2381 , n1124 , n1506 );
nor ( n2382 , n2381 , n1170 );
and ( n2383 , n1010 , n1482 );
nor ( n2384 , n2383 , n1035 );
or ( n2385 , n2384 , n2373 );
nand ( n2386 , n2385 , n1266 );
nor ( n2387 , n1490 , n1241 );
or ( n2388 , n2386 , n2387 );
nand ( n2389 , n2388 , n2371 );
nand ( n2390 , n2376 , n2380 , n2382 , n2389 );
not ( n2391 , n2316 );
nand ( n2392 , n2348 , n2349 , n2390 , n2391 );
not ( n2393 , n1944 );
and ( n2394 , n1706 , n2393 );
not ( n2395 , n1942 );
nor ( n2396 , n2394 , n2395 );
nand ( n2397 , n1651 , n1936 , n2335 );
nand ( n2398 , n2396 , n2397 );
not ( n2399 , n2338 );
and ( n2400 , n2398 , n2399 );
nor ( n2401 , n2400 , n1795 );
nand ( n2402 , n2346 , n2392 , n2401 );
nand ( n2403 , n2019 , n2402 );
nor ( n2404 , n2301 , n2402 );
nor ( n2405 , n2300 , n2292 );
nor ( n2406 , n2404 , n2405 );
nand ( n2407 , n2403 , n2406 );
nand ( n2408 , n2407 , n2029 );
nand ( n2409 , n2315 , n2408 );
nand ( n2410 , n2407 , n2307 );
not ( n2411 , n2300 );
and ( n2412 , n2411 , n744 );
not ( n2413 , n2009 );
and ( n2414 , n2028 , n2413 );
nor ( n2415 , n2412 , n2414 );
nand ( n2416 , n2410 , n2415 );
nor ( n2417 , n2409 , n2416 );
not ( n2418 , n1752 );
nand ( n2419 , n1793 , n1768 );
buf ( n2420 , n2419 );
not ( n2421 , n2420 );
not ( n2422 , n2421 );
not ( n2423 , n2422 );
not ( n2424 , n1768 );
or ( n2425 , n2423 , n2424 );
not ( n2426 , n1724 );
not ( n2427 , n1173 );
nand ( n2428 , n1066 , n1204 , n2427 );
nor ( n2429 , n2428 , n1103 );
nand ( n2430 , n2429 , n1166 );
not ( n2431 , n1696 );
nor ( n2432 , n2430 , n2431 );
nand ( n2433 , n2426 , n2432 );
not ( n2434 , n1754 );
nor ( n2435 , n2433 , n2434 );
not ( n2436 , n1763 );
not ( n2437 , n2436 );
not ( n2438 , n2437 );
nor ( n2439 , n2435 , n2438 );
not ( n2440 , n2439 );
buf ( n2441 , n2420 );
not ( n2442 , n2441 );
nand ( n2443 , n2438 , n2435 );
nand ( n2444 , n2440 , n2442 , n2443 );
nand ( n2445 , n2425 , n2444 );
not ( n2446 , n2445 );
not ( n2447 , n2446 );
or ( n2448 , n2418 , n2447 );
buf ( n2449 , n2421 );
not ( n2450 , n2449 );
and ( n2451 , n2437 , n1791 );
and ( n2452 , n1788 , n2436 );
nor ( n2453 , n2451 , n2452 );
not ( n2454 , n2453 );
not ( n2455 , n2443 );
or ( n2456 , n2454 , n2455 );
or ( n2457 , n2453 , n2443 );
nand ( n2458 , n2456 , n2457 );
not ( n2459 , n2458 );
or ( n2460 , n2450 , n2459 );
buf ( n2461 , n1794 );
buf ( n2462 , n2461 );
not ( n2463 , n2462 );
nand ( n2464 , n2460 , n2463 );
nand ( n2465 , n2464 , n1771 );
nand ( n2466 , n2448 , n2465 );
not ( n2467 , n2466 );
not ( n2468 , n1745 );
not ( n2469 , n1749 );
not ( n2470 , n2449 );
not ( n2471 , n2470 );
or ( n2472 , n2469 , n2471 );
not ( n2473 , n1747 );
not ( n2474 , n2433 );
nor ( n2475 , n2473 , n2474 );
not ( n2476 , n2475 );
not ( n2477 , n2420 );
not ( n2478 , n2477 );
not ( n2479 , n2478 );
nor ( n2480 , n1747 , n2433 );
not ( n2481 , n2480 );
nand ( n2482 , n2476 , n2479 , n2481 );
nand ( n2483 , n2472 , n2482 );
not ( n2484 , n2483 );
nand ( n2485 , n2468 , n2484 );
buf ( n2486 , n1741 );
not ( n2487 , n2486 );
not ( n2488 , n1734 );
not ( n2489 , n2480 );
and ( n2490 , n2488 , n2489 );
and ( n2491 , n1734 , n2480 );
nor ( n2492 , n2490 , n2491 );
and ( n2493 , n2442 , n2492 );
not ( n2494 , n2442 );
not ( n2495 , n1737 );
and ( n2496 , n2494 , n2495 );
or ( n2497 , n2493 , n2496 );
nand ( n2498 , n2487 , n2497 );
nand ( n2499 , n2467 , n2485 , n2498 );
not ( n2500 , n2499 );
not ( n2501 , n2442 );
buf ( n2502 , n2432 );
nand ( n2503 , n2502 , n1669 );
not ( n2504 , n1702 );
nor ( n2505 , n2503 , n2504 );
xor ( n2506 , n2505 , n1686 );
not ( n2507 , n2506 );
or ( n2508 , n2501 , n2507 );
not ( n2509 , n2477 );
not ( n2510 , n1689 );
nand ( n2511 , n2509 , n2510 );
nand ( n2512 , n2508 , n2511 );
nor ( n2513 , n2512 , n1691 );
not ( n2514 , n1704 );
not ( n2515 , n2420 );
not ( n2516 , n2515 );
buf ( n2517 , n2516 );
not ( n2518 , n2517 );
or ( n2519 , n2514 , n2518 );
not ( n2520 , n2504 );
not ( n2521 , n2503 );
nor ( n2522 , n2520 , n2521 );
not ( n2523 , n2522 );
not ( n2524 , n2420 );
buf ( n2525 , n2524 );
not ( n2526 , n2505 );
nand ( n2527 , n2523 , n2525 , n2526 );
nand ( n2528 , n2519 , n2527 );
nor ( n2529 , n2528 , n1694 );
nor ( n2530 , n2513 , n2529 );
not ( n2531 , n2530 );
not ( n2532 , n2441 );
not ( n2533 , n2532 );
not ( n2534 , n1646 );
buf ( n2535 , n1632 );
not ( n2536 , n2535 );
nand ( n2537 , n2536 , n2502 );
not ( n2538 , n2537 );
or ( n2539 , n2534 , n2538 );
or ( n2540 , n1646 , n2537 );
nand ( n2541 , n2539 , n2540 );
not ( n2542 , n2541 );
or ( n2543 , n2533 , n2542 );
not ( n2544 , n1648 );
nand ( n2545 , n2544 , n2516 );
nand ( n2546 , n2543 , n2545 );
nor ( n2547 , n2546 , n1640 );
nor ( n2548 , n2531 , n2547 );
buf ( n2549 , n1634 );
nand ( n2550 , n2549 , n2509 );
not ( n2551 , n2535 );
nor ( n2552 , n2551 , n2502 );
not ( n2553 , n2552 );
nand ( n2554 , n2553 , n2525 , n2537 );
and ( n2555 , n2550 , n2554 );
nand ( n2556 , n1934 , n2555 );
nand ( n2557 , n2500 , n2548 , n2556 );
not ( n2558 , n2557 );
not ( n2559 , n1971 );
not ( n2560 , n2559 );
not ( n2561 , n2509 );
or ( n2562 , n2560 , n2561 );
not ( n2563 , n1907 );
not ( n2564 , n2430 );
not ( n2565 , n2564 );
nand ( n2566 , n2563 , n2565 );
nor ( n2567 , n2565 , n2563 );
not ( n2568 , n2567 );
nand ( n2569 , n2566 , n2477 , n2568 );
nand ( n2570 , n2562 , n2569 );
or ( n2571 , n1900 , n2570 );
buf ( n2572 , n1864 );
not ( n2573 , n2572 );
not ( n2574 , n2441 );
or ( n2575 , n2573 , n2574 );
not ( n2576 , n2564 );
not ( n2577 , n1855 );
nor ( n2578 , n2576 , n2577 );
xnor ( n2579 , n2578 , n2158 );
nand ( n2580 , n2579 , n2477 );
nand ( n2581 , n2575 , n2580 );
nor ( n2582 , n1870 , n2581 );
not ( n2583 , n2564 );
not ( n2584 , n1872 );
nor ( n2585 , n2583 , n2584 );
xnor ( n2586 , n2585 , n1876 );
or ( n2587 , n2422 , n2586 );
buf ( n2588 , n1882 );
nand ( n2589 , n2441 , n2588 );
nand ( n2590 , n2587 , n2589 );
nor ( n2591 , n1888 , n2590 );
nor ( n2592 , n2582 , n2591 );
not ( n2593 , n1929 );
not ( n2594 , n2567 );
not ( n2595 , n1914 );
not ( n2596 , n2595 );
and ( n2597 , n2594 , n2596 );
and ( n2598 , n2595 , n2567 );
nor ( n2599 , n2597 , n2598 );
or ( n2600 , n2517 , n2599 );
nand ( n2601 , n2516 , n1974 );
nand ( n2602 , n2600 , n2601 );
not ( n2603 , n2602 );
nand ( n2604 , n2593 , n2603 );
and ( n2605 , n2571 , n2592 , n2604 );
not ( n2606 , n2422 );
not ( n2607 , n1828 );
not ( n2608 , n1824 );
nor ( n2609 , n2608 , n2430 );
xor ( n2610 , n2607 , n2609 );
and ( n2611 , n2606 , n2610 );
not ( n2612 , n2606 );
and ( n2613 , n2612 , n1955 );
nor ( n2614 , n2611 , n2613 );
not ( n2615 , n2614 );
nand ( n2616 , n2615 , n1956 );
not ( n2617 , n1803 );
not ( n2618 , n1799 );
nor ( n2619 , n2576 , n2618 );
xnor ( n2620 , n2617 , n2619 );
or ( n2621 , n2620 , n2478 );
not ( n2622 , n1805 );
nand ( n2623 , n2622 , n2441 );
nand ( n2624 , n2621 , n2623 );
nor ( n2625 , n1806 , n2624 );
not ( n2626 , n2524 );
not ( n2627 , n1819 );
and ( n2628 , n2626 , n2627 );
not ( n2629 , n2626 );
nand ( n2630 , n2617 , n2609 , n1579 );
xor ( n2631 , n2630 , n1817 );
and ( n2632 , n2629 , n2631 );
nor ( n2633 , n2628 , n2632 );
nor ( n2634 , n1810 , n2633 );
nor ( n2635 , n2625 , n2634 );
not ( n2636 , n1849 );
not ( n2637 , n2449 );
not ( n2638 , n1846 );
and ( n2639 , n2637 , n2638 );
not ( n2640 , n1844 );
nor ( n2641 , n1837 , n2565 );
not ( n2642 , n2641 );
or ( n2643 , n2640 , n2642 );
or ( n2644 , n2641 , n1844 );
nand ( n2645 , n2643 , n2644 );
and ( n2646 , n2525 , n2645 );
nor ( n2647 , n2639 , n2646 );
nand ( n2648 , n2636 , n2647 );
and ( n2649 , n2616 , n2635 , n2648 );
nand ( n2650 , n2558 , n2605 , n2649 );
not ( n2651 , n1181 );
not ( n2652 , n2509 );
or ( n2653 , n2651 , n2652 );
nand ( n2654 , n1175 , n1172 );
nand ( n2655 , n2654 , n2442 , n1208 );
nand ( n2656 , n2653 , n2655 );
not ( n2657 , n2517 );
not ( n2658 , n1209 );
and ( n2659 , n2657 , n2658 );
not ( n2660 , n1209 );
and ( n2661 , n2470 , n2660 );
nor ( n2662 , n2659 , n2661 );
nand ( n2663 , n1202 , n2662 );
nand ( n2664 , n2656 , n1190 , n2663 );
not ( n2665 , n2664 );
not ( n2666 , n2662 );
nand ( n2667 , n1201 , n2666 );
not ( n2668 , n2667 );
or ( n2669 , n2665 , n2668 );
not ( n2670 , n1123 );
not ( n2671 , n2670 );
nor ( n2672 , n2477 , n1110 );
not ( n2673 , n1107 );
nand ( n2674 , n2673 , n2428 );
not ( n2675 , n2429 );
and ( n2676 , n2674 , n2675 , n2515 );
nor ( n2677 , n2672 , n2676 );
nand ( n2678 , n2671 , n2677 );
nand ( n2679 , n2675 , n1163 );
nand ( n2680 , n2679 , n2515 , n2565 );
not ( n2681 , n2680 );
buf ( n2682 , n1169 );
nor ( n2683 , n2477 , n2682 );
nor ( n2684 , n2681 , n2683 );
nand ( n2685 , n1139 , n2684 );
and ( n2686 , n2678 , n2685 );
nand ( n2687 , n2669 , n2686 );
not ( n2688 , n2677 );
nand ( n2689 , n2688 , n2670 , n2685 );
or ( n2690 , n1190 , n2656 );
nand ( n2691 , n2690 , n2686 , n2663 );
not ( n2692 , n2479 );
not ( n2693 , n1034 );
not ( n2694 , n2693 );
or ( n2695 , n2692 , n2694 );
nand ( n2696 , n2470 , n2693 );
nand ( n2697 , n2695 , n2696 );
nor ( n2698 , n2697 , n1017 );
nor ( n2699 , n2691 , n2698 );
not ( n2700 , n1478 );
not ( n2701 , n2470 );
or ( n2702 , n2700 , n2701 );
not ( n2703 , n961 );
nand ( n2704 , n2703 , n950 );
nand ( n2705 , n2606 , n2704 , n1029 );
nand ( n2706 , n2702 , n2705 );
or ( n2707 , n1479 , n2706 );
not ( n2708 , n1240 );
not ( n2709 , n2708 );
not ( n2710 , n2709 );
not ( n2711 , n2517 );
or ( n2712 , n2710 , n2711 );
not ( n2713 , n2168 );
not ( n2714 , n2713 );
nand ( n2715 , n2714 , n1233 );
nand ( n2716 , n2574 , n1242 , n2715 );
nand ( n2717 , n2712 , n2716 );
nor ( n2718 , n1229 , n2717 );
not ( n2719 , n1264 );
not ( n2720 , n1253 );
not ( n2721 , n2720 );
or ( n2722 , n2479 , n2721 );
not ( n2723 , n1242 );
not ( n2724 , n1251 );
or ( n2725 , n2723 , n2724 );
or ( n2726 , n1242 , n1251 );
nand ( n2727 , n2725 , n2726 );
nand ( n2728 , n2449 , n2727 );
nand ( n2729 , n2722 , n2728 );
nor ( n2730 , n2719 , n2729 );
nor ( n2731 , n2718 , n2730 );
not ( n2732 , n1351 );
not ( n2733 , n2732 );
not ( n2734 , n2733 );
not ( n2735 , n2734 );
not ( n2736 , n2735 );
xor ( n2737 , n1328 , n2199 );
or ( n2738 , n2478 , n2737 );
not ( n2739 , n2421 );
nand ( n2740 , n2739 , n1352 );
nand ( n2741 , n2738 , n2740 );
not ( n2742 , n2741 );
or ( n2743 , n2736 , n2742 );
nand ( n2744 , n2743 , n1363 );
not ( n2745 , n1276 );
not ( n2746 , n2745 );
not ( n2747 , n2746 );
not ( n2748 , n2421 );
nand ( n2749 , n2748 , n1297 );
not ( n2750 , n2420 );
not ( n2751 , n1288 );
nand ( n2752 , n2751 , n2230 );
nand ( n2753 , n2750 , n2752 , n1311 );
nand ( n2754 , n2749 , n2753 );
not ( n2755 , n2754 );
and ( n2756 , n2747 , n2755 );
not ( n2757 , n1308 );
not ( n2758 , n2757 );
buf ( n2759 , n1315 );
nor ( n2760 , n2758 , n2759 );
nor ( n2761 , n2756 , n2760 );
nor ( n2762 , n2735 , n2741 );
not ( n2763 , n2762 );
nand ( n2764 , n2744 , n2761 , n2763 );
nor ( n2765 , n1350 , n2762 );
not ( n2766 , n2357 );
nand ( n2767 , n2765 , n2761 , n2766 );
not ( n2768 , n2760 );
nand ( n2769 , n2754 , n2746 , n2768 );
not ( n2770 , n2758 );
not ( n2771 , n2770 );
nand ( n2772 , n2771 , n2759 );
nand ( n2773 , n2764 , n2767 , n2769 , n2772 );
nand ( n2774 , n2699 , n2707 , n2731 , n2773 );
nand ( n2775 , n2687 , n2689 , n2774 );
not ( n2776 , n2691 );
not ( n2777 , n2776 );
not ( n2778 , n2730 );
not ( n2779 , n1229 );
not ( n2780 , n2779 );
nand ( n2781 , n2778 , n2780 , n2717 );
not ( n2782 , n1017 );
not ( n2783 , n2697 );
or ( n2784 , n2782 , n2783 );
nand ( n2785 , n1479 , n2706 );
nand ( n2786 , n2784 , n2785 );
not ( n2787 , n2698 );
nand ( n2788 , n2786 , n2731 , n2787 );
nand ( n2789 , n2719 , n2729 );
nand ( n2790 , n2781 , n2788 , n2789 );
not ( n2791 , n2790 );
or ( n2792 , n2777 , n2791 );
not ( n2793 , n2684 );
nand ( n2794 , n1138 , n2793 );
nand ( n2795 , n2792 , n2794 );
nor ( n2796 , n2775 , n2795 );
or ( n2797 , n2650 , n2796 );
not ( n2798 , n2591 );
nand ( n2799 , n2581 , n1870 , n2798 );
not ( n2800 , n1929 );
not ( n2801 , n2602 );
or ( n2802 , n2800 , n2801 );
nand ( n2803 , n1900 , n2570 );
nand ( n2804 , n2802 , n2803 );
nand ( n2805 , n2804 , n2592 , n2604 );
nand ( n2806 , n1888 , n2590 );
nand ( n2807 , n2799 , n2805 , n2806 );
nand ( n2808 , n2649 , n2807 );
not ( n2809 , n1849 );
not ( n2810 , n2647 );
not ( n2811 , n2810 );
or ( n2812 , n2809 , n2811 );
nand ( n2813 , n2614 , n1822 , n2648 );
nand ( n2814 , n2812 , n2813 );
and ( n2815 , n2635 , n2814 );
not ( n2816 , n2634 );
not ( n2817 , n2816 );
not ( n2818 , n2624 );
nor ( n2819 , n2817 , n2818 , n1807 );
nor ( n2820 , n2815 , n2819 );
nand ( n2821 , n1810 , n2633 );
nand ( n2822 , n2808 , n2820 , n2821 );
not ( n2823 , n2822 );
nor ( n2824 , n2823 , n2557 );
or ( n2825 , n2547 , n1934 , n2555 );
nand ( n2826 , n1640 , n2546 );
nand ( n2827 , n2825 , n2826 );
and ( n2828 , n2530 , n2827 );
not ( n2829 , n2528 );
nor ( n2830 , n2513 , n1695 , n2829 );
not ( n2831 , n2512 );
nor ( n2832 , n2831 , n1692 );
nor ( n2833 , n2828 , n2830 , n2832 );
or ( n2834 , n2833 , n2499 );
and ( n2835 , n2498 , n1745 , n2483 );
not ( n2836 , n2486 );
nor ( n2837 , n2497 , n2836 );
nor ( n2838 , n2835 , n2837 );
or ( n2839 , n2838 , n2466 );
nand ( n2840 , n2445 , n1751 , n2465 );
nand ( n2841 , n2839 , n2840 );
not ( n2842 , n2841 );
not ( n2843 , n2464 );
nand ( n2844 , n2843 , n2069 );
nand ( n2845 , n2834 , n2842 , n2844 );
nor ( n2846 , n2824 , n2845 );
nand ( n2847 , n2797 , n2846 );
or ( n2848 , n2417 , n2847 );
nand ( n2849 , n2408 , n2410 );
not ( n2850 , n2028 );
not ( n2851 , n744 );
or ( n2852 , n2850 , n2851 );
or ( n2853 , n2300 , n2009 );
nand ( n2854 , n2852 , n2853 );
nor ( n2855 , n2849 , n2854 );
not ( n2856 , n2855 );
not ( n2857 , n2315 );
or ( n2858 , n2856 , n2857 );
nand ( n2859 , n2858 , n2847 );
not ( n2860 , n972 );
and ( n2861 , n1000 , n2860 );
not ( n2862 , n1000 );
and ( n2863 , n2862 , n972 );
or ( n2864 , n2861 , n2863 );
nor ( n2865 , n1001 , n2864 );
not ( n2866 , n2865 );
not ( n2867 , n981 );
not ( n2868 , n417 );
not ( n2869 , n2868 );
not ( n2870 , n383 );
or ( n2871 , n2869 , n2870 );
nand ( n2872 , n2871 , n713 );
not ( n2873 , n2872 );
buf ( n2874 , n992 );
nor ( n2875 , n2873 , n2874 );
nand ( n2876 , n2867 , n2875 );
not ( n2877 , n2876 );
not ( n2878 , n2877 );
not ( n2879 , n2875 );
nand ( n2880 , n981 , n2879 );
nand ( n2881 , n2878 , n2880 );
not ( n2882 , n2881 );
not ( n2883 , n2874 );
not ( n2884 , n2872 );
and ( n2885 , n2883 , n2884 );
and ( n2886 , n2874 , n2872 );
nor ( n2887 , n2885 , n2886 );
not ( n2888 , n2887 );
not ( n2889 , n987 );
not ( n2890 , n2876 );
not ( n2891 , n2890 );
or ( n2892 , n2889 , n2891 );
not ( n2893 , n987 );
nand ( n2894 , n2893 , n2876 );
nand ( n2895 , n2892 , n2894 );
nand ( n2896 , n2882 , n2888 , n2895 );
nand ( n2897 , n161 , n2896 );
not ( n2898 , n2022 );
buf ( n2899 , n741 );
not ( n2900 , n2899 );
not ( n2901 , n2900 );
nor ( n2902 , n2866 , n2897 , n2898 , n2901 );
not ( n2903 , n2902 );
nand ( n2904 , n161 , n714 );
nand ( n2905 , n2903 , n158 , n2904 );
nand ( n2906 , n2848 , n2859 , n2905 );
not ( n2907 , n1341 );
not ( n2908 , n1396 );
not ( n2909 , n1464 );
not ( n2910 , n1416 );
nand ( n2911 , n1437 , n2910 );
nor ( n2912 , n2909 , n2911 );
nand ( n2913 , n2908 , n2912 );
nor ( n2914 , n2907 , n2913 );
and ( n2915 , n1351 , n2914 );
nand ( n2916 , n1276 , n2915 );
nor ( n2917 , n2757 , n2916 );
nand ( n2918 , n1479 , n2917 );
not ( n2919 , n2918 );
nand ( n2920 , n1017 , n2919 );
xnor ( n2921 , n2920 , n2779 );
not ( n2922 , n2921 );
not ( n2923 , n2896 );
not ( n2924 , n2923 );
and ( n2925 , n2023 , n2924 );
not ( n2926 , n2306 );
not ( n2927 , n2895 );
not ( n2928 , n2881 );
not ( n2929 , n158 );
not ( n2930 , n2929 );
not ( n2931 , n2888 );
or ( n2932 , n2930 , n2931 );
nand ( n2933 , n158 , n2887 );
nand ( n2934 , n2932 , n2933 );
not ( n2935 , n2934 );
or ( n2936 , n2928 , n2935 );
not ( n2937 , n160 );
nand ( n2938 , n2936 , n2937 );
not ( n2939 , n2938 );
or ( n2940 , n2927 , n2939 );
not ( n2941 , n2895 );
nand ( n2942 , n2882 , n2941 );
nand ( n2943 , n2940 , n2942 );
not ( n2944 , n2888 );
not ( n2945 , n2929 );
not ( n2946 , n2881 );
or ( n2947 , n2945 , n2946 );
nand ( n2948 , n2947 , n2895 );
not ( n2949 , n2948 );
or ( n2950 , n2944 , n2949 );
not ( n2951 , n2933 );
not ( n2952 , n2951 );
not ( n2953 , n2881 );
or ( n2954 , n2952 , n2953 );
not ( n2955 , n159 );
nand ( n2956 , n2954 , n2955 );
nand ( n2957 , n2895 , n2956 );
nand ( n2958 , n2950 , n2957 );
nand ( n2959 , n2943 , n715 , n2958 );
not ( n2960 , n2959 );
and ( n2961 , n2925 , n2926 , n2960 );
not ( n2962 , n2961 );
not ( n2963 , n2962 );
not ( n2964 , n2963 );
not ( n2965 , n2964 );
and ( n2966 , n2922 , n2965 );
and ( n2967 , n2023 , n2924 );
and ( n2968 , n2967 , n740 , n2960 );
not ( n2969 , n2968 );
not ( n2970 , n2969 );
not ( n2971 , n2864 );
not ( n2972 , n2971 );
not ( n2973 , n2693 );
or ( n2974 , n2972 , n2973 );
not ( n2975 , n1429 );
not ( n2976 , n1466 );
nand ( n2977 , n2975 , n2976 );
not ( n2978 , n2977 );
buf ( n2979 , n1349 );
nand ( n2980 , n2978 , n2979 , n1403 );
not ( n2981 , n2980 );
nand ( n2982 , n1352 , n1297 , n2981 );
not ( n2983 , n2982 );
not ( n2984 , n2461 );
nor ( n2985 , n2209 , n2984 );
not ( n2986 , n2985 );
not ( n2987 , n2986 );
nand ( n2988 , n2983 , n2987 );
not ( n2989 , n1315 );
nor ( n2990 , n2988 , n2989 );
nand ( n2991 , n1478 , n2990 );
nor ( n2992 , n2991 , n1034 );
nand ( n2993 , n2709 , n2992 );
not ( n2994 , n2993 );
not ( n2995 , n2721 );
or ( n2996 , n2994 , n2995 );
not ( n2997 , n2993 );
not ( n2998 , n2721 );
and ( n2999 , n2997 , n2998 );
nor ( n3000 , n2999 , n2971 );
nand ( n3001 , n2996 , n3000 );
nand ( n3002 , n2974 , n3001 );
and ( n3003 , n2970 , n3002 );
nor ( n3004 , n2966 , n3003 );
or ( n3005 , n1306 , n1314 );
not ( n3006 , n3005 );
not ( n3007 , n3006 );
not ( n3008 , n2254 );
nand ( n3009 , n3007 , n3008 );
not ( n3010 , n3009 );
not ( n3011 , n2269 );
not ( n3012 , n1327 );
nor ( n3013 , n1393 , n2180 );
not ( n3014 , n3013 );
nand ( n3015 , n3012 , n3014 );
not ( n3016 , n3015 );
nor ( n3017 , n3011 , n3016 );
not ( n3018 , n3017 );
not ( n3019 , n2203 );
not ( n3020 , n1339 );
nand ( n3021 , n3020 , n2196 );
nand ( n3022 , n3019 , n3021 );
not ( n3023 , n3022 );
or ( n3024 , n3018 , n3023 );
not ( n3025 , n3021 );
nand ( n3026 , n3025 , n2203 );
nand ( n3027 , n3024 , n3026 );
and ( n3028 , n1322 , n1330 );
nor ( n3029 , n3028 , n2236 );
not ( n3030 , n2281 );
nand ( n3031 , n1275 , n2229 );
nand ( n3032 , n3030 , n3031 );
not ( n3033 , n3032 );
nor ( n3034 , n3029 , n3033 );
and ( n3035 , n3027 , n3034 );
nand ( n3036 , n3028 , n2236 );
nor ( n3037 , n3036 , n3033 );
nor ( n3038 , n3035 , n3037 );
nand ( n3039 , n2290 , n2185 );
not ( n3040 , n3039 );
not ( n3041 , n1436 );
nor ( n3042 , n3041 , n2209 );
not ( n3043 , n3042 );
not ( n3044 , n1430 );
nor ( n3045 , n3044 , n1458 );
nor ( n3046 , n3043 , n3045 );
not ( n3047 , n1386 );
nor ( n3048 , n3047 , n1467 );
nand ( n3049 , n2285 , n3048 );
nand ( n3050 , n3046 , n3049 );
not ( n3051 , n2285 );
not ( n3052 , n3048 );
nand ( n3053 , n3051 , n3052 );
nand ( n3054 , n3050 , n3053 );
not ( n3055 , n3054 );
or ( n3056 , n3040 , n3055 );
not ( n3057 , n2290 );
not ( n3058 , n2185 );
nand ( n3059 , n3057 , n3058 );
nand ( n3060 , n3056 , n3059 );
not ( n3061 , n3022 );
nor ( n3062 , n3015 , n2269 );
nor ( n3063 , n3061 , n3062 );
and ( n3064 , n3060 , n3063 );
nand ( n3065 , n3064 , n3034 );
not ( n3066 , n3031 );
nand ( n3067 , n3066 , n2281 );
nand ( n3068 , n3038 , n3065 , n3067 );
not ( n3069 , n3068 );
or ( n3070 , n3010 , n3069 );
nand ( n3071 , n3006 , n2254 );
nand ( n3072 , n3070 , n3071 );
not ( n3073 , n3072 );
nand ( n3074 , n1009 , n961 );
not ( n3075 , n3074 );
not ( n3076 , n3075 );
nand ( n3077 , n3076 , n2277 );
not ( n3078 , n3077 );
or ( n3079 , n3073 , n3078 );
nand ( n3080 , n3075 , n2276 );
nand ( n3081 , n3079 , n3080 );
not ( n3082 , n3081 );
not ( n3083 , n3082 );
not ( n3084 , n2273 );
and ( n3085 , n1018 , n3084 );
not ( n3086 , n3085 );
not ( n3087 , n2171 );
and ( n3088 , n3086 , n3087 );
and ( n3089 , n3085 , n2171 );
nor ( n3090 , n3088 , n3089 );
not ( n3091 , n3090 );
not ( n3092 , n3091 );
or ( n3093 , n3083 , n3092 );
and ( n3094 , n3081 , n3090 );
nand ( n3095 , n2021 , n736 );
nand ( n3096 , n2016 , n2305 );
nand ( n3097 , n3095 , n3096 );
nand ( n3098 , n737 , n2306 );
nor ( n3099 , n3097 , n3098 );
nor ( n3100 , n2897 , n2959 );
nand ( n3101 , n3099 , n3100 );
nor ( n3102 , n3094 , n3101 );
nand ( n3103 , n3093 , n3102 );
not ( n3104 , n2780 );
not ( n3105 , n3096 );
and ( n3106 , n727 , n3105 );
not ( n3107 , n3106 );
not ( n3108 , n3100 );
or ( n3109 , n3107 , n3108 );
nor ( n3110 , n2018 , n2306 );
nand ( n3111 , n3110 , n715 , n2924 );
nand ( n3112 , n3109 , n3111 );
not ( n3113 , n3112 );
not ( n3114 , n3113 );
nand ( n3115 , n3104 , n3114 );
not ( n3116 , n61 );
nor ( n3117 , n3116 , n161 );
not ( n3118 , n3117 );
not ( n3119 , n61 );
not ( n3120 , n43 );
nand ( n3121 , n39 , n47 );
not ( n3122 , n3121 );
and ( n3123 , n51 , n3122 );
nand ( n3124 , n35 , n3123 );
nor ( n3125 , n3120 , n3124 );
nand ( n3126 , n59 , n3125 );
not ( n3127 , n3126 );
nand ( n3128 , n3127 , n55 );
not ( n3129 , n3128 );
or ( n3130 , n3119 , n3129 );
or ( n3131 , n61 , n3128 );
nand ( n3132 , n3130 , n3131 );
not ( n3133 , n3097 );
nor ( n3134 , n3133 , n3098 );
nand ( n3135 , n3134 , n3100 );
nand ( n3136 , n3135 , n3101 );
nor ( n3137 , n3136 , n2968 );
nor ( n3138 , n2961 , n3112 );
nand ( n3139 , n3137 , n161 , n3138 );
not ( n3140 , n3139 );
nand ( n3141 , n3132 , n3140 );
not ( n3142 , n1339 );
not ( n3143 , n2266 );
or ( n3144 , n3142 , n3143 );
nand ( n3145 , n3144 , n3021 );
not ( n3146 , n2174 );
not ( n3147 , n1401 );
or ( n3148 , n3146 , n3147 );
nand ( n3149 , n3148 , n3012 );
nand ( n3150 , n3145 , n3149 );
not ( n3151 , n3150 );
not ( n3152 , n3151 );
xor ( n3153 , n1322 , n1330 );
nand ( n3154 , n2197 , n3153 );
not ( n3155 , n3154 );
or ( n3156 , n3152 , n3155 );
not ( n3157 , n2197 );
not ( n3158 , n3153 );
nand ( n3159 , n3157 , n3158 );
nand ( n3160 , n3156 , n3159 );
nor ( n3161 , n2233 , n1293 );
not ( n3162 , n3161 );
nand ( n3163 , n3162 , n3031 );
nor ( n3164 , n2237 , n3163 );
not ( n3165 , n2235 );
not ( n3166 , n1306 );
not ( n3167 , n2255 );
not ( n3168 , n3167 );
or ( n3169 , n3166 , n3168 );
nand ( n3170 , n3169 , n3005 );
nor ( n3171 , n3165 , n3170 );
nor ( n3172 , n3164 , n3171 );
and ( n3173 , n3160 , n3172 );
nand ( n3174 , n2237 , n3163 );
nor ( n3175 , n3174 , n3171 );
nor ( n3176 , n3173 , n3175 );
not ( n3177 , n3154 );
nor ( n3178 , n3145 , n3149 );
nor ( n3179 , n3177 , n3178 );
nand ( n3180 , n1393 , n2180 );
not ( n3181 , n3180 );
nor ( n3182 , n3181 , n3013 );
nand ( n3183 , n1468 , n3182 );
not ( n3184 , n3183 );
nor ( n3185 , n1436 , n1455 );
not ( n3186 , n3185 );
nand ( n3187 , n1455 , n2286 );
nand ( n3188 , n3186 , n3187 );
not ( n3189 , n3188 );
nor ( n3190 , n1455 , n2286 );
nor ( n3191 , n1458 , n2291 );
nor ( n3192 , n3190 , n3191 );
not ( n3193 , n3192 );
or ( n3194 , n3189 , n3193 );
nand ( n3195 , n1460 , n2291 );
nand ( n3196 , n3194 , n3195 );
not ( n3197 , n3196 );
or ( n3198 , n3184 , n3197 );
not ( n3199 , n3182 );
nand ( n3200 , n1469 , n3199 );
nand ( n3201 , n3198 , n3200 );
nand ( n3202 , n3179 , n3201 );
not ( n3203 , n3202 );
nand ( n3204 , n3203 , n3172 );
nand ( n3205 , n3165 , n3170 );
nand ( n3206 , n3176 , n3204 , n3205 );
not ( n3207 , n1479 );
not ( n3208 , n2703 );
or ( n3209 , n3207 , n3208 );
nand ( n3210 , n3209 , n3074 );
not ( n3211 , n3210 );
nand ( n3212 , n2256 , n3211 );
and ( n3213 , n3206 , n3212 );
and ( n3214 , n2259 , n3210 );
nor ( n3215 , n3213 , n3214 );
buf ( n3216 , n2271 );
xor ( n3217 , n1018 , n3084 );
and ( n3218 , n3216 , n3217 );
or ( n3219 , n3215 , n3218 );
not ( n3220 , n3216 );
not ( n3221 , n3217 );
nand ( n3222 , n3220 , n3221 );
nand ( n3223 , n3219 , n3222 );
not ( n3224 , n3223 );
not ( n3225 , n3224 );
not ( n3226 , n2166 );
and ( n3227 , n1228 , n2713 );
not ( n3228 , n1228 );
and ( n3229 , n3228 , n2714 );
nor ( n3230 , n3227 , n3229 );
not ( n3231 , n3230 );
and ( n3232 , n3226 , n3231 );
and ( n3233 , n2166 , n3230 );
nor ( n3234 , n3232 , n3233 );
not ( n3235 , n3234 );
not ( n3236 , n3235 );
or ( n3237 , n3225 , n3236 );
and ( n3238 , n3223 , n3234 );
not ( n3239 , n3135 );
not ( n3240 , n3239 );
nor ( n3241 , n3238 , n3240 );
nand ( n3242 , n3237 , n3241 );
and ( n3243 , n3118 , n3141 , n3242 );
nand ( n3244 , n3004 , n3103 , n3115 , n3243 );
not ( n3245 , n3072 );
not ( n3246 , n3245 );
nand ( n3247 , n3080 , n3077 );
not ( n3248 , n3247 );
or ( n3249 , n3246 , n3248 );
not ( n3250 , n3247 );
and ( n3251 , n3072 , n3250 );
nor ( n3252 , n3251 , n3101 );
nand ( n3253 , n3249 , n3252 );
not ( n3254 , n3215 );
not ( n3255 , n3222 );
nor ( n3256 , n3255 , n3218 );
not ( n3257 , n3256 );
not ( n3258 , n3257 );
or ( n3259 , n3254 , n3258 );
not ( n3260 , n3215 );
and ( n3261 , n3260 , n3256 );
not ( n3262 , n3239 );
nor ( n3263 , n3261 , n3262 );
nand ( n3264 , n3259 , n3263 );
not ( n3265 , n55 );
not ( n3266 , n3126 );
or ( n3267 , n3265 , n3266 );
or ( n3268 , n55 , n3126 );
nand ( n3269 , n3267 , n3268 );
nand ( n3270 , n3269 , n3140 );
and ( n3271 , n3253 , n3264 , n3270 );
nand ( n3272 , n1018 , n3114 );
not ( n3273 , n55 );
nor ( n3274 , n3273 , n161 );
not ( n3275 , n3274 );
and ( n3276 , n2918 , n1017 );
not ( n3277 , n2918 );
and ( n3278 , n3277 , n1018 );
nor ( n3279 , n3276 , n3278 );
not ( n3280 , n3279 );
not ( n3281 , n2962 );
and ( n3282 , n3280 , n3281 );
not ( n3283 , n2971 );
not ( n3284 , n1478 );
or ( n3285 , n3283 , n3284 );
nor ( n3286 , n2709 , n2992 );
not ( n3287 , n3286 );
nand ( n3288 , n3287 , n2993 , n2864 );
nand ( n3289 , n3285 , n3288 );
and ( n3290 , n3289 , n2970 );
nor ( n3291 , n3282 , n3290 );
nand ( n3292 , n3271 , n3272 , n3275 , n3291 );
and ( n3293 , n3059 , n3039 );
not ( n3294 , n3293 );
not ( n3295 , n3054 );
not ( n3296 , n3295 );
or ( n3297 , n3294 , n3296 );
or ( n3298 , n3293 , n3295 );
nand ( n3299 , n3297 , n3298 );
and ( n3300 , n3099 , n3299 );
and ( n3301 , n2022 , n2926 );
and ( n3302 , n2912 , n2908 );
not ( n3303 , n2912 );
not ( n3304 , n2908 );
and ( n3305 , n3303 , n3304 );
nor ( n3306 , n3302 , n3305 );
and ( n3307 , n3301 , n3306 );
nor ( n3308 , n3300 , n3307 );
not ( n3309 , n3308 );
or ( n3310 , n3096 , n2926 );
nand ( n3311 , n3095 , n3310 );
not ( n3312 , n3183 );
not ( n3313 , n3200 );
nor ( n3314 , n3312 , n3313 );
xor ( n3315 , n3314 , n3196 );
nand ( n3316 , n3311 , n3315 );
nand ( n3317 , n3106 , n3304 );
not ( n3318 , n2971 );
buf ( n3319 , n2976 );
not ( n3320 , n3319 );
or ( n3321 , n3318 , n3320 );
buf ( n3322 , n2979 );
not ( n3323 , n3322 );
not ( n3324 , n3323 );
and ( n3325 , n2975 , n2985 );
nand ( n3326 , n3319 , n3325 );
nor ( n3327 , n3326 , n1404 );
not ( n3328 , n3327 );
not ( n3329 , n3328 );
or ( n3330 , n3324 , n3329 );
and ( n3331 , n3322 , n3327 );
nor ( n3332 , n3331 , n2971 );
nand ( n3333 , n3330 , n3332 );
nand ( n3334 , n3321 , n3333 );
nand ( n3335 , n2900 , n3334 );
nand ( n3336 , n3316 , n3317 , n3335 );
nor ( n3337 , n3309 , n3336 );
nor ( n3338 , n714 , n2897 );
not ( n3339 , n3338 );
and ( n3340 , n3096 , n2898 , n3098 );
or ( n3341 , n3339 , n3340 , n2958 , n2943 );
or ( n3342 , n3337 , n3341 );
not ( n3343 , n3341 );
or ( n3344 , n939 , n3343 );
nand ( n3345 , n3342 , n3344 );
not ( n3346 , n2917 );
and ( n3347 , n3346 , n1479 );
not ( n3348 , n3346 );
and ( n3349 , n3348 , n1009 );
nor ( n3350 , n3347 , n3349 );
or ( n3351 , n3350 , n2962 );
not ( n3352 , n161 );
nand ( n3353 , n59 , n3352 );
nand ( n3354 , n3351 , n3353 );
not ( n3355 , n3101 );
not ( n3356 , n3355 );
nand ( n3357 , n3071 , n3009 );
not ( n3358 , n3357 );
not ( n3359 , n3068 );
or ( n3360 , n3358 , n3359 );
or ( n3361 , n3357 , n3068 );
nand ( n3362 , n3360 , n3361 );
not ( n3363 , n3362 );
or ( n3364 , n3356 , n3363 );
not ( n3365 , n3206 );
not ( n3366 , n3214 );
nand ( n3367 , n3366 , n3212 );
not ( n3368 , n3367 );
not ( n3369 , n3368 );
or ( n3370 , n3365 , n3369 );
not ( n3371 , n3206 );
and ( n3372 , n3371 , n3367 );
nor ( n3373 , n3372 , n3135 );
nand ( n3374 , n3370 , n3373 );
nand ( n3375 , n3364 , n3374 );
nor ( n3376 , n3354 , n3375 );
or ( n3377 , n59 , n3125 );
nand ( n3378 , n3377 , n3126 , n3140 );
not ( n3379 , n3113 );
nand ( n3380 , n1009 , n3379 );
not ( n3381 , n2971 );
not ( n3382 , n1315 );
or ( n3383 , n3381 , n3382 );
not ( n3384 , n2992 );
nand ( n3385 , n2991 , n1034 );
nand ( n3386 , n3384 , n3385 , n2864 );
nand ( n3387 , n3383 , n3386 );
nand ( n3388 , n3387 , n2970 );
nand ( n3389 , n3376 , n3378 , n3380 , n3388 );
not ( n3390 , n43 );
nor ( n3391 , n3390 , n161 );
not ( n3392 , n2770 );
not ( n3393 , n3379 );
or ( n3394 , n3392 , n3393 );
not ( n3395 , n3139 );
not ( n3396 , n43 );
nand ( n3397 , n3396 , n3124 );
not ( n3398 , n3125 );
nand ( n3399 , n3395 , n3397 , n3398 );
nand ( n3400 , n3394 , n3399 );
nor ( n3401 , n3391 , n3400 );
not ( n3402 , n3160 );
not ( n3403 , n3402 );
not ( n3404 , n3202 );
or ( n3405 , n3403 , n3404 );
not ( n3406 , n3164 );
nand ( n3407 , n3405 , n3406 );
nand ( n3408 , n3407 , n3174 );
not ( n3409 , n3171 );
and ( n3410 , n3205 , n3409 );
and ( n3411 , n3408 , n3410 );
nor ( n3412 , n3411 , n3240 );
not ( n3413 , n3410 );
not ( n3414 , n3408 );
nand ( n3415 , n3413 , n3414 );
and ( n3416 , n3412 , n3415 );
not ( n3417 , n3027 );
not ( n3418 , n3417 );
not ( n3419 , n3064 );
not ( n3420 , n3419 );
or ( n3421 , n3418 , n3420 );
not ( n3422 , n3029 );
nand ( n3423 , n3421 , n3422 );
nand ( n3424 , n3423 , n3036 );
nand ( n3425 , n3067 , n3032 );
not ( n3426 , n3425 );
and ( n3427 , n3424 , n3426 );
not ( n3428 , n3424 );
and ( n3429 , n3428 , n3425 );
nor ( n3430 , n3427 , n3429 );
and ( n3431 , n3430 , n3355 );
nor ( n3432 , n3416 , n3431 );
not ( n3433 , n2916 );
and ( n3434 , n3433 , n2757 );
not ( n3435 , n3433 );
and ( n3436 , n3435 , n2758 );
nor ( n3437 , n3434 , n3436 );
not ( n3438 , n3437 );
not ( n3439 , n2962 );
and ( n3440 , n3438 , n3439 );
not ( n3441 , n2991 );
not ( n3442 , n966 );
not ( n3443 , n2990 );
not ( n3444 , n3443 );
or ( n3445 , n3442 , n3444 );
nand ( n3446 , n3445 , n2864 );
or ( n3447 , n3441 , n3446 );
not ( n3448 , n1297 );
or ( n3449 , n2864 , n3448 );
nand ( n3450 , n3447 , n3449 );
and ( n3451 , n2970 , n3450 );
nor ( n3452 , n3440 , n3451 );
nand ( n3453 , n3401 , n3432 , n3452 );
not ( n3454 , n52 );
not ( n3455 , n3341 );
or ( n3456 , n3454 , n3455 );
not ( n3457 , n2971 );
buf ( n3458 , n3322 );
not ( n3459 , n3458 );
or ( n3460 , n3457 , n3459 );
not ( n3461 , n3448 );
not ( n3462 , n2986 );
nand ( n3463 , n2981 , n3462 );
nor ( n3464 , n1331 , n3463 );
not ( n3465 , n3464 );
not ( n3466 , n3465 );
or ( n3467 , n3461 , n3466 );
and ( n3468 , n1297 , n3464 );
nor ( n3469 , n3468 , n2971 );
nand ( n3470 , n3467 , n3469 );
nand ( n3471 , n3460 , n3470 );
and ( n3472 , n2900 , n3471 );
and ( n3473 , n2914 , n2733 );
not ( n3474 , n2914 );
and ( n3475 , n3474 , n2732 );
nor ( n3476 , n3473 , n3475 );
and ( n3477 , n3301 , n3476 );
and ( n3478 , n3106 , n2734 );
nor ( n3479 , n3477 , n3478 );
not ( n3480 , n3178 );
not ( n3481 , n3480 );
not ( n3482 , n3201 );
not ( n3483 , n3482 );
not ( n3484 , n3483 );
or ( n3485 , n3481 , n3484 );
not ( n3486 , n3151 );
nand ( n3487 , n3485 , n3486 );
not ( n3488 , n3487 );
nand ( n3489 , n3159 , n3154 );
not ( n3490 , n3489 );
or ( n3491 , n3488 , n3490 );
or ( n3492 , n3487 , n3489 );
nand ( n3493 , n3491 , n3492 );
nand ( n3494 , n3311 , n3493 );
not ( n3495 , n3060 );
not ( n3496 , n3495 );
not ( n3497 , n3062 );
and ( n3498 , n3496 , n3497 );
nor ( n3499 , n3498 , n3017 );
not ( n3500 , n3499 );
and ( n3501 , n3026 , n3022 );
not ( n3502 , n3501 );
or ( n3503 , n3500 , n3502 );
or ( n3504 , n3499 , n3501 );
nand ( n3505 , n3503 , n3504 );
nand ( n3506 , n3099 , n3505 );
nand ( n3507 , n3479 , n3494 , n3506 );
nor ( n3508 , n3472 , n3507 );
or ( n3509 , n3508 , n3341 );
nand ( n3510 , n3456 , n3509 );
not ( n3511 , n50 );
not ( n3512 , n2943 );
not ( n3513 , n2958 );
nor ( n3514 , n3340 , n3513 );
nand ( n3515 , n3512 , n3338 , n3514 );
not ( n3516 , n3515 );
or ( n3517 , n3511 , n3516 );
or ( n3518 , n3508 , n3515 );
nand ( n3519 , n3517 , n3518 );
not ( n3520 , n45 );
and ( n3521 , n3341 , n3520 );
not ( n3522 , n3341 );
not ( n3523 , n2899 );
not ( n3524 , n2971 );
not ( n3525 , n1403 );
or ( n3526 , n3524 , n3525 );
not ( n3527 , n3463 );
nor ( n3528 , n1352 , n3527 );
not ( n3529 , n3528 );
nand ( n3530 , n3529 , n2864 , n3465 );
nand ( n3531 , n3526 , n3530 );
and ( n3532 , n3523 , n3531 );
not ( n3533 , n1341 );
and ( n3534 , n3533 , n2913 );
nor ( n3535 , n3534 , n2914 );
and ( n3536 , n3301 , n3535 );
and ( n3537 , n3106 , n3533 );
nor ( n3538 , n3536 , n3537 );
nand ( n3539 , n3486 , n3480 );
xor ( n3540 , n3482 , n3539 );
nand ( n3541 , n3540 , n3311 );
not ( n3542 , n3017 );
nand ( n3543 , n3542 , n3497 );
xor ( n3544 , n3495 , n3543 );
nand ( n3545 , n3544 , n3099 );
nand ( n3546 , n3538 , n3541 , n3545 );
nor ( n3547 , n3532 , n3546 );
and ( n3548 , n3522 , n3547 );
nor ( n3549 , n3521 , n3548 );
and ( n3550 , n2898 , n740 );
nor ( n3551 , n3550 , n3514 );
not ( n3552 , n2017 );
not ( n3553 , n2926 );
or ( n3554 , n3552 , n3553 );
nand ( n3555 , n3554 , n3512 );
nand ( n3556 , n3551 , n3338 , n3555 );
and ( n3557 , n49 , n3556 );
nand ( n3558 , n3338 , n2943 );
nor ( n3559 , n2958 , n3558 );
nand ( n3560 , n3106 , n3559 );
not ( n3561 , n3560 );
and ( n3562 , n2734 , n3561 );
xor ( n3563 , n51 , n3122 );
not ( n3564 , n3111 );
and ( n3565 , n3563 , n3564 );
nor ( n3566 , n3557 , n3562 , n3565 );
nand ( n3567 , n3301 , n3559 );
not ( n3568 , n3567 );
not ( n3569 , n3476 );
not ( n3570 , n3569 );
and ( n3571 , n3568 , n3570 );
nor ( n3572 , n2958 , n3558 );
and ( n3573 , n3099 , n3572 );
and ( n3574 , n3573 , n3505 );
nor ( n3575 , n3571 , n3574 );
nand ( n3576 , n3134 , n3572 );
not ( n3577 , n3576 );
nand ( n3578 , n3577 , n3493 );
nor ( n3579 , n2898 , n741 );
and ( n3580 , n3579 , n3559 );
nand ( n3581 , n3471 , n3580 );
nand ( n3582 , n3566 , n3575 , n3578 , n3581 );
not ( n3583 , n35 );
not ( n3584 , n3123 );
nand ( n3585 , n3583 , n3584 );
and ( n3586 , n3585 , n3124 , n3140 );
not ( n3587 , n35 );
nor ( n3588 , n3587 , n161 );
nor ( n3589 , n3586 , n3588 );
not ( n3590 , n2746 );
nand ( n3591 , n3590 , n3114 );
nand ( n3592 , n3059 , n3295 );
nand ( n3593 , n3592 , n3063 , n3039 );
nand ( n3594 , n3417 , n3593 );
not ( n3595 , n3594 );
nand ( n3596 , n3036 , n3422 );
not ( n3597 , n3596 );
and ( n3598 , n3595 , n3597 );
and ( n3599 , n3594 , n3596 );
nor ( n3600 , n3598 , n3599 );
nor ( n3601 , n3600 , n3101 );
or ( n3602 , n3313 , n3196 );
not ( n3603 , n3179 );
not ( n3604 , n3183 );
nor ( n3605 , n3603 , n3604 );
nand ( n3606 , n3602 , n3605 );
nand ( n3607 , n3402 , n3606 );
not ( n3608 , n3607 );
and ( n3609 , n3174 , n3406 );
not ( n3610 , n3609 );
or ( n3611 , n3608 , n3610 );
nand ( n3612 , n3611 , n3239 );
nor ( n3613 , n3607 , n3609 );
nor ( n3614 , n3612 , n3613 );
nor ( n3615 , n3601 , n3614 );
not ( n3616 , n2962 );
not ( n3617 , n2915 );
not ( n3618 , n2745 );
and ( n3619 , n3617 , n3618 );
not ( n3620 , n3617 );
and ( n3621 , n3620 , n2745 );
nor ( n3622 , n3619 , n3621 );
not ( n3623 , n3622 );
and ( n3624 , n3616 , n3623 );
not ( n3625 , n2971 );
not ( n3626 , n1352 );
or ( n3627 , n3625 , n3626 );
not ( n3628 , n2988 );
nor ( n3629 , n3628 , n1315 );
not ( n3630 , n3629 );
nand ( n3631 , n3630 , n2864 , n3443 );
nand ( n3632 , n3627 , n3631 );
and ( n3633 , n2970 , n3632 );
nor ( n3634 , n3624 , n3633 );
nand ( n3635 , n3589 , n3591 , n3615 , n3634 );
not ( n3636 , n51 );
nor ( n3637 , n3636 , n161 );
not ( n3638 , n3493 );
or ( n3639 , n3240 , n3638 );
nand ( n3640 , n3355 , n3505 );
nand ( n3641 , n3639 , n3640 );
nor ( n3642 , n3637 , n3641 );
and ( n3643 , n3563 , n3140 );
not ( n3644 , n2735 );
and ( n3645 , n3644 , n3379 );
nor ( n3646 , n3643 , n3645 );
nand ( n3647 , n2963 , n3476 );
nand ( n3648 , n3471 , n2970 );
nand ( n3649 , n3642 , n3646 , n3647 , n3648 );
or ( n3650 , n39 , n47 );
nand ( n3651 , n3650 , n3121 );
not ( n3652 , n3651 );
and ( n3653 , n3652 , n3140 );
not ( n3654 , n3544 );
or ( n3655 , n3654 , n3101 );
not ( n3656 , n3535 );
or ( n3657 , n2962 , n3656 );
nand ( n3658 , n3655 , n3657 );
nor ( n3659 , n3653 , n3658 );
not ( n3660 , n3533 );
not ( n3661 , n3660 );
nand ( n3662 , n3661 , n3114 );
nand ( n3663 , n47 , n3352 );
not ( n3664 , n3540 );
not ( n3665 , n3664 );
not ( n3666 , n3239 );
not ( n3667 , n3666 );
and ( n3668 , n3665 , n3667 );
and ( n3669 , n3531 , n2970 );
nor ( n3670 , n3668 , n3669 );
nand ( n3671 , n3659 , n3662 , n3663 , n3670 );
not ( n3672 , n2971 );
not ( n3673 , n2975 );
not ( n3674 , n3673 );
not ( n3675 , n3674 );
or ( n3676 , n3672 , n3675 );
not ( n3677 , n3326 );
nor ( n3678 , n3677 , n1403 );
not ( n3679 , n3678 );
nand ( n3680 , n3679 , n2864 , n3328 );
nand ( n3681 , n3676 , n3680 );
and ( n3682 , n2900 , n3681 );
not ( n3683 , n2909 );
xnor ( n3684 , n2911 , n3683 );
and ( n3685 , n3301 , n3684 );
not ( n3686 , n3683 );
and ( n3687 , n3106 , n3686 );
nor ( n3688 , n3685 , n3687 );
nand ( n3689 , n3053 , n3049 );
not ( n3690 , n3689 );
not ( n3691 , n3046 );
or ( n3692 , n3690 , n3691 );
or ( n3693 , n3689 , n3046 );
nand ( n3694 , n3692 , n3693 );
and ( n3695 , n3099 , n3694 );
not ( n3696 , n3185 );
not ( n3697 , n3696 );
not ( n3698 , n3190 );
nand ( n3699 , n3697 , n3698 );
nand ( n3700 , n3699 , n3187 );
not ( n3701 , n3191 );
nand ( n3702 , n3195 , n3701 );
not ( n3703 , n3702 );
and ( n3704 , n3700 , n3703 );
not ( n3705 , n3700 );
and ( n3706 , n3705 , n3702 );
nor ( n3707 , n3704 , n3706 );
and ( n3708 , n3311 , n3707 );
nor ( n3709 , n3695 , n3708 );
nand ( n3710 , n3688 , n3709 );
nor ( n3711 , n3682 , n3710 );
or ( n3712 , n3711 , n3341 );
not ( n3713 , n156 );
or ( n3714 , n3713 , n3343 );
nand ( n3715 , n3712 , n3714 );
and ( n3716 , n3299 , n3355 );
and ( n3717 , n3304 , n3379 );
nor ( n3718 , n1279 , n161 );
nor ( n3719 , n3716 , n3717 , n3718 );
and ( n3720 , n1279 , n3140 );
not ( n3721 , n3666 );
and ( n3722 , n3721 , n3315 );
nor ( n3723 , n3720 , n3722 );
nand ( n3724 , n2963 , n3306 );
nand ( n3725 , n2970 , n3334 );
nand ( n3726 , n3719 , n3723 , n3724 , n3725 );
and ( n3727 , n37 , n3556 );
and ( n3728 , n3304 , n3561 );
and ( n3729 , n1279 , n3564 );
nor ( n3730 , n3727 , n3728 , n3729 );
and ( n3731 , n3299 , n3573 );
not ( n3732 , n3567 );
and ( n3733 , n3732 , n3306 );
nor ( n3734 , n3731 , n3733 );
nand ( n3735 , n3577 , n3315 );
nand ( n3736 , n3580 , n3334 );
nand ( n3737 , n3730 , n3734 , n3735 , n3736 );
and ( n3738 , n3686 , n3561 );
and ( n3739 , n3573 , n3694 );
and ( n3740 , n154 , n3564 );
nor ( n3741 , n3738 , n3739 , n3740 );
and ( n3742 , n3684 , n3732 );
and ( n3743 , n155 , n3556 );
nor ( n3744 , n3742 , n3743 );
nand ( n3745 , n3580 , n3681 );
nand ( n3746 , n3577 , n3707 );
nand ( n3747 , n3741 , n3744 , n3745 , n3746 );
and ( n3748 , n3732 , n3535 );
or ( n3749 , n3660 , n3560 );
or ( n3750 , n3651 , n3111 );
nand ( n3751 , n3749 , n3750 );
nor ( n3752 , n3748 , n3751 );
and ( n3753 , n48 , n3556 );
and ( n3754 , n3544 , n3573 );
nor ( n3755 , n3753 , n3754 );
nand ( n3756 , n3540 , n3577 );
nand ( n3757 , n3531 , n3580 );
nand ( n3758 , n3752 , n3755 , n3756 , n3757 );
and ( n3759 , n3686 , n3114 );
and ( n3760 , n3355 , n3694 );
nor ( n3761 , n3759 , n3760 );
and ( n3762 , n3684 , n2963 );
and ( n3763 , n3721 , n3707 );
nor ( n3764 , n3762 , n3763 );
nand ( n3765 , n2970 , n3681 );
nand ( n3766 , n161 , n3139 );
nand ( n3767 , n154 , n3766 );
nand ( n3768 , n3761 , n3764 , n3765 , n3767 );
nor ( n3769 , n3319 , n3325 );
not ( n3770 , n3769 );
nand ( n3771 , n3770 , n3326 , n2864 );
nand ( n3772 , n2971 , n1455 );
nand ( n3773 , n3771 , n3772 );
and ( n3774 , n3523 , n3773 );
not ( n3775 , n3696 );
not ( n3776 , n3187 );
not ( n3777 , n3698 );
nor ( n3778 , n3776 , n3777 );
not ( n3779 , n3778 );
or ( n3780 , n3775 , n3779 );
or ( n3781 , n3696 , n3778 );
nand ( n3782 , n3780 , n3781 );
and ( n3783 , n3311 , n3782 );
not ( n3784 , n3042 );
not ( n3785 , n3045 );
or ( n3786 , n3784 , n3785 );
or ( n3787 , n3042 , n3045 );
nand ( n3788 , n3786 , n3787 );
and ( n3789 , n3099 , n3788 );
nor ( n3790 , n3783 , n3789 );
not ( n3791 , n2910 );
xnor ( n3792 , n3791 , n1437 );
and ( n3793 , n3301 , n3792 );
and ( n3794 , n3106 , n3791 );
nor ( n3795 , n3793 , n3794 );
nand ( n3796 , n3790 , n3795 );
nor ( n3797 , n3774 , n3796 );
or ( n3798 , n3797 , n3341 );
not ( n3799 , n151 );
or ( n3800 , n3799 , n3343 );
nand ( n3801 , n3798 , n3800 );
nor ( n3802 , n3674 , n3462 );
not ( n3803 , n3802 );
not ( n3804 , n3325 );
nand ( n3805 , n3803 , n2864 , n3804 );
or ( n3806 , n2899 , n3805 );
nand ( n3807 , n3099 , n2211 );
nand ( n3808 , n3806 , n3807 );
not ( n3809 , n3311 );
not ( n3810 , n2211 );
or ( n3811 , n3809 , n3810 );
or ( n3812 , n3106 , n3301 );
not ( n3813 , n1437 );
nand ( n3814 , n3812 , n3813 );
nand ( n3815 , n3811 , n3814 );
nor ( n3816 , n3808 , n3815 );
or ( n3817 , n3816 , n3341 );
not ( n3818 , n149 );
or ( n3819 , n3818 , n3343 );
nand ( n3820 , n3817 , n3819 );
not ( n3821 , n148 );
and ( n3822 , n3515 , n3821 );
not ( n3823 , n3515 );
and ( n3824 , n3823 , n3816 );
nor ( n3825 , n3822 , n3824 );
and ( n3826 , n3782 , n3577 );
and ( n3827 , n3573 , n3788 );
not ( n3828 , n150 );
nor ( n3829 , n3828 , n3111 );
nor ( n3830 , n3826 , n3827 , n3829 );
and ( n3831 , n153 , n3556 );
and ( n3832 , n3791 , n3561 );
nor ( n3833 , n3831 , n3832 );
nand ( n3834 , n3792 , n3732 );
nand ( n3835 , n3773 , n3580 );
nand ( n3836 , n3830 , n3833 , n3834 , n3835 );
and ( n3837 , n150 , n3766 );
and ( n3838 , n3791 , n3112 );
nor ( n3839 , n3837 , n3838 );
and ( n3840 , n3782 , n3239 );
and ( n3841 , n3355 , n3788 );
nor ( n3842 , n3840 , n3841 );
not ( n3843 , n2962 );
nand ( n3844 , n3792 , n3843 );
not ( n3845 , n2969 );
nand ( n3846 , n3773 , n3845 );
nand ( n3847 , n3839 , n3842 , n3844 , n3846 );
and ( n3848 , n3573 , n2211 );
and ( n3849 , n146 , n3564 );
nor ( n3850 , n3848 , n3849 );
not ( n3851 , n3576 );
not ( n3852 , n2211 );
not ( n3853 , n3852 );
and ( n3854 , n3851 , n3853 );
nand ( n3855 , n3560 , n3567 );
and ( n3856 , n3813 , n3855 );
nor ( n3857 , n3854 , n3856 );
not ( n3858 , n3805 );
nand ( n3859 , n3580 , n3858 );
nand ( n3860 , n147 , n3556 );
nand ( n3861 , n3850 , n3857 , n3859 , n3860 );
not ( n3862 , n3138 );
nand ( n3863 , n3813 , n3862 );
nand ( n3864 , n3136 , n2211 );
nand ( n3865 , n3845 , n3858 );
nand ( n3866 , n146 , n3766 );
nand ( n3867 , n3863 , n3864 , n3865 , n3866 );
not ( n3868 , n2923 );
nor ( n3869 , n714 , n3868 );
nand ( n3870 , n161 , n3869 );
not ( n3871 , n3870 );
not ( n3872 , n3871 );
buf ( n3873 , n3872 );
not ( n3874 , n3873 );
and ( n3875 , n3874 , n2495 );
not ( n3876 , n3874 );
not ( n3877 , n174 );
and ( n3878 , n3876 , n3877 );
nor ( n3879 , n3875 , n3878 );
not ( n3880 , n2510 );
or ( n3881 , n3873 , n3880 );
not ( n3882 , n175 );
not ( n3883 , n3870 );
not ( n3884 , n3883 );
buf ( n3885 , n3884 );
not ( n3886 , n3885 );
or ( n3887 , n3882 , n3886 );
nand ( n3888 , n3881 , n3887 );
and ( n3889 , n3886 , n1648 );
not ( n3890 , n3886 );
not ( n3891 , n177 );
and ( n3892 , n3890 , n3891 );
nor ( n3893 , n3889 , n3892 );
not ( n3894 , n205 );
and ( n3895 , n3873 , n3894 );
not ( n3896 , n3873 );
and ( n3897 , n3896 , n1769 );
nor ( n3898 , n3895 , n3897 );
or ( n3899 , n3873 , n1748 );
not ( n3900 , n206 );
not ( n3901 , n3872 );
or ( n3902 , n3900 , n3901 );
nand ( n3903 , n3899 , n3902 );
not ( n3904 , n3871 );
buf ( n3905 , n3904 );
not ( n3906 , n2549 );
or ( n3907 , n3905 , n3906 );
not ( n3908 , n178 );
not ( n3909 , n3871 );
not ( n3910 , n3909 );
or ( n3911 , n3908 , n3910 );
nand ( n3912 , n3907 , n3911 );
not ( n3913 , n173 );
and ( n3914 , n3885 , n3913 );
not ( n3915 , n3885 );
not ( n3916 , n2462 );
and ( n3917 , n3915 , n3916 );
nor ( n3918 , n3914 , n3917 );
not ( n3919 , n3884 );
not ( n3920 , n3919 );
or ( n3921 , n3920 , n1705 );
not ( n3922 , n176 );
or ( n3923 , n3922 , n3910 );
nand ( n3924 , n3921 , n3923 );
and ( n3925 , n3886 , n2627 );
not ( n3926 , n3886 );
not ( n3927 , n179 );
and ( n3928 , n3926 , n3927 );
nor ( n3929 , n3925 , n3928 );
not ( n3930 , n210 );
and ( n3931 , n3909 , n3930 );
not ( n3932 , n3909 );
and ( n3933 , n3932 , n2682 );
nor ( n3934 , n3931 , n3933 );
not ( n3935 , n211 );
and ( n3936 , n3905 , n3935 );
not ( n3937 , n3905 );
and ( n3938 , n3937 , n1209 );
nor ( n3939 , n3936 , n3938 );
not ( n3940 , n2720 );
or ( n3941 , n3920 , n3940 );
not ( n3942 , n213 );
or ( n3943 , n3942 , n3910 );
nand ( n3944 , n3941 , n3943 );
not ( n3945 , n218 );
and ( n3946 , n3872 , n3945 );
not ( n3947 , n3872 );
and ( n3948 , n3947 , n1110 );
nor ( n3949 , n3946 , n3948 );
and ( n3950 , n3886 , n1955 );
not ( n3951 , n3886 );
not ( n3952 , n181 );
and ( n3953 , n3951 , n3952 );
nor ( n3954 , n3950 , n3953 );
not ( n3955 , n3871 );
not ( n3956 , n1181 );
or ( n3957 , n3955 , n3956 );
nand ( n3958 , n212 , n3884 );
nand ( n3959 , n3957 , n3958 );
not ( n3960 , n2622 );
or ( n3961 , n3905 , n3960 );
not ( n3962 , n180 );
or ( n3963 , n3962 , n3919 );
nand ( n3964 , n3961 , n3963 );
or ( n3965 , n3873 , n1846 );
not ( n3966 , n203 );
or ( n3967 , n3966 , n3901 );
nand ( n3968 , n3965 , n3967 );
not ( n3969 , n2588 );
or ( n3970 , n3920 , n3969 );
not ( n3971 , n204 );
or ( n3972 , n3971 , n3910 );
nand ( n3973 , n3970 , n3972 );
not ( n3974 , n2572 );
or ( n3975 , n3920 , n3974 );
not ( n3976 , n207 );
or ( n3977 , n3976 , n3910 );
nand ( n3978 , n3975 , n3977 );
or ( n3979 , n3920 , n1919 );
not ( n3980 , n208 );
or ( n3981 , n3980 , n3910 );
nand ( n3982 , n3979 , n3981 );
not ( n3983 , n214 );
not ( n3984 , n3871 );
not ( n3985 , n3984 );
or ( n3986 , n3983 , n3985 );
or ( n3987 , n3909 , n2708 );
nand ( n3988 , n3986 , n3987 );
not ( n3989 , n215 );
not ( n3990 , n3909 );
or ( n3991 , n3989 , n3990 );
or ( n3992 , n3872 , n1034 );
nand ( n3993 , n3991 , n3992 );
or ( n3994 , n3905 , n1971 );
not ( n3995 , n209 );
or ( n3996 , n3995 , n3919 );
nand ( n3997 , n3994 , n3996 );
or ( n3998 , n714 , n737 );
not ( n3999 , n1001 );
or ( n4000 , n3999 , n2971 );
nand ( n4001 , n3998 , n4000 );
not ( n4002 , n3869 );
nand ( n4003 , n4001 , n161 , n4002 );
not ( n4004 , n4003 );
and ( n4005 , n221 , n4004 );
and ( n4006 , n111 , n3352 );
nor ( n4007 , n4005 , n4006 );
not ( n4008 , n1884 );
xor ( n4009 , n110 , n4008 );
not ( n4010 , n113 );
nand ( n4011 , n4010 , n1866 );
not ( n4012 , n122 );
nand ( n4013 , n4012 , n1894 );
not ( n4014 , n4013 );
not ( n4015 , n1923 );
nor ( n4016 , n117 , n4015 );
nor ( n4017 , n4014 , n4016 );
nand ( n4018 , n4011 , n4017 );
not ( n4019 , n4018 );
nor ( n4020 , n79 , n1125 );
not ( n4021 , n4020 );
not ( n4022 , n82 );
nand ( n4023 , n4022 , n1111 );
nand ( n4024 , n4021 , n4023 );
not ( n4025 , n74 );
not ( n4026 , n500 );
nand ( n4027 , n4025 , n4026 );
not ( n4028 , n70 );
not ( n4029 , n1192 );
nand ( n4030 , n4028 , n4029 );
and ( n4031 , n4027 , n4030 );
nor ( n4032 , n63 , n1214 );
not ( n4033 , n1255 );
nor ( n4034 , n66 , n4033 );
nor ( n4035 , n4032 , n4034 );
nand ( n4036 , n58 , n967 );
not ( n4037 , n599 );
nor ( n4038 , n54 , n4037 );
or ( n4039 , n4036 , n4038 );
nand ( n4040 , n54 , n4037 );
nand ( n4041 , n4039 , n4040 );
and ( n4042 , n4035 , n4041 );
nand ( n4043 , n63 , n1214 );
or ( n4044 , n4043 , n4034 );
nand ( n4045 , n66 , n1256 );
nand ( n4046 , n4044 , n4045 );
nor ( n4047 , n4042 , n4046 );
nand ( n4048 , n34 , n1270 );
not ( n4049 , n4048 );
nor ( n4050 , n41 , n626 );
not ( n4051 , n4050 );
and ( n4052 , n4049 , n4051 );
not ( n4053 , n1269 );
nor ( n4054 , n34 , n4053 );
nor ( n4055 , n4054 , n4050 );
and ( n4056 , n46 , n1333 );
not ( n4057 , n4056 );
not ( n4058 , n637 );
or ( n4059 , n50 , n4058 );
not ( n4060 , n4059 );
or ( n4061 , n4057 , n4060 );
nand ( n4062 , n50 , n1318 );
nand ( n4063 , n4061 , n4062 );
and ( n4064 , n4055 , n4063 );
nor ( n4065 , n4052 , n4064 );
nand ( n4066 , n41 , n1299 );
nor ( n4067 , n46 , n1334 );
not ( n4068 , n506 );
or ( n4069 , n38 , n4068 );
nor ( n4070 , n157 , n567 );
nand ( n4071 , n6 , n148 );
not ( n4072 , n4071 );
nand ( n4073 , n4072 , n152 );
not ( n4074 , n152 );
not ( n4075 , n4071 );
or ( n4076 , n4074 , n4075 );
or ( n4077 , n152 , n4071 );
nand ( n4078 , n4076 , n4077 );
nand ( n4079 , n4078 , n650 );
and ( n4080 , n4073 , n4079 );
or ( n4081 , n4070 , n4080 );
nand ( n4082 , n157 , n567 );
nand ( n4083 , n4081 , n4082 );
and ( n4084 , n4069 , n4083 );
not ( n4085 , n506 );
and ( n4086 , n38 , n4085 );
nor ( n4087 , n4084 , n4086 );
nor ( n4088 , n4067 , n4087 );
and ( n4089 , n4059 , n4088 );
nand ( n4090 , n4055 , n4089 );
and ( n4091 , n4065 , n4066 , n4090 );
nor ( n4092 , n58 , n967 );
nor ( n4093 , n4091 , n4092 , n4038 );
nand ( n4094 , n4035 , n4093 );
nand ( n4095 , n4047 , n4094 );
nand ( n4096 , n4031 , n4095 );
nor ( n4097 , n4024 , n4096 );
and ( n4098 , n4019 , n4097 );
not ( n4099 , n4011 );
nand ( n4100 , n122 , n1895 );
or ( n4101 , n4100 , n4016 );
nand ( n4102 , n117 , n1924 );
nand ( n4103 , n4101 , n4102 );
not ( n4104 , n4103 );
or ( n4105 , n4099 , n4104 );
not ( n4106 , n4024 );
and ( n4107 , n74 , n500 );
and ( n4108 , n4107 , n4030 );
not ( n4109 , n70 );
nor ( n4110 , n4109 , n1193 );
nor ( n4111 , n4108 , n4110 );
not ( n4112 , n4111 );
and ( n4113 , n4106 , n4112 );
nand ( n4114 , n82 , n1112 );
or ( n4115 , n4114 , n4020 );
nand ( n4116 , n79 , n1127 );
nand ( n4117 , n4115 , n4116 );
nor ( n4118 , n4113 , n4117 );
or ( n4119 , n4018 , n4118 );
nand ( n4120 , n4105 , n4119 );
not ( n4121 , n113 );
nor ( n4122 , n4121 , n1866 );
nor ( n4123 , n4098 , n4120 , n4122 );
or ( n4124 , n4009 , n4123 );
nand ( n4125 , n4009 , n4123 );
nor ( n4126 , n3999 , n2864 );
or ( n4127 , n738 , n2897 );
nand ( n4128 , n4127 , n2904 );
nand ( n4129 , n4126 , n4128 );
not ( n4130 , n4129 );
nand ( n4131 , n4124 , n4125 , n4130 );
not ( n4132 , n4008 );
not ( n4133 , n4128 );
not ( n4134 , n4133 );
not ( n4135 , n3999 );
nor ( n4136 , n4135 , n2971 );
nand ( n4137 , n4134 , n4136 );
not ( n4138 , n4137 );
nand ( n4139 , n4132 , n4138 );
and ( n4140 , n109 , n4008 );
not ( n4141 , n109 );
and ( n4142 , n4141 , n1884 );
nor ( n4143 , n4140 , n4142 );
not ( n4144 , n4143 );
nor ( n4145 , n112 , n1865 );
not ( n4146 , n4145 );
nor ( n4147 , n121 , n1893 );
nor ( n4148 , n118 , n1922 );
nor ( n4149 , n4147 , n4148 );
nand ( n4150 , n4146 , n4149 );
not ( n4151 , n78 );
nand ( n4152 , n4151 , n707 );
not ( n4153 , n4152 );
nor ( n4154 , n81 , n681 );
nor ( n4155 , n4153 , n4154 );
not ( n4156 , n73 );
nor ( n4157 , n4156 , n4026 );
not ( n4158 , n69 );
nand ( n4159 , n4158 , n695 );
and ( n4160 , n4157 , n4159 );
not ( n4161 , n69 );
nor ( n4162 , n4161 , n695 );
nor ( n4163 , n4160 , n4162 );
not ( n4164 , n4163 );
and ( n4165 , n4155 , n4164 );
and ( n4166 , n81 , n681 );
and ( n4167 , n4166 , n4152 );
not ( n4168 , n78 );
nor ( n4169 , n4168 , n1126 );
nor ( n4170 , n4165 , n4167 , n4169 );
or ( n4171 , n4150 , n4170 );
nand ( n4172 , n121 , n1893 );
or ( n4173 , n4172 , n4148 );
nand ( n4174 , n118 , n1924 );
nand ( n4175 , n4173 , n4174 );
not ( n4176 , n4175 );
or ( n4177 , n4145 , n4176 );
not ( n4178 , n4150 );
or ( n4179 , n73 , n500 );
and ( n4180 , n4179 , n4159 );
nor ( n4181 , n62 , n1214 );
nor ( n4182 , n65 , n667 );
nor ( n4183 , n4181 , n4182 );
nand ( n4184 , n57 , n967 );
nor ( n4185 , n53 , n4037 );
or ( n4186 , n4184 , n4185 );
nand ( n4187 , n53 , n4037 );
nand ( n4188 , n4186 , n4187 );
and ( n4189 , n4183 , n4188 );
nand ( n4190 , n62 , n1214 );
or ( n4191 , n4190 , n4182 );
nand ( n4192 , n65 , n1256 );
nand ( n4193 , n4191 , n4192 );
nor ( n4194 , n4189 , n4193 );
nand ( n4195 , n33 , n1270 );
not ( n4196 , n4195 );
nor ( n4197 , n42 , n626 );
not ( n4198 , n4197 );
and ( n4199 , n4196 , n4198 );
nor ( n4200 , n33 , n525 );
nor ( n4201 , n4200 , n4197 );
not ( n4202 , n637 );
nor ( n4203 , n49 , n4202 );
or ( n4204 , n48 , n1334 );
nand ( n4205 , n942 , n506 );
not ( n4206 , n4205 );
nor ( n4207 , n155 , n567 );
not ( n4208 , n153 );
nand ( n4209 , n6 , n147 );
not ( n4210 , n4209 );
not ( n4211 , n4210 );
or ( n4212 , n4208 , n4211 );
not ( n4213 , n153 );
not ( n4214 , n4209 );
or ( n4215 , n4213 , n4214 );
or ( n4216 , n153 , n4209 );
nand ( n4217 , n4215 , n4216 );
nand ( n4218 , n4217 , n650 );
nand ( n4219 , n4212 , n4218 );
not ( n4220 , n4219 );
or ( n4221 , n4207 , n4220 );
nand ( n4222 , n155 , n567 );
nand ( n4223 , n4221 , n4222 );
not ( n4224 , n4223 );
or ( n4225 , n4206 , n4224 );
nand ( n4226 , n37 , n507 );
nand ( n4227 , n4225 , n4226 );
nand ( n4228 , n4204 , n4227 );
nor ( n4229 , n4203 , n4228 );
and ( n4230 , n4201 , n4229 );
nor ( n4231 , n4199 , n4230 );
nand ( n4232 , n42 , n1299 );
nand ( n4233 , n48 , n1333 );
or ( n4234 , n4233 , n4203 );
nand ( n4235 , n49 , n1318 );
nand ( n4236 , n4234 , n4235 );
nand ( n4237 , n4201 , n4236 );
and ( n4238 , n4231 , n4232 , n4237 );
nor ( n4239 , n57 , n967 );
nor ( n4240 , n4238 , n4239 , n4185 );
nand ( n4241 , n4183 , n4240 );
nand ( n4242 , n4194 , n4241 );
nand ( n4243 , n4180 , n4242 );
not ( n4244 , n4243 );
nand ( n4245 , n4155 , n4244 );
not ( n4246 , n4245 );
and ( n4247 , n4178 , n4246 );
not ( n4248 , n112 );
nor ( n4249 , n4248 , n1866 );
nor ( n4250 , n4247 , n4249 );
nand ( n4251 , n4171 , n4177 , n4250 );
not ( n4252 , n4251 );
or ( n4253 , n4144 , n4252 );
or ( n4254 , n4143 , n4251 );
nand ( n4255 , n4253 , n4254 );
nand ( n4256 , n2865 , n4128 );
not ( n4257 , n4256 );
nand ( n4258 , n4255 , n4257 );
nand ( n4259 , n4007 , n4131 , n4139 , n4258 );
and ( n4260 , n222 , n4004 );
and ( n4261 , n115 , n3352 );
nor ( n4262 , n4260 , n4261 );
not ( n4263 , n4122 );
nand ( n4264 , n4263 , n4011 );
not ( n4265 , n4097 );
nand ( n4266 , n4265 , n4118 );
and ( n4267 , n4017 , n4266 );
nor ( n4268 , n4267 , n4103 );
or ( n4269 , n4264 , n4268 );
nand ( n4270 , n4264 , n4268 );
nand ( n4271 , n4269 , n4270 , n4130 );
not ( n4272 , n1866 );
nand ( n4273 , n4272 , n4138 );
nor ( n4274 , n4249 , n4145 );
not ( n4275 , n4274 );
nand ( n4276 , n4170 , n4245 );
and ( n4277 , n4149 , n4276 );
nor ( n4278 , n4277 , n4175 );
not ( n4279 , n4278 );
or ( n4280 , n4275 , n4279 );
or ( n4281 , n4274 , n4278 );
nand ( n4282 , n4280 , n4281 );
nand ( n4283 , n4282 , n4257 );
nand ( n4284 , n4262 , n4271 , n4273 , n4283 );
and ( n4285 , n223 , n4004 );
and ( n4286 , n119 , n3352 );
nor ( n4287 , n4285 , n4286 );
not ( n4288 , n4102 );
nor ( n4289 , n4288 , n4016 );
not ( n4290 , n4013 );
not ( n4291 , n4266 );
or ( n4292 , n4290 , n4291 );
nand ( n4293 , n4292 , n4100 );
or ( n4294 , n4289 , n4293 );
nand ( n4295 , n4289 , n4293 );
nand ( n4296 , n4294 , n4295 , n4130 );
not ( n4297 , n1925 );
nand ( n4298 , n4297 , n4138 );
not ( n4299 , n4148 );
nand ( n4300 , n4299 , n4174 );
not ( n4301 , n4300 );
not ( n4302 , n4276 );
or ( n4303 , n4147 , n4302 );
nand ( n4304 , n4303 , n4172 );
not ( n4305 , n4304 );
or ( n4306 , n4301 , n4305 );
or ( n4307 , n4300 , n4304 );
nand ( n4308 , n4306 , n4307 );
nand ( n4309 , n4308 , n4257 );
nand ( n4310 , n4287 , n4296 , n4298 , n4309 );
and ( n4311 , n224 , n4004 );
and ( n4312 , n123 , n3352 );
nor ( n4313 , n4311 , n4312 );
and ( n4314 , n4100 , n4013 );
or ( n4315 , n4314 , n4266 );
nand ( n4316 , n4314 , n4266 );
nand ( n4317 , n4315 , n4316 , n4130 );
not ( n4318 , n1896 );
nand ( n4319 , n4318 , n4138 );
not ( n4320 , n4147 );
nand ( n4321 , n4320 , n4172 );
not ( n4322 , n4321 );
not ( n4323 , n4276 );
or ( n4324 , n4322 , n4323 );
or ( n4325 , n4321 , n4276 );
nand ( n4326 , n4324 , n4325 );
nand ( n4327 , n4326 , n4257 );
nand ( n4328 , n4313 , n4317 , n4319 , n4327 );
not ( n4329 , n4169 );
nand ( n4330 , n4329 , n4152 );
not ( n4331 , n4330 );
not ( n4332 , n4154 );
nand ( n4333 , n4332 , n4180 );
or ( n4334 , n4333 , n4241 );
or ( n4335 , n4154 , n4163 );
not ( n4336 , n4333 );
not ( n4337 , n4194 );
and ( n4338 , n4336 , n4337 );
nor ( n4339 , n4338 , n4166 );
nand ( n4340 , n4334 , n4335 , n4339 );
nand ( n4341 , n4331 , n4340 );
not ( n4342 , n4340 );
nand ( n4343 , n4330 , n4342 );
and ( n4344 , n4341 , n4343 , n4257 );
and ( n4345 , n225 , n4004 );
nor ( n4346 , n4344 , n4345 );
not ( n4347 , n1128 );
and ( n4348 , n4347 , n4138 );
and ( n4349 , n77 , n3352 );
nor ( n4350 , n4348 , n4349 );
not ( n4351 , n4020 );
nand ( n4352 , n4351 , n4116 );
not ( n4353 , n4111 );
and ( n4354 , n4023 , n4353 );
nand ( n4355 , n4023 , n4031 );
or ( n4356 , n4355 , n4094 );
nand ( n4357 , n4356 , n4114 );
nor ( n4358 , n4355 , n4047 );
nor ( n4359 , n4354 , n4357 , n4358 );
or ( n4360 , n4352 , n4359 );
nand ( n4361 , n4352 , n4359 );
nand ( n4362 , n4360 , n4361 , n4130 );
nand ( n4363 , n4346 , n4350 , n4362 );
nor ( n4364 , n4166 , n4154 );
nand ( n4365 , n4163 , n4243 );
nand ( n4366 , n4364 , n4365 );
not ( n4367 , n4364 );
not ( n4368 , n4365 );
nand ( n4369 , n4367 , n4368 );
and ( n4370 , n4366 , n4369 , n4257 );
and ( n4371 , n226 , n4004 );
nor ( n4372 , n4370 , n4371 );
not ( n4373 , n1113 );
and ( n4374 , n4373 , n4138 );
and ( n4375 , n83 , n3352 );
nor ( n4376 , n4374 , n4375 );
and ( n4377 , n4114 , n4023 );
nand ( n4378 , n4111 , n4096 );
or ( n4379 , n4377 , n4378 );
nand ( n4380 , n4377 , n4378 );
nand ( n4381 , n4379 , n4380 , n4130 );
nand ( n4382 , n4372 , n4376 , n4381 );
not ( n4383 , n1193 );
and ( n4384 , n4383 , n4138 );
and ( n4385 , n71 , n3352 );
nor ( n4386 , n4384 , n4385 );
not ( n4387 , n4110 );
nand ( n4388 , n4387 , n4030 );
and ( n4389 , n4027 , n4095 );
nor ( n4390 , n4389 , n4107 );
or ( n4391 , n4388 , n4390 );
nand ( n4392 , n4388 , n4390 );
nand ( n4393 , n4391 , n4392 , n4130 );
not ( n4394 , n4162 );
nand ( n4395 , n4394 , n4159 );
and ( n4396 , n4179 , n4242 );
nor ( n4397 , n4396 , n4157 );
or ( n4398 , n4395 , n4397 );
nand ( n4399 , n4395 , n4397 );
nand ( n4400 , n4398 , n4399 , n4257 );
nand ( n4401 , n227 , n4004 );
nand ( n4402 , n4386 , n4393 , n4400 , n4401 );
and ( n4403 , n500 , n4138 );
and ( n4404 , n75 , n3352 );
nor ( n4405 , n4403 , n4404 );
not ( n4406 , n4027 );
nor ( n4407 , n4406 , n4107 );
or ( n4408 , n4407 , n4095 );
nand ( n4409 , n4407 , n4095 );
nand ( n4410 , n4408 , n4409 , n4130 );
not ( n4411 , n4179 );
nor ( n4412 , n4411 , n4157 );
or ( n4413 , n4412 , n4242 );
nand ( n4414 , n4412 , n4242 );
nand ( n4415 , n4413 , n4414 , n4257 );
nand ( n4416 , n228 , n4004 );
nand ( n4417 , n4405 , n4410 , n4415 , n4416 );
and ( n4418 , n1258 , n4138 );
and ( n4419 , n67 , n3352 );
nor ( n4420 , n4418 , n4419 );
not ( n4421 , n4045 );
nor ( n4422 , n4421 , n4034 );
nor ( n4423 , n4041 , n4093 );
or ( n4424 , n4032 , n4423 );
nand ( n4425 , n4424 , n4043 );
or ( n4426 , n4422 , n4425 );
nand ( n4427 , n4422 , n4425 );
nand ( n4428 , n4426 , n4427 , n4130 );
not ( n4429 , n4192 );
nor ( n4430 , n4429 , n4182 );
nor ( n4431 , n4188 , n4240 );
or ( n4432 , n4181 , n4431 );
nand ( n4433 , n4432 , n4190 );
or ( n4434 , n4430 , n4433 );
nand ( n4435 , n4430 , n4433 );
nand ( n4436 , n4434 , n4435 , n4257 );
nand ( n4437 , n229 , n4004 );
nand ( n4438 , n4420 , n4428 , n4436 , n4437 );
not ( n4439 , n1215 );
and ( n4440 , n4439 , n4138 );
nor ( n4441 , n4440 , n3117 );
not ( n4442 , n4032 );
nand ( n4443 , n4442 , n4043 );
or ( n4444 , n4443 , n4423 );
nand ( n4445 , n4443 , n4423 );
nand ( n4446 , n4444 , n4445 , n4130 );
not ( n4447 , n4181 );
nand ( n4448 , n4447 , n4190 );
or ( n4449 , n4448 , n4431 );
nand ( n4450 , n4448 , n4431 );
nand ( n4451 , n4449 , n4450 , n4257 );
nand ( n4452 , n230 , n4004 );
nand ( n4453 , n4441 , n4446 , n4451 , n4452 );
and ( n4454 , n4037 , n4138 );
nor ( n4455 , n4454 , n3274 );
not ( n4456 , n4040 );
nor ( n4457 , n4456 , n4038 );
or ( n4458 , n4092 , n4091 );
nand ( n4459 , n4458 , n4036 );
or ( n4460 , n4457 , n4459 );
nand ( n4461 , n4457 , n4459 );
nand ( n4462 , n4460 , n4461 , n4130 );
not ( n4463 , n4187 );
nor ( n4464 , n4463 , n4185 );
or ( n4465 , n4239 , n4238 );
nand ( n4466 , n4465 , n4184 );
or ( n4467 , n4464 , n4466 );
nand ( n4468 , n4464 , n4466 );
nand ( n4469 , n4467 , n4468 , n4257 );
nand ( n4470 , n231 , n4004 );
nand ( n4471 , n4455 , n4462 , n4469 , n4470 );
and ( n4472 , n967 , n4138 );
not ( n4473 , n3353 );
nor ( n4474 , n4472 , n4473 );
not ( n4475 , n4092 );
nand ( n4476 , n4475 , n4036 );
or ( n4477 , n4476 , n4091 );
nand ( n4478 , n4476 , n4091 );
nand ( n4479 , n4477 , n4478 , n4130 );
not ( n4480 , n4239 );
nand ( n4481 , n4480 , n4184 );
or ( n4482 , n4481 , n4238 );
nand ( n4483 , n4481 , n4238 );
nand ( n4484 , n4482 , n4483 , n4257 );
nand ( n4485 , n232 , n4004 );
nand ( n4486 , n4474 , n4479 , n4484 , n4485 );
and ( n4487 , n233 , n4004 );
nor ( n4488 , n4487 , n3391 );
not ( n4489 , n4066 );
nor ( n4490 , n4489 , n4050 );
nor ( n4491 , n4063 , n4089 );
or ( n4492 , n4054 , n4491 );
nand ( n4493 , n4492 , n4048 );
or ( n4494 , n4490 , n4493 );
nand ( n4495 , n4490 , n4493 );
nand ( n4496 , n4494 , n4495 , n4130 );
not ( n4497 , n1300 );
nand ( n4498 , n4497 , n4138 );
not ( n4499 , n4232 );
nor ( n4500 , n4499 , n4197 );
nor ( n4501 , n4236 , n4229 );
or ( n4502 , n4200 , n4501 );
nand ( n4503 , n4502 , n4195 );
or ( n4504 , n4500 , n4503 );
nand ( n4505 , n4500 , n4503 );
nand ( n4506 , n4504 , n4505 , n4257 );
nand ( n4507 , n4488 , n4496 , n4498 , n4506 );
and ( n4508 , n234 , n4004 );
nor ( n4509 , n4508 , n3588 );
not ( n4510 , n4054 );
nand ( n4511 , n4510 , n4048 );
or ( n4512 , n4511 , n4491 );
nand ( n4513 , n4511 , n4491 );
nand ( n4514 , n4512 , n4513 , n4130 );
nand ( n4515 , n1270 , n4138 );
not ( n4516 , n4195 );
nor ( n4517 , n4516 , n4200 );
not ( n4518 , n4517 );
not ( n4519 , n4501 );
or ( n4520 , n4518 , n4519 );
or ( n4521 , n4517 , n4501 );
nand ( n4522 , n4520 , n4521 );
nand ( n4523 , n4522 , n4257 );
nand ( n4524 , n4509 , n4514 , n4515 , n4523 );
and ( n4525 , n235 , n4004 );
nor ( n4526 , n4525 , n3637 );
nand ( n4527 , n4062 , n4059 );
nor ( n4528 , n4056 , n4088 );
or ( n4529 , n4527 , n4528 );
nand ( n4530 , n4527 , n4528 );
nand ( n4531 , n4529 , n4530 , n4130 );
not ( n4532 , n1319 );
nand ( n4533 , n4532 , n4138 );
not ( n4534 , n4203 );
nand ( n4535 , n4534 , n4235 );
not ( n4536 , n4535 );
nand ( n4537 , n4233 , n4228 );
not ( n4538 , n4537 );
or ( n4539 , n4536 , n4538 );
or ( n4540 , n4535 , n4537 );
nand ( n4541 , n4539 , n4540 );
nand ( n4542 , n4541 , n4257 );
nand ( n4543 , n4526 , n4531 , n4533 , n4542 );
nor ( n4544 , n4056 , n4067 );
not ( n4545 , n4087 );
nand ( n4546 , n4544 , n4545 );
not ( n4547 , n4544 );
nand ( n4548 , n4547 , n4087 );
and ( n4549 , n4546 , n4548 , n4130 );
not ( n4550 , n6 );
and ( n4551 , n147 , n2865 );
and ( n4552 , n148 , n4126 );
nor ( n4553 , n4551 , n4552 );
and ( n4554 , n4550 , n4553 );
not ( n4555 , n6 );
nor ( n4556 , n4555 , n4553 );
nor ( n4557 , n4554 , n4556 , n3870 );
nor ( n4558 , n4549 , n4557 );
nand ( n4559 , n236 , n4004 );
nand ( n4560 , n4233 , n4204 );
not ( n4561 , n4560 );
nand ( n4562 , n4561 , n4227 );
not ( n4563 , n4227 );
nand ( n4564 , n4560 , n4563 );
and ( n4565 , n4562 , n4564 , n4257 );
and ( n4566 , n1334 , n4138 );
nor ( n4567 , n4565 , n4566 );
nand ( n4568 , n4558 , n4559 , n3663 , n4567 );
and ( n4569 , n237 , n4004 );
nor ( n4570 , n4569 , n3718 );
not ( n4571 , n4069 );
nor ( n4572 , n4571 , n4086 );
or ( n4573 , n4572 , n4083 );
nand ( n4574 , n4572 , n4083 );
nand ( n4575 , n4573 , n4574 , n4130 );
not ( n4576 , n1388 );
nand ( n4577 , n4576 , n4138 );
nand ( n4578 , n4226 , n4205 );
not ( n4579 , n4578 );
not ( n4580 , n4223 );
or ( n4581 , n4579 , n4580 );
or ( n4582 , n4578 , n4223 );
nand ( n4583 , n4581 , n4582 );
nand ( n4584 , n4583 , n4257 );
nand ( n4585 , n4570 , n4575 , n4577 , n4584 );
and ( n4586 , n238 , n4004 );
nor ( n4587 , n4586 , n4557 );
not ( n4588 , n4222 );
nor ( n4589 , n4588 , n4207 );
not ( n4590 , n4589 );
nand ( n4591 , n4220 , n4590 );
nand ( n4592 , n4219 , n4589 );
and ( n4593 , n4591 , n4592 , n4257 );
not ( n4594 , n154 );
nor ( n4595 , n4594 , n161 );
nor ( n4596 , n4593 , n4595 );
nand ( n4597 , n567 , n4138 );
not ( n4598 , n4070 );
nand ( n4599 , n4598 , n4082 );
or ( n4600 , n4080 , n4599 );
nand ( n4601 , n4080 , n4599 );
nand ( n4602 , n4600 , n4601 , n4130 );
nand ( n4603 , n4587 , n4596 , n4597 , n4602 );
and ( n4604 , n239 , n4004 );
and ( n4605 , n150 , n3352 );
nor ( n4606 , n4604 , n4605 );
not ( n4607 , n651 );
or ( n4608 , n4078 , n4607 );
nand ( n4609 , n4608 , n4079 , n4130 );
nand ( n4610 , n4607 , n4138 );
or ( n4611 , n4217 , n4607 );
nand ( n4612 , n4611 , n4218 , n4257 );
nand ( n4613 , n4606 , n4609 , n4610 , n4612 );
and ( n4614 , n240 , n4004 );
and ( n4615 , n146 , n3352 );
nor ( n4616 , n4614 , n4615 );
not ( n4617 , n6 );
or ( n4618 , n4617 , n3821 );
or ( n4619 , n6 , n148 );
nand ( n4620 , n4618 , n4619 , n4130 );
nand ( n4621 , n6 , n4138 );
not ( n4622 , n6 );
or ( n4623 , n4622 , n1446 );
or ( n4624 , n6 , n147 );
nand ( n4625 , n4623 , n4624 , n4257 );
nand ( n4626 , n4616 , n4620 , n4621 , n4625 );
or ( n4627 , n3904 , n966 );
not ( n4628 , n3883 );
nand ( n4629 , n216 , n4628 );
nand ( n4630 , n4627 , n4629 );
not ( n4631 , n217 );
not ( n4632 , n3904 );
or ( n4633 , n4631 , n4632 );
or ( n4634 , n3909 , n2989 );
nand ( n4635 , n4633 , n4634 );
not ( n4636 , n3871 );
or ( n4637 , n4636 , n3448 );
nand ( n4638 , n219 , n4628 );
nand ( n4639 , n4637 , n4638 );
not ( n4640 , n3458 );
or ( n4641 , n3904 , n4640 );
nand ( n4642 , n241 , n4628 );
nand ( n4643 , n4641 , n4642 );
or ( n4644 , n4636 , n1404 );
not ( n4645 , n3883 );
nand ( n4646 , n242 , n4645 );
nand ( n4647 , n4644 , n4646 );
not ( n4648 , n3319 );
or ( n4649 , n4636 , n4648 );
nand ( n4650 , n243 , n4628 );
nand ( n4651 , n4649 , n4650 );
or ( n4652 , n4636 , n3673 );
nand ( n4653 , n244 , n4645 );
nand ( n4654 , n4652 , n4653 );
or ( n4655 , n4636 , n2209 );
nand ( n4656 , n245 , n4645 );
nand ( n4657 , n4655 , n4656 );
or ( n4658 , n3904 , n1331 );
not ( n4659 , n3883 );
nand ( n4660 , n220 , n4659 );
nand ( n4661 , n4658 , n4660 );
not ( n4662 , n160 );
not ( n4663 , n3339 );
or ( n4664 , n4662 , n4663 );
nand ( n4665 , n4664 , n3558 );
not ( n4666 , n1510 );
and ( n4667 , n739 , n2924 );
nor ( n4668 , n4667 , n714 );
or ( n4669 , n4666 , n4668 );
nand ( n4670 , n4669 , n161 );
not ( n4671 , n159 );
not ( n4672 , n3339 );
or ( n4673 , n4671 , n4672 );
or ( n4674 , n3339 , n3513 );
nand ( n4675 , n4673 , n4674 );
not ( n4676 , n187 );
not ( n4677 , n3352 );
or ( n4678 , n4676 , n4677 );
not ( n4679 , n835 );
or ( n4680 , n3352 , n4679 );
nand ( n4681 , n4678 , n4680 );
not ( n4682 , n189 );
not ( n4683 , n3352 );
or ( n4684 , n4682 , n4683 );
or ( n4685 , n3352 , n856 );
nand ( n4686 , n4684 , n4685 );
not ( n4687 , n198 );
not ( n4688 , n3352 );
or ( n4689 , n4687 , n4688 );
or ( n4690 , n3352 , n2015 );
nand ( n4691 , n4689 , n4690 );
not ( n4692 , n193 );
not ( n4693 , n3352 );
or ( n4694 , n4692 , n4693 );
or ( n4695 , n3352 , n2874 );
nand ( n4696 , n4694 , n4695 );
not ( n4697 , n188 );
not ( n4698 , n3352 );
or ( n4699 , n4697 , n4698 );
or ( n4700 , n3352 , n2860 );
nand ( n4701 , n4699 , n4700 );
not ( n4702 , n192 );
not ( n4703 , n3352 );
or ( n4704 , n4702 , n4703 );
or ( n4705 , n3352 , n987 );
nand ( n4706 , n4704 , n4705 );
not ( n4707 , n200 );
not ( n4708 , n3352 );
or ( n4709 , n4707 , n4708 );
or ( n4710 , n3352 , n1921 );
nand ( n4711 , n4709 , n4710 );
not ( n4712 , n186 );
not ( n4713 , n3352 );
or ( n4714 , n4712 , n4713 );
or ( n4715 , n3352 , n1257 );
nand ( n4716 , n4714 , n4715 );
not ( n4717 , n182 );
not ( n4718 , n3352 );
or ( n4719 , n4717 , n4718 );
or ( n4720 , n3352 , n1126 );
nand ( n4721 , n4719 , n4720 );
not ( n4722 , n201 );
not ( n4723 , n3352 );
or ( n4724 , n4722 , n4723 );
or ( n4725 , n3352 , n610 );
nand ( n4726 , n4724 , n4725 );
not ( n4727 , n184 );
not ( n4728 , n3352 );
or ( n4729 , n4727 , n4728 );
or ( n4730 , n3352 , n1193 );
nand ( n4731 , n4729 , n4730 );
not ( n4732 , n165 );
not ( n4733 , n3352 );
or ( n4734 , n4732 , n4733 );
or ( n4735 , n3352 , n1300 );
nand ( n4736 , n4734 , n4735 );
not ( n4737 , n183 );
not ( n4738 , n3352 );
or ( n4739 , n4737 , n4738 );
or ( n4740 , n3352 , n1111 );
nand ( n4741 , n4739 , n4740 );
or ( n4742 , n3352 , n4026 );
or ( n4743 , n1182 , n161 );
nand ( n4744 , n4742 , n4743 );
not ( n4745 , n162 );
not ( n4746 , n3352 );
or ( n4747 , n4745 , n4746 );
or ( n4748 , n3352 , n1215 );
nand ( n4749 , n4747 , n4748 );
or ( n4750 , n3352 , n599 );
or ( n4751 , n1015 , n161 );
nand ( n4752 , n4750 , n4751 );
not ( n4753 , n164 );
not ( n4754 , n3352 );
or ( n4755 , n4753 , n4754 );
or ( n4756 , n3352 , n533 );
nand ( n4757 , n4755 , n4756 );
and ( n4758 , n3352 , n190 );
not ( n4759 , n3352 );
and ( n4760 , n4759 , n2868 );
or ( n4761 , n4758 , n4760 );
endmodule
