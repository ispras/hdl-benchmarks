module mul_21_11_11(a, b, c);
  input [20:0] a;
  input [10:0] b;
  output [10:0] c;
  assign c = a * b;
endmodule
