// IWLS benchmark module "MultiplierB_32" printed on Wed May 29 22:12:35 2002
module MultiplierB_32(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \30 , \31 , \32 , \33 , \98 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ;
output
  \98 ;
reg
  \2 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ,
  \67 ,
  \68 ,
  \69 ,
  \70 ,
  \71 ,
  \72 ,
  \73 ,
  \74 ,
  \75 ,
  \76 ,
  \77 ,
  \78 ,
  \79 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ;
wire
  \370 ,
  \371 ,
  \375 ,
  \376 ,
  \377 ,
  \[145] ,
  \383 ,
  \386 ,
  \389 ,
  \[146] ,
  \392 ,
  \395 ,
  \398 ,
  \[147] ,
  \[148] ,
  \[64] ,
  \[149] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \401 ,
  \404 ,
  \407 ,
  \410 ,
  \413 ,
  \416 ,
  \419 ,
  \422 ,
  \425 ,
  \428 ,
  \[150] ,
  \431 ,
  \434 ,
  \437 ,
  \[151] ,
  \440 ,
  \443 ,
  \446 ,
  \449 ,
  \[152] ,
  \452 ,
  \455 ,
  \458 ,
  \[153] ,
  \461 ,
  \464 ,
  \467 ,
  \[154] ,
  \[70] ,
  \470 ,
  \[155] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[78] ,
  \[79] ,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[100] ,
  \[99] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[108] ,
  \[109] ,
  \[110] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \[116] ,
  \[117] ,
  \[118] ,
  \[119] ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \[126] ,
  \[127] ,
  \[128] ,
  \[129] ,
  \226 ,
  \[130] ,
  \230 ,
  \231 ,
  \235 ,
  \236 ,
  \[131] ,
  \240 ,
  \241 ,
  \245 ,
  \246 ,
  \[132] ,
  \250 ,
  \251 ,
  \255 ,
  \256 ,
  \[133] ,
  \260 ,
  \261 ,
  \265 ,
  \266 ,
  \[134] ,
  \270 ,
  \271 ,
  \275 ,
  \276 ,
  \[135] ,
  \280 ,
  \281 ,
  \285 ,
  \286 ,
  \[136] ,
  \290 ,
  \291 ,
  \295 ,
  \296 ,
  \[137] ,
  \[138] ,
  \[139] ,
  \300 ,
  \301 ,
  \305 ,
  \306 ,
  \310 ,
  \311 ,
  \315 ,
  \316 ,
  \320 ,
  \321 ,
  \325 ,
  \326 ,
  \[140] ,
  \330 ,
  \331 ,
  \335 ,
  \336 ,
  \[141] ,
  \340 ,
  \341 ,
  \345 ,
  \346 ,
  \[142] ,
  \350 ,
  \351 ,
  \355 ,
  \356 ,
  \[143] ,
  \360 ,
  \361 ,
  \365 ,
  \366 ,
  \[144] ;
assign
  \370  = (~\366  & \467 ) | (~\467  & \94 ),
  \371  = (~\[155]  & ~\470 ) | (\[155]  & \470 ),
  \375  = (~\371  & \470 ) | (~\470  & \95 ),
  \376  = (~\377  & (\33  & \1 )) | (~\377  & \2 ),
  \377  = \2  & (\33  & \1 ),
  \[145]  = ~\22  | ~\1 ,
  \383  = (~\36  & \66 ) | (\36  & ~\66 ),
  \386  = (~\37  & \67 ) | (\37  & ~\67 ),
  \389  = (~\38  & \68 ) | (\38  & ~\68 ),
  \[146]  = ~\23  | ~\1 ,
  \392  = (~\39  & \69 ) | (\39  & ~\69 ),
  \395  = (~\40  & \70 ) | (\40  & ~\70 ),
  \398  = (~\41  & \71 ) | (\41  & ~\71 ),
  \[147]  = ~\24  | ~\1 ,
  \[148]  = ~\25  | ~\1 ,
  \[64]  = \231 ,
  \[149]  = ~\26  | ~\1 ,
  \[65]  = \236 ,
  \[66]  = \241 ,
  \[67]  = \246 ,
  \[68]  = \251 ,
  \[69]  = \256 ,
  \401  = (~\42  & \72 ) | (\42  & ~\72 ),
  \404  = (~\43  & \73 ) | (\43  & ~\73 ),
  \407  = (~\44  & \74 ) | (\44  & ~\74 ),
  \410  = (~\45  & \75 ) | (\45  & ~\75 ),
  \413  = (~\46  & \76 ) | (\46  & ~\76 ),
  \416  = (~\47  & \77 ) | (\47  & ~\77 ),
  \419  = (~\48  & \78 ) | (\48  & ~\78 ),
  \422  = (~\49  & \79 ) | (\49  & ~\79 ),
  \425  = (~\50  & \80 ) | (\50  & ~\80 ),
  \428  = (~\51  & \81 ) | (\51  & ~\81 ),
  \[150]  = ~\27  | ~\1 ,
  \431  = (~\52  & \82 ) | (\52  & ~\82 ),
  \434  = (~\53  & \83 ) | (\53  & ~\83 ),
  \437  = (~\54  & \84 ) | (\54  & ~\84 ),
  \[151]  = ~\28  | ~\1 ,
  \440  = (~\55  & \85 ) | (\55  & ~\85 ),
  \443  = (~\56  & \86 ) | (\56  & ~\86 ),
  \446  = (~\57  & \87 ) | (\57  & ~\87 ),
  \449  = (~\58  & \88 ) | (\58  & ~\88 ),
  \[152]  = ~\29  | ~\1 ,
  \452  = (~\59  & \89 ) | (\59  & ~\89 ),
  \455  = (~\60  & \90 ) | (\60  & ~\90 ),
  \458  = (~\61  & \91 ) | (\61  & ~\91 ),
  \[153]  = ~\30  | ~\1 ,
  \461  = (~\62  & \92 ) | (\62  & ~\92 ),
  \464  = (~\63  & \93 ) | (\63  & ~\93 ),
  \467  = (~\64  & \94 ) | (\64  & ~\94 ),
  \[154]  = ~\31  | ~\1 ,
  \[70]  = \261 ,
  \470  = (~\65  & \95 ) | (\65  & ~\95 ),
  \[155]  = ~\32  | ~\1 ,
  \[71]  = \266 ,
  \[72]  = \271 ,
  \[73]  = \276 ,
  \[74]  = \281 ,
  \[75]  = \286 ,
  \[76]  = \291 ,
  \[77]  = \296 ,
  \[78]  = \301 ,
  \[79]  = \306 ,
  \[80]  = \311 ,
  \[81]  = \316 ,
  \[82]  = \321 ,
  \[83]  = \326 ,
  \[84]  = \331 ,
  \[85]  = \336 ,
  \[86]  = \341 ,
  \[87]  = \346 ,
  \[88]  = \351 ,
  \[89]  = \356 ,
  \[90]  = \361 ,
  \[91]  = \366 ,
  \[92]  = \371 ,
  \[93]  = \376 ,
  \[94]  = \230 ,
  \[95]  = \235 ,
  \[96]  = \240 ,
  \[97]  = \245 ,
  \[98]  = \250 ,
  \[100]  = \260 ,
  \[99]  = \255 ,
  \[101]  = \265 ,
  \[102]  = \270 ,
  \[103]  = \275 ,
  \98  = \226 ,
  \[104]  = \280 ,
  \[105]  = \285 ,
  \[106]  = \290 ,
  \[107]  = \295 ,
  \[108]  = \300 ,
  \[109]  = \305 ,
  \[110]  = \310 ,
  \[111]  = \315 ,
  \[112]  = \320 ,
  \[113]  = \325 ,
  \[114]  = \330 ,
  \[115]  = \335 ,
  \[116]  = \340 ,
  \[117]  = \345 ,
  \[118]  = \350 ,
  \[119]  = \355 ,
  \[120]  = \360 ,
  \[121]  = \365 ,
  \[122]  = \370 ,
  \[123]  = \375 ,
  \[124]  = \377 ,
  \[126]  = ~\3  | ~\1 ,
  \[127]  = ~\4  | ~\1 ,
  \[128]  = ~\5  | ~\1 ,
  \[129]  = ~\6  | ~\1 ,
  \226  = (~\[126]  & ~\383 ) | (\[126]  & \383 ),
  \[130]  = ~\7  | ~\1 ,
  \230  = (~\226  & \383 ) | (~\383  & \66 ),
  \231  = (~\[127]  & ~\386 ) | (\[127]  & \386 ),
  \235  = (~\231  & \386 ) | (~\386  & \67 ),
  \236  = (~\[128]  & ~\389 ) | (\[128]  & \389 ),
  \[131]  = ~\8  | ~\1 ,
  \240  = (~\236  & \389 ) | (~\389  & \68 ),
  \241  = (~\[129]  & ~\392 ) | (\[129]  & \392 ),
  \245  = (~\241  & \392 ) | (~\392  & \69 ),
  \246  = (~\[130]  & ~\395 ) | (\[130]  & \395 ),
  \[132]  = ~\9  | ~\1 ,
  \250  = (~\246  & \395 ) | (~\395  & \70 ),
  \251  = (~\[131]  & ~\398 ) | (\[131]  & \398 ),
  \255  = (~\251  & \398 ) | (~\398  & \71 ),
  \256  = (~\[132]  & ~\401 ) | (\[132]  & \401 ),
  \[133]  = ~\10  | ~\1 ,
  \260  = (~\256  & \401 ) | (~\401  & \72 ),
  \261  = (~\[133]  & ~\404 ) | (\[133]  & \404 ),
  \265  = (~\261  & \404 ) | (~\404  & \73 ),
  \266  = (~\[134]  & ~\407 ) | (\[134]  & \407 ),
  \[134]  = ~\11  | ~\1 ,
  \270  = (~\266  & \407 ) | (~\407  & \74 ),
  \271  = (~\[135]  & ~\410 ) | (\[135]  & \410 ),
  \275  = (~\271  & \410 ) | (~\410  & \75 ),
  \276  = (~\[136]  & ~\413 ) | (\[136]  & \413 ),
  \[135]  = ~\12  | ~\1 ,
  \280  = (~\276  & \413 ) | (~\413  & \76 ),
  \281  = (~\[137]  & ~\416 ) | (\[137]  & \416 ),
  \285  = (~\281  & \416 ) | (~\416  & \77 ),
  \286  = (~\[138]  & ~\419 ) | (\[138]  & \419 ),
  \[136]  = ~\13  | ~\1 ,
  \290  = (~\286  & \419 ) | (~\419  & \78 ),
  \291  = (~\[139]  & ~\422 ) | (\[139]  & \422 ),
  \295  = (~\291  & \422 ) | (~\422  & \79 ),
  \296  = (~\[140]  & ~\425 ) | (\[140]  & \425 ),
  \[137]  = ~\14  | ~\1 ,
  \[138]  = ~\15  | ~\1 ,
  \[139]  = ~\16  | ~\1 ,
  \300  = (~\296  & \425 ) | (~\425  & \80 ),
  \301  = (~\[141]  & ~\428 ) | (\[141]  & \428 ),
  \305  = (~\301  & \428 ) | (~\428  & \81 ),
  \306  = (~\[142]  & ~\431 ) | (\[142]  & \431 ),
  \310  = (~\306  & \431 ) | (~\431  & \82 ),
  \311  = (~\[143]  & ~\434 ) | (\[143]  & \434 ),
  \315  = (~\311  & \434 ) | (~\434  & \83 ),
  \316  = (~\[144]  & ~\437 ) | (\[144]  & \437 ),
  \320  = (~\316  & \437 ) | (~\437  & \84 ),
  \321  = (~\[145]  & ~\440 ) | (\[145]  & \440 ),
  \325  = (~\321  & \440 ) | (~\440  & \85 ),
  \326  = (~\[146]  & ~\443 ) | (\[146]  & \443 ),
  \[140]  = ~\17  | ~\1 ,
  \330  = (~\326  & \443 ) | (~\443  & \86 ),
  \331  = (~\[147]  & ~\446 ) | (\[147]  & \446 ),
  \335  = (~\331  & \446 ) | (~\446  & \87 ),
  \336  = (~\[148]  & ~\449 ) | (\[148]  & \449 ),
  \[141]  = ~\18  | ~\1 ,
  \340  = (~\336  & \449 ) | (~\449  & \88 ),
  \341  = (~\[149]  & ~\452 ) | (\[149]  & \452 ),
  \345  = (~\341  & \452 ) | (~\452  & \89 ),
  \346  = (~\[150]  & ~\455 ) | (\[150]  & \455 ),
  \[142]  = ~\19  | ~\1 ,
  \350  = (~\346  & \455 ) | (~\455  & \90 ),
  \351  = (~\[151]  & ~\458 ) | (\[151]  & \458 ),
  \355  = (~\351  & \458 ) | (~\458  & \91 ),
  \356  = (~\[152]  & ~\461 ) | (\[152]  & \461 ),
  \[143]  = ~\20  | ~\1 ,
  \360  = (~\356  & \461 ) | (~\461  & \92 ),
  \361  = (~\[153]  & ~\464 ) | (\[153]  & \464 ),
  \365  = (~\361  & \464 ) | (~\464  & \93 ),
  \366  = (~\[154]  & ~\467 ) | (\[154]  & \467 ),
  \[144]  = ~\21  | ~\1 ;
always begin
  \2  = \[64] ;
  \36  = \[65] ;
  \37  = \[66] ;
  \38  = \[67] ;
  \39  = \[68] ;
  \40  = \[69] ;
  \41  = \[70] ;
  \42  = \[71] ;
  \43  = \[72] ;
  \44  = \[73] ;
  \45  = \[74] ;
  \46  = \[75] ;
  \47  = \[76] ;
  \48  = \[77] ;
  \49  = \[78] ;
  \50  = \[79] ;
  \51  = \[80] ;
  \52  = \[81] ;
  \53  = \[82] ;
  \54  = \[83] ;
  \55  = \[84] ;
  \56  = \[85] ;
  \57  = \[86] ;
  \58  = \[87] ;
  \59  = \[88] ;
  \60  = \[89] ;
  \61  = \[90] ;
  \62  = \[91] ;
  \63  = \[92] ;
  \64  = \[93] ;
  \65  = \[94] ;
  \66  = \[95] ;
  \67  = \[96] ;
  \68  = \[97] ;
  \69  = \[98] ;
  \70  = \[99] ;
  \71  = \[100] ;
  \72  = \[101] ;
  \73  = \[102] ;
  \74  = \[103] ;
  \75  = \[104] ;
  \76  = \[105] ;
  \77  = \[106] ;
  \78  = \[107] ;
  \79  = \[108] ;
  \80  = \[109] ;
  \81  = \[110] ;
  \82  = \[111] ;
  \83  = \[112] ;
  \84  = \[113] ;
  \85  = \[114] ;
  \86  = \[115] ;
  \87  = \[116] ;
  \88  = \[117] ;
  \89  = \[118] ;
  \90  = \[119] ;
  \91  = \[120] ;
  \92  = \[121] ;
  \93  = \[122] ;
  \94  = \[123] ;
  \95  = \[124] ;
end
initial begin
  \2  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
  \49  = 0;
  \50  = 0;
  \51  = 0;
  \52  = 0;
  \53  = 0;
  \54  = 0;
  \55  = 0;
  \56  = 0;
  \57  = 0;
  \58  = 0;
  \59  = 0;
  \60  = 0;
  \61  = 0;
  \62  = 0;
  \63  = 0;
  \64  = 0;
  \65  = 0;
  \66  = 0;
  \67  = 0;
  \68  = 0;
  \69  = 0;
  \70  = 0;
  \71  = 0;
  \72  = 0;
  \73  = 0;
  \74  = 0;
  \75  = 0;
  \76  = 0;
  \77  = 0;
  \78  = 0;
  \79  = 0;
  \80  = 0;
  \81  = 0;
  \82  = 0;
  \83  = 0;
  \84  = 0;
  \85  = 0;
  \86  = 0;
  \87  = 0;
  \88  = 0;
  \89  = 0;
  \90  = 0;
  \91  = 0;
  \92  = 0;
  \93  = 0;
  \94  = 0;
  \95  = 0;
end
endmodule

