//NOTE: no-implementation module stub

`define N 0

module DSP_CORE (
    input wire BGn,
    input wire BMSn,
    input wire CLKO,
    input wire [0:0] CMAinx,
    input wire CMSn,
    input wire CM_cs,
    input wire CM_oe,
    input wire [0:0] CM_rd0,
    input wire [0:0] CM_rd1,
    input wire [0:0] CM_rd2,
    input wire [0:0] CM_rd3,
    input wire [0:0] CM_rd4,
    input wire [0:0] CM_rd5,
    input wire [0:0] CM_rd6,
    input wire [0:0] CM_rd7,
    input wire [0:0] CM_rdm,
    input wire [0:0] CM_wd,
    input wire CM_web,
    input wire CMo_cs0,
    input wire CMo_cs1,
    input wire CMo_cs2,
    input wire CMo_cs3,
    input wire CMo_cs4,
    input wire CMo_cs5,
    input wire CMo_cs6,
    input wire CMo_cs7,
    input wire CMo_oe0,
    input wire CMo_oe1,
    input wire CMo_oe2,
    input wire CMo_oe3,
    input wire CMo_oe4,
    input wire CMo_oe5,
    input wire CMo_oe6,
    input wire CMo_oe7,
    input wire DMAinx,
    input wire DMSn,
    input wire DM_cs,
    input wire DM_oe,
    input wire [0:0] DM_rd0,
    input wire [0:0] DM_rd1,
    input wire [0:0] DM_rd2,
    input wire [0:0] DM_rd3,
    input wire [0:0] DM_rd4,
    input wire [0:0] DM_rd5,
    input wire [0:0] DM_rd6,
    input wire [0:0] DM_rd7,
    input wire [0:0] DM_rdm,
    input wire [0:0] DM_wd,
    input wire DMo_cs0,
    input wire DMo_cs1,
    input wire DMo_cs2,
    input wire DMo_cs3,
    input wire DMo_cs4,
    input wire DMo_cs5,
    input wire DMo_cs6,
    input wire DMo_cs7,
    input wire DMo_oe0,
    input wire DMo_oe1,
    input wire DMo_oe2,
    input wire DMo_oe3,
    input wire DMo_oe4,
    input wire DMo_oe5,
    input wire DMo_oe6,
    input wire DMo_oe7,
    input wire DMo_web,
    input wire DSPCLK_cm0,
    input wire DSPCLK_cm1,
    input wire DSPCLK_cm2,
    input wire DSPCLK_dm0,
    input wire DSPCLK_dm1,
    input wire DSPCLK_dm2,
    input wire DSPCLK_pm0,
    input wire DSPCLK_pm1,
    input wire DSPCLK_pm2,
    input wire [0:0] EA_do,
    input wire EA_oe,
    input wire ECMA_EN,
    input wire ECMSn,
    input wire [0:0] ED_do,
    input wire ED_oe_14_8,
    input wire ED_oe_15,
    input wire ED_oe_7_0,
    input wire IACKn,
    input wire [0:0] IAD_do,
    input wire IAD_oe,
    input wire [0:0] IDo,
    input wire IDoe,
    input wire IOSn,
    input wire IRFS0,
    input wire IRFS1,
    input wire ISCLK0,
    input wire ISCLK1,
    input wire ITFS0,
    input wire ITFS1,
    input wire PIO_oe,
    input wire [0:0] PIO_out,
    input wire PMAinx,
    input wire PMSn,
    input wire PM_bdry_sel,
    input wire [0:0] PM_rd0,
    input wire [0:0] PM_rd1,
    input wire [0:0] PM_rd2,
    input wire [0:0] PM_rd3,
    input wire [0:0] PM_rd4,
    input wire [0:0] PM_rd5,
    input wire [0:0] PM_rd6,
    input wire [0:0] PM_rd7,
    input wire [0:0] PM_wd,
    input wire PMo_cs0,
    input wire PMo_cs1,
    input wire PMo_cs2,
    input wire PMo_cs3,
    input wire PMo_cs4,
    input wire PMo_cs5,
    input wire PMo_cs6,
    input wire PMo_cs7,
    input wire PMo_oe0,
    input wire PMo_oe1,
    input wire PMo_oe2,
    input wire PMo_oe3,
    input wire PMo_oe4,
    input wire PMo_oe5,
    input wire PMo_oe6,
    input wire PMo_oe7,
    input wire PMo_web,
    input wire PWDACK,
    input wire RDn,
    input wire RFS0,
    input wire RFS1,
    input wire SCANIN1,
    input wire SCANIN2,
    input wire SCANIN3,
    input wire SCANIN4,
    input wire SCANIN5,
    input wire SCANIN6,
    input wire SCANIN7,
    input wire SCANIN8,
    input wire SCAN_ENABLE,
    input wire SCAN_TEST,
    input wire SCLK0,
    input wire SCLK1,
    input wire [0:0] TD0,
    input wire [0:0] TD1,
    input wire TFS0,
    input wire TFS1,
    input wire T_BMODE,
    input wire T_BRn,
    input wire T_CLKI_OSC,
    input wire T_CLKI_PLL,
    input wire T_EA,
    input wire T_ED,
    input wire T_GOICE,
    input wire T_IAD,
    input wire T_IAL,
    input wire T_ICE_RSTn,
    input wire T_ICK,
    input wire T_ID,
    input wire T_IMS,
    input wire T_IRDn,
    input wire T_IRQ0n,
    input wire T_IRQ1n,
    input wire T_IRQ2n,
    input wire T_IRQE0n,
    input wire T_IRQE1n,
    input wire T_IRQL1n,
    input wire T_ISn,
    input wire T_IWRn,
    input wire T_MMAP,
    input wire T_PIOin,
    input wire T_PWDn,
    input wire [0:0] T_RD0,
    input wire [0:0] T_RD1,
    input wire T_RFS0,
    input wire T_RFS1,
    input wire T_RSTn,
    input wire T_SCLK0,
    input wire T_SCLK1,
    input wire T_Sel_PLL,
    input wire T_TFS0,
    input wire T_TFS1,
    input wire T_TMODE,
    input wire WRn,
    input wire XTALoffn,
    input wire DSPCLK_insert_buf_i,

    output wire DSPCLK_insert_buf_o,
    output wire SCANOUT1,
    output wire SCANOUT2,
    output wire SCANOUT3,
    output wire SCANOUT4,
    output wire SCANOUT5,
    output wire SCANOUT6,
    output wire SCANOUT7,
    output wire SCANOUT8
);

endmodule;
