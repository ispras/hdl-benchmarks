//NOTE: no-implementation module stub

module REG16LC (
    input DSPCLK,
    input MMR_web,
    input TCR_we,
    input [15:0] DMD,
    output [15:0] TCR,
    input T_RST
);
endmodule
