//NOTE: no-implementation module stub

module GtCLK_BUF (
    output Z,
    input A
);

endmodule
