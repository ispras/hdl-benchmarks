module s35932_bench(
  blif_clk_net,
  blif_reset_net,
  DATA_0_31,
  DATA_0_30,
  DATA_0_29,
  DATA_0_28,
  DATA_0_27,
  DATA_0_26,
  DATA_0_25,
  DATA_0_24,
  DATA_0_23,
  DATA_0_22,
  DATA_0_21,
  DATA_0_20,
  DATA_0_19,
  DATA_0_18,
  DATA_0_17,
  DATA_0_16,
  DATA_0_15,
  DATA_0_14,
  DATA_0_13,
  DATA_0_12,
  DATA_0_11,
  DATA_0_10,
  DATA_0_9,
  DATA_0_8,
  DATA_0_7,
  DATA_0_6,
  DATA_0_5,
  DATA_0_4,
  DATA_0_3,
  DATA_0_2,
  DATA_0_1,
  DATA_0_0,
  RESET,
  TM1,
  TM0,
  DATA_9_31,
  DATA_9_30,
  DATA_9_29,
  DATA_9_28,
  DATA_9_27,
  DATA_9_26,
  DATA_9_25,
  DATA_9_24,
  DATA_9_23,
  DATA_9_22,
  DATA_9_21,
  DATA_9_20,
  DATA_9_19,
  DATA_9_18,
  DATA_9_17,
  DATA_9_16,
  DATA_9_15,
  DATA_9_14,
  DATA_9_13,
  DATA_9_12,
  DATA_9_11,
  DATA_9_10,
  DATA_9_9,
  DATA_9_8,
  DATA_9_7,
  DATA_9_6,
  DATA_9_5,
  DATA_9_4,
  DATA_9_3,
  DATA_9_2,
  DATA_9_1,
  DATA_9_0,
  CRC_OUT_9_0,
  CRC_OUT_9_1,
  CRC_OUT_9_2,
  CRC_OUT_9_3,
  CRC_OUT_9_4,
  CRC_OUT_9_5,
  CRC_OUT_9_6,
  CRC_OUT_9_7,
  CRC_OUT_9_8,
  CRC_OUT_9_9,
  CRC_OUT_9_10,
  CRC_OUT_9_11,
  CRC_OUT_9_12,
  CRC_OUT_9_13,
  CRC_OUT_9_14,
  CRC_OUT_9_15,
  CRC_OUT_9_16,
  CRC_OUT_9_17,
  CRC_OUT_9_18,
  CRC_OUT_9_19,
  CRC_OUT_9_20,
  CRC_OUT_9_21,
  CRC_OUT_9_22,
  CRC_OUT_9_23,
  CRC_OUT_9_24,
  CRC_OUT_9_25,
  CRC_OUT_9_26,
  CRC_OUT_9_27,
  CRC_OUT_9_28,
  CRC_OUT_9_29,
  CRC_OUT_9_30,
  CRC_OUT_9_31,
  CRC_OUT_8_0,
  CRC_OUT_8_1,
  CRC_OUT_8_2,
  CRC_OUT_8_3,
  CRC_OUT_8_4,
  CRC_OUT_8_5,
  CRC_OUT_8_6,
  CRC_OUT_8_7,
  CRC_OUT_8_8,
  CRC_OUT_8_9,
  CRC_OUT_8_10,
  CRC_OUT_8_11,
  CRC_OUT_8_12,
  CRC_OUT_8_13,
  CRC_OUT_8_14,
  CRC_OUT_8_15,
  CRC_OUT_8_16,
  CRC_OUT_8_17,
  CRC_OUT_8_18,
  CRC_OUT_8_19,
  CRC_OUT_8_20,
  CRC_OUT_8_21,
  CRC_OUT_8_22,
  CRC_OUT_8_23,
  CRC_OUT_8_24,
  CRC_OUT_8_25,
  CRC_OUT_8_26,
  CRC_OUT_8_27,
  CRC_OUT_8_28,
  CRC_OUT_8_29,
  CRC_OUT_8_30,
  CRC_OUT_8_31,
  CRC_OUT_7_0,
  CRC_OUT_7_1,
  CRC_OUT_7_2,
  CRC_OUT_7_3,
  CRC_OUT_7_4,
  CRC_OUT_7_5,
  CRC_OUT_7_6,
  CRC_OUT_7_7,
  CRC_OUT_7_8,
  CRC_OUT_7_9,
  CRC_OUT_7_10,
  CRC_OUT_7_11,
  CRC_OUT_7_12,
  CRC_OUT_7_13,
  CRC_OUT_7_14,
  CRC_OUT_7_15,
  CRC_OUT_7_16,
  CRC_OUT_7_17,
  CRC_OUT_7_18,
  CRC_OUT_7_19,
  CRC_OUT_7_20,
  CRC_OUT_7_21,
  CRC_OUT_7_22,
  CRC_OUT_7_23,
  CRC_OUT_7_24,
  CRC_OUT_7_25,
  CRC_OUT_7_26,
  CRC_OUT_7_27,
  CRC_OUT_7_28,
  CRC_OUT_7_29,
  CRC_OUT_7_30,
  CRC_OUT_7_31,
  CRC_OUT_6_0,
  CRC_OUT_6_1,
  CRC_OUT_6_2,
  CRC_OUT_6_3,
  CRC_OUT_6_4,
  CRC_OUT_6_5,
  CRC_OUT_6_6,
  CRC_OUT_6_7,
  CRC_OUT_6_8,
  CRC_OUT_6_9,
  CRC_OUT_6_10,
  CRC_OUT_6_11,
  CRC_OUT_6_12,
  CRC_OUT_6_13,
  CRC_OUT_6_14,
  CRC_OUT_6_15,
  CRC_OUT_6_16,
  CRC_OUT_6_17,
  CRC_OUT_6_18,
  CRC_OUT_6_19,
  CRC_OUT_6_20,
  CRC_OUT_6_21,
  CRC_OUT_6_22,
  CRC_OUT_6_23,
  CRC_OUT_6_24,
  CRC_OUT_6_25,
  CRC_OUT_6_26,
  CRC_OUT_6_27,
  CRC_OUT_6_28,
  CRC_OUT_6_29,
  CRC_OUT_6_30,
  CRC_OUT_6_31,
  CRC_OUT_5_0,
  CRC_OUT_5_1,
  CRC_OUT_5_2,
  CRC_OUT_5_3,
  CRC_OUT_5_4,
  CRC_OUT_5_5,
  CRC_OUT_5_6,
  CRC_OUT_5_7,
  CRC_OUT_5_8,
  CRC_OUT_5_9,
  CRC_OUT_5_10,
  CRC_OUT_5_11,
  CRC_OUT_5_12,
  CRC_OUT_5_13,
  CRC_OUT_5_14,
  CRC_OUT_5_15,
  CRC_OUT_5_16,
  CRC_OUT_5_17,
  CRC_OUT_5_18,
  CRC_OUT_5_19,
  CRC_OUT_5_20,
  CRC_OUT_5_21,
  CRC_OUT_5_22,
  CRC_OUT_5_23,
  CRC_OUT_5_24,
  CRC_OUT_5_25,
  CRC_OUT_5_26,
  CRC_OUT_5_27,
  CRC_OUT_5_28,
  CRC_OUT_5_29,
  CRC_OUT_5_30,
  CRC_OUT_5_31,
  CRC_OUT_4_0,
  CRC_OUT_4_1,
  CRC_OUT_4_2,
  CRC_OUT_4_3,
  CRC_OUT_4_4,
  CRC_OUT_4_5,
  CRC_OUT_4_6,
  CRC_OUT_4_7,
  CRC_OUT_4_8,
  CRC_OUT_4_9,
  CRC_OUT_4_10,
  CRC_OUT_4_11,
  CRC_OUT_4_12,
  CRC_OUT_4_13,
  CRC_OUT_4_14,
  CRC_OUT_4_15,
  CRC_OUT_4_16,
  CRC_OUT_4_17,
  CRC_OUT_4_18,
  CRC_OUT_4_19,
  CRC_OUT_4_20,
  CRC_OUT_4_21,
  CRC_OUT_4_22,
  CRC_OUT_4_23,
  CRC_OUT_4_24,
  CRC_OUT_4_25,
  CRC_OUT_4_26,
  CRC_OUT_4_27,
  CRC_OUT_4_28,
  CRC_OUT_4_29,
  CRC_OUT_4_30,
  CRC_OUT_4_31,
  CRC_OUT_3_0,
  CRC_OUT_3_1,
  CRC_OUT_3_2,
  CRC_OUT_3_3,
  CRC_OUT_3_4,
  CRC_OUT_3_5,
  CRC_OUT_3_6,
  CRC_OUT_3_7,
  CRC_OUT_3_8,
  CRC_OUT_3_9,
  CRC_OUT_3_10,
  CRC_OUT_3_11,
  CRC_OUT_3_12,
  CRC_OUT_3_13,
  CRC_OUT_3_14,
  CRC_OUT_3_15,
  CRC_OUT_3_16,
  CRC_OUT_3_17,
  CRC_OUT_3_18,
  CRC_OUT_3_19,
  CRC_OUT_3_20,
  CRC_OUT_3_21,
  CRC_OUT_3_22,
  CRC_OUT_3_23,
  CRC_OUT_3_24,
  CRC_OUT_3_25,
  CRC_OUT_3_26,
  CRC_OUT_3_27,
  CRC_OUT_3_28,
  CRC_OUT_3_29,
  CRC_OUT_3_30,
  CRC_OUT_3_31,
  CRC_OUT_2_0,
  CRC_OUT_2_1,
  CRC_OUT_2_2,
  CRC_OUT_2_3,
  CRC_OUT_2_4,
  CRC_OUT_2_5,
  CRC_OUT_2_6,
  CRC_OUT_2_7,
  CRC_OUT_2_8,
  CRC_OUT_2_9,
  CRC_OUT_2_10,
  CRC_OUT_2_11,
  CRC_OUT_2_12,
  CRC_OUT_2_13,
  CRC_OUT_2_14,
  CRC_OUT_2_15,
  CRC_OUT_2_16,
  CRC_OUT_2_17,
  CRC_OUT_2_18,
  CRC_OUT_2_19,
  CRC_OUT_2_20,
  CRC_OUT_2_21,
  CRC_OUT_2_22,
  CRC_OUT_2_23,
  CRC_OUT_2_24,
  CRC_OUT_2_25,
  CRC_OUT_2_26,
  CRC_OUT_2_27,
  CRC_OUT_2_28,
  CRC_OUT_2_29,
  CRC_OUT_2_30,
  CRC_OUT_2_31,
  CRC_OUT_1_0,
  CRC_OUT_1_1,
  CRC_OUT_1_2,
  CRC_OUT_1_3,
  CRC_OUT_1_4,
  CRC_OUT_1_5,
  CRC_OUT_1_6,
  CRC_OUT_1_7,
  CRC_OUT_1_8,
  CRC_OUT_1_9,
  CRC_OUT_1_10,
  CRC_OUT_1_11,
  CRC_OUT_1_12,
  CRC_OUT_1_13,
  CRC_OUT_1_14,
  CRC_OUT_1_15,
  CRC_OUT_1_16,
  CRC_OUT_1_17,
  CRC_OUT_1_18,
  CRC_OUT_1_19,
  CRC_OUT_1_20,
  CRC_OUT_1_21,
  CRC_OUT_1_22,
  CRC_OUT_1_23,
  CRC_OUT_1_24,
  CRC_OUT_1_25,
  CRC_OUT_1_26,
  CRC_OUT_1_27,
  CRC_OUT_1_28,
  CRC_OUT_1_29,
  CRC_OUT_1_30,
  CRC_OUT_1_31);
input blif_clk_net;
input blif_reset_net;
input DATA_0_31;
input DATA_0_30;
input DATA_0_29;
input DATA_0_28;
input DATA_0_27;
input DATA_0_26;
input DATA_0_25;
input DATA_0_24;
input DATA_0_23;
input DATA_0_22;
input DATA_0_21;
input DATA_0_20;
input DATA_0_19;
input DATA_0_18;
input DATA_0_17;
input DATA_0_16;
input DATA_0_15;
input DATA_0_14;
input DATA_0_13;
input DATA_0_12;
input DATA_0_11;
input DATA_0_10;
input DATA_0_9;
input DATA_0_8;
input DATA_0_7;
input DATA_0_6;
input DATA_0_5;
input DATA_0_4;
input DATA_0_3;
input DATA_0_2;
input DATA_0_1;
input DATA_0_0;
input RESET;
input TM1;
input TM0;
output DATA_9_31;
output DATA_9_30;
output DATA_9_29;
output DATA_9_28;
output DATA_9_27;
output DATA_9_26;
output DATA_9_25;
output DATA_9_24;
output DATA_9_23;
output DATA_9_22;
output DATA_9_21;
output DATA_9_20;
output DATA_9_19;
output DATA_9_18;
output DATA_9_17;
output DATA_9_16;
output DATA_9_15;
output DATA_9_14;
output DATA_9_13;
output DATA_9_12;
output DATA_9_11;
output DATA_9_10;
output DATA_9_9;
output DATA_9_8;
output DATA_9_7;
output DATA_9_6;
output DATA_9_5;
output DATA_9_4;
output DATA_9_3;
output DATA_9_2;
output DATA_9_1;
output DATA_9_0;
output CRC_OUT_9_0;
output CRC_OUT_9_1;
output CRC_OUT_9_2;
output CRC_OUT_9_3;
output CRC_OUT_9_4;
output CRC_OUT_9_5;
output CRC_OUT_9_6;
output CRC_OUT_9_7;
output CRC_OUT_9_8;
output CRC_OUT_9_9;
output CRC_OUT_9_10;
output CRC_OUT_9_11;
output CRC_OUT_9_12;
output CRC_OUT_9_13;
output CRC_OUT_9_14;
output CRC_OUT_9_15;
output CRC_OUT_9_16;
output CRC_OUT_9_17;
output CRC_OUT_9_18;
output CRC_OUT_9_19;
output CRC_OUT_9_20;
output CRC_OUT_9_21;
output CRC_OUT_9_22;
output CRC_OUT_9_23;
output CRC_OUT_9_24;
output CRC_OUT_9_25;
output CRC_OUT_9_26;
output CRC_OUT_9_27;
output CRC_OUT_9_28;
output CRC_OUT_9_29;
output CRC_OUT_9_30;
output CRC_OUT_9_31;
output CRC_OUT_8_0;
output CRC_OUT_8_1;
output CRC_OUT_8_2;
output CRC_OUT_8_3;
output CRC_OUT_8_4;
output CRC_OUT_8_5;
output CRC_OUT_8_6;
output CRC_OUT_8_7;
output CRC_OUT_8_8;
output CRC_OUT_8_9;
output CRC_OUT_8_10;
output CRC_OUT_8_11;
output CRC_OUT_8_12;
output CRC_OUT_8_13;
output CRC_OUT_8_14;
output CRC_OUT_8_15;
output CRC_OUT_8_16;
output CRC_OUT_8_17;
output CRC_OUT_8_18;
output CRC_OUT_8_19;
output CRC_OUT_8_20;
output CRC_OUT_8_21;
output CRC_OUT_8_22;
output CRC_OUT_8_23;
output CRC_OUT_8_24;
output CRC_OUT_8_25;
output CRC_OUT_8_26;
output CRC_OUT_8_27;
output CRC_OUT_8_28;
output CRC_OUT_8_29;
output CRC_OUT_8_30;
output CRC_OUT_8_31;
output CRC_OUT_7_0;
output CRC_OUT_7_1;
output CRC_OUT_7_2;
output CRC_OUT_7_3;
output CRC_OUT_7_4;
output CRC_OUT_7_5;
output CRC_OUT_7_6;
output CRC_OUT_7_7;
output CRC_OUT_7_8;
output CRC_OUT_7_9;
output CRC_OUT_7_10;
output CRC_OUT_7_11;
output CRC_OUT_7_12;
output CRC_OUT_7_13;
output CRC_OUT_7_14;
output CRC_OUT_7_15;
output CRC_OUT_7_16;
output CRC_OUT_7_17;
output CRC_OUT_7_18;
output CRC_OUT_7_19;
output CRC_OUT_7_20;
output CRC_OUT_7_21;
output CRC_OUT_7_22;
output CRC_OUT_7_23;
output CRC_OUT_7_24;
output CRC_OUT_7_25;
output CRC_OUT_7_26;
output CRC_OUT_7_27;
output CRC_OUT_7_28;
output CRC_OUT_7_29;
output CRC_OUT_7_30;
output CRC_OUT_7_31;
output CRC_OUT_6_0;
output CRC_OUT_6_1;
output CRC_OUT_6_2;
output CRC_OUT_6_3;
output CRC_OUT_6_4;
output CRC_OUT_6_5;
output CRC_OUT_6_6;
output CRC_OUT_6_7;
output CRC_OUT_6_8;
output CRC_OUT_6_9;
output CRC_OUT_6_10;
output CRC_OUT_6_11;
output CRC_OUT_6_12;
output CRC_OUT_6_13;
output CRC_OUT_6_14;
output CRC_OUT_6_15;
output CRC_OUT_6_16;
output CRC_OUT_6_17;
output CRC_OUT_6_18;
output CRC_OUT_6_19;
output CRC_OUT_6_20;
output CRC_OUT_6_21;
output CRC_OUT_6_22;
output CRC_OUT_6_23;
output CRC_OUT_6_24;
output CRC_OUT_6_25;
output CRC_OUT_6_26;
output CRC_OUT_6_27;
output CRC_OUT_6_28;
output CRC_OUT_6_29;
output CRC_OUT_6_30;
output CRC_OUT_6_31;
output CRC_OUT_5_0;
output CRC_OUT_5_1;
output CRC_OUT_5_2;
output CRC_OUT_5_3;
output CRC_OUT_5_4;
output CRC_OUT_5_5;
output CRC_OUT_5_6;
output CRC_OUT_5_7;
output CRC_OUT_5_8;
output CRC_OUT_5_9;
output CRC_OUT_5_10;
output CRC_OUT_5_11;
output CRC_OUT_5_12;
output CRC_OUT_5_13;
output CRC_OUT_5_14;
output CRC_OUT_5_15;
output CRC_OUT_5_16;
output CRC_OUT_5_17;
output CRC_OUT_5_18;
output CRC_OUT_5_19;
output CRC_OUT_5_20;
output CRC_OUT_5_21;
output CRC_OUT_5_22;
output CRC_OUT_5_23;
output CRC_OUT_5_24;
output CRC_OUT_5_25;
output CRC_OUT_5_26;
output CRC_OUT_5_27;
output CRC_OUT_5_28;
output CRC_OUT_5_29;
output CRC_OUT_5_30;
output CRC_OUT_5_31;
output CRC_OUT_4_0;
output CRC_OUT_4_1;
output CRC_OUT_4_2;
output CRC_OUT_4_3;
output CRC_OUT_4_4;
output CRC_OUT_4_5;
output CRC_OUT_4_6;
output CRC_OUT_4_7;
output CRC_OUT_4_8;
output CRC_OUT_4_9;
output CRC_OUT_4_10;
output CRC_OUT_4_11;
output CRC_OUT_4_12;
output CRC_OUT_4_13;
output CRC_OUT_4_14;
output CRC_OUT_4_15;
output CRC_OUT_4_16;
output CRC_OUT_4_17;
output CRC_OUT_4_18;
output CRC_OUT_4_19;
output CRC_OUT_4_20;
output CRC_OUT_4_21;
output CRC_OUT_4_22;
output CRC_OUT_4_23;
output CRC_OUT_4_24;
output CRC_OUT_4_25;
output CRC_OUT_4_26;
output CRC_OUT_4_27;
output CRC_OUT_4_28;
output CRC_OUT_4_29;
output CRC_OUT_4_30;
output CRC_OUT_4_31;
output CRC_OUT_3_0;
output CRC_OUT_3_1;
output CRC_OUT_3_2;
output CRC_OUT_3_3;
output CRC_OUT_3_4;
output CRC_OUT_3_5;
output CRC_OUT_3_6;
output CRC_OUT_3_7;
output CRC_OUT_3_8;
output CRC_OUT_3_9;
output CRC_OUT_3_10;
output CRC_OUT_3_11;
output CRC_OUT_3_12;
output CRC_OUT_3_13;
output CRC_OUT_3_14;
output CRC_OUT_3_15;
output CRC_OUT_3_16;
output CRC_OUT_3_17;
output CRC_OUT_3_18;
output CRC_OUT_3_19;
output CRC_OUT_3_20;
output CRC_OUT_3_21;
output CRC_OUT_3_22;
output CRC_OUT_3_23;
output CRC_OUT_3_24;
output CRC_OUT_3_25;
output CRC_OUT_3_26;
output CRC_OUT_3_27;
output CRC_OUT_3_28;
output CRC_OUT_3_29;
output CRC_OUT_3_30;
output CRC_OUT_3_31;
output CRC_OUT_2_0;
output CRC_OUT_2_1;
output CRC_OUT_2_2;
output CRC_OUT_2_3;
output CRC_OUT_2_4;
output CRC_OUT_2_5;
output CRC_OUT_2_6;
output CRC_OUT_2_7;
output CRC_OUT_2_8;
output CRC_OUT_2_9;
output CRC_OUT_2_10;
output CRC_OUT_2_11;
output CRC_OUT_2_12;
output CRC_OUT_2_13;
output CRC_OUT_2_14;
output CRC_OUT_2_15;
output CRC_OUT_2_16;
output CRC_OUT_2_17;
output CRC_OUT_2_18;
output CRC_OUT_2_19;
output CRC_OUT_2_20;
output CRC_OUT_2_21;
output CRC_OUT_2_22;
output CRC_OUT_2_23;
output CRC_OUT_2_24;
output CRC_OUT_2_25;
output CRC_OUT_2_26;
output CRC_OUT_2_27;
output CRC_OUT_2_28;
output CRC_OUT_2_29;
output CRC_OUT_2_30;
output CRC_OUT_2_31;
output CRC_OUT_1_0;
output CRC_OUT_1_1;
output CRC_OUT_1_2;
output CRC_OUT_1_3;
output CRC_OUT_1_4;
output CRC_OUT_1_5;
output CRC_OUT_1_6;
output CRC_OUT_1_7;
output CRC_OUT_1_8;
output CRC_OUT_1_9;
output CRC_OUT_1_10;
output CRC_OUT_1_11;
output CRC_OUT_1_12;
output CRC_OUT_1_13;
output CRC_OUT_1_14;
output CRC_OUT_1_15;
output CRC_OUT_1_16;
output CRC_OUT_1_17;
output CRC_OUT_1_18;
output CRC_OUT_1_19;
output CRC_OUT_1_20;
output CRC_OUT_1_21;
output CRC_OUT_1_22;
output CRC_OUT_1_23;
output CRC_OUT_1_24;
output CRC_OUT_1_25;
output CRC_OUT_1_26;
output CRC_OUT_1_27;
output CRC_OUT_1_28;
output CRC_OUT_1_29;
output CRC_OUT_1_30;
output CRC_OUT_1_31;
reg WX485;
reg WX487;
reg WX489;
reg WX491;
reg WX493;
reg WX495;
reg WX497;
reg WX499;
reg WX501;
reg WX503;
reg WX505;
reg WX507;
reg WX509;
reg WX511;
reg WX513;
reg WX515;
reg WX517;
reg WX519;
reg WX521;
reg WX523;
reg WX525;
reg WX527;
reg WX529;
reg WX531;
reg WX533;
reg WX535;
reg WX537;
reg WX539;
reg WX541;
reg WX543;
reg WX545;
reg WX547;
reg WX645;
reg WX647;
reg WX649;
reg WX651;
reg WX653;
reg WX655;
reg WX657;
reg WX659;
reg WX661;
reg WX663;
reg WX665;
reg WX667;
reg WX669;
reg WX671;
reg WX673;
reg WX675;
reg WX677;
reg WX679;
reg WX681;
reg WX683;
reg WX685;
reg WX687;
reg WX689;
reg WX691;
reg WX693;
reg WX695;
reg WX697;
reg WX699;
reg WX701;
reg WX703;
reg WX705;
reg WX707;
reg WX709;
reg WX711;
reg WX713;
reg WX715;
reg WX717;
reg WX719;
reg WX721;
reg WX723;
reg WX725;
reg WX727;
reg WX729;
reg WX731;
reg WX733;
reg WX735;
reg WX737;
reg WX739;
reg WX741;
reg WX743;
reg WX745;
reg WX747;
reg WX749;
reg WX751;
reg WX753;
reg WX755;
reg WX757;
reg WX759;
reg WX761;
reg WX763;
reg WX765;
reg WX767;
reg WX769;
reg WX771;
reg WX773;
reg WX775;
reg WX777;
reg WX779;
reg WX781;
reg WX783;
reg WX785;
reg WX787;
reg WX789;
reg WX791;
reg WX793;
reg WX795;
reg WX797;
reg WX799;
reg WX801;
reg WX803;
reg WX805;
reg WX807;
reg WX809;
reg WX811;
reg WX813;
reg WX815;
reg WX817;
reg WX819;
reg WX821;
reg WX823;
reg WX825;
reg WX827;
reg WX829;
reg WX831;
reg WX833;
reg WX835;
reg WX837;
reg WX839;
reg WX841;
reg WX843;
reg WX845;
reg WX847;
reg WX849;
reg WX851;
reg WX853;
reg WX855;
reg WX857;
reg WX859;
reg WX861;
reg WX863;
reg WX865;
reg WX867;
reg WX869;
reg WX871;
reg WX873;
reg WX875;
reg WX877;
reg WX879;
reg WX881;
reg WX883;
reg WX885;
reg WX887;
reg WX889;
reg WX891;
reg WX893;
reg WX895;
reg WX897;
reg WX899;
reg _2077_;
reg _2078_;
reg _2079_;
reg _2080_;
reg _2081_;
reg _2082_;
reg _2083_;
reg _2084_;
reg _2085_;
reg _2086_;
reg _2087_;
reg _2088_;
reg _2089_;
reg _2090_;
reg _2091_;
reg _2092_;
reg _2093_;
reg _2094_;
reg _2095_;
reg _2096_;
reg _2097_;
reg _2098_;
reg _2099_;
reg _2100_;
reg _2101_;
reg _2102_;
reg _2103_;
reg _2104_;
reg _2105_;
reg _2106_;
reg _2107_;
reg _2108_;
reg WX1778;
reg WX1780;
reg WX1782;
reg WX1784;
reg WX1786;
reg WX1788;
reg WX1790;
reg WX1792;
reg WX1794;
reg WX1796;
reg WX1798;
reg WX1800;
reg WX1802;
reg WX1804;
reg WX1806;
reg WX1808;
reg WX1810;
reg WX1812;
reg WX1814;
reg WX1816;
reg WX1818;
reg WX1820;
reg WX1822;
reg WX1824;
reg WX1826;
reg WX1828;
reg WX1830;
reg WX1832;
reg WX1834;
reg WX1836;
reg WX1838;
reg WX1840;
reg WX1938;
reg WX1940;
reg WX1942;
reg WX1944;
reg WX1946;
reg WX1948;
reg WX1950;
reg WX1952;
reg WX1954;
reg WX1956;
reg WX1958;
reg WX1960;
reg WX1962;
reg WX1964;
reg WX1966;
reg WX1968;
reg WX1970;
reg WX1972;
reg WX1974;
reg WX1976;
reg WX1978;
reg WX1980;
reg WX1982;
reg WX1984;
reg WX1986;
reg WX1988;
reg WX1990;
reg WX1992;
reg WX1994;
reg WX1996;
reg WX1998;
reg WX2000;
reg WX2002;
reg WX2004;
reg WX2006;
reg WX2008;
reg WX2010;
reg WX2012;
reg WX2014;
reg WX2016;
reg WX2018;
reg WX2020;
reg WX2022;
reg WX2024;
reg WX2026;
reg WX2028;
reg WX2030;
reg WX2032;
reg WX2034;
reg WX2036;
reg WX2038;
reg WX2040;
reg WX2042;
reg WX2044;
reg WX2046;
reg WX2048;
reg WX2050;
reg WX2052;
reg WX2054;
reg WX2056;
reg WX2058;
reg WX2060;
reg WX2062;
reg WX2064;
reg WX2066;
reg WX2068;
reg WX2070;
reg WX2072;
reg WX2074;
reg WX2076;
reg WX2078;
reg WX2080;
reg WX2082;
reg WX2084;
reg WX2086;
reg WX2088;
reg WX2090;
reg WX2092;
reg WX2094;
reg WX2096;
reg WX2098;
reg WX2100;
reg WX2102;
reg WX2104;
reg WX2106;
reg WX2108;
reg WX2110;
reg WX2112;
reg WX2114;
reg WX2116;
reg WX2118;
reg WX2120;
reg WX2122;
reg WX2124;
reg WX2126;
reg WX2128;
reg WX2130;
reg WX2132;
reg WX2134;
reg WX2136;
reg WX2138;
reg WX2140;
reg WX2142;
reg WX2144;
reg WX2146;
reg WX2148;
reg WX2150;
reg WX2152;
reg WX2154;
reg WX2156;
reg WX2158;
reg WX2160;
reg WX2162;
reg WX2164;
reg WX2166;
reg WX2168;
reg WX2170;
reg WX2172;
reg WX2174;
reg WX2176;
reg WX2178;
reg WX2180;
reg WX2182;
reg WX2184;
reg WX2186;
reg WX2188;
reg WX2190;
reg WX2192;
reg _2109_;
reg _2110_;
reg _2111_;
reg _2112_;
reg _2113_;
reg _2114_;
reg _2115_;
reg _2116_;
reg _2117_;
reg _2118_;
reg _2119_;
reg _2120_;
reg _2121_;
reg _2122_;
reg _2123_;
reg _2124_;
reg _2125_;
reg _2126_;
reg _2127_;
reg _2128_;
reg _2129_;
reg _2130_;
reg _2131_;
reg _2132_;
reg _2133_;
reg _2134_;
reg _2135_;
reg _2136_;
reg _2137_;
reg _2138_;
reg _2139_;
reg _2140_;
reg WX3071;
reg WX3073;
reg WX3075;
reg WX3077;
reg WX3079;
reg WX3081;
reg WX3083;
reg WX3085;
reg WX3087;
reg WX3089;
reg WX3091;
reg WX3093;
reg WX3095;
reg WX3097;
reg WX3099;
reg WX3101;
reg WX3103;
reg WX3105;
reg WX3107;
reg WX3109;
reg WX3111;
reg WX3113;
reg WX3115;
reg WX3117;
reg WX3119;
reg WX3121;
reg WX3123;
reg WX3125;
reg WX3127;
reg WX3129;
reg WX3131;
reg WX3133;
reg WX3231;
reg WX3233;
reg WX3235;
reg WX3237;
reg WX3239;
reg WX3241;
reg WX3243;
reg WX3245;
reg WX3247;
reg WX3249;
reg WX3251;
reg WX3253;
reg WX3255;
reg WX3257;
reg WX3259;
reg WX3261;
reg WX3263;
reg WX3265;
reg WX3267;
reg WX3269;
reg WX3271;
reg WX3273;
reg WX3275;
reg WX3277;
reg WX3279;
reg WX3281;
reg WX3283;
reg WX3285;
reg WX3287;
reg WX3289;
reg WX3291;
reg WX3293;
reg WX3295;
reg WX3297;
reg WX3299;
reg WX3301;
reg WX3303;
reg WX3305;
reg WX3307;
reg WX3309;
reg WX3311;
reg WX3313;
reg WX3315;
reg WX3317;
reg WX3319;
reg WX3321;
reg WX3323;
reg WX3325;
reg WX3327;
reg WX3329;
reg WX3331;
reg WX3333;
reg WX3335;
reg WX3337;
reg WX3339;
reg WX3341;
reg WX3343;
reg WX3345;
reg WX3347;
reg WX3349;
reg WX3351;
reg WX3353;
reg WX3355;
reg WX3357;
reg WX3359;
reg WX3361;
reg WX3363;
reg WX3365;
reg WX3367;
reg WX3369;
reg WX3371;
reg WX3373;
reg WX3375;
reg WX3377;
reg WX3379;
reg WX3381;
reg WX3383;
reg WX3385;
reg WX3387;
reg WX3389;
reg WX3391;
reg WX3393;
reg WX3395;
reg WX3397;
reg WX3399;
reg WX3401;
reg WX3403;
reg WX3405;
reg WX3407;
reg WX3409;
reg WX3411;
reg WX3413;
reg WX3415;
reg WX3417;
reg WX3419;
reg WX3421;
reg WX3423;
reg WX3425;
reg WX3427;
reg WX3429;
reg WX3431;
reg WX3433;
reg WX3435;
reg WX3437;
reg WX3439;
reg WX3441;
reg WX3443;
reg WX3445;
reg WX3447;
reg WX3449;
reg WX3451;
reg WX3453;
reg WX3455;
reg WX3457;
reg WX3459;
reg WX3461;
reg WX3463;
reg WX3465;
reg WX3467;
reg WX3469;
reg WX3471;
reg WX3473;
reg WX3475;
reg WX3477;
reg WX3479;
reg WX3481;
reg WX3483;
reg WX3485;
reg _2141_;
reg _2142_;
reg _2143_;
reg _2144_;
reg _2145_;
reg _2146_;
reg _2147_;
reg _2148_;
reg _2149_;
reg _2150_;
reg _2151_;
reg _2152_;
reg _2153_;
reg _2154_;
reg _2155_;
reg _2156_;
reg _2157_;
reg _2158_;
reg _2159_;
reg _2160_;
reg _2161_;
reg _2162_;
reg _2163_;
reg _2164_;
reg _2165_;
reg _2166_;
reg _2167_;
reg _2168_;
reg _2169_;
reg _2170_;
reg _2171_;
reg _2172_;
reg WX4364;
reg WX4366;
reg WX4368;
reg WX4370;
reg WX4372;
reg WX4374;
reg WX4376;
reg WX4378;
reg WX4380;
reg WX4382;
reg WX4384;
reg WX4386;
reg WX4388;
reg WX4390;
reg WX4392;
reg WX4394;
reg WX4396;
reg WX4398;
reg WX4400;
reg WX4402;
reg WX4404;
reg WX4406;
reg WX4408;
reg WX4410;
reg WX4412;
reg WX4414;
reg WX4416;
reg WX4418;
reg WX4420;
reg WX4422;
reg WX4424;
reg WX4426;
reg WX4524;
reg WX4526;
reg WX4528;
reg WX4530;
reg WX4532;
reg WX4534;
reg WX4536;
reg WX4538;
reg WX4540;
reg WX4542;
reg WX4544;
reg WX4546;
reg WX4548;
reg WX4550;
reg WX4552;
reg WX4554;
reg WX4556;
reg WX4558;
reg WX4560;
reg WX4562;
reg WX4564;
reg WX4566;
reg WX4568;
reg WX4570;
reg WX4572;
reg WX4574;
reg WX4576;
reg WX4578;
reg WX4580;
reg WX4582;
reg WX4584;
reg WX4586;
reg WX4588;
reg WX4590;
reg WX4592;
reg WX4594;
reg WX4596;
reg WX4598;
reg WX4600;
reg WX4602;
reg WX4604;
reg WX4606;
reg WX4608;
reg WX4610;
reg WX4612;
reg WX4614;
reg WX4616;
reg WX4618;
reg WX4620;
reg WX4622;
reg WX4624;
reg WX4626;
reg WX4628;
reg WX4630;
reg WX4632;
reg WX4634;
reg WX4636;
reg WX4638;
reg WX4640;
reg WX4642;
reg WX4644;
reg WX4646;
reg WX4648;
reg WX4650;
reg WX4652;
reg WX4654;
reg WX4656;
reg WX4658;
reg WX4660;
reg WX4662;
reg WX4664;
reg WX4666;
reg WX4668;
reg WX4670;
reg WX4672;
reg WX4674;
reg WX4676;
reg WX4678;
reg WX4680;
reg WX4682;
reg WX4684;
reg WX4686;
reg WX4688;
reg WX4690;
reg WX4692;
reg WX4694;
reg WX4696;
reg WX4698;
reg WX4700;
reg WX4702;
reg WX4704;
reg WX4706;
reg WX4708;
reg WX4710;
reg WX4712;
reg WX4714;
reg WX4716;
reg WX4718;
reg WX4720;
reg WX4722;
reg WX4724;
reg WX4726;
reg WX4728;
reg WX4730;
reg WX4732;
reg WX4734;
reg WX4736;
reg WX4738;
reg WX4740;
reg WX4742;
reg WX4744;
reg WX4746;
reg WX4748;
reg WX4750;
reg WX4752;
reg WX4754;
reg WX4756;
reg WX4758;
reg WX4760;
reg WX4762;
reg WX4764;
reg WX4766;
reg WX4768;
reg WX4770;
reg WX4772;
reg WX4774;
reg WX4776;
reg WX4778;
reg _2173_;
reg _2174_;
reg _2175_;
reg _2176_;
reg _2177_;
reg _2178_;
reg _2179_;
reg _2180_;
reg _2181_;
reg _2182_;
reg _2183_;
reg _2184_;
reg _2185_;
reg _2186_;
reg _2187_;
reg _2188_;
reg _2189_;
reg _2190_;
reg _2191_;
reg _2192_;
reg _2193_;
reg _2194_;
reg _2195_;
reg _2196_;
reg _2197_;
reg _2198_;
reg _2199_;
reg _2200_;
reg _2201_;
reg _2202_;
reg _2203_;
reg _2204_;
reg WX5657;
reg WX5659;
reg WX5661;
reg WX5663;
reg WX5665;
reg WX5667;
reg WX5669;
reg WX5671;
reg WX5673;
reg WX5675;
reg WX5677;
reg WX5679;
reg WX5681;
reg WX5683;
reg WX5685;
reg WX5687;
reg WX5689;
reg WX5691;
reg WX5693;
reg WX5695;
reg WX5697;
reg WX5699;
reg WX5701;
reg WX5703;
reg WX5705;
reg WX5707;
reg WX5709;
reg WX5711;
reg WX5713;
reg WX5715;
reg WX5717;
reg WX5719;
reg WX5817;
reg WX5819;
reg WX5821;
reg WX5823;
reg WX5825;
reg WX5827;
reg WX5829;
reg WX5831;
reg WX5833;
reg WX5835;
reg WX5837;
reg WX5839;
reg WX5841;
reg WX5843;
reg WX5845;
reg WX5847;
reg WX5849;
reg WX5851;
reg WX5853;
reg WX5855;
reg WX5857;
reg WX5859;
reg WX5861;
reg WX5863;
reg WX5865;
reg WX5867;
reg WX5869;
reg WX5871;
reg WX5873;
reg WX5875;
reg WX5877;
reg WX5879;
reg WX5881;
reg WX5883;
reg WX5885;
reg WX5887;
reg WX5889;
reg WX5891;
reg WX5893;
reg WX5895;
reg WX5897;
reg WX5899;
reg WX5901;
reg WX5903;
reg WX5905;
reg WX5907;
reg WX5909;
reg WX5911;
reg WX5913;
reg WX5915;
reg WX5917;
reg WX5919;
reg WX5921;
reg WX5923;
reg WX5925;
reg WX5927;
reg WX5929;
reg WX5931;
reg WX5933;
reg WX5935;
reg WX5937;
reg WX5939;
reg WX5941;
reg WX5943;
reg WX5945;
reg WX5947;
reg WX5949;
reg WX5951;
reg WX5953;
reg WX5955;
reg WX5957;
reg WX5959;
reg WX5961;
reg WX5963;
reg WX5965;
reg WX5967;
reg WX5969;
reg WX5971;
reg WX5973;
reg WX5975;
reg WX5977;
reg WX5979;
reg WX5981;
reg WX5983;
reg WX5985;
reg WX5987;
reg WX5989;
reg WX5991;
reg WX5993;
reg WX5995;
reg WX5997;
reg WX5999;
reg WX6001;
reg WX6003;
reg WX6005;
reg WX6007;
reg WX6009;
reg WX6011;
reg WX6013;
reg WX6015;
reg WX6017;
reg WX6019;
reg WX6021;
reg WX6023;
reg WX6025;
reg WX6027;
reg WX6029;
reg WX6031;
reg WX6033;
reg WX6035;
reg WX6037;
reg WX6039;
reg WX6041;
reg WX6043;
reg WX6045;
reg WX6047;
reg WX6049;
reg WX6051;
reg WX6053;
reg WX6055;
reg WX6057;
reg WX6059;
reg WX6061;
reg WX6063;
reg WX6065;
reg WX6067;
reg WX6069;
reg WX6071;
reg _2205_;
reg _2206_;
reg _2207_;
reg _2208_;
reg _2209_;
reg _2210_;
reg _2211_;
reg _2212_;
reg _2213_;
reg _2214_;
reg _2215_;
reg _2216_;
reg _2217_;
reg _2218_;
reg _2219_;
reg _2220_;
reg _2221_;
reg _2222_;
reg _2223_;
reg _2224_;
reg _2225_;
reg _2226_;
reg _2227_;
reg _2228_;
reg _2229_;
reg _2230_;
reg _2231_;
reg _2232_;
reg _2233_;
reg _2234_;
reg _2235_;
reg _2236_;
reg WX6950;
reg WX6952;
reg WX6954;
reg WX6956;
reg WX6958;
reg WX6960;
reg WX6962;
reg WX6964;
reg WX6966;
reg WX6968;
reg WX6970;
reg WX6972;
reg WX6974;
reg WX6976;
reg WX6978;
reg WX6980;
reg WX6982;
reg WX6984;
reg WX6986;
reg WX6988;
reg WX6990;
reg WX6992;
reg WX6994;
reg WX6996;
reg WX6998;
reg WX7000;
reg WX7002;
reg WX7004;
reg WX7006;
reg WX7008;
reg WX7010;
reg WX7012;
reg WX7110;
reg WX7112;
reg WX7114;
reg WX7116;
reg WX7118;
reg WX7120;
reg WX7122;
reg WX7124;
reg WX7126;
reg WX7128;
reg WX7130;
reg WX7132;
reg WX7134;
reg WX7136;
reg WX7138;
reg WX7140;
reg WX7142;
reg WX7144;
reg WX7146;
reg WX7148;
reg WX7150;
reg WX7152;
reg WX7154;
reg WX7156;
reg WX7158;
reg WX7160;
reg WX7162;
reg WX7164;
reg WX7166;
reg WX7168;
reg WX7170;
reg WX7172;
reg WX7174;
reg WX7176;
reg WX7178;
reg WX7180;
reg WX7182;
reg WX7184;
reg WX7186;
reg WX7188;
reg WX7190;
reg WX7192;
reg WX7194;
reg WX7196;
reg WX7198;
reg WX7200;
reg WX7202;
reg WX7204;
reg WX7206;
reg WX7208;
reg WX7210;
reg WX7212;
reg WX7214;
reg WX7216;
reg WX7218;
reg WX7220;
reg WX7222;
reg WX7224;
reg WX7226;
reg WX7228;
reg WX7230;
reg WX7232;
reg WX7234;
reg WX7236;
reg WX7238;
reg WX7240;
reg WX7242;
reg WX7244;
reg WX7246;
reg WX7248;
reg WX7250;
reg WX7252;
reg WX7254;
reg WX7256;
reg WX7258;
reg WX7260;
reg WX7262;
reg WX7264;
reg WX7266;
reg WX7268;
reg WX7270;
reg WX7272;
reg WX7274;
reg WX7276;
reg WX7278;
reg WX7280;
reg WX7282;
reg WX7284;
reg WX7286;
reg WX7288;
reg WX7290;
reg WX7292;
reg WX7294;
reg WX7296;
reg WX7298;
reg WX7300;
reg WX7302;
reg WX7304;
reg WX7306;
reg WX7308;
reg WX7310;
reg WX7312;
reg WX7314;
reg WX7316;
reg WX7318;
reg WX7320;
reg WX7322;
reg WX7324;
reg WX7326;
reg WX7328;
reg WX7330;
reg WX7332;
reg WX7334;
reg WX7336;
reg WX7338;
reg WX7340;
reg WX7342;
reg WX7344;
reg WX7346;
reg WX7348;
reg WX7350;
reg WX7352;
reg WX7354;
reg WX7356;
reg WX7358;
reg WX7360;
reg WX7362;
reg WX7364;
reg _2237_;
reg _2238_;
reg _2239_;
reg _2240_;
reg _2241_;
reg _2242_;
reg _2243_;
reg _2244_;
reg _2245_;
reg _2246_;
reg _2247_;
reg _2248_;
reg _2249_;
reg _2250_;
reg _2251_;
reg _2252_;
reg _2253_;
reg _2254_;
reg _2255_;
reg _2256_;
reg _2257_;
reg _2258_;
reg _2259_;
reg _2260_;
reg _2261_;
reg _2262_;
reg _2263_;
reg _2264_;
reg _2265_;
reg _2266_;
reg _2267_;
reg _2268_;
reg WX8243;
reg WX8245;
reg WX8247;
reg WX8249;
reg WX8251;
reg WX8253;
reg WX8255;
reg WX8257;
reg WX8259;
reg WX8261;
reg WX8263;
reg WX8265;
reg WX8267;
reg WX8269;
reg WX8271;
reg WX8273;
reg WX8275;
reg WX8277;
reg WX8279;
reg WX8281;
reg WX8283;
reg WX8285;
reg WX8287;
reg WX8289;
reg WX8291;
reg WX8293;
reg WX8295;
reg WX8297;
reg WX8299;
reg WX8301;
reg WX8303;
reg WX8305;
reg WX8403;
reg WX8405;
reg WX8407;
reg WX8409;
reg WX8411;
reg WX8413;
reg WX8415;
reg WX8417;
reg WX8419;
reg WX8421;
reg WX8423;
reg WX8425;
reg WX8427;
reg WX8429;
reg WX8431;
reg WX8433;
reg WX8435;
reg WX8437;
reg WX8439;
reg WX8441;
reg WX8443;
reg WX8445;
reg WX8447;
reg WX8449;
reg WX8451;
reg WX8453;
reg WX8455;
reg WX8457;
reg WX8459;
reg WX8461;
reg WX8463;
reg WX8465;
reg WX8467;
reg WX8469;
reg WX8471;
reg WX8473;
reg WX8475;
reg WX8477;
reg WX8479;
reg WX8481;
reg WX8483;
reg WX8485;
reg WX8487;
reg WX8489;
reg WX8491;
reg WX8493;
reg WX8495;
reg WX8497;
reg WX8499;
reg WX8501;
reg WX8503;
reg WX8505;
reg WX8507;
reg WX8509;
reg WX8511;
reg WX8513;
reg WX8515;
reg WX8517;
reg WX8519;
reg WX8521;
reg WX8523;
reg WX8525;
reg WX8527;
reg WX8529;
reg WX8531;
reg WX8533;
reg WX8535;
reg WX8537;
reg WX8539;
reg WX8541;
reg WX8543;
reg WX8545;
reg WX8547;
reg WX8549;
reg WX8551;
reg WX8553;
reg WX8555;
reg WX8557;
reg WX8559;
reg WX8561;
reg WX8563;
reg WX8565;
reg WX8567;
reg WX8569;
reg WX8571;
reg WX8573;
reg WX8575;
reg WX8577;
reg WX8579;
reg WX8581;
reg WX8583;
reg WX8585;
reg WX8587;
reg WX8589;
reg WX8591;
reg WX8593;
reg WX8595;
reg WX8597;
reg WX8599;
reg WX8601;
reg WX8603;
reg WX8605;
reg WX8607;
reg WX8609;
reg WX8611;
reg WX8613;
reg WX8615;
reg WX8617;
reg WX8619;
reg WX8621;
reg WX8623;
reg WX8625;
reg WX8627;
reg WX8629;
reg WX8631;
reg WX8633;
reg WX8635;
reg WX8637;
reg WX8639;
reg WX8641;
reg WX8643;
reg WX8645;
reg WX8647;
reg WX8649;
reg WX8651;
reg WX8653;
reg WX8655;
reg WX8657;
reg _2269_;
reg _2270_;
reg _2271_;
reg _2272_;
reg _2273_;
reg _2274_;
reg _2275_;
reg _2276_;
reg _2277_;
reg _2278_;
reg _2279_;
reg _2280_;
reg _2281_;
reg _2282_;
reg _2283_;
reg _2284_;
reg _2285_;
reg _2286_;
reg _2287_;
reg _2288_;
reg _2289_;
reg _2290_;
reg _2291_;
reg _2292_;
reg _2293_;
reg _2294_;
reg _2295_;
reg _2296_;
reg _2297_;
reg _2298_;
reg _2299_;
reg _2300_;
reg WX9536;
reg WX9538;
reg WX9540;
reg WX9542;
reg WX9544;
reg WX9546;
reg WX9548;
reg WX9550;
reg WX9552;
reg WX9554;
reg WX9556;
reg WX9558;
reg WX9560;
reg WX9562;
reg WX9564;
reg WX9566;
reg WX9568;
reg WX9570;
reg WX9572;
reg WX9574;
reg WX9576;
reg WX9578;
reg WX9580;
reg WX9582;
reg WX9584;
reg WX9586;
reg WX9588;
reg WX9590;
reg WX9592;
reg WX9594;
reg WX9596;
reg WX9598;
reg WX9696;
reg WX9698;
reg WX9700;
reg WX9702;
reg WX9704;
reg WX9706;
reg WX9708;
reg WX9710;
reg WX9712;
reg WX9714;
reg WX9716;
reg WX9718;
reg WX9720;
reg WX9722;
reg WX9724;
reg WX9726;
reg WX9728;
reg WX9730;
reg WX9732;
reg WX9734;
reg WX9736;
reg WX9738;
reg WX9740;
reg WX9742;
reg WX9744;
reg WX9746;
reg WX9748;
reg WX9750;
reg WX9752;
reg WX9754;
reg WX9756;
reg WX9758;
reg WX9760;
reg WX9762;
reg WX9764;
reg WX9766;
reg WX9768;
reg WX9770;
reg WX9772;
reg WX9774;
reg WX9776;
reg WX9778;
reg WX9780;
reg WX9782;
reg WX9784;
reg WX9786;
reg WX9788;
reg WX9790;
reg WX9792;
reg WX9794;
reg WX9796;
reg WX9798;
reg WX9800;
reg WX9802;
reg WX9804;
reg WX9806;
reg WX9808;
reg WX9810;
reg WX9812;
reg WX9814;
reg WX9816;
reg WX9818;
reg WX9820;
reg WX9822;
reg WX9824;
reg WX9826;
reg WX9828;
reg WX9830;
reg WX9832;
reg WX9834;
reg WX9836;
reg WX9838;
reg WX9840;
reg WX9842;
reg WX9844;
reg WX9846;
reg WX9848;
reg WX9850;
reg WX9852;
reg WX9854;
reg WX9856;
reg WX9858;
reg WX9860;
reg WX9862;
reg WX9864;
reg WX9866;
reg WX9868;
reg WX9870;
reg WX9872;
reg WX9874;
reg WX9876;
reg WX9878;
reg WX9880;
reg WX9882;
reg WX9884;
reg WX9886;
reg WX9888;
reg WX9890;
reg WX9892;
reg WX9894;
reg WX9896;
reg WX9898;
reg WX9900;
reg WX9902;
reg WX9904;
reg WX9906;
reg WX9908;
reg WX9910;
reg WX9912;
reg WX9914;
reg WX9916;
reg WX9918;
reg WX9920;
reg WX9922;
reg WX9924;
reg WX9926;
reg WX9928;
reg WX9930;
reg WX9932;
reg WX9934;
reg WX9936;
reg WX9938;
reg WX9940;
reg WX9942;
reg WX9944;
reg WX9946;
reg WX9948;
reg WX9950;
reg _2301_;
reg _2302_;
reg _2303_;
reg _2304_;
reg _2305_;
reg _2306_;
reg _2307_;
reg _2308_;
reg _2309_;
reg _2310_;
reg _2311_;
reg _2312_;
reg _2313_;
reg _2314_;
reg _2315_;
reg _2316_;
reg _2317_;
reg _2318_;
reg _2319_;
reg _2320_;
reg _2321_;
reg _2322_;
reg _2323_;
reg _2324_;
reg _2325_;
reg _2326_;
reg _2327_;
reg _2328_;
reg _2329_;
reg _2330_;
reg _2331_;
reg _2332_;
reg WX10829;
reg WX10831;
reg WX10833;
reg WX10835;
reg WX10837;
reg WX10839;
reg WX10841;
reg WX10843;
reg WX10845;
reg WX10847;
reg WX10849;
reg WX10851;
reg WX10853;
reg WX10855;
reg WX10857;
reg WX10859;
reg WX10861;
reg WX10863;
reg WX10865;
reg WX10867;
reg WX10869;
reg WX10871;
reg WX10873;
reg WX10875;
reg WX10877;
reg WX10879;
reg WX10881;
reg WX10883;
reg WX10885;
reg WX10887;
reg WX10889;
reg WX10891;
reg WX10989;
reg WX10991;
reg WX10993;
reg WX10995;
reg WX10997;
reg WX10999;
reg WX11001;
reg WX11003;
reg WX11005;
reg WX11007;
reg WX11009;
reg WX11011;
reg WX11013;
reg WX11015;
reg WX11017;
reg WX11019;
reg WX11021;
reg WX11023;
reg WX11025;
reg WX11027;
reg WX11029;
reg WX11031;
reg WX11033;
reg WX11035;
reg WX11037;
reg WX11039;
reg WX11041;
reg WX11043;
reg WX11045;
reg WX11047;
reg WX11049;
reg WX11051;
reg WX11053;
reg WX11055;
reg WX11057;
reg WX11059;
reg WX11061;
reg WX11063;
reg WX11065;
reg WX11067;
reg WX11069;
reg WX11071;
reg WX11073;
reg WX11075;
reg WX11077;
reg WX11079;
reg WX11081;
reg WX11083;
reg WX11085;
reg WX11087;
reg WX11089;
reg WX11091;
reg WX11093;
reg WX11095;
reg WX11097;
reg WX11099;
reg WX11101;
reg WX11103;
reg WX11105;
reg WX11107;
reg WX11109;
reg WX11111;
reg WX11113;
reg WX11115;
reg WX11117;
reg WX11119;
reg WX11121;
reg WX11123;
reg WX11125;
reg WX11127;
reg WX11129;
reg WX11131;
reg WX11133;
reg WX11135;
reg WX11137;
reg WX11139;
reg WX11141;
reg WX11143;
reg WX11145;
reg WX11147;
reg WX11149;
reg WX11151;
reg WX11153;
reg WX11155;
reg WX11157;
reg WX11159;
reg WX11161;
reg WX11163;
reg WX11165;
reg WX11167;
reg WX11169;
reg WX11171;
reg WX11173;
reg WX11175;
reg WX11177;
reg WX11179;
reg WX11181;
reg WX11183;
reg WX11185;
reg WX11187;
reg WX11189;
reg WX11191;
reg WX11193;
reg WX11195;
reg WX11197;
reg WX11199;
reg WX11201;
reg WX11203;
reg WX11205;
reg WX11207;
reg WX11209;
reg WX11211;
reg WX11213;
reg WX11215;
reg WX11217;
reg WX11219;
reg WX11221;
reg WX11223;
reg WX11225;
reg WX11227;
reg WX11229;
reg WX11231;
reg WX11233;
reg WX11235;
reg WX11237;
reg WX11239;
reg WX11241;
reg WX11243;
reg _2333_;
reg _2334_;
reg _2335_;
reg _2336_;
reg _2337_;
reg _2338_;
reg _2339_;
reg _2340_;
reg _2341_;
reg _2342_;
reg _2343_;
reg _2344_;
reg _2345_;
reg _2346_;
reg _2347_;
reg _2348_;
reg _2349_;
reg _2350_;
reg _2351_;
reg _2352_;
reg _2353_;
reg _2354_;
reg _2355_;
reg _2356_;
reg _2357_;
reg _2358_;
reg _2359_;
reg _2360_;
reg _2361_;
reg _2362_;
reg _2363_;
reg _2364_;
wire II26071;
wire WX6414;
wire WX9613;
wire WX7987;
wire WX2450;
wire II2229;
wire II30149;
wire II2963;
wire WX8188;
wire WX3931;
wire WX7670;
wire WX6302;
wire II22919;
wire WX6164;
wire WX239;
wire WX330;
wire II3642;
wire II26018;
wire II15405;
wire II15147;
wire WX2904;
wire WX8882;
wire WX5365;
wire WX8975;
wire WX5343;
wire II14615;
wire WX3563;
wire WX8062;
wire II14260;
wire WX1525;
wire WX1406;
wire II10585;
wire WX11054;
wire II34796;
wire WX4953;
wire II2499;
wire II1988;
wire II26172;
wire II26856;
wire II26252;
wire II30929;
wire WX2627;
wire WX4973;
wire II34098;
wire WX11574;
wire WX11360;
wire WX2993;
wire WX11558;
wire II26791;
wire WX10544;
wire WX9283;
wire WX10599;
wire WX4974;
wire II18597;
wire WX5460;
wire WX8768;
wire WX11251;
wire II11517;
wire II35012;
wire WX3416;
wire II34750;
wire WX6728;
wire WX929;
wire WX10790;
wire WX5064;
wire II18100;
wire WX5449;
wire WX11506;
wire WX5280;
wire WX8596;
wire WX5285;
wire II23455;
wire WX2773;
wire WX555;
wire II30288;
wire WX3489;
wire WX2358;
wire II2801;
wire II11440;
wire WX4831;
wire II18830;
wire WX11342;
wire WX6651;
wire WX7488;
wire WX8391;
wire WX3548;
wire WX2055;
wire II34818;
wire WX11012;
wire II22850;
wire WX9078;
wire WX10766;
wire WX101;
wire II34928;
wire II30781;
wire WX5348;
wire WX2693;
wire II10883;
wire II18254;
wire WX800;
wire WX10138;
wire II30379;
wire WX9691;
wire WX3662;
wire II6735;
wire II6615;
wire II10029;
wire WX8250;
wire II11427;
wire WX2565;
wire WX8089;
wire II23667;
wire II30759;
wire WX404;
wire II2011;
wire WX7621;
wire II23645;
wire WX6095;
wire II19577;
wire WX4242;
wire WX10193;
wire WX6026;
wire WX1941;
wire II2064;
wire WX2230;
wire WX10644;
wire WX6599;
wire WX550;
wire WX2922;
wire WX3450;
wire II23569;
wire WX4873;
wire II18915;
wire WX2543;
wire WX7809;
wire WX4172;
wire WX8268;
wire II30118;
wire WX591;
wire WX901;
wire II7072;
wire WX918;
wire WX10014;
wire II35687;
wire II15314;
wire II30643;
wire WX6696;
wire II23583;
wire WX7061;
wire WX1708;
wire WX971;
wire WX10687;
wire II23207;
wire WX5086;
wire WX954;
wire II15486;
wire WX7007;
wire II30505;
wire WX11092;
wire WX10051;
wire WX7723;
wire WX8614;
wire WX10888;
wire WX10237;
wire WX1383;
wire II6009;
wire II2808;
wire WX7887;
wire II15711;
wire II3691;
wire WX10173;
wire II3444;
wire WX7817;
wire WX1050;
wire WX9695;
wire WX10524;
wire II23736;
wire II14284;
wire WX8963;
wire II18797;
wire WX3178;
wire II6901;
wire WX3175;
wire II19542;
wire II18883;
wire WX3722;
wire II14893;
wire WX2709;
wire WX8899;
wire II7695;
wire II6643;
wire WX8025;
wire WX3366;
wire WX838;
wire WX5473;
wire WX10951;
wire WX627;
wire WX4993;
wire WX3227;
wire II18273;
wire II2451;
wire WX6720;
wire II19111;
wire WX1663;
wire II27515;
wire WX11596;
wire WX7880;
wire II19730;
wire WX1553;
wire WX4297;
wire II18232;
wire II6922;
wire WX4575;
wire WX8692;
wire II30706;
wire WX631;
wire II30474;
wire II11495;
wire WX6654;
wire WX9579;
wire II30805;
wire II27290;
wire WX5316;
wire WX4350;
wire II2136;
wire II2811;
wire II14506;
wire WX5179;
wire II31563;
wire WX6741;
wire WX6365;
wire II10244;
wire WX5816;
wire WX1640;
wire II6861;
wire WX4919;
wire WX3537;
wire WX9849;
wire II3487;
wire II34980;
wire II34771;
wire II30424;
wire WX3681;
wire WX10690;
wire II14057;
wire WX508;
wire II34510;
wire WX4216;
wire WX6378;
wire WX10019;
wire WX10499;
wire WX1680;
wire WX339;
wire II31614;
wire WX8294;
wire WX2941;
wire WX936;
wire II2034;
wire WX6042;
wire WX399;
wire WX6814;
wire WX1359;
wire WX36;
wire II14359;
wire WX8670;
wire WX10471;
wire WX2497;
wire WX4328;
wire WX10669;
wire WX9036;
wire WX4613;
wire II31689;
wire WX8772;
wire WX5910;
wire II18759;
wire WX378;
wire WX8474;
wire II6225;
wire II10470;
wire II22749;
wire II10485;
wire WX10925;
wire WX5264;
wire WX5760;
wire WX4438;
wire WX2909;
wire II26157;
wire II10341;
wire II22476;
wire WX9355;
wire WX1334;
wire II10834;
wire II31193;
wire II18750;
wire WX9547;
wire WX6749;
wire WX6434;
wire WX5559;
wire II27109;
wire WX10549;
wire WX7415;
wire WX5199;
wire WX10492;
wire II18008;
wire II31670;
wire II18285;
wire WX8892;
wire WX4899;
wire II2654;
wire WX6868;
wire WX6527;
wire II22680;
wire II6156;
wire WX10093;
wire WX7837;
wire II31256;
wire WX225;
wire WX8376;
wire WX7195;
wire WX7800;
wire II3485;
wire II18211;
wire WX8973;
wire WX8855;
wire WX10272;
wire WX4603;
wire II22423;
wire II30316;
wire WX3207;
wire WX6977;
wire WX6926;
wire WX2093;
wire II6031;
wire WX5121;
wire WX4781;
wire II18567;
wire WX9913;
wire II11337;
wire WX9227;
wire II34686;
wire II26692;
wire WX2732;
wire WX6243;
wire II19412;
wire WX6078;
wire II27553;
wire WX4894;
wire WX1807;
wire WX605;
wire WX10386;
wire WX4854;
wire WX3033;
wire WX597;
wire II10184;
wire II26733;
wire WX164;
wire II18481;
wire II26822;
wire II14159;
wire II19660;
wire WX6252;
wire II10647;
wire WX6153;
wire II3131;
wire WX10295;
wire II18192;
wire WX11482;
wire WX6730;
wire II18373;
wire WX8805;
wire WX7591;
wire II27186;
wire WX5572;
wire WX4317;
wire WX3797;
wire II35094;
wire WX998;
wire II18502;
wire II2142;
wire WX5020;
wire WX8246;
wire II2793;
wire WX11531;
wire II10292;
wire WX7669;
wire WX4944;
wire WX11529;
wire II10269;
wire WX3482;
wire II2422;
wire II30898;
wire II27714;
wire WX11326;
wire WX11369;
wire WX5982;
wire WX9741;
wire WX3074;
wire II22045;
wire WX9412;
wire II19556;
wire WX9382;
wire WX2729;
wire WX844;
wire II19074;
wire II22113;
wire WX2787;
wire WX5104;
wire WX10041;
wire WX4117;
wire II14747;
wire WX10907;
wire WX7942;
wire WX10446;
wire WX9131;
wire II22697;
wire WX10146;
wire WX5832;
wire WX9115;
wire WX7971;
wire WX4579;
wire WX6789;
wire WX6197;
wire II10604;
wire WX416;
wire WX397;
wire WX4994;
wire WX6791;
wire WX5552;
wire WX10239;
wire II35548;
wire II34136;
wire II10363;
wire WX4109;
wire II14522;
wire WX9501;
wire II7554;
wire II27587;
wire II34989;
wire WX4933;
wire WX4033;
wire II22538;
wire WX10734;
wire WX6384;
wire WX5737;
wire WX1910;
wire WX9797;
wire WX90;
wire WX2005;
wire WX6577;
wire WX6326;
wire II35432;
wire II6325;
wire WX328;
wire WX2391;
wire II31738;
wire WX1843;
wire WX9260;
wire WX10990;
wire II19449;
wire WX8988;
wire WX11287;
wire II3521;
wire II15629;
wire WX6371;
wire WX2511;
wire WX5938;
wire WX4663;
wire II18921;
wire WX4122;
wire II18195;
wire WX8086;
wire WX7293;
wire WX1148;
wire WX6422;
wire WX1697;
wire WX6348;
wire WX5185;
wire WX266;
wire WX9313;
wire WX7852;
wire WX8028;
wire II23118;
wire WX5797;
wire WX850;
wire II7633;
wire WX3754;
wire II22616;
wire WX6508;
wire II30533;
wire WX8852;
wire WX10264;
wire WX5425;
wire II10666;
wire WX10065;
wire WX234;
wire WX3691;
wire II23378;
wire WX6101;
wire WX5794;
wire WX5588;
wire WX9026;
wire WX10116;
wire WX3940;
wire WX8494;
wire WX2364;
wire II35132;
wire WX4451;
wire II14807;
wire WX3996;
wire II10695;
wire II22190;
wire WX11605;
wire II10919;
wire II34275;
wire WX2294;
wire II27615;
wire II6566;
wire WX435;
wire WX5662;
wire II3704;
wire WX5765;
wire WX74;
wire WX8146;
wire WX1204;
wire II27121;
wire WX6260;
wire WX5755;
wire II23517;
wire II34739;
wire WX1935;
wire WX6130;
wire II15340;
wire II18993;
wire II3514;
wire II2865;
wire WX9214;
wire II14236;
wire WX4826;
wire WX1496;
wire II22129;
wire WX4807;
wire WX10945;
wire WX3598;
wire WX7921;
wire II26391;
wire WX5044;
wire WX1254;
wire WX1961;
wire II18929;
wire WX5924;
wire II7682;
wire WX8220;
wire WX7522;
wire WX2141;
wire WX6622;
wire WX9979;
wire II11496;
wire II31115;
wire WX1388;
wire WX11242;
wire II10115;
wire WX3787;
wire WX1931;
wire WX7231;
wire II11713;
wire WX6294;
wire II22965;
wire WX4811;
wire WX5173;
wire WX3613;
wire II26330;
wire WX10830;
wire WX1629;
wire WX7451;
wire WX5750;
wire WX2370;
wire II10772;
wire WX5227;
wire WX1506;
wire WX9460;
wire II10223;
wire WX10968;
wire II26698;
wire WX226;
wire WX10828;
wire WX643;
wire WX6442;
wire WX3864;
wire WX287;
wire WX2896;
wire II22874;
wire II15367;
wire WX3214;
wire II30350;
wire WX7439;
wire II34911;
wire II14328;
wire WX4336;
wire WX7253;
wire II6528;
wire WX3532;
wire II26195;
wire II10633;
wire II7703;
wire WX3751;
wire WX11086;
wire II22036;
wire WX2378;
wire WX9262;
wire WX2546;
wire WX9470;
wire II22600;
wire II6589;
wire II14631;
wire WX11459;
wire WX10567;
wire WX6677;
wire WX10808;
wire WX7794;
wire II34221;
wire II7332;
wire WX5729;
wire II30187;
wire WX1021;
wire WX7299;
wire II2043;
wire II22316;
wire II26352;
wire WX2765;
wire II26412;
wire II18444;
wire WX6490;
wire WX1431;
wire II26702;
wire WX4519;
wire II34082;
wire WX7039;
wire WX7032;
wire II26574;
wire II14962;
wire WX10778;
wire II19514;
wire WX1573;
wire WX3236;
wire II18099;
wire II2343;
wire II2104;
wire WX6234;
wire II2328;
wire II22307;
wire II2873;
wire WX315;
wire WX4516;
wire II30580;
wire WX10651;
wire II11323;
wire WX10219;
wire WX10323;
wire II34293;
wire II11244;
wire II35223;
wire WX5492;
wire II34057;
wire WX3670;
wire II30658;
wire WX8956;
wire WX9208;
wire II34463;
wire II26629;
wire II15419;
wire II18425;
wire WX8715;
wire II2368;
wire WX7391;
wire WX4761;
wire II6234;
wire II18939;
wire II10973;
wire II22810;
wire WX1227;
wire WX64;
wire II26313;
wire II10308;
wire II2266;
wire WX4204;
wire WX5331;
wire WX9181;
wire WX2466;
wire II15275;
wire II6366;
wire WX11351;
wire WX11308;
wire II30542;
wire WX11006;
wire WX6672;
wire II6971;
wire WX8915;
wire WX3648;
wire II26531;
wire II14392;
wire II27265;
wire II3470;
wire WX6183;
wire WX1053;
wire II3365;
wire WX2246;
wire II26265;
wire II18388;
wire WX138;
wire WX11512;
wire WX420;
wire WX4870;
wire II34631;
wire WX8139;
wire WX10425;
wire II19690;
wire WX9524;
wire WX4152;
wire II6124;
wire WX1905;
wire WX2899;
wire WX1712;
wire WX11614;
wire WX10899;
wire WX4683;
wire WX2782;
wire WX7603;
wire WX6887;
wire II14149;
wire WX6686;
wire WX2745;
wire II34724;
wire II14538;
wire II2647;
wire WX9100;
wire WX2273;
wire WX9370;
wire II15509;
wire II35554;
wire II30628;
wire II18087;
wire II30598;
wire WX1483;
wire WX4129;
wire WX6224;
wire WX4545;
wire WX1069;
wire WX1111;
wire II22941;
wire WX7090;
wire WX8204;
wire II10021;
wire WX11156;
wire WX8618;
wire II34197;
wire WX10642;
wire WX2930;
wire WX602;
wire II22935;
wire II6025;
wire II35315;
wire II11453;
wire WX534;
wire WX2482;
wire II3416;
wire II18403;
wire WX11277;
wire II11596;
wire II2787;
wire II10678;
wire WX10467;
wire II22711;
wire II19498;
wire WX2663;
wire WX2925;
wire II34399;
wire II26994;
wire II18409;
wire II18402;
wire II6281;
wire WX7481;
wire WX6246;
wire WX4843;
wire II14785;
wire II35276;
wire WX2495;
wire WX10285;
wire WX10404;
wire WX1514;
wire WX2469;
wire WX5900;
wire II7647;
wire WX7775;
wire WX6955;
wire WX6540;
wire II6467;
wire II31386;
wire WX9425;
wire WX2657;
wire II14647;
wire WX6896;
wire WX1894;
wire II34811;
wire WX3096;
wire WX2978;
wire WX10788;
wire II22322;
wire II19085;
wire II34400;
wire WX2413;
wire WX656;
wire WX10616;
wire WX5475;
wire WX2224;
wire WX458;
wire WX9432;
wire WX8466;
wire II31477;
wire II30908;
wire WX2428;
wire WX9670;
wire WX5069;
wire II34959;
wire II26779;
wire WX3009;
wire WX3908;
wire II26877;
wire WX7375;
wire WX9389;
wire II18575;
wire II27560;
wire II35575;
wire WX9342;
wire II19112;
wire WX6291;
wire WX8252;
wire WX3542;
wire WX6715;
wire II30457;
wire WX7519;
wire WX1031;
wire WX1165;
wire WX5743;
wire II31724;
wire II6522;
wire WX2271;
wire WX1324;
wire II18535;
wire II6209;
wire WX5095;
wire WX251;
wire WX4332;
wire II6575;
wire WX9960;
wire WX4199;
wire WX10636;
wire II3655;
wire WX465;
wire II10279;
wire WX9633;
wire II31426;
wire WX471;
wire WX6946;
wire WX6820;
wire WX3318;
wire WX7568;
wire WX7097;
wire WX6526;
wire II7241;
wire WX8919;
wire II18496;
wire II2661;
wire WX10561;
wire WX1936;
wire II10129;
wire II26027;
wire WX10078;
wire II26841;
wire WX10769;
wire WX8438;
wire WX6796;
wire WX7995;
wire II10384;
wire WX1633;
wire WX11473;
wire WX1501;
wire WX3266;
wire WX8229;
wire WX5676;
wire WX10157;
wire WX366;
wire II22571;
wire WX85;
wire WX7370;
wire II19529;
wire WX6333;
wire WX5377;
wire WX6583;
wire WX3604;
wire WX8564;
wire WX8214;
wire WX6492;
wire WX9320;
wire WX6173;
wire II18595;
wire WX337;
wire WX6930;
wire II30211;
wire WX3610;
wire WX4014;
wire II30621;
wire WX3964;
wire WX5457;
wire WX3852;
wire WX9553;
wire WX5878;
wire WX4256;
wire WX7653;
wire WX11030;
wire II14794;
wire WX2460;
wire WX1987;
wire II18413;
wire WX5242;
wire II10270;
wire WX7675;
wire WX10988;
wire WX7108;
wire WX108;
wire II10237;
wire II35497;
wire II35237;
wire II34160;
wire WX6763;
wire WX7606;
wire WX9705;
wire WX7755;
wire II18893;
wire II22077;
wire II14382;
wire II26988;
wire WX5232;
wire WX6281;
wire WX4924;
wire II22300;
wire WX114;
wire II2374;
wire WX2671;
wire WX7711;
wire WX648;
wire II35340;
wire II14321;
wire II31348;
wire WX2137;
wire II2840;
wire II18488;
wire WX9254;
wire II30674;
wire WX6129;
wire WX2593;
wire II22586;
wire WX8053;
wire WX5169;
wire II14924;
wire WX265;
wire II22170;
wire II18527;
wire WX7045;
wire WX5531;
wire WX9595;
wire WX3042;
wire WX2928;
wire WX9988;
wire WX961;
wire WX4922;
wire II31154;
wire WX666;
wire WX10554;
wire II31114;
wire II26367;
wire II2555;
wire WX4984;
wire WX7181;
wire WX9621;
wire II19191;
wire WX6605;
wire II34678;
wire II19385;
wire II31205;
wire II27565;
wire WX4541;
wire WX2798;
wire WX3636;
wire II10323;
wire WX2912;
wire WX6702;
wire WX5602;
wire WX4880;
wire WX10288;
wire WX10045;
wire WX7803;
wire II10557;
wire WX5624;
wire WX3066;
wire WX856;
wire WX2705;
wire II14507;
wire II10013;
wire WX10211;
wire WX9379;
wire WX10897;
wire WX2916;
wire WX9688;
wire II26826;
wire II26807;
wire WX2717;
wire WX4276;
wire II26933;
wire II31543;
wire WX8389;
wire II7436;
wire WX7468;
wire WX9374;
wire II23195;
wire II34579;
wire II14754;
wire WX2194;
wire II18511;
wire WX2252;
wire WX5019;
wire WX4062;
wire II26033;
wire II18109;
wire WX11164;
wire WX4343;
wire II6674;
wire II22291;
wire WX6609;
wire II7653;
wire WX9673;
wire WX924;
wire WX5370;
wire WX2523;
wire WX2959;
wire WX9873;
wire WX175;
wire II6010;
wire WX564;
wire II11651;
wire WX2288;
wire II34765;
wire WX2815;
wire WX411;
wire WX10962;
wire II14373;
wire WX2524;
wire WX2557;
wire WX2647;
wire II35003;
wire WX2823;
wire II23456;
wire II6784;
wire WX10513;
wire II15669;
wire II30161;
wire II34556;
wire WX3556;
wire WX8552;
wire WX1476;
wire WX10813;
wire WX4965;
wire WX3937;
wire WX7161;
wire II6550;
wire II30342;
wire II10222;
wire WX6568;
wire II11272;
wire WX6563;
wire WX11450;
wire WX2689;
wire II6217;
wire WX4002;
wire II18799;
wire II14500;
wire II35561;
wire WX1286;
wire WX7496;
wire WX8094;
wire WX1116;
wire WX4132;
wire WX3723;
wire II26647;
wire II27003;
wire WX7627;
wire II22083;
wire II10161;
wire II2399;
wire WX7872;
wire WX5894;
wire II34455;
wire WX987;
wire II3208;
wire WX3841;
wire WX6767;
wire WX3185;
wire WX3571;
wire WX2457;
wire II6512;
wire II6350;
wire WX4487;
wire II34508;
wire II22773;
wire WX7612;
wire WX978;
wire WX1811;
wire II14413;
wire WX2368;
wire WX11116;
wire WX557;
wire WX11210;
wire II6535;
wire WX2234;
wire WX1537;
wire II14606;
wire WX1105;
wire WX10932;
wire WX1464;
wire II26916;
wire II26769;
wire WX613;
wire II31399;
wire II26383;
wire WX5522;
wire WX5070;
wire II22137;
wire WX1542;
wire II22446;
wire II6800;
wire WX4467;
wire II14120;
wire WX3657;
wire WX6818;
wire WX5350;
wire WX6832;
wire II22981;
wire II30069;
wire II10331;
wire WX2198;
wire WX514;
wire WX5297;
wire II2351;
wire WX5453;
wire WX2699;
wire II30285;
wire II23482;
wire WX11310;
wire WX9271;
wire WX5397;
wire WX2999;
wire II10619;
wire WX10347;
wire WX6668;
wire WX3412;
wire WX4961;
wire WX6304;
wire WX8339;
wire WX4937;
wire WX9647;
wire WX3491;
wire WX8994;
wire II26165;
wire II3507;
wire II2274;
wire WX1398;
wire II35262;
wire WX3478;
wire WX6709;
wire WX9512;
wire WX5011;
wire WX8366;
wire WX7553;
wire WX7862;
wire II15705;
wire WX8662;
wire WX2109;
wire II31745;
wire II11311;
wire II10317;
wire II26228;
wire II31282;
wire WX332;
wire II34998;
wire WX10764;
wire WX7631;
wire WX11337;
wire WX1565;
wire WX2589;
wire II34151;
wire WX10529;
wire WX1459;
wire WX6426;
wire WX11258;
wire WX8578;
wire WX3927;
wire II23144;
wire WX8902;
wire WX7464;
wire WX9721;
wire II30769;
wire WX10399;
wire WX9937;
wire WX6484;
wire WX10634;
wire II14096;
wire WX3406;
wire II6473;
wire WX1602;
wire WX2308;
wire WX9094;
wire WX11273;
wire WX6627;
wire WX7508;
wire WX1260;
wire II14979;
wire WX5860;
wire WX6801;
wire WX6517;
wire II19347;
wire II6978;
wire WX10682;
wire II14909;
wire WX4407;
wire WX6775;
wire WX9250;
wire WX674;
wire II26717;
wire WX8000;
wire WX10292;
wire WX7578;
wire WX9452;
wire WX7087;
wire WX8244;
wire WX7586;
wire WX7529;
wire II19371;
wire WX1599;
wire WX4253;
wire II2849;
wire II6240;
wire WX2756;
wire II10263;
wire WX10530;
wire WX10928;
wire WX6134;
wire WX11028;
wire WX2214;
wire WX794;
wire II14724;
wire WX3703;
wire WX6482;
wire II14466;
wire II26142;
wire WX212;
wire WX8009;
wire II2429;
wire WX3979;
wire II6398;
wire WX5646;
wire WX9504;
wire WX431;
wire WX931;
wire WX2189;
wire WX3221;
wire II34269;
wire II18745;
wire WX5776;
wire WX9687;
wire II30362;
wire II27082;
wire WX8516;
wire II22469;
wire WX5392;
wire II22864;
wire WX2869;
wire WX9220;
wire II2114;
wire II3183;
wire II30813;
wire II30426;
wire II34982;
wire WX5055;
wire II14414;
wire WX7647;
wire WX7189;
wire WX3982;
wire WX690;
wire WX4042;
wire WX98;
wire II10347;
wire WX1475;
wire II35541;
wire WX9583;
wire WX3442;
wire II10137;
wire II35171;
wire WX6880;
wire II2252;
wire WX4104;
wire WX2320;
wire II31453;
wire WX5805;
wire II26887;
wire WX8406;
wire WX10757;
wire WX279;
wire II35737;
wire WX6353;
wire WX10061;
wire WX4221;
wire II18630;
wire II6002;
wire WX4036;
wire II34618;
wire WX10713;
wire II30433;
wire WX10392;
wire II34827;
wire WX3330;
wire WX10660;
wire WX10184;
wire II35510;
wire WX11404;
wire WX9005;
wire II30047;
wire WX8817;
wire WX11489;
wire WX5642;
wire WX1687;
wire II30386;
wire II22523;
wire WX2800;
wire II6560;
wire WX5544;
wire WX8330;
wire II7618;
wire II18660;
wire II3549;
wire WX7664;
wire II3492;
wire WX9144;
wire II6715;
wire II19648;
wire WX7442;
wire II15470;
wire WX7215;
wire II35584;
wire II18853;
wire II19124;
wire WX1795;
wire WX4324;
wire WX635;
wire WX5561;
wire WX8171;
wire II10051;
wire WX4301;
wire WX2504;
wire WX4245;
wire WX1679;
wire WX10355;
wire II18240;
wire WX4759;
wire II7675;
wire II26135;
wire WX8742;
wire II23728;
wire II31640;
wire WX8340;
wire WX6315;
wire WX8620;
wire II15069;
wire WX4076;
wire WX1249;
wire II10354;
wire WX10906;
wire II30325;
wire WX572;
wire II34803;
wire WX9563;
wire WX8382;
wire II31296;
wire WX9340;
wire WX8198;
wire WX1883;
wire II18667;
wire WX4563;
wire II30186;
wire WX2636;
wire WX9735;
wire II15459;
wire WX4454;
wire WX3744;
wire II14313;
wire II10874;
wire WX10103;
wire II6954;
wire II2501;
wire WX10536;
wire WX6515;
wire WX1502;
wire WX2579;
wire II23644;
wire WX45;
wire WX2919;
wire II18248;
wire II34384;
wire II18440;
wire II14258;
wire II18156;
wire II14933;
wire WX1643;
wire II22841;
wire II11630;
wire II26895;
wire WX3717;
wire WX1736;
wire WX5920;
wire II11361;
wire II14150;
wire II26304;
wire II7575;
wire II26056;
wire WX9867;
wire WX10576;
wire II22657;
wire WX894;
wire WX10121;
wire WX9316;
wire II30704;
wire WX6084;
wire II14353;
wire WX4983;
wire WX230;
wire WX4235;
wire WX9173;
wire WX5111;
wire WX8574;
wire II3633;
wire II10570;
wire II3417;
wire WX10976;
wire II19269;
wire WX308;
wire WX3201;
wire WX6081;
wire II10609;
wire II6286;
wire II30961;
wire II26113;
wire WX7473;
wire II22330;
wire WX8942;
wire II10596;
wire WX4095;
wire II22463;
wire WX2937;
wire WX3626;
wire WX1170;
wire WX3171;
wire WX9096;
wire WX68;
wire WX9895;
wire II34748;
wire II5995;
wire II35710;
wire WX4186;
wire II31529;
wire WX10692;
wire WX2059;
wire WX1004;
wire WX5321;
wire WX11455;
wire WX10466;
wire II14172;
wire WX1995;
wire WX1837;
wire WX1919;
wire WX3010;
wire WX3621;
wire WX2673;
wire WX5032;
wire WX6585;
wire II18588;
wire WX10672;
wire WX4423;
wire WX1716;
wire WX3136;
wire II6962;
wire WX8778;
wire WX10281;
wire WX134;
wire II26321;
wire WX2720;
wire II3592;
wire WX3920;
wire WX2812;
wire WX6637;
wire II30395;
wire WX4507;
wire II14436;
wire II2203;
wire WX354;
wire II10741;
wire WX2776;
wire WX10154;
wire WX10009;
wire WX6468;
wire II14872;
wire WX9543;
wire II23497;
wire II3338;
wire II2514;
wire II35158;
wire II26295;
wire II31635;
wire WX2849;
wire WX221;
wire WX9194;
wire II34525;
wire WX3878;
wire WX834;
wire WX9971;
wire WX8178;
wire II30077;
wire II7540;
wire WX1758;
wire WX11148;
wire WX1744;
wire II26058;
wire WX1771;
wire WX9403;
wire WX53;
wire WX10656;
wire II35694;
wire WX9475;
wire WX1370;
wire II2854;
wire WX7078;
wire II30869;
wire WX9223;
wire WX5555;
wire II6899;
wire WX8706;
wire WX8325;
wire II22378;
wire II18812;
wire WX9292;
wire II27608;
wire WX5653;
wire WX4472;
wire II3234;
wire WX10199;
wire WX1582;
wire WX8920;
wire WX8760;
wire II30502;
wire II30201;
wire WX8132;
wire WX5410;
wire II6506;
wire II27670;
wire WX9466;
wire WX6758;
wire WX4903;
wire II35626;
wire WX7843;
wire WX9193;
wire II2059;
wire II6497;
wire WX4510;
wire WX6983;
wire WX3595;
wire WX9186;
wire II30874;
wire WX3007;
wire II2065;
wire WX10451;
wire WX1077;
wire II26584;
wire II14397;
wire WX2877;
wire WX9959;
wire II18187;
wire II14800;
wire WX8484;
wire II26452;
wire II18130;
wire II10920;
wire WX6368;
wire II7689;
wire II22122;
wire II19255;
wire II10030;
wire WX6337;
wire II22989;
wire II30798;
wire WX8656;
wire WX2473;
wire WX2349;
wire WX10622;
wire II6116;
wire II30070;
wire WX3696;
wire II34662;
wire II6374;
wire WX8239;
wire WX5043;
wire WX7865;
wire WX1487;
wire II22817;
wire WX8066;
wire WX1167;
wire WX2621;
wire WX3634;
wire WX1906;
wire II27331;
wire II2586;
wire WX10220;
wire WX3191;
wire WX8354;
wire WX6751;
wire II3529;
wire WX8879;
wire WX5733;
wire II18055;
wire WX1650;
wire WX242;
wire II22518;
wire WX2393;
wire II15354;
wire WX11415;
wire II2439;
wire WX1821;
wire WX184;
wire WX7702;
wire II26505;
wire II7356;
wire WX323;
wire WX3803;
wire II6892;
wire II7371;
wire WX1393;
wire WX8602;
wire WX9243;
wire WX6846;
wire WX2965;
wire WX4955;
wire WX994;
wire WX8161;
wire WX9435;
wire WX2768;
wire II18117;
wire II2824;
wire WX10134;
wire II6457;
wire II18327;
wire WX6912;
wire WX2229;
wire WX5882;
wire WX6878;
wire WX10089;
wire WX6454;
wire WX5284;
wire II3558;
wire WX140;
wire WX5161;
wire II30738;
wire II2889;
wire WX346;
wire II31558;
wire WX131;
wire II30962;
wire II26398;
wire WX4649;
wire WX10161;
wire WX6157;
wire WX3120;
wire WX6444;
wire II35652;
wire II19319;
wire II3261;
wire WX10255;
wire WX9992;
wire II22764;
wire II10371;
wire WX11299;
wire II14776;
wire WX8168;
wire II30233;
wire II18332;
wire WX9483;
wire II18613;
wire II18227;
wire II27473;
wire WX5824;
wire WX7075;
wire WX447;
wire WX10311;
wire II7228;
wire II6708;
wire WX2550;
wire WX4727;
wire WX2445;
wire WX5251;
wire II2530;
wire WX2035;
wire II6938;
wire WX1242;
wire II6806;
wire WX10315;
wire WX5290;
wire II22740;
wire II14563;
wire II27200;
wire II34492;
wire WX6214;
wire II26282;
wire WX7369;
wire WX197;
wire II14290;
wire II2746;
wire II30951;
wire WX4801;
wire II10108;
wire WX7856;
wire II34336;
wire WX2437;
wire WX348;
wire WX1352;
wire WX4415;
wire II18234;
wire WX5289;
wire WX3727;
wire WX1891;
wire II27657;
wire WX9322;
wire WX3386;
wire WX6219;
wire WX272;
wire WX9108;
wire WX2342;
wire WX81;
wire WX11424;
wire II22206;
wire II10152;
wire II22346;
wire WX9332;
wire WX1150;
wire WX9156;
wire II14064;
wire II27097;
wire WX8811;
wire II10062;
wire WX5195;
wire WX6347;
wire WX7543;
wire II2398;
wire WX2408;
wire II10671;
wire WX5134;
wire WX2503;
wire WX1010;
wire WX8669;
wire WX577;
wire WX4460;
wire WX5007;
wire II15650;
wire WX1235;
wire WX4192;
wire WX2748;
wire WX1094;
wire II6854;
wire WX1929;
wire WX3108;
wire WX10872;
wire WX6969;
wire II2576;
wire WX3581;
wire II18846;
wire II22950;
wire WX1886;
wire WX10754;
wire II10432;
wire II18673;
wire II14663;
wire WX3619;
wire WX7913;
wire WX1752;
wire WX6450;
wire II6420;
wire II2591;
wire WX9954;
wire WX7071;
wire WX4399;
wire II27663;
wire WX4687;
wire II14042;
wire WX7396;
wire II18960;
wire WX5246;
wire II2640;
wire II30349;
wire WX4877;
wire WX5631;
wire II14950;
wire WX11586;
wire II15301;
wire II23091;
wire WX1060;
wire II19436;
wire II23639;
wire WX2853;
wire WX1212;
wire WX4142;
wire II6054;
wire WX7691;
wire WX6267;
wire II30254;
wire WX5089;
wire WX11184;
wire WX7938;
wire WX9302;
wire WX3023;
wire II14847;
wire II2617;
wire WX7698;
wire II26608;
wire II22759;
wire WX1198;
wire WX6785;
wire WX3936;
wire WX1136;
wire WX9571;
wire WX1300;
wire WX8968;
wire WX11549;
wire WX1877;
wire WX10723;
wire II30791;
wire II34212;
wire WX7135;
wire WX384;
wire II30194;
wire II34206;
wire II26978;
wire WX1797;
wire WX3156;
wire WX2886;
wire II35289;
wire II6141;
wire WX6230;
wire WX2803;
wire WX7456;
wire II30087;
wire II30177;
wire WX3028;
wire II22898;
wire II34708;
wire WX3145;
wire WX5507;
wire II22387;
wire WX5052;
wire WX293;
wire WX3833;
wire WX4363;
wire WX6645;
wire WX8420;
wire WX7743;
wire WX11463;
wire II14089;
wire II35184;
wire II35680;
wire II35752;
wire WX3342;
wire WX776;
wire II2088;
wire II14142;
wire WX5489;
wire WX9016;
wire WX11062;
wire II22090;
wire WX4669;
wire II11233;
wire WX9062;
wire WX7333;
wire II18490;
wire II7482;
wire WX4857;
wire II34874;
wire II30518;
wire WX10965;
wire WX980;
wire II18945;
wire WX10596;
wire WX6022;
wire II2415;
wire WX3522;
wire WX1762;
wire WX9357;
wire WX7727;
wire WX4084;
wire WX598;
wire WX6549;
wire WX3732;
wire WX3494;
wire WX9235;
wire WX8032;
wire II7149;
wire II14011;
wire WX11246;
wire WX4149;
wire WX5517;
wire II23540;
wire II6428;
wire WX10708;
wire II14018;
wire II30993;
wire II10899;
wire WX6827;
wire WX11302;
wire II18683;
wire WX9667;
wire WX5638;
wire WX4695;
wire II7161;
wire II3661;
wire WX718;
wire WX9967;
wire II14544;
wire II34973;
wire II30417;
wire WX5300;
wire WX8073;
wire WX6202;
wire WX3529;
wire II30272;
wire WX5635;
wire WX8108;
wire WX6893;
wire WX4294;
wire WX5502;
wire II14740;
wire WX8844;
wire II2313;
wire WX5327;
wire WX4050;
wire II23660;
wire WX5952;
wire WX8191;
wire WX5210;
wire WX5512;
wire WX2335;
wire II31513;
wire WX8058;
wire II26838;
wire II22624;
wire WX2216;
wire WX3679;
wire II35353;
wire II22215;
wire WX6538;
wire WX3784;
wire WX2831;
wire II27110;
wire II2547;
wire WX4308;
wire WX11449;
wire WX2401;
wire WX5593;
wire II34026;
wire II14049;
wire WX10031;
wire WX3322;
wire II35611;
wire WX8351;
wire II30937;
wire WX10958;
wire II30519;
wire WX10785;
wire WX2973;
wire WX4539;
wire WX1348;
wire WX3580;
wire WX8900;
wire II18969;
wire II18163;
wire II18737;
wire II7507;
wire WX11375;
wire WX10504;
wire WX5239;
wire WX4890;
wire II15328;
wire WX6280;
wire II26817;
wire II34941;
wire II34433;
wire WX8151;
wire WX1427;
wire WX1509;
wire WX9532;
wire II14127;
wire WX1016;
wire WX4267;
wire II14337;
wire WX9032;
wire WX10073;
wire WX8298;
wire WX2642;
wire WX7163;
wire WX4281;
wire WX4915;
wire WX3654;
wire II7096;
wire WX4250;
wire II35209;
wire WX10475;
wire II22718;
wire WX8398;
wire WX1889;
wire WX8276;
wire II14253;
wire II23652;
wire WX3012;
wire II34755;
wire WX39;
wire WX3628;
wire II30868;
wire WX4786;
wire WX10737;
wire II18179;
wire WX6573;
wire WX8759;
wire II14190;
wire WX8082;
wire II2500;
wire WX5842;
wire WX10496;
wire WX6256;
wire II14105;
wire II2934;
wire WX6614;
wire II22500;
wire WX5498;
wire II18451;
wire WX8085;
wire II23429;
wire WX8044;
wire WX11202;
wire WX7974;
wire WX6821;
wire II6606;
wire WX6148;
wire II26066;
wire WX9110;
wire II23259;
wire II15641;
wire WX6923;
wire II23504;
wire II14367;
wire WX8022;
wire WX10040;
wire WX255;
wire WX309;
wire II26497;
wire WX5742;
wire WX2448;
wire WX154;
wire WX6920;
wire II27149;
wire II23196;
wire II14250;
wire WX466;
wire WX6839;
wire II2561;
wire WX6192;
wire WX4913;
wire WX4493;
wire II30039;
wire WX7907;
wire II9996;
wire WX10718;
wire WX7093;
wire WX4026;
wire WX10631;
wire WX2850;
wire WX7381;
wire II3586;
wire II18936;
wire WX7380;
wire WX10994;
wire WX10126;
wire II18792;
wire WX6318;
wire WX7976;
wire II30032;
wire II30304;
wire WX2725;
wire WX7423;
wire II34779;
wire WX9346;
wire WX10964;
wire WX8931;
wire II6845;
wire II2151;
wire II22787;
wire WX6973;
wire WX10442;
wire WX6176;
wire WX10755;
wire II15643;
wire WX6744;
wire WX311;
wire WX8938;
wire WX2839;
wire WX7371;
wire WX10389;
wire WX4850;
wire WX7595;
wire WX7924;
wire II10759;
wire II34276;
wire WX8860;
wire II14027;
wire II22415;
wire WX3203;
wire WX670;
wire II22786;
wire WX7418;
wire WX848;
wire II26763;
wire WX9119;
wire II30333;
wire II6969;
wire WX1368;
wire WX4228;
wire WX6987;
wire WX2001;
wire WX5100;
wire II30883;
wire WX4793;
wire WX3002;
wire II22811;
wire WX5431;
wire II14311;
wire WX3946;
wire WX4260;
wire II14422;
wire II7396;
wire WX11477;
wire WX8965;
wire WX9398;
wire WX2161;
wire WX8047;
wire II11063;
wire WX2764;
wire WX706;
wire WX1685;
wire WX3559;
wire II6233;
wire II2560;
wire WX10415;
wire WX2631;
wire WX1100;
wire WX3774;
wire WX790;
wire WX6593;
wire WX9134;
wire WX10018;
wire WX5219;
wire II3157;
wire WX9976;
wire WX4599;
wire WX3950;
wire II26373;
wire II11582;
wire WX4553;
wire WX6309;
wire WX4703;
wire WX3163;
wire II30527;
wire WX1920;
wire WX4930;
wire WX7665;
wire II18754;
wire II10859;
wire WX5986;
wire II22152;
wire II26335;
wire II34477;
wire WX2538;
wire WX8801;
wire WX3668;
wire WX2375;
wire WX1316;
wire WX9557;
wire II6527;
wire II23695;
wire II22641;
wire WX10794;
wire WX7657;
wire WX2043;
wire WX5836;
wire WX9883;
wire WX3793;
wire II35645;
wire WX6344;
wire WX6795;
wire WX1020;
wire WX8195;
wire WX6075;
wire WX2619;
wire II14678;
wire II34367;
wire WX7869;
wire II23546;
wire WX11538;
wire II6766;
wire WX6030;
wire WX5772;
wire WX4861;
wire WX6028;
wire WX3078;
wire WX816;
wire WX9276;
wire WX7823;
wire WX8540;
wire II14717;
wire WX11554;
wire WX4211;
wire WX9386;
wire WX8796;
wire II15678;
wire WX6375;
wire WX4313;
wire WX4354;
wire WX3685;
wire WX3993;
wire WX5362;
wire WX10741;
wire WX6776;
wire II10944;
wire II11193;
wire II18024;
wire WX8470;
wire II27532;
wire WX610;
wire II6303;
wire II2158;
wire II30760;
wire WX11364;
wire WX8809;
wire II34538;
wire II6736;
wire WX6724;
wire WX7890;
wire WX1521;
wire WX5966;
wire WX9757;
wire II10579;
wire II14761;
wire WX6504;
wire WX7735;
wire II14531;
wire WX7683;
wire II23182;
wire II2942;
wire WX7349;
wire WX105;
wire II11487;
wire WX8610;
wire II14407;
wire II6134;
wire II14485;
wire WX5047;
wire II26924;
wire WX11100;
wire WX2319;
wire WX1030;
wire WX11590;
wire WX10519;
wire II34337;
wire II18310;
wire II34680;
wire WX5496;
wire II18317;
wire II18544;
wire WX10935;
wire II31218;
wire WX569;
wire WX3090;
wire II18335;
wire WX4979;
wire II34353;
wire WX162;
wire WX5528;
wire WX9070;
wire WX5081;
wire II11154;
wire WX6328;
wire II35013;
wire II18506;
wire WX5476;
wire WX3799;
wire WX8752;
wire II11206;
wire II26884;
wire II30765;
wire II14900;
wire WX2431;
wire WX7957;
wire WX3804;
wire II15573;
wire WX2297;
wire II14113;
wire WX3159;
wire WX9017;
wire II34106;
wire WX5340;
wire WX7100;
wire WX1074;
wire II18869;
wire II30052;
wire WX9444;
wire WX4443;
wire WX2794;
wire WX2537;
wire WX8142;
wire II6165;
wire II11686;
wire II34484;
wire II31244;
wire II2220;
wire WX5191;
wire WX10979;
wire II3696;
wire II6580;
wire WX10507;
wire WX10060;
wire WX3591;
wire II30381;
wire II2406;
wire WX4239;
wire WX453;
wire II22640;
wire WX7637;
wire II11666;
wire WX6091;
wire WX7883;
wire II10201;
wire II3570;
wire WX8784;
wire WX551;
wire WX11486;
wire II14624;
wire WX5345;
wire WX6169;
wire WX10299;
wire II30924;
wire WX3302;
wire WX2713;
wire WX2926;
wire WX1579;
wire II34260;
wire II19633;
wire WX394;
wire II27292;
wire II26299;
wire WX913;
wire II18564;
wire WX10177;
wire WX6275;
wire WX4848;
wire II14733;
wire WX11222;
wire WX1029;
wire WX2177;
wire II15664;
wire WX1556;
wire II30946;
wire II15648;
wire II27162;
wire WX4000;
wire WX7946;
wire WX6393;
wire WX7003;
wire WX3747;
wire WX8506;
wire WX4257;
wire II15095;
wire WX926;
wire WX7950;
wire WX6658;
wire WX750;
wire WX4359;
wire WX10683;
wire WX7607;
wire WX10382;
wire II30247;
wire WX2561;
wire II14833;
wire WX9287;
wire WX9622;
wire WX5996;
wire II2307;
wire II18016;
wire WX3430;
wire WX4023;
wire WX9056;
wire WX10422;
wire WX9201;
wire II18216;
wire II30939;
wire WX4827;
wire II6839;
wire WX11050;
wire II14818;
wire WX1909;
wire II27733;
wire WX10227;
wire II10385;
wire WX1646;
wire WX10233;
wire WX4431;
wire II22107;
wire WX10894;
wire WX1454;
wire II26274;
wire WX6160;
wire II26901;
wire II26190;
wire II18692;
wire WX1401;
wire WX3058;
wire WX8184;
wire II22392;
wire II14578;
wire II10580;
wire WX483;
wire WX6361;
wire II7422;
wire II34245;
wire II6661;
wire II2748;
wire II31401;
wire WX5464;
wire II22068;
wire WX2149;
wire WX8361;
wire II6318;
wire WX2750;
wire WX4970;
wire WX802;
wire II26528;
wire WX1437;
wire II18278;
wire WX10779;
wire II22633;
wire II14591;
wire WX1528;
wire WX7897;
wire II10617;
wire II30558;
wire II19653;
wire II23715;
wire WX3332;
wire II7057;
wire WX9853;
wire II26591;
wire WX4280;
wire WX9837;
wire II11553;
wire WX9326;
wire WX3543;
wire WX5813;
wire II23273;
wire WX2799;
wire WX3910;
wire WX9575;
wire II34524;
wire WX1246;
wire II34330;
wire WX8681;
wire II6646;
wire II26358;
wire WX2454;
wire WX5702;
wire WX11630;
wire WX11520;
wire WX3960;
wire WX6959;
wire WX8462;
wire WX7751;
wire WX1160;
wire II18961;
wire II26243;
wire WX1898;
wire II31626;
wire WX3046;
wire WX6343;
wire II31528;
wire WX1338;
wire II6629;
wire WX7679;
wire II18806;
wire WX11152;
wire II6914;
wire II26544;
wire II22671;
wire II22579;
wire WX10858;
wire II10843;
wire WX2021;
wire II30983;
wire WX9634;
wire WX6221;
wire WX3528;
wire WX5904;
wire WX3495;
wire II10031;
wire II18627;
wire II2827;
wire WX4482;
wire WX5028;
wire WX4195;
wire WX9162;
wire WX1065;
wire II3577;
wire WX3350;
wire II26088;
wire II26786;
wire WX123;
wire WX5267;
wire WX10612;
wire WX9637;
wire WX6228;
wire WX1610;
wire II18139;
wire WX5125;
wire WX159;
wire WX6522;
wire II35105;
wire II31490;
wire II30975;
wire II7498;
wire II30572;
wire II30269;
wire II18642;
wire WX6937;
wire WX1461;
wire II6614;
wire WX10036;
wire WX8122;
wire WX9267;
wire II18906;
wire WX11397;
wire II6101;
wire WX6824;
wire WX9964;
wire WX3260;
wire WX5235;
wire II34546;
wire II30613;
wire II14880;
wire WX5613;
wire WX7787;
wire WX9279;
wire WX4434;
wire WX2667;
wire WX7935;
wire II14887;
wire II23235;
wire WX8307;
wire WX5944;
wire WX1099;
wire II19476;
wire II19576;
wire II26683;
wire WX7963;
wire WX4889;
wire II15501;
wire II14917;
wire II22259;
wire WX8560;
wire WX4950;
wire WX4291;
wire WX5781;
wire WX3890;
wire II10465;
wire WX203;
wire WX5155;
wire WX10484;
wire II2485;
wire II30682;
wire WX419;
wire II30689;
wire WX6942;
wire II11336;
wire WX764;
wire II35354;
wire II22905;
wire WX2277;
wire WX652;
wire WX10598;
wire WX2700;
wire II23603;
wire II34717;
wire II10275;
wire WX5090;
wire WX7133;
wire WX3726;
wire II15276;
wire WX8114;
wire II10756;
wire WX1636;
wire WX1039;
wire WX6554;
wire WX5358;
wire II26483;
wire WX1157;
wire II30877;
wire II31633;
wire II10037;
wire WX878;
wire II34648;
wire WX6290;
wire WX8786;
wire WX10020;
wire II22750;
wire WX5315;
wire WX3740;
wire WX6571;
wire II7568;
wire WX10940;
wire II30108;
wire WX2623;
wire II34633;
wire WX3179;
wire II26104;
wire II26971;
wire WX6578;
wire WX11446;
wire II22073;
wire WX7781;
wire WX4305;
wire WX2540;
wire II2606;
wire II11540;
wire II31725;
wire II2741;
wire WX3600;
wire II2663;
wire WX1859;
wire II23638;
wire WX9541;
wire II14499;
wire II11610;
wire WX11620;
wire WX3140;
wire WX3262;
wire II22252;
wire WX2331;
wire II34710;
wire WX7327;
wire WX4927;
wire WX4165;
wire WX2133;
wire II14335;
wire II18689;
wire II6591;
wire WX1767;
wire WX10359;
wire WX6655;
wire WX3643;
wire WX5780;
wire WX1417;
wire II22881;
wire II10424;
wire WX11468;
wire II2677;
wire WX4018;
wire II6797;
wire WX8921;
wire WX3695;
wire II23597;
wire II7535;
wire WX4617;
wire WX2507;
wire II10811;
wire WX7056;
wire WX5207;
wire WX7535;
wire WX247;
wire WX11597;
wire WX10677;
wire WX10984;
wire WX5385;
wire WX2808;
wire II30758;
wire II6336;
wire II2423;
wire II7624;
wire WX4876;
wire WX3152;
wire WX5025;
wire II14390;
wire II22663;
wire WX8984;
wire II11526;
wire II34588;
wire WX11018;
wire WX2980;
wire WX7994;
wire WX6010;
wire WX3771;
wire II19591;
wire WX6858;
wire II34137;
wire WX6032;
wire WX1819;
wire II34864;
wire WX864;
wire WX3587;
wire II15606;
wire II10417;
wire WX7563;
wire WX7518;
wire WX110;
wire II2609;
wire WX1220;
wire II35618;
wire WX2783;
wire WX2490;
wire II35673;
wire II15684;
wire WX7771;
wire II18304;
wire WX11102;
wire WX5277;
wire WX9809;
wire WX5258;
wire WX5928;
wire II22998;
wire WX222;
wire WX3708;
wire II34898;
wire II26125;
wire II11075;
wire II18320;
wire II6115;
wire II10393;
wire WX6634;
wire WX11436;
wire WX3769;
wire II14081;
wire WX5535;
wire II6945;
wire WX8136;
wire WX7101;
wire II15593;
wire WX1186;
wire II7596;
wire II18118;
wire WX333;
wire II6930;
wire WX9781;
wire II3710;
wire WX8386;
wire WX10139;
wire WX8747;
wire II22827;
wire II22253;
wire WX5761;
wire II22834;
wire WX9677;
wire WX10069;
wire WX4126;
wire II22619;
wire II6435;
wire II19562;
wire II27227;
wire WX7229;
wire WX6322;
wire WX6287;
wire WX1856;
wire WX9521;
wire II34130;
wire WX2354;
wire WX9211;
wire II15185;
wire II7176;
wire WX5138;
wire II6193;
wire II2903;
wire II6170;
wire WX78;
wire II22159;
wire II26319;
wire II34694;
wire WX1203;
wire WX3758;
wire WX3828;
wire WX1151;
wire II3092;
wire WX10253;
wire WX7257;
wire II19703;
wire II6131;
wire WX2960;
wire WX2416;
wire II11608;
wire WX1690;
wire WX1043;
wire WX8225;
wire II35145;
wire II2765;
wire II30913;
wire WX8098;
wire WX2977;
wire II31414;
wire II26150;
wire WX7952;
wire II14764;
wire II35198;
wire II19606;
wire WX1241;
wire II30023;
wire WX9204;
wire II18053;
wire WX8109;
wire WX9141;
wire II22996;
wire II14809;
wire WX283;
wire WX448;
wire WX4815;
wire II7135;
wire WX7836;
wire II31100;
wire II18854;
wire WX10939;
wire WX7235;
wire WX2318;
wire II2058;
wire WX8091;
wire WX1517;
wire II18845;
wire WX10819;
wire WX10258;
wire II3499;
wire II26870;
wire WX1983;
wire II23338;
wire WX1250;
wire II35639;
wire II19243;
wire WX3448;
wire WX11322;
wire WX5754;
wire II34321;
wire WX4822;
wire WX3218;
wire II23723;
wire II22594;
wire II14181;
wire II26171;
wire WX8233;
wire II19569;
wire WX5722;
wire II7292;
wire II30202;
wire WX10918;
wire WX9601;
wire WX10647;
wire WX6752;
wire WX1703;
wire II10795;
wire WX2330;
wire WX8758;
wire WX6864;
wire WX1442;
wire WX955;
wire WX2652;
wire WX9528;
wire WX8911;
wire WX5790;
wire WX2498;
wire WX3674;
wire II34965;
wire II30409;
wire WX2011;
wire WX11002;
wire II14281;
wire II15692;
wire II22361;
wire II10689;
wire II22991;
wire WX10834;
wire II27278;
wire WX5990;
wire II6258;
wire II35632;
wire WX11418;
wire II3626;
wire WX2741;
wire II26290;
wire II2910;
wire WX6860;
wire II22780;
wire WX2238;
wire WX6673;
wire WX5469;
wire WX8859;
wire WX10812;
wire II22859;
wire WX8856;
wire II23616;
wire WX2950;
wire WX9314;
wire II3275;
wire WX6771;
wire WX10433;
wire II35722;
wire II2003;
wire WX1667;
wire II15172;
wire WX10920;
wire WX9711;
wire WX8679;
wire II26405;
wire II22913;
wire WX11048;
wire II27607;
wire WX10166;
wire WX6105;
wire WX7036;
wire II26578;
wire II14655;
wire WX8719;
wire II30827;
wire II34734;
wire WX5226;
wire II15516;
wire II6405;
wire II6373;
wire WX7857;
wire WX11265;
wire WX6683;
wire II2856;
wire II10454;
wire II26568;
wire II26699;
wire II22355;
wire WX1390;
wire WX10327;
wire WX2381;
wire WX1492;
wire WX2865;
wire WX9014;
wire WX2893;
wire II31006;
wire WX968;
wire WX8711;
wire II10642;
wire WX11347;
wire WX367;
wire II19604;
wire WX5421;
wire WX7221;
wire II10780;
wire II2198;
wire WX424;
wire WX4177;
wire WX11304;
wire II26639;
wire II11466;
wire WX7799;
wire II2182;
wire II22368;
wire WX10143;
wire WX11495;
wire WX60;
wire WX10207;
wire WX8674;
wire II34601;
wire WX1371;
wire WX7581;
wire II2259;
wire WX2881;
wire WX351;
wire II31598;
wire II6243;
wire II18583;
wire II14904;
wire WX6154;
wire II6596;
wire WX5747;
wire II10518;
wire WX8015;
wire II34207;
wire WX7917;
wire II14322;
wire II18821;
wire II10680;
wire WX7660;
wire WX7547;
wire WX1057;
wire WX911;
wire WX7643;
wire II7477;
wire II7521;
wire WX1737;
wire II30278;
wire WX7504;
wire WX1001;
wire WX2071;
wire WX11072;
wire II31677;
wire II10649;
wire WX7868;
wire WX4118;
wire WX7057;
wire WX4521;
wire II30635;
wire WX9863;
wire II18955;
wire II15262;
wire WX5378;
wire WX11120;
wire II5993;
wire WX7747;
wire II30225;
wire WX11545;
wire WX2441;
wire II2770;
wire II2460;
wire WX4111;
wire WX786;
wire WX7191;
wire WX3712;
wire WX5320;
wire II10911;
wire II18606;
wire WX8584;
wire WX9381;
wire WX1915;
wire WX2346;
wire II18699;
wire WX11066;
wire WX11390;
wire II31230;
wire II14036;
wire WX8725;
wire WX2515;
wire II34936;
wire WX1008;
wire II2129;
wire WX379;
wire WX11372;
wire II2338;
wire II31362;
wire II22687;
wire WX5114;
wire WX9040;
wire WX5540;
wire WX702;
wire WX4101;
wire WX952;
wire WX2397;
wire WX10606;
wire WX8369;
wire II26237;
wire II2469;
wire II27580;
wire II3544;
wire II19462;
wire II6187;
wire WX95;
wire WX4290;
wire II34446;
wire WX9001;
wire WX10663;
wire II7318;
wire WX5806;
wire II34656;
wire WX3846;
wire WX5649;
wire II31535;
wire WX6141;
wire WX3739;
wire WX3961;
wire WX2185;
wire WX7313;
wire WX10396;
wire WX1547;
wire II10044;
wire WX1413;
wire WX1378;
wire II27740;
wire WX3116;
wire WX9539;
wire II14219;
wire II2291;
wire II34712;
wire WX2280;
wire WX7574;
wire WX4141;
wire II2538;
wire II6412;
wire WX7689;
wire II11482;
wire WX9655;
wire II18363;
wire WX8723;
wire WX9656;
wire II35443;
wire WX5801;
wire II3145;
wire II10711;
wire II23555;
wire WX10242;
wire WX6436;
wire WX7477;
wire WX959;
wire WX10487;
wire WX1833;
wire II11609;
wire WX1609;
wire WX48;
wire II27524;
wire WX576;
wire WX2145;
wire II10789;
wire II30449;
wire WX6819;
wire II10091;
wire WX4046;
wire WX1446;
wire WX2324;
wire II6001;
wire WX7411;
wire WX2099;
wire WX2527;
wire WX6138;
wire WX10021;
wire II11479;
wire WX1174;
wire WX6902;
wire WX10180;
wire WX7374;
wire WX9418;
wire WX4884;
wire II3670;
wire WX4091;
wire II2546;
wire WX1675;
wire II18859;
wire II6326;
wire WX10601;
wire WX9148;
wire WX8624;
wire WX9825;
wire WX2489;
wire WX2633;
wire II22104;
wire WX1533;
wire II18471;
wire II10369;
wire WX6179;
wire WX7808;
wire II22604;
wire WX3535;
wire II26361;
wire WX9899;
wire II34340;
wire WX608;
wire WX581;
wire WX252;
wire WX2830;
wire WX5629;
wire II18769;
wire II18480;
wire WX7463;
wire II23286;
wire II34409;
wire WX3498;
wire WX8344;
wire WX9166;
wire WX5708;
wire II14856;
wire II10370;
wire WX5872;
wire II23261;
wire WX10462;
wire II18263;
wire WX10972;
wire WX7853;
wire II30650;
wire II19667;
wire II34169;
wire WX8241;
wire WX4182;
wire WX4567;
wire II6395;
wire WX4072;
wire WX10509;
wire WX496;
wire WX9496;
wire WX10001;
wire WX6087;
wire WX71;
wire WX2571;
wire II34347;
wire WX329;
wire WX1078;
wire WX6589;
wire II14687;
wire WX8311;
wire WX6080;
wire II3493;
wire WX5107;
wire II6038;
wire WX10198;
wire WX3800;
wire II10440;
wire WX5759;
wire II2446;
wire WX7157;
wire WX4939;
wire WX6805;
wire WX6358;
wire WX7026;
wire II3105;
wire II3117;
wire WX7812;
wire WX6284;
wire WX4947;
wire II14446;
wire WX4185;
wire WX3625;
wire WX5612;
wire II34431;
wire WX7083;
wire WX10106;
wire WX1848;
wire II2330;
wire II31336;
wire WX10005;
wire II6846;
wire II19717;
wire WX11315;
wire WX3975;
wire WX373;
wire WX216;
wire II19710;
wire II23403;
wire WX5547;
wire WX8688;
wire WX6000;
wire II22797;
wire WX9662;
wire WX4099;
wire WX10550;
wire II6690;
wire WX2739;
wire II10898;
wire WX10557;
wire II14346;
wire II2863;
wire II6907;
wire WX7982;
wire WX3420;
wire WX3917;
wire WX7283;
wire WX8918;
wire II26445;
wire WX5075;
wire WX6601;
wire II35716;
wire WX5151;
wire WX9947;
wire WX7933;
wire WX10480;
wire II18574;
wire WX3812;
wire WX3894;
wire WX4006;
wire II14670;
wire WX7720;
wire WX8336;
wire WX8698;
wire II10214;
wire WX1774;
wire WX1670;
wire WX3062;
wire WX11454;
wire WX3472;
wire II18180;
wire WX9605;
wire II2167;
wire II11671;
wire II27136;
wire WX1777;
wire WX11548;
wire WX6351;
wire II27644;
wire WX7267;
wire II11706;
wire II26438;
wire WX8341;
wire WX5625;
wire WX8288;
wire II11650;
wire II27593;
wire II26474;
wire WX5353;
wire II22331;
wire II35483;
wire II31087;
wire WX4387;
wire II10170;
wire II19190;
wire WX8350;
wire WX11356;
wire WX5940;
wire II30440;
wire WX11412;
wire II10656;
wire WX7650;
wire WX3575;
wire II14575;
wire WX1073;
wire WX5620;
wire WX1868;
wire II22562;
wire II22222;
wire II11166;
wire WX908;
wire WX1999;
wire WX2685;
wire WX1133;
wire II30486;
wire WX6567;
wire WX7877;
wire WX3552;
wire II22199;
wire WX1719;
wire WX10110;
wire WX3811;
wire WX6272;
wire WX10695;
wire II10565;
wire WX41;
wire II27433;
wire WX1562;
wire WX6755;
wire WX8634;
wire II14700;
wire WX2819;
wire WX3126;
wire II18341;
wire WX3972;
wire WX1850;
wire II35518;
wire WX9669;
wire WX10862;
wire II31607;
wire WX9231;
wire II18202;
wire WX11333;
wire WX10279;
wire WX3051;
wire WX5336;
wire WX4960;
wire WX9644;
wire WX947;
wire II27572;
wire WX5018;
wire WX7532;
wire WX2039;
wire WX8592;
wire II2523;
wire II10558;
wire WX11214;
wire WX4272;
wire WX11293;
wire WX7828;
wire WX7876;
wire WX10449;
wire WX8737;
wire WX1576;
wire WX730;
wire WX8189;
wire II14987;
wire WX1730;
wire WX6618;
wire WX617;
wire WX3314;
wire WX6661;
wire II27539;
wire WX8887;
wire II3479;
wire WX10587;
wire WX8872;
wire WX10421;
wire WX7492;
wire WX6066;
wire WX2882;
wire WX4800;
wire WX5440;
wire WX5954;
wire II34122;
wire II10293;
wire WX974;
wire WX11563;
wire II19152;
wire WX614;
wire WX10804;
wire WX8906;
wire WX2287;
wire WX11176;
wire WX10510;
wire WX10774;
wire II7582;
wire WX3821;
wire II34243;
wire WX8928;
wire II14863;
wire WX11234;
wire WX1341;
wire II10046;
wire WX3181;
wire II23156;
wire WX8825;
wire II14298;
wire WX4066;
wire WX4207;
wire WX11284;
wire WX4200;
wire WX6427;
wire WX9415;
wire WX2644;
wire II34935;
wire WX3222;
wire WX1109;
wire II10929;
wire II10589;
wire WX11218;
wire WX9120;
wire WX2265;
wire WX7514;
wire WX4452;
wire II7548;
wire WX5382;
wire II10199;
wire II2468;
wire WX7173;
wire II2430;
wire WX9440;
wire WX3513;
wire WX11606;
wire WX1569;
wire II22285;
wire WX132;
wire II34154;
wire WX1468;
wire WX4836;
wire WX3082;
wire WX5273;
wire WX3464;
wire WX8147;
wire WX10428;
wire II23363;
wire II31206;
wire WX10760;
wire II34236;
wire II11297;
wire WX4723;
wire WX9643;
wire WX5389;
wire WX10525;
wire WX7539;
wire II34966;
wire II11568;
wire WX2528;
wire WX4969;
wire II31167;
wire II18223;
wire WX9104;
wire WX5726;
wire II15133;
wire II2414;
wire WX4089;
wire II11617;
wire II2096;
wire II14072;
wire II10523;
wire WX2857;
wire II22554;
wire II18526;
wire II14079;
wire WX10750;
wire WX8665;
wire II3455;
wire WX8370;
wire WX9152;
wire WX3736;
wire WX10056;
wire II18170;
wire WX6781;
wire II15379;
wire II34665;
wire WX10591;
wire II27720;
wire WX7452;
wire II26653;
wire II22588;
wire WX5015;
wire II7513;
wire WX1722;
wire II2700;
wire WX1092;
wire WX10520;
wire WX8424;
wire WX9455;
wire WX1036;
wire WX4039;
wire WX2654;
wire II34112;
wire WX11206;
wire WX9727;
wire WX6249;
wire II7111;
wire II2870;
wire II3537;
wire WX3836;
wire II10501;
wire II6218;
wire II18682;
wire WX7526;
wire WX9068;
wire WX4864;
wire II30776;
wire II10868;
wire II10626;
wire WX7460;
wire WX2195;
wire II31452;
wire II11271;
wire WX436;
wire WX9306;
wire WX5436;
wire II34943;
wire WX6122;
wire WX6693;
wire WX5375;
wire WX6263;
wire WX11634;
wire WX5503;
wire WX2757;
wire WX4032;
wire II10804;
wire II2926;
wire II19215;
wire WX10929;
wire II22532;
wire II7462;
wire WX5597;
wire WX11438;
wire WX9138;
wire II30992;
wire WX1489;
wire WX4497;
wire II26345;
wire WX3818;
wire WX7351;
wire WX7117;
wire II18218;
wire WX1873;
wire WX4263;
wire WX2019;
wire II18775;
wire II3067;
wire II2028;
wire II10826;
wire WX6208;
wire WX10301;
wire WX10781;
wire WX3666;
wire WX4146;
wire WX5078;
wire WX7014;
wire WX4637;
wire II27317;
wire II7715;
wire II7617;
wire II34216;
wire WX3027;
wire II30102;
wire II10192;
wire WX3966;
wire WX1761;
wire WX5056;
wire II27719;
wire WX5516;
wire II22383;
wire WX2761;
wire WX11603;
wire WX6474;
wire WX5293;
wire WX1874;
wire II11623;
wire WX10913;
wire WX9587;
wire II35534;
wire II14585;
wire II34370;
wire WX10308;
wire II26025;
wire WX297;
wire II18084;
wire WX380;
wire II22231;
wire WX1257;
wire WX5639;
wire WX6511;
wire II23686;
wire II22120;
wire II14213;
wire WX4232;
wire WX3568;
wire WX3141;
wire WX3352;
wire WX10547;
wire II7666;
wire WX5238;
wire WX3780;
wire WX1823;
wire WX10701;
wire II2708;
wire II2833;
wire WX2995;
wire WX9955;
wire WX3743;
wire II14638;
wire WX10817;
wire II22492;
wire WX2404;
wire WX4989;
wire WX7893;
wire II26630;
wire II10402;
wire WX462;
wire II2734;
wire II27705;
wire WX2085;
wire II34879;
wire WX4659;
wire WX6207;
wire WX5323;
wire WX7848;
wire WX8175;
wire WX5484;
wire WX1298;
wire II2105;
wire II7148;
wire WX1959;
wire WX7337;
wire II22098;
wire II22175;
wire II14955;
wire WX8155;
wire WX8104;
wire WX623;
wire WX7509;
wire WX10187;
wire WX3196;
wire WX1664;
wire WX6706;
wire WX2201;
wire II2235;
wire II23247;
wire WX11384;
wire WX9422;
wire WX6546;
wire WX8849;
wire II26466;
wire WX8039;
wire II10477;
wire II18785;
wire WX8840;
wire WX11188;
wire II7499;
wire WX5369;
wire WX8208;
wire WX4464;
wire II6280;
wire WX2113;
wire II22432;
wire WX5214;
wire WX2948;
wire WX2835;
wire WX8035;
wire WX7042;
wire WX7435;
wire II22462;
wire II2361;
wire II26249;
wire WX4904;
wire WX4287;
wire II18134;
wire WX2240;
wire WX6534;
wire II11400;
wire WX10625;
wire II31578;
wire II27499;
wire WX7674;
wire II6622;
wire II6093;
wire WX6535;
wire II15431;
wire WX772;
wire II19725;
wire WX303;
wire II26590;
wire II3352;
wire WX8734;
wire WX10113;
wire WX8685;
wire II30605;
wire WX6768;
wire WX4428;
wire II22890;
wire II31504;
wire WX5061;
wire WX5000;
wire WX10876;
wire WX3016;
wire II10409;
wire II31322;
wire II2947;
wire WX6502;
wire II2312;
wire II11322;
wire WX7499;
wire WX4477;
wire WX7074;
wire II26522;
wire II10089;
wire II18875;
wire WX4139;
wire WX4057;
wire II19549;
wire WX2845;
wire WX1586;
wire WX58;
wire WX7928;
wire WX2427;
wire II19583;
wire II7702;
wire WX11640;
wire WX2433;
wire WX11510;
wire II30843;
wire WX7706;
wire WX8704;
wire WX11508;
wire WX2828;
wire WX4737;
wire WX3688;
wire WX8792;
wire WX5581;
wire II34339;
wire WX144;
wire WX3924;
wire II35738;
wire WX9296;
wire II2925;
wire II31613;
wire WX1654;
wire WX4178;
wire WX9517;
wire WX10247;
wire WX3943;
wire WX1467;
wire II18723;
wire WX8695;
wire WX10214;
wire II10403;
wire WX2661;
wire II18837;
wire II27213;
wire II30852;
wire II22820;
wire II18356;
wire II11114;
wire WX1973;
wire WX6188;
wire II2083;
wire WX4509;
wire WX4959;
wire WX6109;
wire WX358;
wire WX4169;
wire WX2508;
wire II14166;
wire WX8764;
wire II23311;
wire WX6390;
wire WX9407;
wire WX5414;
wire II34190;
wire WX9479;
wire WX5403;
wire II26745;
wire WX126;
wire WX1193;
wire WX11458;
wire WX4502;
wire WX2772;
wire II30665;
wire II18518;
wire WX9508;
wire WX1699;
wire II30567;
wire WX2779;
wire WX56;
wire II19372;
wire II6720;
wire WX7365;
wire WX8126;
wire WX9197;
wire II30722;
wire II15538;
wire WX8480;
wire WX10652;
wire II23351;
wire WX343;
wire II26624;
wire WX9366;
wire WX4940;
wire WX9091;
wire WX10212;
wire II34050;
wire II6637;
wire II34851;
wire II23350;
wire WX5445;
wire WX2477;
wire WX832;
wire II31001;
wire WX310;
wire WX5165;
wire WX9246;
wire II27394;
wire WX11666;
wire WX2474;
wire WX7446;
wire II34307;
wire WX5491;
wire WX9350;
wire WX2676;
wire WX5255;
wire WX2969;
wire II30889;
wire II34887;
wire WX3639;
wire II15698;
wire WX9616;
wire WX9439;
wire WX992;
wire II30131;
wire II30955;
wire II6830;
wire WX5129;
wire WX1236;
wire WX8836;
wire II3508;
wire WX3630;
wire WX8172;
wire WX2379;
wire II26280;
wire WX6133;
wire WX233;
wire WX892;
wire WX10269;
wire II30551;
wire WX7427;
wire WX4707;
wire II26707;
wire WX8953;
wire II7490;
wire WX8998;
wire WX6873;
wire WX5886;
wire II27501;
wire WX1434;
wire WX3390;
wire WX3504;
wire WX180;
wire WX11096;
wire WX5482;
wire II7150;
wire WX7739;
wire WX7599;
wire WX3699;
wire WX2249;
wire II6776;
wire WX1219;
wire II35598;
wire II3366;
wire WX5428;
wire II30579;
wire II3404;
wire WX10456;
wire WX3827;
wire WX11515;
wire II22455;
wire II6364;
wire II22166;
wire II2679;
wire II34960;
wire II30404;
wire WX6916;
wire WX5260;
wire WX10085;
wire II7590;
wire II18441;
wire WX5307;
wire WX8946;
wire WX2388;
wire WX4949;
wire WX11656;
wire II34719;
wire II19178;
wire WX9625;
wire WX6842;
wire WX3902;
wire WX5568;
wire WX8875;
wire WX884;
wire WX9996;
wire WX8388;
wire WX7400;
wire II6953;
wire WX6118;
wire WX3518;
wire WX11420;
wire WX1729;
wire WX7243;
wire II6761;
wire WX4805;
wire WX2173;
wire II19359;
wire WX2870;
wire WX320;
wire WX1743;
wire WX276;
wire WX10132;
wire WX8029;
wire WX1276;
wire II2630;
wire WX9209;
wire II10672;
wire WX9707;
wire WX8716;
wire II23169;
wire II31308;
wire WX1892;
wire WX5413;
wire II34894;
wire WX10846;
wire WX10914;
wire WX5261;
wire II27459;
wire II2027;
wire WX4206;
wire WX4825;
wire WX9434;
wire WX7225;
wire WX5388;
wire WX10477;
wire WX11178;
wire WX3697;
wire WX9763;
wire II35352;
wire II10849;
wire WX1209;
wire WX1396;
wire WX5130;
wire WX1757;
wire II31310;
wire II30154;
wire WX3183;
wire WX5274;
wire II27396;
wire WX10621;
wire WX1934;
wire WX245;
wire WX10827;
wire II10665;
wire WX2446;
wire II6179;
wire WX1930;
wire WX8092;
wire II14559;
wire WX7604;
wire WX8127;
wire II10224;
wire II34502;
wire II14941;
wire WX4814;
wire II30208;
wire II6937;
wire II34222;
wire WX3786;
wire WX4498;
wire WX3765;
wire WX10946;
wire II34858;
wire II22879;
wire II22014;
wire WX8192;
wire WX5686;
wire WX1207;
wire II7344;
wire II10603;
wire WX11410;
wire WX3802;
wire WX6170;
wire WX1189;
wire II14786;
wire WX10609;
wire WX9219;
wire WX82;
wire WX4956;
wire II18196;
wire WX6550;
wire WX1621;
wire WX4123;
wire II15106;
wire WX7583;
wire II34509;
wire WX1827;
wire WX6448;
wire II22352;
wire II10740;
wire WX6222;
wire II14862;
wire II2885;
wire II22929;
wire WX2679;
wire WX10066;
wire II22617;
wire WX375;
wire WX10775;
wire WX6100;
wire WX4011;
wire WX8430;
wire II35653;
wire II19563;
wire WX5534;
wire WX7104;
wire WX5456;
wire WX2314;
wire WX1969;
wire WX8530;
wire WX235;
wire WX10254;
wire WX9785;
wire II3093;
wire II18342;
wire WX130;
wire WX11270;
wire WX360;
wire WX281;
wire WX2553;
wire II23246;
wire II30541;
wire WX4439;
wire II22037;
wire II18719;
wire II10100;
wire II7688;
wire II10967;
wire WX1226;
wire WX6383;
wire II26314;
wire II14291;
wire WX8528;
wire II10547;
wire WX2467;
wire WX8916;
wire WX8955;
wire II15236;
wire II11715;
wire II31605;
wire II30657;
wire II22681;
wire II15250;
wire WX1745;
wire WX6867;
wire II19676;
wire WX6566;
wire WX6888;
wire WX4054;
wire II18458;
wire WX754;
wire II10007;
wire WX11350;
wire WX7311;
wire WX306;
wire WX8854;
wire WX1628;
wire WX3649;
wire WX2651;
wire II14437;
wire WX8743;
wire II34464;
wire II22973;
wire II26729;
wire WX2781;
wire II30534;
wire WX11479;
wire II30851;
wire WX10412;
wire WX11425;
wire WX9463;
wire WX3138;
wire II6119;
wire II18007;
wire WX9192;
wire WX5249;
wire II27199;
wire II18712;
wire II31683;
wire II14005;
wire II14438;
wire WX286;
wire II11673;
wire WX2898;
wire II27264;
wire WX9715;
wire II27342;
wire II11257;
wire WX11106;
wire WX1272;
wire WX7203;
wire II2529;
wire II34316;
wire WX4518;
wire WX10538;
wire II30675;
wire II18753;
wire II34083;
wire II26351;
wire II14167;
wire II31584;
wire II31718;
wire WX2434;
wire II26096;
wire WX4679;
wire II7331;
wire WX11521;
wire WX11407;
wire WX8812;
wire WX5250;
wire WX6377;
wire WX9228;
wire II6265;
wire II23377;
wire II14383;
wire WX1515;
wire WX1182;
wire WX10218;
wire WX3006;
wire II14873;
wire WX1041;
wire II18048;
wire WX50;
wire WX4485;
wire II34362;
wire WX4459;
wire II2382;
wire WX10711;
wire WX10659;
wire WX9345;
wire II26413;
wire WX1895;
wire WX57;
wire WX8671;
wire WX9474;
wire WX4210;
wire II35589;
wire II34290;
wire WX2533;
wire WX8326;
wire II27500;
wire WX858;
wire WX9010;
wire WX10564;
wire II2113;
wire II34159;
wire WX2954;
wire WX9044;
wire WX3462;
wire II15225;
wire WX8394;
wire II35418;
wire WX2157;
wire WX10493;
wire II35640;
wire WX962;
wire II2699;
wire WX2500;
wire II14964;
wire WX6537;
wire WX7376;
wire WX3043;
wire WX3935;
wire II2072;
wire WX6559;
wire WX2429;
wire II34299;
wire WX192;
wire II26778;
wire WX6438;
wire WX10724;
wire WX7459;
wire WX5746;
wire II18077;
wire WX5864;
wire WX1296;
wire WX2270;
wire II31648;
wire WX200;
wire WX4753;
wire WX7107;
wire II15608;
wire WX3521;
wire WX10439;
wire WX2282;
wire WX2970;
wire II11502;
wire II31191;
wire II3249;
wire II34593;
wire WX2279;
wire WX3640;
wire WX459;
wire II35638;
wire II6868;
wire WX6947;
wire WX1614;
wire WX8052;
wire WX2083;
wire II30193;
wire II10285;
wire II26327;
wire II14143;
wire II30232;
wire WX7845;
wire II18426;
wire II26981;
wire WX1444;
wire WX9371;
wire II30309;
wire WX9631;
wire II26840;
wire II31243;
wire II15433;
wire WX9236;
wire WX7478;
wire WX1482;
wire II3312;
wire WX259;
wire II14305;
wire WX1594;
wire WX6678;
wire II6062;
wire WX4531;
wire WX4085;
wire WX250;
wire WX2272;
wire WX10807;
wire WX3162;
wire WX6407;
wire WX10705;
wire II7215;
wire WX8400;
wire II18992;
wire WX4203;
wire WX11301;
wire II6753;
wire II19425;
wire WX4844;
wire WX2235;
wire II15446;
wire II7408;
wire WX7914;
wire II23443;
wire II3662;
wire WX1532;
wire WX1587;
wire II34895;
wire WX4285;
wire II30300;
wire II10906;
wire II2786;
wire WX4721;
wire II23509;
wire II34562;
wire WX5326;
wire WX6121;
wire II22666;
wire WX2461;
wire WX7046;
wire WX1326;
wire WX7654;
wire II26808;
wire WX3148;
wire WX9632;
wire II14043;
wire WX3860;
wire II2470;
wire II19334;
wire WX7615;
wire WX6266;
wire WX8095;
wire WX100;
wire II6201;
wire WX470;
wire II18598;
wire WX11464;
wire WX4191;
wire WX9164;
wire WX8945;
wire II27134;
wire WX10234;
wire WX7609;
wire WX6282;
wire WX4344;
wire II18404;
wire II11720;
wire WX10032;
wire WX10167;
wire WX5570;
wire WX2363;
wire II27329;
wire II27544;
wire WX10365;
wire II15636;
wire WX1477;
wire WX2747;
wire II6683;
wire WX9893;
wire WX988;
wire WX4362;
wire II2601;
wire WX2856;
wire WX642;
wire II34422;
wire WX9022;
wire WX7967;
wire II27545;
wire WX7431;
wire WX5211;
wire WX4921;
wire II2314;
wire WX260;
wire WX9987;
wire WX8067;
wire WX10054;
wire II34709;
wire WX6648;
wire II35406;
wire WX11020;
wire WX6933;
wire II2662;
wire WX7866;
wire WX3292;
wire WX1500;
wire WX7562;
wire WX969;
wire WX2105;
wire WX1130;
wire WX9980;
wire WX6110;
wire II27686;
wire WX4871;
wire WX1312;
wire WX4711;
wire WX7695;
wire WX6963;
wire WX6574;
wire WX387;
wire II18736;
wire WX6014;
wire WX3618;
wire WX10090;
wire II30712;
wire WX1705;
wire WX5053;
wire WX7397;
wire II34052;
wire WX9689;
wire II30388;
wire II2871;
wire WX1763;
wire II18070;
wire WX10405;
wire II18596;
wire WX9305;
wire II23679;
wire II30356;
wire WX8228;
wire II10981;
wire II6885;
wire II2358;
wire WX7716;
wire II2608;
wire WX11084;
wire II26166;
wire WX9488;
wire WX9454;
wire WX443;
wire WX6953;
wire II34958;
wire WX5088;
wire WX1331;
wire II18412;
wire WX11228;
wire II30068;
wire II2761;
wire WX8240;
wire WX2362;
wire WX11224;
wire II18552;
wire WX3824;
wire II30226;
wire II11664;
wire WX1801;
wire WX2412;
wire II22076;
wire II30378;
wire WX9690;
wire WX3122;
wire WX2686;
wire WX9392;
wire WX11610;
wire WX1947;
wire WX125;
wire II1987;
wire WX5189;
wire WX639;
wire WX11550;
wire WX10761;
wire II23454;
wire WX5472;
wire II34500;
wire WX3745;
wire II2584;
wire WX11343;
wire II22851;
wire WX6652;
wire II34819;
wire WX7630;
wire WX612;
wire WX3874;
wire II14429;
wire II26120;
wire II14408;
wire II10028;
wire II22526;
wire II22315;
wire II30218;
wire II26669;
wire WX830;
wire WX7171;
wire II30030;
wire WX979;
wire WX1456;
wire WX1369;
wire WX8987;
wire WX3990;
wire II10720;
wire II22084;
wire II6542;
wire II10022;
wire II18115;
wire II2320;
wire WX8976;
wire WX4839;
wire WX8302;
wire WX8804;
wire II7605;
wire WX2350;
wire II30806;
wire WX3658;
wire WX6708;
wire II31599;
wire WX3135;
wire WX575;
wire II35120;
wire II26660;
wire II15522;
wire II23092;
wire WX6729;
wire WX3570;
wire WX2905;
wire WX11398;
wire WX2790;
wire II34121;
wire WX8063;
wire II19256;
wire II2686;
wire WX8883;
wire II2477;
wire WX6413;
wire WX4792;
wire WX2902;
wire II34826;
wire II10912;
wire II30751;
wire WX8234;
wire WX6721;
wire II18650;
wire II7317;
wire II2710;
wire II14616;
wire WX1058;
wire II34804;
wire WX3438;
wire II19683;
wire WX3564;
wire WX2419;
wire WX1333;
wire WX6181;
wire WX726;
wire WX4992;
wire II30286;
wire WX8363;
wire WX9747;
wire WX5288;
wire II18798;
wire WX10822;
wire II23735;
wire II14739;
wire WX7888;
wire WX8767;
wire II3585;
wire II26753;
wire II10586;
wire WX8898;
wire WX3932;
wire II34507;
wire II22742;
wire II23155;
wire WX10130;
wire WX1384;
wire WX4975;
wire WX7829;
wire WX8568;
wire WX2458;
wire II18420;
wire WX10419;
wire WX5775;
wire II19599;
wire II11179;
wire WX10786;
wire WX8482;
wire II6642;
wire WX8964;
wire II30348;
wire WX5461;
wire WX8105;
wire WX9052;
wire WX5067;
wire WX2704;
wire WX2315;
wire WX3424;
wire WX912;
wire II2393;
wire WX10714;
wire WX2357;
wire WX7626;
wire II10074;
wire WX1524;
wire WX11524;
wire II26536;
wire II10146;
wire II22795;
wire WX6247;
wire WX405;
wire WX568;
wire II23415;
wire WX684;
wire WX10589;
wire II15173;
wire WX2556;
wire WX4022;
wire II10895;
wire WX951;
wire WX6312;
wire WX10980;
wire WX10201;
wire II10348;
wire WX9833;
wire WX10643;
wire WX7659;
wire WX10514;
wire WX8939;
wire II18916;
wire II35703;
wire II31204;
wire II6908;
wire II35517;
wire WX10010;
wire II14459;
wire WX1405;
wire WX1839;
wire WX3008;
wire II6296;
wire WX909;
wire WX3832;
wire II2019;
wire WX2613;
wire II6870;
wire WX3226;
wire WX6119;
wire II26917;
wire WX6740;
wire WX2646;
wire WX1630;
wire WX1294;
wire II3478;
wire WX11391;
wire WX6046;
wire II30238;
wire WX5349;
wire II3118;
wire II10850;
wire II30341;
wire WX8930;
wire WX3304;
wire WX2015;
wire WX5143;
wire WX3689;
wire II18534;
wire II30466;
wire WX8180;
wire WX6225;
wire WX5621;
wire WX2025;
wire II2306;
wire WX401;
wire WX3650;
wire II22385;
wire WX2754;
wire II30037;
wire II14825;
wire WX11192;
wire WX6598;
wire WX4065;
wire II34105;
wire II30146;
wire WX10898;
wire II2817;
wire WX5736;
wire WX4747;
wire II3572;
wire II34687;
wire II10556;
wire WX590;
wire WX10610;
wire II34795;
wire II3690;
wire WX3553;
wire II3405;
wire II34237;
wire WX6098;
wire WX7069;
wire WX6591;
wire WX4797;
wire WX558;
wire WX7444;
wire WX5085;
wire WX1353;
wire WX3547;
wire WX7590;
wire WX2716;
wire WX8794;
wire WX3001;
wire WX8755;
wire II26908;
wire II30642;
wire II11588;
wire WX1360;
wire II2672;
wire WX5603;
wire II27407;
wire WX1104;
wire II18419;
wire WX9694;
wire WX2656;
wire II26955;
wire II18791;
wire II2794;
wire WX5523;
wire WX920;
wire WX93;
wire WX2795;
wire II19386;
wire II2623;
wire WX9602;
wire WX826;
wire II34572;
wire II10882;
wire WX4154;
wire II23582;
wire II2544;
wire WX10176;
wire WX6165;
wire II14289;
wire WX8524;
wire II3469;
wire II26853;
wire WX596;
wire WX46;
wire WX9114;
wire II14173;
wire II18954;
wire WX73;
wire WX7949;
wire II10461;
wire WX6924;
wire WX7199;
wire II14352;
wire II23222;
wire WX10094;
wire II14492;
wire WX4591;
wire WX3376;
wire II23469;
wire II15550;
wire WX7838;
wire WX876;
wire II18410;
wire WX3296;
wire II23533;
wire WX4789;
wire WX7979;
wire WX3065;
wire WX1171;
wire WX2392;
wire II35119;
wire WX4893;
wire WX9323;
wire WX6699;
wire WX9855;
wire II10726;
wire II14475;
wire WX8974;
wire WX6885;
wire WX1123;
wire WX10696;
wire II30317;
wire WX5110;
wire WX5810;
wire II19411;
wire WX6079;
wire WX5122;
wire II10775;
wire WX8057;
wire II23609;
wire WX6825;
wire WX546;
wire WX1389;
wire WX5758;
wire WX6850;
wire WX391;
wire WX10129;
wire II34398;
wire WX2247;
wire WX6927;
wire II23511;
wire II11296;
wire WX1176;
wire WX165;
wire II18482;
wire II2141;
wire WX4918;
wire WX10454;
wire WX4865;
wire WX3661;
wire WX10998;
wire II30734;
wire II35211;
wire WX9535;
wire WX4215;
wire WX9505;
wire II26716;
wire WX4003;
wire WX4323;
wire II15499;
wire WX2908;
wire WX10472;
wire WX2836;
wire II26691;
wire II27600;
wire II14715;
wire WX9416;
wire WX6370;
wire II11594;
wire WX7729;
wire WX1662;
wire WX150;
wire WX4557;
wire II34951;
wire II34770;
wire WX3627;
wire II22290;
wire WX5890;
wire WX1916;
wire WX11517;
wire WX10049;
wire II2282;
wire WX7895;
wire WX11591;
wire WX10027;
wire WX10293;
wire WX10926;
wire II7696;
wire WX10108;
wire II18443;
wire WX9523;
wire II19668;
wire II6327;
wire WX7941;
wire WX6835;
wire II3054;
wire WX7970;
wire II7576;
wire II19555;
wire II19550;
wire WX10385;
wire WX6137;
wire II14314;
wire WX3246;
wire WX620;
wire WX9139;
wire WX3167;
wire WX10573;
wire WX10331;
wire II6442;
wire WX7576;
wire WX11283;
wire II6487;
wire WX6212;
wire WX6237;
wire WX3665;
wire WX398;
wire WX10836;
wire WX6500;
wire II23285;
wire WX10798;
wire II14568;
wire WX10732;
wire WX11366;
wire WX9589;
wire II26561;
wire II10802;
wire II3635;
wire WX7646;
wire WX6325;
wire WX1781;
wire WX1924;
wire WX7956;
wire II7619;
wire WX10977;
wire WX7386;
wire II26732;
wire WX3596;
wire II18730;
wire II31551;
wire WX8068;
wire WX2169;
wire WX7016;
wire II26516;
wire WX6659;
wire WX3647;
wire WX11361;
wire WX3778;
wire II7555;
wire WX8371;
wire WX1014;
wire II27421;
wire II6963;
wire WX6387;
wire WX1591;
wire II6645;
wire WX3680;
wire II26359;
wire WX2510;
wire WX768;
wire II26236;
wire WX4171;
wire WX1377;
wire WX10145;
wire II35093;
wire II3299;
wire II19125;
wire II22593;
wire WX8980;
wire II14244;
wire II14196;
wire II14058;
wire WX6800;
wire WX8087;
wire II26203;
wire II2585;
wire WX990;
wire WX1490;
wire II18635;
wire WX6349;
wire WX1554;
wire WX6553;
wire WX2721;
wire II31309;
wire WX7009;
wire II18372;
wire WX3456;
wire WX5021;
wire WX4911;
wire II30890;
wire WX11593;
wire WX8008;
wire WX3997;
wire WX1023;
wire WX10905;
wire WX9961;
wire WX3170;
wire WX6152;
wire WX4254;
wire WX7981;
wire II18697;
wire WX3796;
wire WX3026;
wire WX4318;
wire WX7577;
wire II34385;
wire WX7959;
wire II22402;
wire II31732;
wire II18659;
wire II10316;
wire WX9008;
wire II19073;
wire WX6016;
wire II35682;
wire WX2213;
wire II23730;
wire WX2545;
wire WX5874;
wire WX4522;
wire WX2635;
wire WX7361;
wire II30969;
wire WX11327;
wire II34758;
wire WX3354;
wire II31295;
wire II31439;
wire WX211;
wire II14725;
wire WX2309;
wire II26040;
wire II22694;
wire WX10745;
wire WX7661;
wire II6707;
wire WX3192;
wire II27616;
wire II26268;
wire II35625;
wire WX7412;
wire II34584;
wire WX11000;
wire II22966;
wire WX4383;
wire II30310;
wire II2484;
wire II6481;
wire II26273;
wire II26305;
wire II14398;
wire WX10966;
wire II18614;
wire WX2666;
wire II23581;
wire II2369;
wire WX1649;
wire WX11460;
wire WX423;
wire WX6682;
wire WX2874;
wire WX6845;
wire II18978;
wire WX4653;
wire WX1907;
wire II30464;
wire WX227;
wire II30799;
wire II30071;
wire WX10050;
wire II15380;
wire WX316;
wire II31684;
wire WX1486;
wire II26910;
wire WX77;
wire WX1217;
wire II34663;
wire WX9974;
wire II34639;
wire WX5585;
wire II23524;
wire II10162;
wire II22704;
wire WX6316;
wire WX7019;
wire WX4902;
wire WX7712;
wire II10496;
wire II34283;
wire WX3635;
wire WX1195;
wire WX822;
wire WX9951;
wire II35391;
wire WX4504;
wire WX5241;
wire II22688;
wire WX2377;
wire II26397;
wire WX2813;
wire WX1651;
wire WX9293;
wire II34526;
wire II23659;
wire WX8814;
wire WX4153;
wire II2112;
wire II27609;
wire WX4573;
wire II10749;
wire WX3197;
wire WX10500;
wire II10075;
wire WX4391;
wire WX4765;
wire WX11513;
wire II18351;
wire II2383;
wire II19522;
wire WX4194;
wire WX9404;
wire WX9499;
wire WX3785;
wire II6891;
wire WX2974;
wire WX886;
wire WX9999;
wire WX10919;
wire II35159;
wire WX9312;
wire WX11646;
wire WX11298;
wire WX624;
wire II10805;
wire WX3282;
wire II14832;
wire WX4473;
wire WX6215;
wire II30750;
wire WX10443;
wire WX10310;
wire II26390;
wire II34268;
wire II22284;
wire WX11652;
wire WX9354;
wire WX10162;
wire WX8113;
wire WX6218;
wire WX6881;
wire WX10314;
wire WX8884;
wire WX2423;
wire II34619;
wire II7227;
wire WX7733;
wire WX1243;
wire WX1385;
wire WX9362;
wire II10431;
wire II34254;
wire WX67;
wire WX3728;
wire II18333;
wire WX7849;
wire II10107;
wire II10926;
wire WX5423;
wire II22741;
wire II22207;
wire II35736;
wire WX5395;
wire WX4411;
wire WX2609;
wire II14063;
wire WX7050;
wire II18497;
wire WX5228;
wire WX10930;
wire WX271;
wire WX1728;
wire WX2981;
wire II18123;
wire WX7043;
wire WX9217;
wire WX347;
wire WX7919;
wire WX6849;
wire WX9991;
wire WX11443;
wire II14823;
wire II7631;
wire WX5291;
wire II26250;
wire WX278;
wire II2522;
wire WX11430;
wire WX1149;
wire II2431;
wire WX2478;
wire WX2744;
wire WX7263;
wire WX9241;
wire WX9813;
wire WX4348;
wire WX3358;
wire WX4427;
wire II10153;
wire WX10265;
wire II27460;
wire II2920;
wire II22580;
wire WX6194;
wire II11415;
wire WX7701;
wire WX2534;
wire WX1158;
wire II3106;
wire II15564;
wire WX185;
wire WX1817;
wire WX10546;
wire II3557;
wire II3378;
wire II26482;
wire II6273;
wire WX4333;
wire WX8143;
wire II30086;
wire II15523;
wire WX5424;
wire WX8160;
wire WX9793;
wire WX10379;
wire WX7149;
wire II30176;
wire WX9179;
wire WX4080;
wire II31128;
wire WX89;
wire WX385;
wire II34655;
wire II10651;
wire II7681;
wire II18983;
wire II3260;
wire WX7610;
wire WX6466;
wire WX2487;
wire WX2221;
wire II6728;
wire WX10133;
wire WX11138;
wire WX2261;
wire II2646;
wire WX5556;
wire WX345;
wire II18924;
wire WX5448;
wire WX4166;
wire WX9461;
wire II10372;
wire II3705;
wire WX1253;
wire II26506;
wire WX4405;
wire WX1572;
wire II34772;
wire WX6394;
wire II30882;
wire WX4277;
wire WX262;
wire WX6999;
wire WX3849;
wire WX3953;
wire WX2400;
wire II10610;
wire II10332;
wire WX7929;
wire WX1693;
wire WX5632;
wire II30595;
wire II14795;
wire II19438;
wire II26970;
wire WX7307;
wire WX3022;
wire WX6764;
wire WX10753;
wire WX6530;
wire II23548;
wire WX199;
wire WX5511;
wire WX10059;
wire II34391;
wire WX3605;
wire II18379;
wire II30790;
wire II11194;
wire II6140;
wire WX6782;
wire WX8428;
wire WX7357;
wire WX6108;
wire WX3731;
wire WX1190;
wire II34548;
wire WX355;
wire WX4314;
wire WX3840;
wire WX1234;
wire WX8588;
wire WX2045;
wire WX5101;
wire II7252;
wire II11601;
wire II18489;
wire WX1870;
wire WX8991;
wire WX2802;
wire WX4943;
wire WX1452;
wire II23467;
wire WX6523;
wire II10875;
wire II14707;
wire WX3586;
wire WX11254;
wire II34602;
wire WX9257;
wire WX4176;
wire WX1095;
wire II34873;
wire II30517;
wire WX8960;
wire WX7996;
wire WX2407;
wire II2575;
wire II30719;
wire WX5721;
wire WX9885;
wire WX1928;
wire WX9333;
wire II27664;
wire WX4478;
wire WX8213;
wire II2176;
wire II26461;
wire II22942;
wire II19597;
wire II10771;
wire WX8833;
wire WX5844;
wire WX6582;
wire II19397;
wire II22051;
wire WX806;
wire WX782;
wire WX1764;
wire WX5006;
wire WX10650;
wire II23631;
wire WX2846;
wire II27621;
wire WX7690;
wire WX6828;
wire WX7903;
wire WX5964;
wire WX7070;
wire II2901;
wire II18257;
wire II10679;
wire WX862;
wire WX10789;
wire WX4878;
wire WX6623;
wire II14033;
wire WX8839;
wire WX6541;
wire II2048;
wire WX4058;
wire II14646;
wire II22726;
wire II19360;
wire WX9968;
wire WX117;
wire II23702;
wire II26049;
wire II6436;
wire WX4607;
wire II2359;
wire WX484;
wire WX4513;
wire WX5092;
wire WX8845;
wire II22471;
wire WX4743;
wire II10230;
wire WX10434;
wire II34812;
wire II14848;
wire WX6289;
wire II34417;
wire II14552;
wire WX10571;
wire II2579;
wire WX9431;
wire II27635;
wire WX585;
wire II22091;
wire II11645;
wire WX4777;
wire WX6815;
wire WX6737;
wire WX8075;
wire WX5334;
wire WX5501;
wire II2269;
wire II34119;
wire II22454;
wire WX1887;
wire II15614;
wire WX8199;
wire WX7863;
wire WX1340;
wire WX2117;
wire WX6128;
wire II22214;
wire II22595;
wire II19086;
wire WX1955;
wire WX11474;
wire WX1425;
wire WX7301;
wire II35458;
wire II14329;
wire II30458;
wire II34929;
wire II30986;
wire WX4133;
wire WX1032;
wire II22988;
wire II10813;
wire WX1161;
wire WX710;
wire WX9427;
wire II3457;
wire II22502;
wire II14515;
wire WX6716;
wire WX1443;
wire WX4858;
wire II30273;
wire WX9356;
wire WX8203;
wire WX748;
wire WX8030;
wire II26196;
wire WX8120;
wire WX3015;
wire WX7851;
wire WX4148;
wire WX11245;
wire II30471;
wire WX10505;
wire WX10700;
wire II6653;
wire WX4483;
wire II23694;
wire WX2944;
wire WX6292;
wire WX2933;
wire WX2139;
wire WX9136;
wire II6149;
wire II34181;
wire WX10602;
wire II11452;
wire WX2253;
wire WX11388;
wire II34058;
wire II26283;
wire II18626;
wire WX3031;
wire II34306;
wire WX1066;
wire WX5303;
wire WX5636;
wire WX549;
wire II2894;
wire WX9238;
wire II22934;
wire II30169;
wire WX8072;
wire II6429;
wire II26771;
wire II31113;
wire WX1270;
wire II35631;
wire WX7678;
wire WX10569;
wire II18878;
wire II14111;
wire WX10543;
wire WX7467;
wire II10245;
wire WX9426;
wire WX6204;
wire WX10196;
wire II34027;
wire WX8150;
wire WX6114;
wire WX4135;
wire II18884;
wire WX7908;
wire WX9142;
wire II14849;
wire WX9680;
wire WX5771;
wire II7266;
wire WX11541;
wire II11636;
wire WX2824;
wire II2956;
wire WX7490;
wire WX2917;
wire WX4373;
wire II1995;
wire WX3476;
wire WX9666;
wire II6675;
wire II7447;
wire II10539;
wire WX6894;
wire II22849;
wire WX4351;
wire WX10814;
wire II18557;
wire WX7824;
wire WX2289;
wire WX8352;
wire WX3328;
wire WX10931;
wire II2005;
wire WX8730;
wire II31537;
wire II10945;
wire WX2962;
wire WX1545;
wire WX7021;
wire WX8722;
wire II30240;
wire WX6608;
wire WX10276;
wire WX10170;
wire WX3177;
wire WX6562;
wire WX2207;
wire WX3884;
wire II34044;
wire WX11569;
wire II6380;
wire WX9943;
wire WX601;
wire WX11374;
wire II10138;
wire WX7325;
wire II3563;
wire WX5652;
wire WX3980;
wire II2777;
wire WX4585;
wire WX7345;
wire WX8969;
wire II27677;
wire II18852;
wire WX10555;
wire WX7273;
wire WX7986;
wire WX6701;
wire WX2990;
wire WX11405;
wire II34843;
wire II11488;
wire II26366;
wire WX3036;
wire II14732;
wire II22325;
wire II18691;
wire WX7064;
wire II14802;
wire II10526;
wire II18255;
wire WX2712;
wire WX7546;
wire WX981;
wire WX7505;
wire WX8691;
wire WX11267;
wire WX6695;
wire II34030;
wire WX11583;
wire WX6332;
wire WX8347;
wire WX2266;
wire II10324;
wire WX9145;
wire WX7624;
wire WX6203;
wire II26423;
wire WX174;
wire WX2258;
wire II6046;
wire WX254;
wire II27698;
wire WX2542;
wire II19626;
wire WX2197;
wire WX9927;
wire II30559;
wire II10392;
wire II34677;
wire WX915;
wire WX972;
wire II15580;
wire WX4985;
wire II30899;
wire II7123;
wire WX4488;
wire II30528;
wire WX9360;
wire WX4936;
wire II34972;
wire WX10523;
wire WX4733;
wire WX6604;
wire WX7511;
wire WX6366;
wire WX1178;
wire WX5529;
wire WX6425;
wire WX4441;
wire WX7636;
wire WX8338;
wire II27586;
wire WX7489;
wire II26034;
wire II19661;
wire WX3057;
wire II10889;
wire WX3088;
wire II18860;
wire II26932;
wire II22517;
wire WX10463;
wire WX696;
wire II34168;
wire WX6193;
wire II2275;
wire WX11336;
wire WX6062;
wire WX7500;
wire II35261;
wire WX450;
wire WX4282;
wire II15725;
wire WX8795;
wire II34740;
wire WX7482;
wire II11205;
wire WX3132;
wire WX840;
wire WX3510;
wire II30178;
wire II26701;
wire II7504;
wire WX6665;
wire WX7465;
wire WX8314;
wire WX11216;
wire WX1564;
wire II3648;
wire WX1362;
wire II10169;
wire II19543;
wire WX4268;
wire II30619;
wire WX3500;
wire II18124;
wire WX5010;
wire WX1713;
wire WX11257;
wire WX4964;
wire WX11358;
wire WX2697;
wire WX7125;
wire WX8901;
wire WX9097;
wire WX1397;
wire WX2913;
wire II11494;
wire WX9640;
wire WX8861;
wire WX7611;
wire II7306;
wire WX11662;
wire II6449;
wire WX5564;
wire WX2451;
wire WX5071;
wire WX11320;
wire WX4785;
wire II30148;
wire WX8185;
wire II22774;
wire II2964;
wire II34555;
wire II10782;
wire II6351;
wire WX11562;
wire WX7315;
wire WX2887;
wire WX3270;
wire II14110;
wire WX2123;
wire II10930;
wire WX6177;
wire II19490;
wire WX6810;
wire WX8736;
wire WX9101;
wire II27357;
wire WX8821;
wire WX9480;
wire WX5339;
wire II10750;
wire WX4804;
wire WX2522;
wire WX734;
wire WX2735;
wire II34176;
wire WX9282;
wire WX10584;
wire WX5351;
wire II2165;
wire II6769;
wire WX1860;
wire WX2583;
wire II31544;
wire WX4715;
wire WX4466;
wire II19639;
wire WX8590;
wire WX3186;
wire WX6613;
wire WX11311;
wire II26857;
wire II26792;
wire WX7684;
wire II30363;
wire II35542;
wire WX4962;
wire WX6004;
wire WX4049;
wire II2553;
wire WX4094;
wire WX1392;
wire WX8446;
wire II35170;
wire WX3981;
wire II35549;
wire WX7572;
wire WX6498;
wire WX9221;
wire WX10304;
wire II15392;
wire WX5270;
wire WX4041;
wire II14894;
wire WX2191;
wire WX6400;
wire II10696;
wire WX11475;
wire WX3805;
wire WX2575;
wire WX953;
wire II14971;
wire II30960;
wire WX99;
wire WX5898;
wire WX1844;
wire WX5802;
wire II10864;
wire WX6628;
wire WX11381;
wire WX1911;
wire WX10671;
wire II2120;
wire WX10391;
wire WX8626;
wire II2219;
wire WX4241;
wire II2405;
wire II10310;
wire II22540;
wire WX5641;
wire WX10949;
wire WX6253;
wire II34990;
wire II30434;
wire WX3599;
wire WX9652;
wire II35511;
wire II30387;
wire II18900;
wire WX9109;
wire II7610;
wire II31641;
wire II22338;
wire II14134;
wire II6925;
wire WX5796;
wire WX5972;
wire WX10733;
wire II19346;
wire WX995;
wire WX6276;
wire II18604;
wire WX5645;
wire WX8373;
wire WX1603;
wire II14470;
wire II6474;
wire WX1678;
wire WX3577;
wire WX9157;
wire WX6856;
wire II10950;
wire WX10044;
wire II34066;
wire II34415;
wire II2376;
wire II23300;
wire II31505;
wire WX6774;
wire II31696;
wire II6249;
wire WX1367;
wire II11581;
wire II26762;
wire WX1070;
wire WX4597;
wire II6511;
wire WX1536;
wire WX5571;
wire II6697;
wire WX10635;
wire WX9185;
wire WX10406;
wire II6620;
wire WX4145;
wire WX249;
wire WX6514;
wire WX6830;
wire WX5541;
wire II22044;
wire II34836;
wire WX7177;
wire II10268;
wire WX6636;
wire WX10535;
wire WX430;
wire WX2067;
wire WX6352;
wire II6242;
wire II7569;
wire WX7898;
wire WX6478;
wire II26925;
wire II14097;
wire II18092;
wire WX8729;
wire II6458;
wire WX11427;
wire WX5856;
wire WX6516;
wire WX6877;
wire WX1598;
wire WX2936;
wire WX942;
wire WX4549;
wire WX7722;
wire WX4189;
wire WX2866;
wire II26507;
wire WX1735;
wire WX5371;
wire WX5791;
wire WX3338;
wire WX6410;
wire II14683;
wire WX9443;
wire WX10280;
wire WX4187;
wire WX3718;
wire WX7474;
wire II30814;
wire II18905;
wire WX5310;
wire II27691;
wire II23512;
wire WX10120;
wire WX307;
wire WX4830;
wire II14342;
wire WX4784;
wire II11659;
wire WX5553;
wire WX1003;
wire II30114;
wire II22487;
wire II7528;
wire WX8652;
wire II26825;
wire II30295;
wire WX10868;
wire WX6240;
wire WX4855;
wire WX7813;
wire II22889;
wire II5994;
wire WX3208;
wire II34749;
wire WX10485;
wire II30612;
wire WX6584;
wire WX5031;
wire WX8282;
wire WX9829;
wire II34460;
wire WX2505;
wire II10098;
wire WX10183;
wire WX7089;
wire WX1865;
wire II31521;
wire II10160;
wire WX11286;
wire WX10668;
wire II30040;
wire II34786;
wire WX7443;
wire WX1264;
wire II3593;
wire WX137;
wire WX313;
wire WX2641;
wire II7570;
wire WX11581;
wire WX9383;
wire WX7088;
wire II14017;
wire WX3507;
wire II6785;
wire II15120;
wire WX4077;
wire II7674;
wire II30867;
wire WX4455;
wire II6573;
wire II10713;
wire WX42;
wire II30473;
wire WX8381;
wire WX9127;
wire WX9163;
wire II10340;
wire II18247;
wire II19611;
wire II7267;
wire WX5549;
wire II19165;
wire WX8940;
wire WX3629;
wire WX9272;
wire WX8458;
wire II7083;
wire WX758;
wire II14175;
wire II31141;
wire II10842;
wire WX2300;
wire II22709;
wire WX5770;
wire WX6809;
wire II19640;
wire WX1503;
wire II27650;
wire WX2097;
wire WX2630;
wire II7654;
wire WX9672;
wire WX7844;
wire WX8377;
wire WX8893;
wire WX10287;
wire WX10954;
wire WX933;
wire WX6769;
wire WX7640;
wire WX5922;
wire II23604;
wire WX9232;
wire WX3939;
wire II30696;
wire II26429;
wire WX129;
wire WX374;
wire WX8110;
wire II34352;
wire WX204;
wire WX10429;
wire WX10970;
wire WX3346;
wire WX6907;
wire II35610;
wire II15502;
wire II30737;
wire WX2338;
wire II34547;
wire II2353;
wire WX10675;
wire WX10803;
wire WX6617;
wire WX4463;
wire WX6943;
wire WX8196;
wire WX9984;
wire II14692;
wire WX4840;
wire WX10632;
wire WX6533;
wire WX7964;
wire WX2029;
wire WX6543;
wire WX2179;
wire WX6430;
wire WX324;
wire II30326;
wire WX196;
wire II26404;
wire II2362;
wire WX7434;
wire II26182;
wire WX5725;
wire II10418;
wire WX4757;
wire WX5098;
wire II34091;
wire WX10852;
wire II6915;
wire WX5786;
wire WX9593;
wire WX1644;
wire II35570;
wire II2196;
wire WX9189;
wire II14708;
wire II23729;
wire II30672;
wire II22345;
wire II27643;
wire WX4219;
wire WX9153;
wire WX9520;
wire WX3706;
wire WX3166;
wire WX5283;
wire WX10800;
wire II3523;
wire II34603;
wire II22578;
wire II22294;
wire WX10590;
wire II26189;
wire WX8970;
wire WX5764;
wire WX10033;
wire WX10702;
wire WX2807;
wire WX2901;
wire WX1673;
wire WX2758;
wire WX2239;
wire II18807;
wire WX2660;
wire II34693;
wire II6288;
wire II19536;
wire II22662;
wire WX6692;
wire II35660;
wire II6110;
wire WX9636;
wire II6878;
wire WX905;
wire WX9266;
wire WX4569;
wire WX5614;
wire II26211;
wire WX1422;
wire WX4007;
wire WX3047;
wire II2842;
wire WX8101;
wire II7345;
wire II6751;
wire WX6936;
wire WX10097;
wire II7497;
wire WX870;
wire II10812;
wire WX7779;
wire II35533;
wire II34051;
wire WX8099;
wire II26739;
wire WX7761;
wire WX965;
wire II22384;
wire II18030;
wire WX10782;
wire II3235;
wire WX9773;
wire II18676;
wire II34423;
wire WX9484;
wire WX4998;
wire II15683;
wire II34191;
wire WX4395;
wire WX1902;
wire WX1322;
wire WX10394;
wire WX10985;
wire WX9395;
wire WX810;
wire II27201;
wire WX2339;
wire WX7143;
wire WX9132;
wire WX2276;
wire II26607;
wire WX338;
wire WX1481;
wire WX5079;
wire WX5618;
wire II18395;
wire II10276;
wire WX8218;
wire WX7183;
wire II30789;
wire WX1698;
wire WX6168;
wire II15635;
wire WX10508;
wire II6581;
wire WX3617;
wire II35674;
wire II7625;
wire II10061;
wire WX6719;
wire WX10361;
wire II14082;
wire II14918;
wire WX9599;
wire WX7055;
wire II14306;
wire WX1223;
wire WX6857;
wire WX1637;
wire WX8851;
wire II35183;
wire II14136;
wire II6754;
wire WX4310;
wire WX7455;
wire WX4377;
wire WX6957;
wire WX2250;
wire WX5215;
wire II11220;
wire WX6792;
wire II3392;
wire II10083;
wire WX10850;
wire II19592;
wire WX11262;
wire WX9084;
wire WX408;
wire WX10153;
wire II14623;
wire WX8785;
wire II10027;
wire WX3486;
wire WX5057;
wire WX8434;
wire WX2491;
wire WX3741;
wire WX2762;
wire WX1851;
wire II31726;
wire WX6125;
wire WX3394;
wire II34632;
wire WX7700;
wire WX9309;
wire II30775;
wire WX3212;
wire II2207;
wire WX11448;
wire WX3584;
wire II22765;
wire WX3956;
wire II18847;
wire II34647;
wire II14498;
wire II30263;
wire II18289;
wire WX3144;
wire WX7692;
wire WX9518;
wire WX7789;
wire II30713;
wire II18505;
wire II30428;
wire WX3759;
wire II6055;
wire WX10511;
wire II6816;
wire II26947;
wire II14234;
wire WX6233;
wire II18239;
wire WX714;
wire II22254;
wire II34725;
wire WX4098;
wire II15620;
wire WX8636;
wire II26950;
wire WX6104;
wire WX3951;
wire WX5384;
wire WX321;
wire WX589;
wire WX7673;
wire WX11323;
wire WX2389;
wire II18836;
wire WX5159;
wire WX7536;
wire WX10455;
wire WX1857;
wire WX3519;
wire WX8224;
wire WX580;
wire II6365;
wire WX2442;
wire WX10655;
wire WX9478;
wire II26311;
wire WX5254;
wire WX2415;
wire II6102;
wire WX4127;
wire II6047;
wire WX1740;
wire WX4449;
wire WX7033;
wire II22758;
wire II19202;
wire II26993;
wire WX2293;
wire WX6470;
wire II30125;
wire II2057;
wire WX11394;
wire II35597;
wire WX7096;
wire WX7420;
wire WX5769;
wire II31425;
wire WX10026;
wire WX3362;
wire WX3987;
wire II27356;
wire WX5538;
wire II30024;
wire WX9205;
wire WX3768;
wire II23326;
wire II26151;
wire WX8876;
wire WX9743;
wire II27381;
wire II3104;
wire WX6418;
wire II14716;
wire WX10595;
wire II27173;
wire WX4773;
wire WX6712;
wire WX2892;
wire WX3770;
wire WX11516;
wire WX1347;
wire II31654;
wire WX7510;
wire WX8894;
wire II31000;
wire WX1120;
wire WX5223;
wire WX9789;
wire WX8355;
wire WX2675;
wire WX5133;
wire WX6038;
wire WX1625;
wire II30688;
wire WX9438;
wire WX10605;
wire WX10351;
wire WX8490;
wire II23142;
wire WX10149;
wire II6777;
wire WX11457;
wire II2911;
wire II15353;
wire WX7858;
wire II26141;
wire WX4349;
wire WX1129;
wire WX10624;
wire WX10414;
wire II22139;
wire II27472;
wire WX11421;
wire WX8450;
wire WX1256;
wire WX7113;
wire WX3678;
wire WX10266;
wire II15186;
wire II15592;
wire WX8133;
wire WX59;
wire II10827;
wire WX5682;
wire WX2049;
wire WX334;
wire WX9242;
wire WX11016;
wire WX6633;
wire WX2597;
wire WX7587;
wire II15472;
wire WX11439;
wire WX3829;
wire II10744;
wire WX9975;
wire WX8678;
wire II23183;
wire WX6503;
wire II26435;
wire II26374;
wire WX5147;
wire WX9450;
wire WX446;
wire WX11587;
wire WX4494;
wire WX5452;
wire WX2394;
wire II14327;
wire WX11628;
wire II2002;
wire WX8021;
wire WX6391;
wire WX5499;
wire II6498;
wire II26631;
wire II34865;
wire II22679;
wire II11115;
wire WX11266;
wire WX7207;
wire WX7717;
wire II18930;
wire WX2786;
wire WX158;
wire WX11318;
wire II22160;
wire WX4515;
wire II5992;
wire WX10206;
wire II14562;
wire WX6147;
wire WX8790;
wire II31217;
wire WX1051;
wire II22185;
wire II22356;
wire WX5058;
wire II35222;
wire WX6187;
wire WX5670;
wire WX7497;
wire WX9467;
wire WX4157;
wire II27573;
wire WX8410;
wire WX1141;
wire WX10055;
wire II26035;
wire WX8675;
wire II19605;
wire WX9367;
wire WX958;
wire WX9349;
wire II23494;
wire WX282;
wire WX526;
wire WX2862;
wire WX7403;
wire WX9196;
wire WX11496;
wire II30681;
wire II11467;
wire II27485;
wire WX368;
wire II19505;
wire WX1168;
wire II2197;
wire WX2895;
wire WX8935;
wire WX5417;
wire WX7798;
wire II3274;
wire WX8390;
wire WX7797;
wire WX3896;
wire WX10895;
wire II18537;
wire II14336;
wire II14491;
wire II14182;
wire WX2653;
wire WX2374;
wire WX2063;
wire WX10648;
wire II6017;
wire II10681;
wire II14103;
wire II35444;
wire II2508;
wire WX4821;
wire WX11419;
wire WX11618;
wire WX9527;
wire II15302;
wire WX469;
wire WX2262;
wire WX10910;
wire WX2322;
wire II15697;
wire WX8912;
wire II34088;
wire WX7594;
wire WX1185;
wire II23131;
wire WX8397;
wire II22920;
wire II6250;
wire II7291;
wire WX5278;
wire WX11144;
wire WX1704;
wire II11587;
wire II18449;
wire WX9265;
wire WX9459;
wire WX8934;
wire WX9397;
wire WX4435;
wire II26606;
wire WX3725;
wire WX2961;
wire II6162;
wire II2918;
wire WX4675;
wire II7716;
wire WX363;
wire WX11078;
wire WX6779;
wire II14275;
wire II34733;
wire II2730;
wire WX11525;
wire WX10450;
wire II27277;
wire II22572;
wire WX10248;
wire WX10842;
wire WX5140;
wire II14547;
wire WX6863;
wire WX3104;
wire WX2958;
wire WX6288;
wire II34253;
wire II11708;
wire WX3921;
wire WX3382;
wire II6255;
wire II26065;
wire WX8858;
wire II14779;
wire II7240;
wire WX5245;
wire WX9719;
wire WX3608;
wire II30255;
wire WX3773;
wire WX6229;
wire II34430;
wire II6713;
wire WX5409;
wire WX6074;
wire WX395;
wire II26112;
wire WX6829;
wire WX7975;
wire II35569;
wire II14461;
wire WX504;
wire II10144;
wire WX10125;
wire II10399;
wire II10058;
wire WX5594;
wire WX4025;
wire WX2829;
wire WX7382;
wire WX8256;
wire II34150;
wire WX10086;
wire WX1666;
wire WX5668;
wire II22735;
wire II18288;
wire II30828;
wire II30846;
wire II3656;
wire II23672;
wire WX2921;
wire II27741;
wire II18459;
wire WX8687;
wire WX4140;
wire II30279;
wire WX10957;
wire II10441;
wire II15642;
wire WX4492;
wire II34833;
wire II22479;
wire WX6380;
wire II2816;
wire II7639;
wire II34376;
wire II19716;
wire WX4912;
wire WX10388;
wire WX1081;
wire WX3684;
wire WX6854;
wire II15082;
wire WX10409;
wire WX290;
wire WX1593;
wire WX4633;
wire II15670;
wire WX6321;
wire WX3242;
wire II2537;
wire WX6921;
wire WX472;
wire WX4322;
wire II14243;
wire II2159;
wire II34905;
wire WX312;
wire WX2449;
wire WX3372;
wire WX6140;
wire II31668;
wire WX9531;
wire WX5366;
wire WX3957;
wire II14838;
wire WX9859;
wire II10284;
wire WX4914;
wire II2754;
wire II10183;
wire WX7811;
wire WX10973;
wire WX10381;
wire WX4623;
wire II6875;
wire WX9113;
wire II23714;
wire II6952;
wire WX8048;
wire WX9699;
wire II27161;
wire II7214;
wire WX11577;
wire WX1426;
wire WX4832;
wire II7097;
wire WX10577;
wire WX3782;
wire WX9617;
wire WX1518;
wire WX409;
wire WX3815;
wire II10368;
wire WX5113;
wire WX9327;
wire WX10476;
wire II22029;
wire II23651;
wire WX4997;
wire WX8868;
wire WX4289;
wire WX8395;
wire WX1015;
wire WX5479;
wire II34368;
wire II22501;
wire II34805;
wire WX7973;
wire WX9803;
wire WX10884;
wire WX6257;
wire II11128;
wire II7435;
wire II34414;
wire II3484;
wire WX49;
wire WX3240;
wire WX6745;
wire WX8083;
wire II30270;
wire WX7642;
wire WX10230;
wire WX8043;
wire WX11575;
wire II31705;
wire WX2939;
wire WX1912;
wire II14026;
wire WX9154;
wire WX6629;
wire WX6831;
wire WX7805;
wire WX9419;
wire II3516;
wire WX1435;
wire WX1018;
wire II6210;
wire WX2367;
wire WX7951;
wire WX10278;
wire WX5934;
wire WX6374;
wire WX6345;
wire II26258;
wire WX1373;
wire WX11150;
wire II34447;
wire WX4102;
wire WX5268;
wire II9997;
wire II18279;
wire II11699;
wire WX10902;
wire II2222;
wire WX5049;
wire II22897;
wire II31387;
wire WX5108;
wire WX4818;
wire WX104;
wire II26512;
wire II31733;
wire WX1849;
wire WX632;
wire II23547;
wire II6482;
wire II18735;
wire WX10666;
wire WX7573;
wire II18549;
wire WX9567;
wire II11064;
wire WX2101;
wire WX9701;
wire WX10290;
wire II6815;
wire II3600;
wire II6022;
wire WX7911;
wire WX10938;
wire WX11500;
wire II22161;
wire WX6804;
wire II2377;
wire WX215;
wire II7687;
wire II14684;
wire II6186;
wire WX3005;
wire II10262;
wire II22495;
wire WX3622;
wire WX10400;
wire WX8966;
wire II23534;
wire WX3592;
wire WX7841;
wire WX9277;
wire WX11493;
wire II14203;
wire WX8064;
wire II15545;
wire WX1263;
wire II18874;
wire WX2329;
wire WX9118;
wire II18464;
wire II18605;
wire II14569;
wire II22369;
wire WX1175;
wire WX5576;
wire II7071;
wire II10968;
wire WX11478;
wire WX6928;
wire II34493;
wire II7280;
wire II2718;
wire WX6592;
wire WX9135;
wire WX4110;
wire II26133;
wire II14755;
wire II2933;
wire II11512;
wire WX2353;
wire II10857;
wire WX1785;
wire II34408;
wire WX11280;
wire II19345;
wire II2562;
wire II22362;
wire WX7791;
wire WX1108;
wire II10487;
wire WX2643;
wire WX4828;
wire II22407;
wire WX439;
wire II2329;
wire WX3574;
wire II18868;
wire WX7556;
wire II18146;
wire II14592;
wire II6310;
wire II10337;
wire WX9915;
wire II18303;
wire WX11174;
wire II14280;
wire WX4389;
wire II35470;
wire WX8983;
wire II30364;
wire II22123;
wire II11685;
wire WX11414;
wire WX7634;
wire WX9004;
wire WX9074;
wire II34200;
wire WX4158;
wire WX6271;
wire WX4442;
wire II10571;
wire WX7884;
wire WX3086;
wire II14415;
wire II11665;
wire WX11553;
wire II30053;
wire II3698;
wire II34624;
wire WX3928;
wire WX10566;
wire II14901;
wire II15607;
wire WX6991;
wire WX10072;
wire II30139;
wire WX9965;
wire WX4086;
wire WX3286;
wire II22376;
wire WX10112;
wire WX11036;
wire II31153;
wire WX9614;
wire WX2639;
wire WX1965;
wire WX10163;
wire WX3870;
wire II10890;
wire II30155;
wire WX10941;
wire WX616;
wire WX11365;
wire WX2204;
wire WX4709;
wire II6821;
wire WX1520;
wire WX7020;
wire II6739;
wire II6536;
wire WX948;
wire II14530;
wire II34042;
wire II10471;
wire WX6262;
wire II31577;
wire WX5557;
wire II7384;
wire WX1409;
wire WX2769;
wire WX6725;
wire WX1330;
wire WX8979;
wire WX4105;
wire WX8808;
wire WX2311;
wire WX3762;
wire WX5732;
wire II6691;
wire II10186;
wire II34123;
wire II11481;
wire WX3276;
wire WX5443;
wire II18316;
wire II34153;
wire WX10171;
wire WX8826;
wire II30727;
wire II19293;
wire WX11598;
wire WX1380;
wire WX11168;
wire II30588;
wire WX163;
wire WX4667;
wire WX3536;
wire WX7515;
wire WX5550;
wire WX4780;
wire WX7484;
wire II34681;
wire WX4246;
wire II34036;
wire WX6505;
wire WX6656;
wire WX6911;
wire WX11196;
wire WX4525;
wire II14404;
wire WX5080;
wire WX5497;
wire II14529;
wire WX2585;
wire WX559;
wire II22447;
wire II27538;
wire WX11114;
wire II31557;
wire II34324;
wire II22649;
wire II15146;
wire WX2539;
wire II23079;
wire WX5381;
wire WX8042;
wire WX10528;
wire WX9089;
wire II22634;
wire II11101;
wire II34523;
wire II6521;
wire WX9843;
wire WX1400;
wire WX6967;
wire II23234;
wire WX3050;
wire WX932;
wire WX4069;
wire WX11535;
wire II22393;
wire WX1550;
wire WX11570;
wire WX2296;
wire WX5465;
wire WX8260;
wire WX9018;
wire WX6198;
wire WX2530;
wire WX4971;
wire II26592;
wire II30441;
wire WX3217;
wire WX1527;
wire WX5040;
wire II35301;
wire WX4292;
wire II22914;
wire WX11551;
wire WX1290;
wire WX8230;
wire WX10343;
wire WX5361;
wire II31258;
wire WX10015;
wire II6852;
wire WX10226;
wire WX4214;
wire II23716;
wire II10921;
wire WX4035;
wire II31536;
wire WX646;
wire WX5312;
wire WX168;
wire II3339;
wire WX8306;
wire II30860;
wire II15303;
wire WX7153;
wire II18226;
wire WX8236;
wire II3675;
wire WX7629;
wire WX2775;
wire WX4796;
wire II11552;
wire II2152;
wire II6660;
wire WX6705;
wire WX2996;
wire II2772;
wire WX7945;
wire WX3434;
wire WX6161;
wire II30930;
wire II27672;
wire WX8897;
wire WX1337;
wire WX7065;
wire WX1805;
wire WX5026;
wire WX11274;
wire WX4689;
wire WX11292;
wire WX2682;
wire WX561;
wire WX1578;
wire II10961;
wire II15094;
wire WX1773;
wire WX3308;
wire II26940;
wire WX8520;
wire WX10205;
wire WX6094;
wire WX8468;
wire WX1557;
wire WX680;
wire II26646;
wire WX1943;
wire II30893;
wire II26543;
wire WX854;
wire II34061;
wire II31676;
wire II2455;
wire WX7448;
wire WX975;
wire II30334;
wire II26529;
wire WX1901;
wire WX6369;
wire II34471;
wire WX8024;
wire WX4273;
wire II6202;
wire WX6462;
wire WX10048;
wire II22648;
wire II35004;
wire WX4869;
wire WX8910;
wire II10036;
wire WX7804;
wire WX8345;
wire WX6746;
wire WX9606;
wire WX1497;
wire II14197;
wire WX4909;
wire II27370;
wire WX3061;
wire WX7013;
wire WX2424;
wire II2082;
wire WX10300;
wire WX1488;
wire II22880;
wire WX3256;
wire WX6209;
wire II35689;
wire WX5119;
wire WX8841;
wire WX11385;
wire WX9180;
wire WX1618;
wire WX1344;
wire WX5515;
wire WX5236;
wire II10330;
wire WX7840;
wire WX6200;
wire II11401;
wire II26636;
wire II2694;
wire II18072;
wire II10766;
wire WX11250;
wire WX6295;
wire II7122;
wire WX3019;
wire WX5294;
wire II26082;
wire II18774;
wire WX5003;
wire II34476;
wire II34215;
wire II6194;
wire II15579;
wire WX9919;
wire WX6770;
wire WX113;
wire II22533;
wire II31520;
wire WX6421;
wire II10650;
wire II27383;
wire II22099;
wire WX9683;
wire II26078;
wire II11616;
wire WX4031;
wire WX7566;
wire II26833;
wire II15558;
wire WX5437;
wire WX3601;
wire II22601;
wire WX11540;
wire II11575;
wire WX3418;
wire WX11532;
wire WX8512;
wire II15432;
wire II2656;
wire II2097;
wire II30982;
wire WX1939;
wire II14073;
wire WX10539;
wire II18890;
wire WX7991;
wire WX3612;
wire WX2403;
wire WX267;
wire WX3735;
wire II18270;
wire WX6115;
wire WX8546;
wire WX6159;
wire WX2591;
wire II22781;
wire WX10490;
wire WX6641;
wire WX2626;
wire WX4367;
wire WX7757;
wire II7474;
wire II10625;
wire WX7139;
wire II2709;
wire WX2334;
wire II11285;
wire WX11400;
wire II6270;
wire II26654;
wire WX8905;
wire WX342;
wire II14963;
wire WX6915;
wire WX2310;
wire WX8924;
wire WX1471;
wire WX8600;
wire WX7024;
wire II34113;
wire WX6995;
wire II35695;
wire WX7582;
wire II2234;
wire II2927;
wire WX1132;
wire WX2455;
wire II14266;
wire II30976;
wire WX7832;
wire II18666;
wire II18364;
wire WX5330;
wire WX11180;
wire WX8079;
wire WX4299;
wire WX475;
wire WX147;
wire WX3094;
wire WX7894;
wire II14886;
wire WX2241;
wire WX7392;
wire WX5598;
wire II35617;
wire WX2202;
wire II19654;
wire WX9956;
wire WX1062;
wire II2265;
wire II2346;
wire WX10921;
wire II15368;
wire WX6872;
wire WX4988;
wire II34920;
wire II19477;
wire WX5848;
wire WX4691;
wire WX6406;
wire WX7651;
wire WX10915;
wire WX5916;
wire WX6733;
wire II30998;
wire II6862;
wire WX4897;
wire II10492;
wire WX5096;
wire WX8835;
wire II22239;
wire WX4288;
wire II15585;
wire WX10497;
wire II30083;
wire WX6340;
wire II27700;
wire WX744;
wire WX5962;
wire WX10222;
wire WX8731;
wire WX5091;
wire WX7825;
wire WX8036;
wire WX8076;
wire WX8033;
wire WX3149;
wire WX8950;
wire II3353;
wire II35576;
wire II2515;
wire WX3606;
wire II22626;
wire II2570;
wire II26600;
wire WX11539;
wire II22888;
wire II11560;
wire WX9400;
wire II14792;
wire II26128;
wire WX9753;
wire WX149;
wire WX2820;
wire II30179;
wire WX2966;
wire II10509;
wire WX2670;
wire WX4231;
wire WX3748;
wire II22896;
wire II11335;
wire WX10142;
wire WX9168;
wire WX8995;
wire II26560;
wire WX2940;
wire WX3837;
wire WX9739;
wire WX2284;
wire II19281;
wire II18968;
wire II18805;
wire WX4896;
wire II27446;
wire WX5485;
wire WX6979;
wire II34198;
wire WX463;
wire II6426;
wire II14375;
wire WX11453;
wire WX6760;
wire II26242;
wire WX4888;
wire II7667;
wire WX8154;
wire WX5690;
wire WX2281;
wire WX8773;
wire II26987;
wire WX5257;
wire WX9492;
wire II2020;
wire II27706;
wire WX8174;
wire WX3193;
wire WX1611;
wire WX417;
wire WX3506;
wire II18031;
wire II18705;
wire II3286;
wire II22725;
wire II27636;
wire II3262;
wire WX10726;
wire WX8123;
wire II18728;
wire II14001;
wire WX9408;
wire WX294;
wire WX9158;
wire WX5930;
wire II14600;
wire II2183;
wire WX10217;
wire WX9624;
wire WX11580;
wire WX2516;
wire II10238;
wire WX1211;
wire WX5580;
wire WX9970;
wire WX5483;
wire WX11348;
wire II18643;
wire II10307;
wire WX3631;
wire WX8800;
wire WX1143;
wire II15406;
wire WX10037;
wire WX9210;
wire WX8694;
wire II19358;
wire WX5306;
wire II3711;
wire WX5506;
wire II23312;
wire II22585;
wire WX246;
wire WX427;
wire WX3673;
wire II23567;
wire WX10077;
wire WX6301;
wire II26623;
wire WX8701;
wire WX662;
wire WX4503;
wire WX4136;
wire WX8666;
wire II30666;
wire WX7407;
wire II26158;
wire II14630;
wire II10299;
wire II10796;
wire WX7447;
wire II15316;
wire WX5420;
wire WX492;
wire WX3944;
wire II19373;
wire WX2771;
wire II34184;
wire WX11379;
wire WX6841;
wire WX2985;
wire WX2165;
wire WX11098;
wire WX8707;
wire II27212;
wire WX9995;
wire II26119;
wire WX5405;
wire II18387;
wire WX7079;
wire WX10131;
wire II34889;
wire WX8642;
wire II22232;
wire II18816;
wire WX9901;
wire II22067;
wire II34944;
wire II22927;
wire II18294;
wire II10751;
wire WX9149;
wire WX11433;
wire WX10307;
wire WX5828;
wire II22828;
wire II14430;
wire II14607;
wire II31628;
wire II31321;
wire II19242;
wire II34888;
wire WX9285;
wire II26344;
wire WX2953;
wire WX9297;
wire WX3560;
wire WX7927;
wire WX11382;
wire II22910;
wire WX2382;
wire II10510;
wire WX3324;
wire II19137;
wire WX2740;
wire II26585;
wire II10447;
wire WX8791;
wire II26810;
wire II27721;
wire II30355;
wire II30552;
wire II26450;
wire II11140;
wire WX350;
wire WX1655;
wire II31612;
wire II6387;
wire WX9817;
wire WX2878;
wire II14652;
wire II15341;
wire WX6900;
wire WX3139;
wire WX3692;
wire WX9799;
wire WX86;
wire WX1046;
wire WX8763;
wire II19702;
wire II2904;
wire II23617;
wire WX275;
wire WX63;
wire WX11442;
wire WX5664;
wire II10114;
wire II27509;
wire WX7438;
wire II26678;
wire WX5398;
wire II26722;
wire II2973;
wire WX5782;
wire II34615;
wire II18164;
wire II2965;
wire II23352;
wire II19177;
wire WX352;
wire WX7567;
wire WX4078;
wire II22262;
wire II3500;
wire WX11134;
wire II22020;
wire II2701;
wire WX7366;
wire WX9769;
wire WX6398;
wire WX1154;
wire II14188;
wire WX4948;
wire WX8880;
wire WX6808;
wire II22835;
wire WX2871;
wire WX1971;
wire WX4419;
wire WX10637;
wire II6503;
wire WX8658;
wire II6760;
wire WX2605;
wire II6844;
wire WX10375;
wire WX188;
wire II23105;
wire WX10710;
wire WX9725;
wire II7175;
wire II10595;
wire WX223;
wire WX1721;
wire II22974;
wire II14811;
wire WX11238;
wire WX181;
wire II19499;
wire II30132;
wire WX9253;
wire WX2475;
wire II34329;
wire WX3250;
wire WX9175;
wire WX5126;
wire WX8013;
wire WX1755;
wire II15119;
wire WX8952;
wire WX7287;
wire II6831;
wire II34331;
wire II30403;
wire WX2483;
wire II2878;
wire II2723;
wire WX993;
wire WX6239;
wire II6721;
wire II6026;
wire II10937;
wire WX3503;
wire II18041;
wire II31627;
wire WX8117;
wire WX10468;
wire WX4337;
wire WX5444;
wire II6332;
wire II34262;
wire WX10617;
wire WX8164;
wire WX8746;
wire WX6132;
wire WX1511;
wire II30838;
wire II34075;
wire WX2325;
wire WX5137;
wire WX4645;
wire WX1239;
wire WX2225;
wire WX9338;
wire II35365;
wire II26360;
wire WX8454;
wire WX798;
wire II26567;
wire WX1306;
wire WX4862;
wire WX10719;
wire II2251;
wire WX8262;
wire WX2851;
wire WX4090;
wire WX11024;
wire II30720;
wire WX11373;
wire WX7666;
wire II14454;
wire WX866;
wire WX4045;
wire II2848;
wire II18937;
wire WX8051;
wire WX11505;
wire II3144;
wire WX9777;
wire WX1412;
wire II10781;
wire WX7419;
wire WX8227;
wire II34711;
wire II26964;
wire WX10395;
wire WX1546;
wire WX5391;
wire WX4474;
wire II6071;
wire II10362;
wire WX9657;
wire II18022;
wire II22418;
wire II2289;
wire WX2842;
wire II15494;
wire II3543;
wire WX4851;
wire WX10481;
wire WX8137;
wire WX9387;
wire WX4161;
wire WX1429;
wire WX7084;
wire WX5567;
wire II6084;
wire WX7918;
wire II30171;
wire WX4225;
wire WX6308;
wire WX8004;
wire II2010;
wire WX7047;
wire WX1247;
wire II3156;
wire WX1561;
wire WX3809;
wire WX7121;
wire II18347;
wire II2258;
wire WX10160;
wire WX678;
wire WX10262;
wire WX5432;
wire II23709;
wire WX5712;
wire WX5716;
wire WX5948;
wire WX2269;
wire WX2210;
wire WX3644;
wire II27305;
wire WX1991;
wire WX11042;
wire WX1674;
wire II18178;
wire II31661;
wire WX5852;
wire WX3232;
wire WX8740;
wire WX8100;
wire WX3048;
wire II6597;
wire WX5379;
wire WX9502;
wire II35482;
wire WX10791;
wire II35668;
wire WX5201;
wire WX1218;
wire WX641;
wire II10517;
wire WX5354;
wire WX8534;
wire WX1684;
wire WX9048;
wire II14746;
wire WX4719;
wire WX1304;
wire WX8739;
wire II26748;
wire II34107;
wire WX7552;
wire WX6085;
wire WX9092;
wire II19718;
wire WX3174;
wire WX11411;
wire WX1268;
wire WX3398;
wire WX480;
wire WX10107;
wire WX7705;
wire WX4183;
wire WX7658;
wire WX4073;
wire WX94;
wire WX9881;
wire WX2219;
wire II6916;
wire II6394;
wire WX8181;
wire WX2343;
wire WX70;
wire WX6088;
wire WX9376;
wire WX10501;
wire WX5807;
wire WX6588;
wire WX9167;
wire II18722;
wire WX1606;
wire WX4184;
wire WX8646;
wire WX5304;
wire WX3490;
wire II2420;
wire WX4355;
wire WX898;
wire WX4938;
wire WX3994;
wire II22803;
wire II6411;
wire II22198;
wire WX6211;
wire II14158;
wire II10712;
wire WX10006;
wire WX4298;
wire WX2033;
wire WX6754;
wire WX7085;
wire WX10002;
wire WX9009;
wire WX3707;
wire WX5548;
wire WX6357;
wire WX5060;
wire WX7493;
wire WX4304;
wire II18023;
wire WX5519;
wire II35525;
wire WX3497;
wire II19627;
wire WX11314;
wire WX2077;
wire WX3976;
wire WX7833;
wire WX7649;
wire WX10744;
wire II10059;
wire WX6319;
wire II7527;
wire WX157;
wire WX4327;
wire WX478;
wire WX3204;
wire WX10022;
wire WX7321;
wire II18909;
wire WX11307;
wire II6289;
wire II18822;
wire WX10570;
wire II19308;
wire II35417;
wire II26864;
wire WX7726;
wire WX1112;
wire WX8016;
wire II31606;
wire WX9447;
wire WX6250;
wire WX6311;
wire WX1447;
wire WX6008;
wire WX11249;
wire WX9509;
wire WX5976;
wire II18582;
wire WX9123;
wire II14126;
wire WX10488;
wire WX10284;
wire WX6811;
wire II27523;
wire WX10243;
wire WX2509;
wire WX1580;
wire WX3653;
wire WX5402;
wire II6627;
wire WX10182;
wire WX4883;
wire WX6903;
wire WX6143;
wire WX8464;
wire WX8385;
wire WX5674;
wire II18472;
wire II10480;
wire II7189;
wire WX11074;
wire WX1869;
wire WX5036;
wire WX3402;
wire II22244;
wire WX10950;
wire II23402;
wire WX937;
wire II22717;
wire II22710;
wire WX8570;
wire II3607;
wire II14251;
wire II18110;
wire WX3713;
wire II15613;
wire WX2304;
wire WX9676;
wire II26498;
wire WX3721;
wire WX10335;
wire II26051;
wire WX10969;
wire WX11568;
wire WX4581;
wire II15718;
wire WX8818;
wire II18015;
wire II14576;
wire II11363;
wire II10356;
wire II18149;
wire WX9684;
wire WX178;
wire II6704;
wire II23574;
wire WX10192;
wire WX6581;
wire II30412;
wire II31126;
wire WX7902;
wire WX1658;
wire WX5607;
wire WX3428;
wire WX8608;
wire II34988;
wire II10213;
wire II22221;
wire II14283;
wire II34485;
wire WX208;
wire II2173;
wire II7421;
wire WX8830;
wire II10478;
wire II10957;
wire II10177;
wire II22339;
wire WX2708;
wire II11658;
wire WX11607;
wire WX4980;
wire WX7167;
wire WX11332;
wire WX3364;
wire WX173;
wire II19724;
wire WX8865;
wire II30063;
wire II14609;
wire WX3845;
wire WX2151;
wire WX4849;
wire II14701;
wire WX1199;
wire WX10294;
wire WX2988;
wire II19634;
wire WX3817;
wire WX919;
wire II26800;
wire II18565;
wire II35603;
wire WX8310;
wire II15212;
wire WX9877;
wire II6341;
wire II11707;
wire II6302;
wire WX914;
wire WX9105;
wire WX3761;
wire II35484;
wire WX7932;
wire WX7211;
wire II15134;
wire WX6600;
wire WX3781;
wire II19620;
wire WX738;
wire WX8684;
wire WX4907;
wire WX5359;
wire WX5076;
wire WX7820;
wire WX3882;
wire WX10686;
wire WX1568;
wire II6039;
wire WX11295;
wire WX3468;
wire II30636;
wire WX8319;
wire WX4264;
wire II10632;
wire II7395;
wire II10502;
wire WX10818;
wire WX3225;
wire II22903;
wire WX902;
wire II6822;
wire II27679;
wire II22321;
wire II22177;
wire WX35;
wire WX10271;
wire II7084;
wire II31572;
wire II23722;
wire II22276;
wire WX8781;
wire WX5626;
wire WX8335;
wire WX1472;
wire II18568;
wire WX4340;
wire WX9495;
wire WX6350;
wire II11672;
wire WX6058;
wire II35717;
wire II26437;
wire WX8360;
wire WX9423;
wire II34539;
wire WX10188;
wire WX3068;
wire WX9923;
wire WX7620;
wire II14839;
wire II10534;
wire WX1282;
wire WX3888;
wire WX8780;
wire II14956;
wire WX4432;
wire II30915;
wire WX10169;
wire II6746;
wire WX9170;
wire WX6362;
wire WX11546;
wire WX722;
wire II31710;
wire WX7060;
wire II14229;
wire WX1363;
wire II7549;
wire WX5656;
wire WX3514;
wire WX11357;
wire WX10082;
wire II2749;
wire II27434;
wire WX454;
wire II19451;
wire WX604;
wire WX4968;
wire II2467;
wire WX3947;
wire II26087;
wire WX532;
wire II2337;
wire WX692;
wire WX556;
wire II6613;
wire WX3561;
wire WX2366;
wire II34934;
wire WX5698;
wire II18101;
wire WX510;
wire WX5739;
wire WX4453;
wire WX3268;
wire II30604;
wire WX7277;
wire WX7027;
wire II23103;
wire WX1088;
wire II23274;
wire WX8148;
wire WX11128;
wire WX10597;
wire II10253;
wire WX8556;
wire WX381;
wire II10540;
wire WX6669;
wire II6798;
wire II6301;
wire WX10371;
wire II30216;
wire WX1093;
wire WX560;
wire WX9645;
wire WX2690;
wire WX7319;
wire WX11483;
wire WX3967;
wire WX2731;
wire WX1541;
wire II19695;
wire II11692;
wire II18209;
wire WX5455;
wire II31512;
wire WX6052;
wire WX3032;
wire WX7051;
wire II34144;
wire II14299;
wire WX5014;
wire WX2883;
wire WX1438;
wire WX5525;
wire II34787;
wire WX925;
wire II18201;
wire II14067;
wire WX7341;
wire WX7461;
wire II14453;
wire WX8873;
wire II22509;
wire WX7891;
wire WX1575;
wire WX3189;
wire WX2196;
wire WX2420;
wire WX9286;
wire WX1460;
wire II30768;
wire WX3822;
wire II10865;
wire II34129;
wire WX10588;
wire II19151;
wire II26017;
wire WX11566;
wire II11631;
wire WX7687;
wire II10122;
wire WX1899;
wire II11679;
wire II22106;
wire II2498;
wire WX2526;
wire WX8927;
wire II23623;
wire WX2053;
wire WX1455;
wire II11153;
wire II15457;
wire WX5372;
wire II22635;
wire II30109;
wire II26885;
wire WX3182;
wire II18782;
wire II3614;
wire WX3053;
wire WX10772;
wire II22507;
wire II6147;
wire II22128;
wire II26918;
wire II30497;
wire WX2888;
wire II15655;
wire II19689;
wire II22743;
wire WX4303;
wire WX10189;
wire WX3340;
wire WX2459;
wire WX5710;
wire II2018;
wire WX9060;
wire WX9021;
wire WX615;
wire II2144;
wire II34120;
wire WX1732;
wire II2492;
wire WX516;
wire WX1466;
wire WX11312;
wire WX4905;
wire WX7523;
wire WX2751;
wire WX1607;
wire II34743;
wire WX9603;
wire II19294;
wire II19696;
wire II30287;
wire II30045;
wire WX3734;
wire WX8364;
wire II14826;
wire II14222;
wire II10239;
wire WX628;
wire WX8837;
wire WX268;
wire II19682;
wire II10315;
wire II30248;
wire II7562;
wire WX8313;
wire WX8793;
wire WX388;
wire II15587;
wire II27699;
wire WX7501;
wire WX153;
wire WX10618;
wire WX7151;
wire II2436;
wire II34975;
wire II30419;
wire WX5271;
wire WX4967;
wire II18093;
wire II34167;
wire WX3030;
wire II2685;
wire WX5407;
wire II34214;
wire WX3659;
wire II30280;
wire WX5451;
wire II2214;
wire WX1581;
wire II18658;
wire WX10418;
wire WX4489;
wire II26259;
wire WX6424;
wire WX9273;
wire II3509;
wire WX3714;
wire WX5524;
wire WX1457;
wire II10587;
wire II2624;
wire WX11256;
wire WX6356;
wire WX10762;
wire WX3825;
wire WX7677;
wire WX2361;
wire II30954;
wire II18743;
wire II35702;
wire II19099;
wire WX6816;
wire II34780;
wire WX6698;
wire WX1560;
wire WX9931;
wire II10936;
wire WX7864;
wire WX7129;
wire II2276;
wire II7109;
wire WX3962;
wire WX7279;
wire WX11600;
wire WX11294;
wire WX241;
wire WX6396;
wire WX6662;
wire WX10168;
wire WX1604;
wire WX456;
wire WX1539;
wire II11545;
wire WX5651;
wire II22176;
wire WX7424;
wire WX5338;
wire II1990;
wire WX10934;
wire WX6335;
wire II30489;
wire WX5072;
wire WX7873;
wire WX5013;
wire II26700;
wire WX5212;
wire WX10080;
wire II15720;
wire WX4838;
wire II26668;
wire WX8488;
wire WX1714;
wire II22314;
wire WX989;
wire II3119;
wire WX8904;
wire II34308;
wire II6543;
wire WX3742;
wire II18171;
wire WX3511;
wire II30170;
wire WX1567;
wire II19570;
wire II18651;
wire WX991;
wire II30831;
wire WX11377;
wire II18208;
wire WX4872;
wire WX11118;
wire II23701;
wire II7475;
wire II22541;
wire II27623;
wire WX2796;
wire WX5622;
wire II30411;
wire II34238;
wire WX1428;
wire WX2715;
wire WX10670;
wire WX11335;
wire WX4739;
wire WX8582;
wire WX1284;
wire WX9897;
wire WX10152;
wire WX5826;
wire WX2914;
wire II18533;
wire II35563;
wire WX7625;
wire WX9102;
wire WX7295;
wire II30490;
wire WX3991;
wire II18186;
wire WX4986;
wire WX3810;
wire WX5604;
wire II15288;
wire II35005;
wire WX10213;
wire WX565;
wire WX11282;
wire II19489;
wire WX8756;
wire WX3064;
wire II22461;
wire WX3080;
wire WX7445;
wire WX1739;
wire WX6561;
wire II2895;
wire WX536;
wire WX9361;
wire WX171;
wire II22431;
wire II14051;
wire WX10558;
wire WX6607;
wire II10951;
wire WX522;
wire WX6136;
wire WX4341;
wire WX1354;
wire WX9949;
wire II19669;
wire II18581;
wire WX6757;
wire II34991;
wire II30435;
wire WX2521;
wire II27368;
wire WX3440;
wire WX5171;
wire WX3848;
wire II26451;
wire WX2125;
wire WX2187;
wire WX3502;
wire II2166;
wire WX2703;
wire II14965;
wire WX3567;
wire II30340;
wire WX10860;
wire WX6838;
wire WX7022;
wire WX9751;
wire II22796;
wire WX8286;
wire II34741;
wire WX11300;
wire WX10551;
wire II14762;
wire II10175;
wire II6219;
wire II27252;
wire WX10200;
wire WX1638;
wire II10217;
wire WX5116;
wire II15211;
wire WX4278;
wire WX10100;
wire II30565;
wire WX10981;
wire II30145;
wire WX1478;
wire WX10063;
wire WX11543;
wire WX177;
wire WX2687;
wire II27304;
wire II2615;
wire II11270;
wire WX4004;
wire II34540;
wire II14351;
wire WX2910;
wire WX6739;
wire WX1631;
wire WX7598;
wire WX2825;
wire II30394;
wire WX10697;
wire II26490;
wire WX2426;
wire II6682;
wire II15067;
wire WX2645;
wire WX922;
wire WX7713;
wire WX3777;
wire WX1776;
wire II11388;
wire WX8728;
wire WX10101;
wire II35577;
wire WX8380;
wire II14855;
wire II27001;
wire WX10840;
wire WX1835;
wire WX3530;
wire WX10000;
wire WX9650;
wire WX11359;
wire II3605;
wire II23510;
wire II34801;
wire WX8056;
wire WX4589;
wire II7577;
wire WX5589;
wire II11414;
wire II31642;
wire II19512;
wire WX5030;
wire II34453;
wire WX3715;
wire WX6313;
wire II26754;
wire WX8342;
wire II3477;
wire II11524;
wire II22508;
wire WX8735;
wire WX570;
wire II14854;
wire WX10537;
wire WX8207;
wire II22804;
wire WX4074;
wire WX896;
wire WX4456;
wire WX10447;
wire II3564;
wire II11714;
wire II14315;
wire WX1042;
wire WX4887;
wire II34950;
wire WX10240;
wire WX4561;
wire WX9129;
wire II14931;
wire II10053;
wire II31232;
wire II22192;
wire WX5542;
wire WX6510;
wire II2762;
wire WX621;
wire WX9675;
wire WX1861;
wire II34291;
wire II34696;
wire II14034;
wire WX7896;
wire WX8223;
wire II14745;
wire II18721;
wire II2493;
wire WX8011;
wire II34346;
wire II35313;
wire II27692;
wire II22216;
wire II18766;
wire WX1237;
wire WX1734;
wire II2250;
wire II2461;
wire WX10286;
wire WX3719;
wire WX10464;
wire WX1917;
wire II14532;
wire II18783;
wire WX8387;
wire II23532;
wire WX9498;
wire WX9413;
wire WX3017;
wire WX6086;
wire WX8337;
wire WX9126;
wire WX4537;
wire WX4693;
wire WX1531;
wire II10958;
wire II34386;
wire II26430;
wire II22655;
wire WX1177;
wire WX8744;
wire WX1620;
wire WX2248;
wire WX10574;
wire II10206;
wire WX1006;
wire WX7015;
wire WX9146;
wire WX10978;
wire II10168;
wire WX11130;
wire WX9514;
wire II19126;
wire WX8576;
wire WX7810;
wire II14174;
wire II10446;
wire WX8508;
wire WX1540;
wire WX10123;
wire WX7801;
wire WX9171;
wire WX2935;
wire WX10431;
wire II34182;
wire II30815;
wire WX5906;
wire WX1448;
wire WX6780;
wire WX10662;
wire II27601;
wire II18636;
wire WX9581;
wire WX6519;
wire II18698;
wire WX11026;
wire WX2722;
wire II30721;
wire WX7980;
wire WX3876;
wire WX9962;
wire II22957;
wire WX4106;
wire WX83;
wire WX8703;
wire WX11582;
wire WX792;
wire WX1007;
wire WX1862;
wire II27316;
wire II31360;
wire WX11271;
wire WX5932;
wire II6349;
wire II22278;
wire II26546;
wire WX413;
wire WX8007;
wire II6598;
wire II34825;
wire II30891;
wire WX2212;
wire II6241;
wire WX3998;
wire II11622;
wire WX210;
wire II22247;
wire II18348;
wire II22531;
wire II18953;
wire WX6625;
wire WX10680;
wire WX10532;
wire WX1695;
wire WX5560;
wire WX5757;
wire II7520;
wire II10090;
wire WX9909;
wire WX2844;
wire II6139;
wire WX4523;
wire WX5808;
wire WX1597;
wire WX7931;
wire WX5355;
wire WX5648;
wire WX8954;
wire WX10799;
wire WX6486;
wire WX10752;
wire WX2267;
wire WX9372;
wire WX10748;
wire II14094;
wire WX9871;
wire II3634;
wire II10709;
wire WX7269;
wire II14228;
wire WX1923;
wire WX4479;
wire WX7830;
wire II30209;
wire WX7575;
wire II30985;
wire WX1549;
wire II22866;
wire II26235;
wire WX1118;
wire II18908;
wire WX4476;
wire WX7080;
wire WX6798;
wire WX3664;
wire WX2867;
wire II10913;
wire WX10515;
wire WX4044;
wire WX7662;
wire II35666;
wire WX8130;
wire WX4543;
wire II6085;
wire WX5644;
wire WX1000;
wire II6263;
wire II10703;
wire II26537;
wire II26350;
wire WX7251;
wire WX7645;
wire WX244;
wire WX10620;
wire WX1689;
wire II30611;
wire WX1498;
wire WX1395;
wire WX6886;
wire WX672;
wire WX10911;
wire WX5978;
wire WX1411;
wire II7701;
wire WX5582;
wire II6488;
wire II22548;
wire WX8372;
wire WX860;
wire WX4223;
wire WX5946;
wire WX10821;
wire WX10486;
wire II10702;
wire WX4385;
wire WX9653;
wire WX7704;
wire II18325;
wire II22686;
wire II35654;
wire II15524;
wire WX10608;
wire WX3258;
wire WX4082;
wire II18309;
wire WX6355;
wire WX1278;
wire WX9994;
wire II31519;
wire II26219;
wire WX9007;
wire WX4957;
wire WX10148;
wire WX5157;
wire II26218;
wire II2971;
wire WX10257;
wire WX2447;
wire II3556;
wire II34175;
wire II14769;
wire II26174;
wire WX10815;
wire WX11408;
wire II2413;
wire WX8414;
wire WX8163;
wire II35681;
wire WX5262;
wire WX10136;
wire WX10585;
wire WX5302;
wire II31166;
wire WX6446;
wire II6940;
wire WX4946;
wire WX418;
wire II27712;
wire II14816;
wire WX5412;
wire II30357;
wire II26204;
wire II27343;
wire II10673;
wire WX2552;
wire II22013;
wire WX4783;
wire WX5480;
wire WX2208;
wire WX10317;
wire II10294;
wire II18619;
wire WX186;
wire WX6844;
wire WX1346;
wire WX10313;
wire WX11658;
wire WX6456;
wire WX4647;
wire WX10478;
wire WX9353;
wire WX3900;
wire II19217;
wire WX6876;
wire WX5554;
wire II26421;
wire II22022;
wire II14129;
wire WX9298;
wire II31550;
wire WX3157;
wire II18046;
wire II6730;
wire WX2452;
wire II10430;
wire WX6213;
wire WX7040;
wire II27395;
wire WX5002;
wire WX996;
wire II23688;
wire WX9249;
wire II23168;
wire II22145;
wire II31506;
wire II34918;
wire WX3184;
wire WX9334;
wire WX2810;
wire II31719;
wire II14940;
wire WX7187;
wire II6178;
wire WX4499;
wire II3430;
wire II6706;
wire WX9336;
wire II10154;
wire II30736;
wire II31466;
wire II34594;
wire II22821;
wire WX10731;
wire WX1893;
wire WX579;
wire WX2422;
wire WX5136;
wire WX4055;
wire II18010;
wire WX7433;
wire WX8996;
wire II7200;
wire WX5163;
wire WX4417;
wire WX8193;
wire WX7559;
wire II10207;
wire WX4505;
wire II11574;
wire WX6376;
wire II18258;
wire II18752;
wire II18814;
wire WX2435;
wire II2205;
wire II18513;
wire WX1756;
wire II35392;
wire WX2514;
wire II31178;
wire WX5149;
wire WX7584;
wire WX4508;
wire II18172;
wire II14583;
wire WX206;
wire WX7618;
wire II3535;
wire WX51;
wire II10563;
wire WX4775;
wire WX1727;
wire II10076;
wire WX11426;
wire WX2957;
wire WX9229;
wire II2886;
wire WX11642;
wire WX386;
wire WX9473;
wire WX3977;
wire WX8813;
wire WX1720;
wire WX8448;
wire WX5505;
wire WX2286;
wire II6651;
wire II19333;
wire WX10197;
wire WX6339;
wire WX8774;
wire WX9627;
wire II2631;
wire II7460;
wire WX10658;
wire WX2847;
wire WX3388;
wire WX4866;
wire II19282;
wire WX11146;
wire II7542;
wire WX4729;
wire II26144;
wire II14949;
wire WX8697;
wire WX9464;
wire WX11636;
wire WX1485;
wire WX10923;
wire II10658;
wire II23313;
wire WX1071;
wire II2213;
wire II34267;
wire II14439;
wire WX945;
wire II26081;
wire II6894;
wire WX8272;
wire WX1214;
wire II7717;
wire II18877;
wire WX9184;
wire II18713;
wire WX8422;
wire II26289;
wire II18006;
wire II15251;
wire II6064;
wire II31682;
wire WX8832;
wire II14087;
wire II14144;
wire II2090;
wire WX6848;
wire II26205;
wire II18457;
wire II31585;
wire II35715;
wire WX518;
wire WX7839;
wire WX9405;
wire II27551;
wire II26622;
wire WX7018;
wire WX1216;
wire WX2650;
wire II26848;
wire WX7867;
wire WX3280;
wire II6118;
wire II10725;
wire II2949;
wire WX8604;
wire II34616;
wire WX9191;
wire WX10297;
wire WX10453;
wire WX8034;
wire II22819;
wire WX148;
wire II26980;
wire II2909;
wire II10439;
wire II34284;
wire WX5605;
wire WX2678;
wire WX6408;
wire WX8789;
wire II19491;
wire WX9165;
wire WX133;
wire WX6547;
wire II34926;
wire WX7846;
wire WX4361;
wire WX3801;
wire WX9290;
wire WX10956;
wire II10301;
wire WX5599;
wire WX305;
wire WX6097;
wire II31334;
wire WX3554;
wire WX6700;
wire WX668;
wire II15381;
wire II34872;
wire WX8153;
wire WX7430;
wire WX7479;
wire II6628;
wire WX9237;
wire WX5591;
wire WX11328;
wire WX8838;
wire WX1445;
wire WX774;
wire WX5510;
wire II7660;
wire WX9823;
wire WX11068;
wire WX7025;
wire II22059;
wire WX11389;
wire WX451;
wire II7484;
wire II26615;
wire WX3524;
wire WX9561;
wire II26553;
wire WX429;
wire II27558;
wire WX4393;
wire WX2326;
wire WX5193;
wire II10015;
wire II14304;
wire WX11090;
wire WX445;
wire II22602;
wire WX6310;
wire WX10706;
wire II23442;
wire II11349;
wire WX8119;
wire II3663;
wire II30301;
wire WX10594;
wire WX8106;
wire II10120;
wire WX2971;
wire WX8944;
wire WX146;
wire WX6145;
wire II7163;
wire WX583;
wire WX10502;
wire WX6904;
wire II31740;
wire II35419;
wire WX712;
wire II26288;
wire II18047;
wire WX880;
wire WX5325;
wire WX8177;
wire II22625;
wire II34305;
wire WX836;
wire WX9661;
wire II22043;
wire WX7241;
wire II22983;
wire WX191;
wire WX4470;
wire WX10494;
wire II22213;
wire WX8158;
wire II6148;
wire WX982;
wire II7278;
wire WX740;
wire WX1450;
wire WX8846;
wire WX5500;
wire WX10787;
wire II30590;
wire II27546;
wire II26469;
wire II18068;
wire II11700;
wire WX3702;
wire WX9421;
wire WX10703;
wire WX2283;
wire II23339;
wire WX9545;
wire WX1085;
wire II34608;
wire WX882;
wire II7505;
wire WX7854;
wire WX3320;
wire II11503;
wire II27707;
wire II6095;
wire WX7193;
wire II10525;
wire WX9453;
wire WX9150;
wire WX7398;
wire II26064;
wire II6425;
wire WX10627;
wire WX7561;
wire II2227;
wire WX7545;
wire WX10874;
wire WX9218;
wire WX9087;
wire WX9515;
wire WX2501;
wire II15160;
wire WX1880;
wire WX8667;
wire II22563;
wire II14074;
wire WX3014;
wire WX4879;
wire II2593;
wire WX7696;
wire WX3509;
wire II19424;
wire WX2254;
wire WX7137;
wire WX5590;
wire II22430;
wire II19398;
wire WX9668;
wire II10572;
wire WX7904;
wire II18078;
wire WX325;
wire WX6558;
wire II26931;
wire II26048;
wire WX3847;
wire WX5005;
wire WX9681;
wire WX9304;
wire WX7548;
wire WX341;
wire WX7915;
wire WX7179;
wire WX9489;
wire II18688;
wire WX11386;
wire WX5295;
wire WX11584;
wire WX6205;
wire WX1750;
wire II3223;
wire WX6575;
wire II30512;
wire WX1584;
wire II14841;
wire WX442;
wire WX4401;
wire WX8074;
wire WX11297;
wire II34585;
wire WX4512;
wire WX6265;
wire WX11182;
wire II10198;
wire WX10235;
wire WX10053;
wire II14330;
wire WX10542;
wire II22727;
wire II14469;
wire WX872;
wire II34701;
wire II5991;
wire WX3147;
wire WX11465;
wire II7110;
wire WX10572;
wire WX10111;
wire WX4892;
wire II30690;
wire II26444;
wire WX636;
wire II6884;
wire WX1875;
wire WX9534;
wire WX2680;
wire WX7213;
wire II22852;
wire WX4657;
wire WX2805;
wire II2668;
wire II22555;
wire WX8550;
wire WX5009;
wire WX6300;
wire WX6783;
wire WX8006;
wire WX1196;
wire WX9506;
wire WX6647;
wire II31649;
wire II18133;
wire WX6694;
wire WX9368;
wire WX4190;
wire II11181;
wire II27135;
wire II2238;
wire II18256;
wire WX1799;
wire WX7458;
wire WX3070;
wire WX9391;
wire WX4130;
wire II26475;
wire II35250;
wire II6869;
wire WX7353;
wire WX5102;
wire WX8128;
wire WX3021;
wire WX11490;
wire II26109;
wire II14428;
wire II6832;
wire II10069;
wire WX9573;
wire WX2007;
wire WX1615;
wire II34857;
wire WX11340;
wire WX2855;
wire WX261;
wire II26343;
wire WX10303;
wire WX7063;
wire WX3055;
wire II14731;
wire II18790;
wire II3442;
wire WX1027;
wire WX10195;
wire II18947;
wire II15713;
wire II30645;
wire WX6024;
wire WX4798;
wire WX402;
wire WX8211;
wire WX4244;
wire WX520;
wire WX6717;
wire WX8235;
wire WX11248;
wire WX11344;
wire WX1555;
wire WX8348;
wire WX3370;
wire WX8690;
wire WX5818;
wire II2539;
wire II31698;
wire WX3835;
wire II26709;
wire WX5724;
wire II2004;
wire II26422;
wire II11539;
wire WX10016;
wire II30944;
wire WX10721;
wire WX8308;
wire WX593;
wire WX10689;
wire WX10417;
wire WX7944;
wire WX2920;
wire WX4791;
wire WX5814;
wire WX7029;
wire WX6367;
wire WX3557;
wire WX916;
wire WX9693;
wire WX4155;
wire II27408;
wire WX6186;
wire WX11268;
wire II23665;
wire II11533;
wire WX6162;
wire II14749;
wire WX4279;
wire WX8612;
wire WX7623;
wire II34570;
wire II11721;
wire II10246;
wire WX6597;
wire WX2301;
wire WX3484;
wire WX8504;
wire WX5735;
wire II10554;
wire II2778;
wire II18885;
wire WX7005;
wire WX6747;
wire WX8961;
wire II22061;
wire WX2640;
wire WX6120;
wire II14980;
wire II10942;
wire II6381;
wire WX3040;
wire II11088;
wire WX625;
wire WX1336;
wire WX6073;
wire WX8822;
wire II10339;
wire WX5471;
wire II7059;
wire II7070;
wire II14593;
wire WX9011;
wire WX4052;
wire II14676;
wire II26902;
wire WX10522;
wire WX3229;
wire WX2963;
wire II22848;
wire WX600;
wire WX9665;
wire II2128;
wire WX5660;
wire WX538;
wire WX6241;
wire WX8278;
wire II2134;
wire II27160;
wire WX4352;
wire WX3452;
wire WX5318;
wire WX10275;
wire II14801;
wire II34045;
wire II26761;
wire WX8913;
wire II1996;
wire II30862;
wire WX4175;
wire II34532;
wire WX2711;
wire WX6320;
wire II30331;
wire WX6386;
wire II34461;
wire WX5508;
wire II2392;
wire WX11396;
wire II7305;
wire WX5142;
wire II34842;
wire II34554;
wire WX6416;
wire WX6090;
wire WX11321;
wire WX3683;
wire WX4009;
wire WX3985;
wire II15572;
wire WX5950;
wire WX7685;
wire II11376;
wire WX5367;
wire WX7985;
wire II34228;
wire WX2057;
wire II7434;
wire WX9745;
wire WX8986;
wire WX2903;
wire II35495;
wire II26815;
wire WX4803;
wire WX6269;
wire II30147;
wire WX4951;
wire WX198;
wire II34569;
wire WX4583;
wire WX6710;
wire II34392;
wire WX5494;
wire II7448;
wire II22223;
wire WX4447;
wire WX2259;
wire II6667;
wire WX7169;
wire WX9982;
wire II14221;
wire WX2991;
wire WX9038;
wire WX3546;
wire WX4167;
wire II6305;
wire II2803;
wire WX5341;
wire WX5287;
wire II6768;
wire WX11367;
wire WX6506;
wire WX7512;
wire WX11638;
wire II26715;
wire WX10028;
wire II3640;
wire II15571;
wire II10881;
wire WX8766;
wire II6227;
wire WX9529;
wire II26793;
wire II11489;
wire II30093;
wire II10728;
wire II14361;
wire WX2694;
wire II3314;
wire II35568;
wire II22516;
wire WX903;
wire WX6635;
wire WX1523;
wire WX7635;
wire WX3300;
wire WX5048;
wire WX3056;
wire II30241;
wire WX4330;
wire WX3414;
wire WX5282;
wire WX8977;
wire WX7885;
wire II15600;
wire II6549;
wire WX552;
wire II14947;
wire II15277;
wire II27531;
wire II30920;
wire WX5346;
wire II22115;
wire II14661;
wire II3613;
wire WX9911;
wire WX2727;
wire WX5029;
wire WX5694;
wire II2818;
wire II22525;
wire II15662;
wire II22324;
wire WX10613;
wire II18543;
wire WX5408;
wire WX103;
wire WX11056;
wire WX122;
wire II6737;
wire II30054;
wire II26784;
wire WX6726;
wire WX9076;
wire II2454;
wire WX8327;
wire WX820;
wire WX943;
wire WX9259;
wire II15726;
wire II10145;
wire II30581;
wire II22399;
wire WX1361;
wire WX3790;
wire II11519;
wire WX2316;
wire WX956;
wire WX6273;
wire II11580;
wire II2795;
wire WX3792;
wire II22478;
wire WX1590;
wire WX10043;
wire WX8266;
wire WX2079;
wire II34849;
wire WX2809;
wire II18381;
wire WX6395;
wire WX4144;
wire II2424;
wire WX1087;
wire WX10128;
wire WX11220;
wire II30968;
wire WX7905;
wire WX9887;
wire WX6552;
wire WX5980;
wire II26234;
wire WX10109;
wire II15107;
wire WX6855;
wire II23560;
wire WX3072;
wire WX10384;
wire II3080;
wire II22401;
wire WX10826;
wire II26041;
wire II22394;
wire II6188;
wire II19072;
wire II6459;
wire WX11533;
wire WX4357;
wire II6790;
wire WX4625;
wire II6698;
wire WX6151;
wire WX4081;
wire WX10407;
wire WX8374;
wire WX8476;
wire WX7517;
wire II19641;
wire WX11469;
wire WX8320;
wire WX1493;
wire WX10444;
wire II6211;
wire II7680;
wire II19410;
wire II10835;
wire WX1381;
wire WX818;
wire II27629;
wire WX10175;
wire II34378;
wire WX1416;
wire WX2982;
wire II14080;
wire WX4685;
wire II18435;
wire II27279;
wire WX10953;
wire WX7571;
wire II22337;
wire WX4639;
wire II34371;
wire II30626;
wire II2475;
wire II14265;
wire WX9410;
wire WX5998;
wire WX4935;
wire WX7044;
wire WX6419;
wire WX11124;
wire WX4115;
wire WX8023;
wire II10493;
wire II15627;
wire WX1845;
wire WX8807;
wire WX10792;
wire WX6579;
wire WX5360;
wire WX11076;
wire II35118;
wire II7556;
wire II31140;
wire WX5830;
wire WX10736;
wire WX11264;
wire WX4021;
wire II11298;
wire WX2833;
wire II10602;
wire II10983;
wire WX5795;
wire WX3110;
wire II27188;
wire WX10795;
wire II11402;
wire II35527;
wire WX2541;
wire II15657;
wire WX2356;
wire II23272;
wire WX6195;
wire WX11616;
wire II7611;
wire WX8542;
wire II35210;
wire II30807;
wire WX9324;
wire WX4311;
wire II6924;
wire WX7387;
wire II34161;
wire II34479;
wire II19176;
wire WX4295;
wire WX8046;
wire II30472;
wire WX4326;
wire II22353;
wire WX8049;
wire WX5988;
wire WX4218;
wire WX7821;
wire WX2710;
wire WX6631;
wire II2296;
wire WX6040;
wire II10425;
wire WX11578;
wire II34757;
wire WX4910;
wire II30821;
wire II18350;
wire WX7920;
wire II34067;
wire WX8292;
wire II30397;
wire WX934;
wire WX1034;
wire II31697;
wire WX10252;
wire WX1357;
wire II18637;
wire WX3806;
wire II34470;
wire II2283;
wire WX1240;
wire II30800;
wire II31731;
wire WX10095;
wire WX8452;
wire II6033;
wire WX4061;
wire WX43;
wire WX11514;
wire WX9433;
wire WX1179;
wire WX1612;
wire WX1372;
wire II19612;
wire WX7655;
wire WX3539;
wire II7098;
wire II19732;
wire II14714;
wire WX9289;
wire WX11576;
wire II14405;
wire WX6925;
wire II22928;
wire WX1122;
wire WX5041;
wire WX390;
wire WX3527;
wire WX1420;
wire WX1516;
wire II6668;
wire WX6595;
wire WX11413;
wire II11129;
wire II2067;
wire II18154;
wire II34773;
wire WX5579;
wire II30164;
wire WX9615;
wire WX9522;
wire WX7721;
wire WX10339;
wire II19619;
wire WX7197;
wire II18177;
wire WX7413;
wire II3584;
wire II23221;
wire WX3209;
wire WX11285;
wire WX5595;
wire II14020;
wire WX3520;
wire II2189;
wire II22030;
wire WX3916;
wire II15530;
wire WX10629;
wire WX7955;
wire WX392;
wire II30318;
wire WX9446;
wire WX2091;
wire WX9969;
wire II2188;
wire WX6254;
wire WX3593;
wire WX8460;
wire WX4265;
wire II26824;
wire WX8896;
wire WX4856;
wire WX8084;
wire II14787;
wire WX5311;
wire II14622;
wire WX1013;
wire WX6529;
wire WX1789;
wire WX4283;
wire WX10667;
wire II35092;
wire II10758;
wire II27420;
wire WX1701;
wire WX1623;
wire WX10203;
wire WX6679;
wire II2483;
wire WX5741;
wire II2111;
wire WX1993;
wire WX7796;
wire WX2384;
wire II15691;
wire WX11444;
wire II26267;
wire WX9177;
wire WX8870;
wire WX9472;
wire WX8958;
wire II22229;
wire WX11170;
wire WX8949;
wire WX8712;
wire II34089;
wire II23589;
wire II26197;
wire WX9199;
wire WX8815;
wire WX361;
wire WX11522;
wire II22990;
wire WX6185;
wire WX4514;
wire WX11088;
wire II15599;
wire WX11519;
wire II7330;
wire WX8378;
wire WX10357;
wire II2384;
wire II11644;
wire II2600;
wire WX7233;
wire WX8680;
wire II14368;
wire II14831;
wire II11258;
wire WX7037;
wire WX1645;
wire WX7537;
wire WX2143;
wire WX3602;
wire WX7030;
wire WX1225;
wire WX1571;
wire WX2864;
wire II10806;
wire WX5792;
wire WX2726;
wire II14554;
wire WX6236;
wire WX11527;
wire II18521;
wire II27225;
wire WX2791;
wire II10966;
wire II22183;
wire WX4763;
wire WX3234;
wire WX1055;
wire II23595;
wire II30743;
wire WX6889;
wire II10976;
wire WX6681;
wire WX8717;
wire WX1648;
wire II22309;
wire II23324;
wire II10410;
wire WX8616;
wire WX2464;
wire WX422;
wire WX280;
wire WX5244;
wire WX66;
wire WX7816;
wire II14639;
wire WX7405;
wire II18977;
wire WX2327;
wire WX4258;
wire II10975;
wire II34732;
wire II18397;
wire WX7530;
wire WX2544;
wire WX11353;
wire II23525;
wire WX2398;
wire II14002;
wire WX7011;
wire WX136;
wire WX2743;
wire WX4484;
wire WX6674;
wire WX8753;
wire WX3408;
wire II6232;
wire WX2780;
wire II27461;
wire WX5167;
wire WX9183;
wire WX11253;
wire II31479;
wire II30535;
wire WX9630;
wire WX4097;
wire WX7889;
wire II11077;
wire WX1202;
wire II30905;
wire II18923;
wire WX2535;
wire II10462;
wire WX1188;
wire II34835;
wire WX8242;
wire WX8144;
wire WX5803;
wire II35146;
wire II23116;
wire II2444;
wire II10888;
wire WX8393;
wire II14926;
wire II3379;
wire II30332;
wire WX8496;
wire WX1252;
wire II27486;
wire WX38;
wire WX7753;
wire WX5533;
wire WX7850;
wire II26926;
wire WX9462;
wire II22976;
wire WX2975;
wire II26575;
wire II18193;
wire II18371;
wire WX236;
wire II26298;
wire WX4120;
wire WX5753;
wire II19229;
wire II35274;
wire II14645;
wire WX4809;
wire II7640;
wire II3248;
wire WX5275;
wire WX5422;
wire II35675;
wire II14780;
wire WX5536;
wire II15445;
wire WX10458;
wire II34726;
wire WX11428;
wire WX6777;
wire WX8672;
wire WX7769;
wire II30115;
wire WX8885;
wire II26872;
wire WX9080;
wire WX1230;
wire WX1386;
wire WX3752;
wire WX6429;
wire WX8112;
wire II10697;
wire WX1933;
wire II11511;
wire II11602;
wire II19675;
wire WX11435;
wire WX5926;
wire II26328;
wire WX10411;
wire II10851;
wire II3221;
wire II23632;
wire II22511;
wire II30380;
wire II30180;
wire WX7141;
wire WX205;
wire II22263;
wire II30021;
wire WX1504;
wire WX10229;
wire WX2418;
wire WX5394;
wire WX5183;
wire WX842;
wire WX4334;
wire WX9216;
wire WX9240;
wire WX3641;
wire WX9206;
wire II30311;
wire WX7527;
wire WX762;
wire WX4824;
wire WX9363;
wire WX8404;
wire WX11240;
wire WX76;
wire II6956;
wire WX1854;
wire II23519;
wire II23428;
wire WX1049;
wire II30550;
wire WX5586;
wire II2916;
wire WX6440;
wire WX4671;
wire WX9610;
wire WX11480;
wire WX289;
wire WX7247;
wire II10386;
wire WX371;
wire WX2376;
wire WX8212;
wire WX11561;
wire WX10603;
wire WX10640;
wire II23480;
wire WX7968;
wire II11629;
wire WX9264;
wire II6752;
wire WX10563;
wire WX3368;
wire II35249;
wire WX9137;
wire WX5209;
wire WX11491;
wire WX3264;
wire WX3161;
wire WX10806;
wire WX4794;
wire II14384;
wire WX9555;
wire II35405;
wire II7409;
wire II27508;
wire II14421;
wire WX4469;
wire WX8862;
wire WX1765;
wire WX6146;
wire WX7993;
wire II6689;
wire WX2291;
wire II26102;
wire WX2232;
wire II10618;
wire WX9028;
wire WX9989;
wire WX4059;
wire WX5678;
wire WX8562;
wire WX9481;
wire WX7106;
wire WX2131;
wire WX3854;
wire WX2738;
wire WX6765;
wire WX8677;
wire WX4015;
wire WX4991;
wire II6403;
wire WX6103;
wire WX3954;
wire WX10178;
wire WX963;
wire WX7923;
wire II34866;
wire II6828;
wire II34059;
wire WX9178;
wire WX1846;
wire WX7608;
wire II2052;
wire II22609;
wire WX1989;
wire WX8660;
wire II18378;
wire II7612;
wire WX6127;
wire WX11622;
wire WX10159;
wire WX8010;
wire II30239;
wire II26407;
wire WX9597;
wire WX8850;
wire II2880;
wire WX6111;
wire WX1669;
wire WX4926;
wire WX8060;
wire WX4315;
wire II26598;
wire II15199;
wire WX433;
wire WX10423;
wire WX4345;
wire WX116;
wire WX3585;
wire WX2785;
wire WX10232;
wire WX1945;
wire WX263;
wire WX4619;
wire WX10649;
wire WX6524;
wire WX9917;
wire II22136;
wire WX9428;
wire WX2430;
wire II6312;
wire WX6852;
wire WX467;
wire II23503;
wire II7174;
wire WX5419;
wire WX9256;
wire WX11275;
wire WX4813;
wire II15507;
wire WX1787;
wire WX3298;
wire WX4209;
wire WX6688;
wire II14514;
wire WX3039;
wire II10277;
wire WX9239;
wire WX7773;
wire WX5763;
wire WX8202;
wire WX4202;
wire WX5123;
wire WX6939;
wire WX2947;
wire WX4029;
wire II2785;
wire II10325;
wire II34402;
wire II26684;
wire WX2484;
wire II7491;
wire WX1067;
wire WX3098;
wire II35107;
wire WX5902;
wire WX5109;
wire II22959;
wire II26996;
wire WX5462;
wire II23693;
wire WX2932;
wire II34577;
wire WX2821;
wire WX5265;
wire WX5333;
wire WX2629;
wire WX10074;
wire WX2659;
wire WX10127;
wire II30906;
wire WX7709;
wire WX257;
wire II34688;
wire WX10298;
wire WX10469;
wire II30099;
wire WX4845;
wire WX6226;
wire WX7103;
wire II11218;
wire WX5093;
wire WX10321;
wire WX1896;
wire WX1415;
wire WX7437;
wire II2268;
wire WX584;
wire II7382;
wire WX6244;
wire WX1692;
wire WX7961;
wire II3712;
wire II31219;
wire II10463;
wire II35196;
wire WX2222;
wire WX2665;
wire WX6624;
wire WX6941;
wire WX6542;
wire WX9635;
wire WX11204;
wire WX2159;
wire WX6736;
wire WX2411;
wire WX8096;
wire WX8418;
wire WX3764;
wire WX6616;
wire WX1320;
wire WX1424;
wire II2610;
wire WX6975;
wire WX2275;
wire WX6822;
wire II26460;
wire WX6948;
wire WX6174;
wire WX7428;
wire II10286;
wire WX10398;
wire WX6539;
wire WX5578;
wire WX2894;
wire WX6521;
wire II6552;
wire WX11399;
wire WX658;
wire WX4867;
wire II18558;
wire II11509;
wire II34763;
wire WX10856;
wire II26777;
wire WX3316;
wire II2073;
wire II6605;
wire II30459;
wire II35556;
wire WX3866;
wire WX3623;
wire WX1519;
wire II14151;
wire WX473;
wire WX9122;
wire WX8941;
wire WX4886;
wire WX6270;
wire WX4697;
wire WX6735;
wire WX5545;
wire WX4180;
wire II2507;
wire II22728;
wire WX587;
wire II14685;
wire WX10244;
wire WX3458;
wire WX5868;
wire WX3550;
wire II3668;
wire II31669;
wire II34407;
wire WX10730;
wire WX5575;
wire WX10974;
wire WX574;
wire II22449;
wire II23553;
wire II30652;
wire II6807;
wire WX2638;
wire WX4425;
wire II34099;
wire WX8622;
wire WX1686;
wire WX5640;
wire WX6336;
wire WX8654;
wire WX6513;
wire WX5401;
wire WX1440;
wire WX10489;
wire WX10901;
wire WX8869;
wire II14668;
wire II22028;
wire WX11470;
wire II27330;
wire WX4068;
wire II26770;
wire WX2832;
wire WX2321;
wire II27656;
wire WX6258;
wire WX8332;
wire WX6870;
wire WX7806;
wire WX10720;
wire WX6199;
wire WX10578;
wire II35743;
wire WX498;
wire WX6750;
wire WX11422;
wire WX1997;
wire WX6853;
wire WX7485;
wire WX6002;
wire II14242;
wire WX4124;
wire WX10534;
wire II11232;
wire II26381;
wire WX4565;
wire WX9319;
wire II2847;
wire WX10007;
wire WX5039;
wire WX7558;
wire II7673;
wire WX8346;
wire II3169;
wire II15327;
wire WX1677;
wire II3528;
wire WX8686;
wire WX5035;
wire II14934;
wire II35300;
wire WX4113;
wire WX6389;
wire WX10460;
wire II31165;
wire WX5609;
wire II26723;
wire WX9494;
wire WX4093;
wire WX302;
wire WX1793;
wire WX3973;
wire II27574;
wire II14476;
wire WX7466;
wire II22245;
wire II14010;
wire WX3925;
wire WX11317;
wire II30271;
wire WX6082;
wire WX5566;
wire WX957;
wire WX10104;
wire II18473;
wire II3301;
wire II18707;
wire II34832;
wire WX6089;
wire WX5610;
wire WX10283;
wire WX5063;
wire II19320;
wire WX2263;
wire WX10023;
wire WX2073;
wire II10232;
wire WX1080;
wire WX1831;
wire II6419;
wire II31690;
wire WX7859;
wire WX11160;
wire II18760;
wire WX10003;
wire WX1172;
wire II6714;
wire WX4269;
wire II22377;
wire WX6156;
wire WX7834;
wire WX2268;
wire WX9865;
wire WX5077;
wire WX5779;
wire WX8384;
wire WX11494;
wire II6692;
wire II34671;
wire II26552;
wire WX4143;
wire WX10306;
wire WX10401;
wire WX4547;
wire WX619;
wire WX9966;
wire WX3153;
wire WX1262;
wire II35287;
wire II26847;
wire WX11370;
wire WX11158;
wire WX4381;
wire WX5749;
wire WX1113;
wire II31271;
wire II14902;
wire II18116;
wire II31675;
wire II6248;
wire WX8017;
wire II10952;
wire II6504;
wire WX9125;
wire WX6640;
wire WX1473;
wire WX369;
wire WX1210;
wire WX9003;
wire II2336;
wire II6947;
wire WX2573;
wire II14460;
wire WX7506;
wire II2174;
wire II10261;
wire II14521;
wire WX9679;
wire II30596;
wire WX7641;
wire WX9685;
wire WX9143;
wire WX6480;
wire II14204;
wire II14653;
wire II34092;
wire WX5059;
wire WX9458;
wire WX4103;
wire WX9503;
wire II3143;
wire WX10693;
wire II23673;
wire WX7870;
wire II7265;
wire WX1866;
wire WX2517;
wire II2554;
wire II18382;
wire WX3906;
wire WX1583;
wire II7659;
wire WX1927;
wire II15671;
wire WX3533;
wire II6079;
wire WX4247;
wire II22734;
wire II3683;
wire WX5942;
wire WX2559;
wire WX7265;
wire II11480;
wire II31388;
wire WX4817;
wire II34904;
wire WX5390;
wire WX7331;
wire WX3114;
wire WX10665;
wire WX1097;
wire II2035;
wire WX9658;
wire WX4371;
wire WX700;
wire WX4859;
wire II14119;
wire WX3783;
wire II35445;
wire WX10291;
wire II27382;
wire II6410;
wire WX11080;
wire WX8819;
wire II27148;
wire II3542;
wire II18242;
wire II14098;
wire WX10482;
wire II6814;
wire WX10185;
wire WX4307;
wire WX5563;
wire II30728;
wire II6519;
wire II14135;
wire WX9106;
wire II6745;
wire II26485;
wire WX10904;
wire WX976;
wire WX4048;
wire WX5558;
wire WX10942;
wire II2747;
wire II26939;
wire WX8632;
wire WX8926;
wire WX2285;
wire WX6663;
wire II6451;
wire WX3143;
wire WX8367;
wire II19150;
wire WX633;
wire II7547;
wire II34143;
wire II34043;
wire WX2406;
wire WX8594;
wire WX2037;
wire II31600;
wire II14296;
wire WX9064;
wire WX7516;
wire WX11212;
wire WX270;
wire WX3858;
wire WX10715;
wire II11547;
wire WX8827;
wire II7085;
wire WX6910;
wire WX2438;
wire WX4802;
wire II3236;
wire II27537;
wire II31101;
wire II34323;
wire II6537;
wire WX11291;
wire WX2884;
wire WX5442;
wire II34531;
wire WX6064;
wire WX7520;
wire II22448;
wire WX3573;
wire WX4981;
wire WX9364;
wire WX7131;
wire WX5896;
wire WX562;
wire WX5956;
wire WX11565;
wire WX5380;
wire II34037;
wire WX7372;
wire II31269;
wire II10927;
wire WX2569;
wire WX9442;
wire WX9526;
wire II10247;
wire WX1463;
wire WX3515;
wire WX906;
wire II34060;
wire WX5520;
wire WX10527;
wire II26614;
wire II26226;
wire II11566;
wire WX9648;
wire WX4963;
wire WX7303;
wire II22283;
wire II10346;
wire WX9935;
wire WX7028;
wire WX7826;
wire WX6420;
wire II10338;
wire WX10512;
wire II19723;
wire WX1107;
wire WX6919;
wire WX9905;
wire WX5870;
wire II11428;
wire WX7633;
wire II6356;
wire II31139;
wire WX1751;
wire WX172;
wire WX5356;
wire II26111;
wire WX6666;
wire WX4051;
wire II34625;
wire WX10164;
wire II10106;
wire WX9641;
wire WX3984;
wire WX5438;
wire WX6704;
wire WX11339;
wire WX3493;
wire II11348;
wire WX11608;
wire WX5787;
wire WX9485;
wire WX2340;
wire WX8908;
wire II6782;
wire WX9771;
wire WX7155;
wire II22703;
wire II26050;
wire II7162;
wire II10254;
wire WX3134;
wire WX9098;
wire WX5822;
wire WX1710;
wire II30931;
wire II26443;
wire II14709;
wire WX10047;
wire II14344;
wire WX2778;
wire II15264;
wire II6087;
wire WX923;
wire WX10580;
wire WX2649;
wire II6635;
wire WX7291;
wire WX5728;
wire WX5017;
wire WX2683;
wire II23721;
wire II27678;
wire WX6603;
wire II27567;
wire II6397;
wire II26453;
wire WX7081;
wire WX228;
wire WX11008;
wire WX9945;
wire II34028;
wire WX1135;
wire WX10556;
wire II26645;
wire II6976;
wire II14444;
wire II27595;
wire II6676;
wire WX1535;
wire WX4274;
wire WX7281;
wire II34703;
wire WX11070;
wire WX7549;
wire WX4197;
wire II7253;
wire II34996;
wire WX2518;
wire WX7937;
wire WX2997;
wire WX3060;
wire II10479;
wire WX2525;
wire WX804;
wire WX1772;
wire WX4008;
wire WX7068;
wire II23298;
wire II7201;
wire WX8334;
wire WX10067;
wire WX1197;
wire WX4300;
wire WX6331;
wire WX7555;
wire WX4627;
wire WX9607;
wire WX8318;
wire II2548;
wire WX8586;
wire II2725;
wire WX5778;
wire II22293;
wire II14482;
wire II27642;
wire WX542;
wire WX7059;
wire II10216;
wire II3598;
wire II26839;
wire II30504;
wire WX3838;
wire WX10810;
wire II11168;
wire II19618;
wire WX11452;
wire II14360;
wire II18302;
wire WX9377;
wire WX11354;
wire WX5655;
wire II27084;
wire WX10204;
wire II6520;
wire WX11567;
wire II26428;
wire WX11331;
wire WX7449;
wire II27435;
wire II31089;
wire WX10345;
wire WX5627;
wire II18946;
wire WX10560;
wire WX11461;
wire WX940;
wire WX5313;
wire II3647;
wire WX5153;
wire II22867;
wire II26057;
wire WX3892;
wire WX3814;
wire WX3844;
wire WX3444;
wire II11637;
wire WX2706;
wire II19590;
wire WX1717;
wire WX107;
wire II10176;
wire WX4293;
wire II2110;
wire II31152;
wire WX9224;
wire II3391;
wire WX6565;
wire II23541;
wire WX9761;
wire II35339;
wire II22494;
wire WX11383;
wire WX4188;
wire WX5633;
wire WX7217;
wire WX10545;
wire WX11456;
wire II22724;
wire WX6116;
wire WX1350;
wire WX8732;
wire II10400;
wire WX8951;
wire WX4238;
wire II18086;
wire II2940;
wire II14374;
wire II26264;
wire WX8157;
wire WX8357;
wire II31180;
wire WX5486;
wire WX3198;
wire II18621;
wire WX4397;
wire WX2023;
wire II23417;
wire WX6544;
wire II11389;
wire II7514;
wire WX11560;
wire WX9409;
wire II7668;
wire II14235;
wire II22757;
wire WX7899;
wire WX6778;
wire II6877;
wire II14561;
wire II30256;
wire II34259;
wire II6890;
wire II10620;
wire II18612;
wire WX9620;
wire WX1715;
wire II19535;
wire II14778;
wire II6287;
wire II30697;
wire WX9384;
wire II34309;
wire WX8071;
wire WX10034;
wire II6551;
wire WX6882;
wire II2080;
wire WX1259;
wire WX8102;
wire II10533;
wire WX9359;
wire II14546;
wire WX9233;
wire WX4605;
wire WX7718;
wire WX8775;
wire II14249;
wire II3669;
wire II19307;
wire WX8316;
wire WX1128;
wire WX1672;
wire II34912;
wire WX195;
wire WX9827;
wire WX788;
wire WX10674;
wire WX949;
wire WX2337;
wire WX2425;
wire WX3505;
wire WX10393;
wire WX770;
wire WX8842;
wire WX9530;
wire WX8217;
wire WX128;
wire II26863;
wire WX2242;
wire WX8486;
wire II30999;
wire WX8201;
wire II15471;
wire WX4908;
wire WX8037;
wire II6837;
wire II30124;
wire WX441;
wire WX9308;
wire WX5888;
wire WX3106;
wire WX7672;
wire WX10115;
wire WX10438;
wire WX5099;
wire WX1884;
wire II18620;
wire WX8078;
wire WX2003;
wire II23078;
wire WX2513;
wire WX8834;
wire WX5298;
wire WX1233;
wire WX11324;
wire II10012;
wire II31619;
wire II30138;
wire WX6908;
wire II18225;
wire WX8683;
wire WX6532;
wire WX9375;
wire WX10289;
wire WX2244;
wire WX8888;
wire WX11186;
wire WX4725;
wire WX169;
wire II30084;
wire WX3970;
wire WX11208;
wire II6475;
wire WX8663;
wire II14118;
wire WX9729;
wire WX2989;
wire II22486;
wire WX11447;
wire WX6587;
wire WX9303;
wire WX5583;
wire II2578;
wire WX11261;
wire II30774;
wire WX3018;
wire WX4087;
wire WX9401;
wire WX2549;
wire WX1724;
wire WX10058;
wire WX7900;
wire WX6124;
wire WX438;
wire WX2840;
wire II14508;
wire WX6793;
wire II14879;
wire II30100;
wire II34810;
wire WX7999;
wire II6271;
wire II10503;
wire II19521;
wire WX10062;
wire WX3583;
wire II10682;
wire WX6630;
wire WX3738;
wire II6056;
wire WX9759;
wire WX3470;
wire WX2859;
wire WX6261;
wire II15621;
wire WX9420;
wire WX5434;
wire II30262;
wire II10743;
wire WX6691;
wire WX9629;
wire II19585;
wire WX2205;
wire WX9585;
wire II6048;
wire WX5216;
wire WX1090;
wire II26655;
wire II15492;
wire II10734;
wire II10082;
wire WX6297;
wire WX6401;
wire WX1957;
wire II22952;
wire II30481;
wire II10387;
wire II35582;
wire II30223;
wire WX9066;
wire WX4038;
wire II35532;
wire WX11094;
wire WX5514;
wire WX7693;
wire WX11487;
wire WX984;
wire WX6201;
wire II19189;
wire WX412;
wire WX10870;
wire WX11232;
wire II18675;
wire WX356;
wire WX4261;
wire II22238;
wire II31127;
wire II6181;
wire II26738;
wire WX11588;
wire WX4222;
wire WX10866;
wire WX2347;
wire II22153;
wire II2081;
wire WX7454;
wire WX5054;
wire II22944;
wire II34781;
wire WX9133;
wire WX7741;
wire WX2599;
wire II18566;
wire II30876;
wire WX6890;
wire WX8002;
wire WX2256;
wire WX10783;
wire WX460;
wire WX1746;
wire WX2479;
wire WX11378;
wire WX4229;
wire II6722;
wire WX7115;
wire WX1878;
wire WX2875;
wire WX9957;
wire II22556;
wire WX7367;
wire WX3025;
wire WX8375;
wire II6317;
wire II6274;
wire II30564;
wire WX11660;
wire WX2183;
wire WX8356;
wire WX4942;
wire II6559;
wire II15727;
wire II6729;
wire WX189;
wire II31655;
wire II2702;
wire II35326;
wire WX7759;
wire II34881;
wire II3184;
wire WX6452;
wire WX5222;
wire WX4705;
wire II14608;
wire II6612;
wire II26140;
wire WX8134;
wire WX1432;
wire WX2755;
wire II27239;
wire II3551;
wire WX219;
wire WX182;
wire II2841;
wire WX9437;
wire II27095;
wire WX2395;
wire WX10465;
wire WX3904;
wire II35729;
wire WX10087;
wire WX1376;
wire II10828;
wire WX3677;
wire WX7614;
wire WX6307;
wire WX5447;
wire II9998;
wire WX9511;
wire II2731;
wire WX8167;
wire II30231;
wire WX2470;
wire WX2203;
wire WX11503;
wire WX716;
wire WX6840;
wire WX10267;
wire II34114;
wire WX1741;
wire WX588;
wire WX322;
wire WX5253;
wire WX6766;
wire II26794;
wire WX7588;
wire WX11654;
wire WX2443;
wire WX7737;
wire WX6871;
wire WX4448;
wire II2532;
wire WX3952;
wire II2237;
wire WX1871;
wire WX7926;
wire WX2872;
wire WX6417;
wire WX5399;
wire WX5309;
wire WX9549;
wire II23526;
wire II18161;
wire WX2171;
wire WX10581;
wire WX8798;
wire WX10249;
wire II7358;
wire II18394;
wire II26605;
wire WX6803;
wire WX9990;
wire WX571;
wire II34516;
wire II23130;
wire II14988;
wire II10377;
wire WX9330;
wire WX8426;
wire WX9245;
wire II31620;
wire II35457;
wire WX8770;
wire II35731;
wire WX4137;
wire WX1979;
wire II35596;
wire WX7119;
wire II6955;
wire II34949;
wire WX4835;
wire WX6713;
wire WX298;
wire WX1726;
wire WX1600;
wire WX8877;
wire II3621;
wire WX8828;
wire WX9270;
wire WX3988;
wire WX231;
wire WX2386;
wire WX3729;
wire II27355;
wire II14066;
wire WX2371;
wire WX8186;
wire II23194;
wire WX5132;
wire WX4475;
wire II14125;
wire II10434;
wire WX8708;
wire II26020;
wire WX10156;
wire WX7076;
wire WX5248;
wire WX9339;
wire WX8659;
wire WX1115;
wire WX7239;
wire II27665;
wire WX1037;
wire II2717;
wire WX6107;
wire WX2816;
wire II30845;
wire II18295;
wire WX4462;
wire II30442;
wire WX4735;
wire WX9188;
wire II18358;
wire II30660;
wire II14274;
wire WX9477;
wire WX7402;
wire WX1913;
wire II22200;
wire II6163;
wire II10068;
wire WX1423;
wire II22826;
wire II19138;
wire II31704;
wire WX143;
wire II6388;
wire WX1656;
wire WX5478;
wire WX9476;
wire WX5804;
wire WX9952;
wire WX3938;
wire WX6216;
wire II22268;
wire II14501;
wire WX3609;
wire WX8933;
wire II34145;
wire II23658;
wire WX4079;
wire WX7708;
wire II23576;
wire WX2567;
wire WX3211;
wire WX7498;
wire WX9294;
wire II30078;
wire WX1142;
wire WX4641;
wire WX1052;
wire II22053;
wire II22678;
wire WX3922;
wire WX10098;
wire WX3637;
wire WX6834;
wire WX9468;
wire WX8762;
wire II11116;
wire II26640;
wire WX3941;
wire WX4495;
wire WX10654;
wire WX8936;
wire II30796;
wire WX3579;
wire WX9195;
wire WX97;
wire WX2723;
wire WX5740;
wire WX9608;
wire WX10878;
wire WX54;
wire WX2129;
wire WX4901;
wire II6604;
wire WX4500;
wire WX291;
wire II26740;
wire II35624;
wire WX10927;
wire II18938;
wire II11362;
wire II3065;
wire WX4771;
wire WX8721;
wire II22370;
wire WX6472;
wire II35709;
wire II31465;
wire WX10604;
wire II30667;
wire WX5416;
wire II23495;
wire WX10260;
wire WX1169;
wire WX6989;
wire WX8197;
wire II15536;
wire II19506;
wire WX5433;
wire WX814;
wire II18433;
wire WX7954;
wire II22306;
wire II22363;
wire WX4028;
wire WX10231;
wire WX640;
wire WX8003;
wire WX1102;
wire WX3410;
wire II30207;
wire WX752;
wire II31591;
wire WX10743;
wire II26375;
wire WX6131;
wire WX8116;
wire WX3645;
wire WX4226;
wire WX6093;
wire WX6985;
wire WX2766;
wire WX4996;
wire II6155;
wire WX7593;
wire WX1975;
wire II2408;
wire WX5050;
wire WX4749;
wire WX3795;
wire WX7048;
wire WX2163;
wire WX9396;
wire WX11594;
wire WX5984;
wire WX5022;
wire WX846;
wire WX7881;
wire WX1238;
wire II35341;
wire WX11289;
wire II14391;
wire WX3772;
wire II22105;
wire II30402;
wire WX4932;
wire WX396;
wire II11497;
wire WX5493;
wire WX10611;
wire WX5084;
wire WX766;
wire WX8170;
wire WX9559;
wire WX11664;
wire II6343;
wire II3170;
wire WX7725;
wire WX3000;
wire II3364;
wire II6203;
wire II10664;
wire WX6797;
wire II34820;
wire WX2843;
wire II26677;
wire II14972;
wire II26094;
wire WX9274;
wire II18411;
wire WX335;
wire WX2617;
wire WX434;
wire II3606;
wire WX8027;
wire II23220;
wire WX4108;
wire WX8050;
wire II6023;
wire WX2041;
wire II18465;
wire WX6859;
wire WX11032;
wire WX11670;
wire II26948;
wire WX2218;
wire WX6373;
wire WX2531;
wire WX10796;
wire WX3541;
wire II10123;
wire II35647;
wire II3078;
wire WX8379;
wire WX11362;
wire WX5799;
wire WX2938;
wire WX6012;
wire WX1526;
wire WX7031;
wire II26513;
wire WX9328;
wire WX1022;
wire WX8803;
wire WX3076;
wire WX6557;
wire II6072;
wire WX8069;
wire WX4213;
wire WX1841;
wire II10818;
wire II15676;
wire II30659;
wire II18986;
wire WX8226;
wire II26941;
wire WX8498;
wire II26965;
wire II22168;
wire WX5834;
wire WX3290;
wire WX6235;
wire II10361;
wire WX9998;
wire WX8948;
wire II34292;
wire WX8866;
wire II18280;
wire WX10473;
wire WX2155;
wire WX5811;
wire II34794;
wire II2298;
wire II10000;
wire II2864;
wire WX1404;
wire II35604;
wire II15145;
wire WX5045;
wire WX8779;
wire WX6812;
wire WX6612;
wire WX9847;
wire II27602;
wire WX4681;
wire WX4917;
wire WX477;
wire WX119;
wire WX4812;
wire WX6251;
wire WX10083;
wire II26854;
wire WX3652;
wire WX2852;
wire WX6142;
wire WX8020;
wire II10640;
wire II15407;
wire WX9321;
wire II14157;
wire II10858;
wire II22275;
wire WX2305;
wire WX6929;
wire WX11200;
wire WX6077;
wire WX1616;
wire WX9117;
wire WX2352;
wire WX4788;
wire WX5474;
wire II3340;
wire II26909;
wire II2563;
wire II14537;
wire II14528;
wire WX1588;
wire WX11592;
wire WX10124;
wire WX1017;
wire II22873;
wire WX8296;
wire WX4852;
wire WX481;
wire WX6509;
wire WX8041;
wire WX2226;
wire WX8442;
wire WX1592;
wire WX2480;
wire II34068;
wire II30548;
wire WX3205;
wire II22789;
wire II2932;
wire WX7940;
wire WX3934;
wire WX890;
wire WX7219;
wire WX7383;
wire WX11052;
wire WX10270;
wire II7489;
wire WX4577;
wire WX1191;
wire WX156;
wire WX124;
wire WX7551;
wire WX3049;
wire WX7329;
wire II14840;
wire II15704;
wire II26747;
wire II22089;
wire II26180;
wire WX8080;
wire WX10387;
wire WX1144;
wire II30365;
wire WX595;
wire WX11626;
wire II10797;
wire II22169;
wire II35524;
wire WX1661;
wire II23129;
wire WX1507;
wire II10448;
wire II18287;
wire WX938;
wire WX1244;
wire II26118;
wire WX7421;
wire II35224;
wire WX4491;
wire WX8971;
wire WX5127;
wire WX7910;
wire WX7978;
wire WX8702;
wire II34274;
wire II6295;
wire II22417;
wire WX166;
wire II14237;
wire WX6742;
wire WX1696;
wire WX2837;
wire II26159;
wire WX10459;
wire WX5838;
wire II26187;
wire WX10380;
wire WX3035;
wire WX2563;
wire WX9618;
wire II30302;
wire WX1809;
wire WX7470;
wire WX6897;
wire WX1491;
wire II2300;
wire II11245;
wire II2732;
wire II15517;
wire II6644;
wire WX6891;
wire WX2967;
wire WX2702;
wire WX3632;
wire WX1366;
wire WX7819;
wire II27369;
wire WX4906;
wire WX5574;
wire II26547;
wire WX10685;
wire WX9388;
wire II18690;
wire WX8782;
wire WX3216;
wire WX3069;
wire WX3432;
wire WX1683;
wire WX1652;
wire WX1967;
wire WX3749;
wire WX3831;
wire II14376;
wire WX3566;
wire WX3760;
wire II34073;
wire WX4240;
wire WX8231;
wire II30373;
wire II27735;
wire II6658;
wire II23233;
wire WX5840;
wire WX3480;
wire II14957;
wire WX1558;
wire WX2365;
wire WX6048;
wire II31662;
wire II2079;
wire WX2111;
wire II15393;
wire II34494;
wire II30335;
wire WX7667;
wire II22695;
wire WX7416;
wire II6859;
wire WX6182;
wire WX7948;
wire WX9058;
wire II23575;
wire WX7001;
wire WX9020;
wire WX4433;
wire II26499;
wire II30953;
wire WX1314;
wire WX8538;
wire WX5774;
wire WX7542;
wire WX10191;
wire WX8518;
wire WX3173;
wire WX540;
wire WX9577;
wire II18148;
wire WX8182;
wire WX3816;
wire WX6935;
wire WX5466;
wire II19464;
wire II34522;
wire WX1063;
wire WX7393;
wire WX4829;
wire II35471;
wire II22631;
wire WX607;
wire WX1659;
wire WX4159;
wire II2042;
wire WX11571;
wire WX7688;
wire II14632;
wire II19655;
wire WX4234;
wire II26593;
wire II2670;
wire WX7619;
wire II14282;
wire WX2707;
wire II11615;
wire WX11632;
wire WX10011;
wire WX5608;
wire WX5731;
wire II2951;
wire WX1551;
wire II26801;
wire WX928;
wire WX11556;
wire WX2906;
wire WX4150;
wire WX4795;
wire WX6363;
wire WX11552;
wire WX7165;
wire II6823;
wire II18271;
wire WX1439;
wire II3676;
wire II6367;
wire WX1903;
wire II2839;
wire WX3334;
wire II15223;
wire II2321;
wire WX5068;
wire WX3995;
wire II3472;
wire II22012;
wire WX8472;
wire WX5454;
wire II26962;
wire II34501;
wire WX7054;
wire WX7681;
wire WX2414;
wire II6738;
wire II30922;
wire II18319;
wire II26671;
wire II10472;
wire WX4819;
wire II6582;
wire II30217;
wire WX10440;
wire II2622;
wire WX10071;
wire WX10517;
wire II30603;
wire WX5968;
wire WX5526;
wire II10541;
wire II6863;
wire WX7989;
wire WX7892;
wire II18898;
wire WX6167;
wire II34515;
wire II6077;
wire II34231;
wire II22647;
wire WX4198;
wire WX160;
wire II18102;
wire II19519;
wire WX8982;
wire II27579;
wire WX6639;
wire II18536;
wire WX11504;
wire WX3958;
wire II26832;
wire II34128;
wire II26886;
wire II6568;
wire II10020;
wire II14452;
wire WX2312;
wire WX2601;
wire II14895;
wire WX6722;
wire WX11599;
wire WX4976;
wire WX11244;
wire II26016;
wire WX10179;
wire II6132;
wire II27108;
wire II2958;
wire WX209;
wire II3502;
wire II18528;
wire WX455;
wire WX10771;
wire WX11401;
wire WX8323;
wire II3579;
wire WX8248;
wire WX4551;
wire WX9939;
wire WX11278;
wire II6443;
wire II22408;
wire II18504;
wire WX3487;
wire II30629;
wire II30641;
wire WX10119;
wire II30767;
wire II26127;
wire WX8237;
wire II2437;
wire WX8221;
wire WX11557;
wire II23181;
wire II22144;
wire II18141;
wire II22790;
wire WX2924;
wire WX4445;
wire II2245;
wire II10182;
wire II31571;
wire II11441;
wire WX2734;
wire WX6190;
wire WX553;
wire WX11484;
wire WX6381;
wire WX2691;
wire WX7639;
wire II26731;
wire WX382;
wire II34035;
wire II10548;
wire WX3948;
wire WX8140;
wire II2026;
wire WX7565;
wire WX5994;
wire II26977;
wire II30914;
wire II34817;
wire WX10864;
wire WX9344;
wire WX6494;
wire II22075;
wire WX7099;
wire II18738;
wire II19646;
wire WX364;
wire II7710;
wire WX7997;
wire II10960;
wire II7137;
wire II27447;
wire WX2492;
wire II18891;
wire II14267;
wire II18365;
wire II30900;
wire WX3165;
wire WX3823;
wire II2879;
wire WX10892;
wire WX1852;
wire WX4012;
wire II6490;
wire II30782;
wire II27516;
wire WX2299;
wire WX4929;
wire WX8788;
wire II34957;
wire WX1419;
wire WX10767;
wire WX10645;
wire WX9261;
wire WX4019;
wire II26212;
wire II34987;
wire WX10809;
wire WX8923;
wire II11561;
wire WX2625;
wire II15628;
wire WX2333;
wire WX7992;
wire WX1634;
wire WX8093;
wire WX5105;
wire WX10091;
wire WX9088;
wire II15197;
wire WX6761;
wire II2607;
wire II26879;
wire WX5509;
wire WX3052;
wire WX1480;
wire WX2986;
wire II31373;
wire II3684;
wire II14878;
wire II26662;
wire WX6520;
wire WX10776;
wire WX10435;
wire II23365;
wire WX87;
wire WX8014;
wire II34586;
wire WX5083;
wire II10787;
wire II10415;
wire WX9986;
wire II6799;
wire II26337;
wire WX4920;
wire II27685;
wire WX5738;
wire WX10325;
wire II34247;
wire II23077;
wire WX6034;
wire II23390;
wire II14756;
wire II22197;
wire WX11110;
wire WX2806;
wire WX3150;
wire WX8909;
wire WX4116;
wire WX4841;
wire WX6786;
wire II22895;
wire WX4205;
wire II6195;
wire WX9869;
wire WX10740;
wire WX10426;
wire WX5205;
wire WX10679;
wire WX999;
wire WX4898;
wire II34438;
wire WX407;
wire WX2462;
wire WX11046;
wire WX6971;
wire II14198;
wire WX6096;
wire WX4874;
wire WX10076;
wire II10306;
wire WX3160;
wire II35236;
wire WX9929;
wire WX7440;
wire II11102;
wire WX112;
wire WX3919;
wire WX1126;
wire WX4895;
wire WX10676;
wire WX10727;
wire II27727;
wire WX5197;
wire WX10948;
wire WX9281;
wire WX9807;
wire II18967;
wire II11426;
wire WX9731;
wire WX3705;
wire II18040;
wire II18427;
wire WX9169;
wire II14793;
wire WX6341;
wire WX6944;
wire WX224;
wire II30062;
wire WX9394;
wire WX1162;
wire II19280;
wire II34469;
wire II30859;
wire II14693;
wire WX1512;
wire WX9160;
wire WX1343;
wire WX9491;
wire WX2292;
wire II10896;
wire WX3294;
wire WX4251;
wire II26986;
wire II3287;
wire WX8401;
wire WX10959;
wire WX9311;
wire WX8890;
wire II18704;
wire II34152;
wire II30705;
wire WX6223;
wire WX9301;
wire II2228;
wire WX8124;
wire II19564;
wire WX4631;
wire II34925;
wire II23376;
wire II31564;
wire WX9791;
wire WX10038;
wire II2825;
wire WX5317;
wire II6921;
wire II34199;
wire II11454;
wire WX11526;
wire WX9269;
wire II2638;
wire WX7969;
wire WX4665;
wire WX4480;
wire WX9424;
wire WX2089;
wire WX9537;
wire WX1403;
wire WX5783;
wire II19164;
wire WX6431;
wire II22439;
wire WX1619;
wire WX3607;
wire II35590;
wire WX1768;
wire WX2236;
wire WX6620;
wire II26685;
wire II14919;
wire II15237;
wire WX7965;
wire WX3615;
wire WX7377;
wire II34486;
wire II14885;
wire II19578;
wire II18079;
wire II15634;
wire WX5233;
wire II10710;
wire WX9639;
wire II18038;
wire WX3312;
wire II11284;
wire WX5619;
wire WX10251;
wire WX2943;
wire WX9983;
wire WX10491;
wire WX10498;
wire WX2669;
wire WX11471;
wire WX10802;
wire WX1985;
wire WX6296;
wire WX8055;
wire WX7984;
wire WX7092;
wire II10131;
wire WX1627;
wire II15559;
wire WX4882;
wire WX9839;
wire WX5097;
wire II19528;
wire WX6732;
wire WX7255;
wire II30455;
wire WX654;
wire II15578;
wire WX3526;
wire WX6158;
wire II30094;
wire II3132;
wire WX11395;
wire WX9019;
wire WX6826;
wire II11693;
wire II7561;
wire WX9703;
wire II10005;
wire WX10141;
wire WX5752;
wire II2305;
wire WX6932;
wire WX1641;
wire II2191;
wire II18009;
wire WX1355;
wire WX6385;
wire WX5240;
wire WX10922;
wire II22926;
wire II30676;
wire WX852;
wire II34135;
wire II22771;
wire WX6644;
wire II22539;
wire WX11004;
wire WX4436;
wire WX1155;
wire II30543;
wire II14025;
wire WX10565;
wire WX10225;
wire II3195;
wire II22610;
wire WX3238;
wire WX6232;
wire WX10832;
wire II26957;
wire II10456;
wire II34563;
wire II3196;
wire II2206;
wire II2345;
wire II22911;
wire II35431;
wire WX327;
wire II22299;
wire WX3720;
wire WX7034;
wire II18456;
wire II18714;
wire WX6901;
wire II31008;
wire II34448;
wire WX5427;
wire WX5459;
wire II35172;
wire II6108;
wire II11090;
wire II18644;
wire WX5118;
wire WX2979;
wire II22066;
wire II22573;
wire WX8799;
wire WX6675;
wire WX403;
wire II34360;
wire WX5615;
wire II18061;
wire II15485;
wire II2792;
wire II26149;
wire WX2390;
wire II26637;
wire WX6670;
wire WX11497;
wire WX62;
wire II22857;
wire WX2952;
wire II23618;
wire WX10430;
wire WX6685;
wire WX10540;
wire II6126;
wire II34369;
wire WX6773;
wire II35724;
wire II3325;
wire II2919;
wire WX11349;
wire WX2863;
wire WX3693;
wire WX2891;
wire WX4356;
wire II14187;
wire WX3672;
wire WX5768;
wire WX10916;
wire WX1754;
wire WX4810;
wire II14910;
wire WX6379;
wire WX3687;
wire WX6285;
wire WX3044;
wire WX7406;
wire II6016;
wire II22673;
wire II22182;
wire WX1748;
wire WX6862;
wire WX9159;
wire II35380;
wire II6630;
wire II2858;
wire II22836;
wire WX11306;
wire WX1494;
wire WX10209;
wire WX2860;
wire WX7409;
wire II6460;
wire WX317;
wire II23708;
wire WX8500;
wire WX7601;
wire II10687;
wire WX3843;
wire WX5530;
wire WX7592;
wire II6224;
wire WX7223;
wire II34185;
wire II10093;
wire WX1206;
wire II15342;
wire WX2147;
wire II10648;
wire II35378;
wire WX3767;
wire II22975;
wire WX4070;
wire WX1059;
wire II10594;
wire WX3789;
wire WX3187;
wire WX9252;
wire WX1146;
wire WX3989;
wire WX8138;
wire WX10137;
wire II10904;
wire WX11434;
wire II6333;
wire WX9174;
wire II30025;
wire WX5537;
wire WX9765;
wire WX6412;
wire WX4820;
wire WX11154;
wire II7188;
wire II6932;
wire WX7765;
wire WX5329;
wire WX8745;
wire WX121;
wire WX3756;
wire WX9213;
wire II2281;
wire WX8713;
wire II34076;
wire II30549;
wire WX6238;
wire WX4338;
wire II23590;
wire II6334;
wire II30977;
wire II10516;
wire II18843;
wire WX5279;
wire WX4677;
wire WX10402;
wire II34896;
wire II35393;
wire WX5387;
wire WX9034;
wire WX4335;
wire II35131;
wire WX6883;
wire II34223;
wire WX11431;
wire WX4621;
wire WX10614;
wire II30830;
wire II30820;
wire II26312;
wire WX5286;
wire II3628;
wire II18829;
wire WX1045;
wire WX10992;
wire WX1624;
wire WX5404;
wire WX3755;
wire WX9202;
wire WX5217;
wire II3501;
wire WX2555;
wire WX426;
wire II2693;
wire WX7533;
wire WX9978;
wire WX7785;
wire II34641;
wire WX6277;
wire WX6403;
wire WX2383;
wire WX7237;
wire WX2496;
wire WX5745;
wire II3530;
wire WX10824;
wire WX8321;
wire WX3538;
wire WX1184;
wire WX285;
wire WX6866;
wire WX11392;
wire II27742;
wire WX8881;
wire WX1153;
wire II7604;
wire II10229;
wire II34355;
wire WX8408;
wire WX3180;
wire WX6399;
wire II31412;
wire II26173;
wire II10113;
wire WX950;
wire II27122;
wire WX4767;
wire WX10638;
wire WX4162;
wire II14771;
wire WX10943;
wire WX9430;
wire WX6875;
wire II26392;
wire WX8848;
wire WX7521;
wire II26281;
wire II30984;
wire WX6428;
wire WX7249;
wire WX7390;
wire WX1139;
wire WX6476;
wire WX9819;
wire WX141;
wire II26894;
wire II10773;
wire WX10975;
wire WX3158;
wire WX5892;
wire II18823;
wire WX10312;
wire WX2453;
wire II14227;
wire WX10140;
wire WX5332;
wire WX2607;
wire WX486;
wire II2344;
wire WX5784;
wire WX9337;
wire II2756;
wire WX3690;
wire WX2421;
wire WX2061;
wire WX11288;
wire WX2402;
wire WX9352;
wire II18396;
wire WX349;
wire WX9215;
wire WX7569;
wire WX11472;
wire WX2200;
wire II34600;
wire WX8165;
wire II7370;
wire WX1048;
wire WX997;
wire WX11650;
wire II11603;
wire WX5259;
wire WX2303;
wire WX2811;
wire WX9335;
wire WX1351;
wire II19704;
wire II27552;
wire WX10628;
wire II34617;
wire WX9172;
wire II19423;
wire WX3215;
wire WX11432;
wire WX2964;
wire WX10309;
wire WX10908;
wire WX1125;
wire WX7703;
wire WX11441;
wire II27559;
wire WX5488;
wire WX1863;
wire II14377;
wire WX8145;
wire WX2472;
wire II2390;
wire WX7289;
wire WX9611;
wire II2524;
wire II6382;
wire II6208;
wire II22228;
wire II18922;
wire II2715;
wire WX3356;
wire II19087;
wire II31711;
wire WX5266;
wire II26175;
wire WX4444;
wire II30076;
wire II35751;
wire II7512;
wire WX7855;
wire II26266;
wire WX8005;
wire WX5305;
wire WX6847;
wire WX2485;
wire WX10135;
wire II30745;
wire WX10117;
wire WX8162;
wire WX11604;
wire WX8179;
wire II14601;
wire WX10457;
wire WX4450;
wire WX10228;
wire II2826;
wire WX10263;
wire WX2344;
wire II31179;
wire II6567;
wire II10790;
wire II22696;
wire WX5481;
wire WX1694;
wire II2639;
wire WX4945;
wire WX6279;
wire WX11136;
wire II11259;
wire WX6210;
wire II2872;
wire II19513;
wire WX10099;
wire WX2223;
wire II27614;
wire II22936;
wire II34919;
wire WX4160;
wire WX5692;
wire WX10820;
wire II10657;
wire WX10092;
wire II15418;
wire WX9626;
wire II6893;
wire II22191;
wire II26420;
wire II35591;
wire WX3326;
wire II15566;
wire II2462;
wire II10694;
wire WX7404;
wire II26436;
wire WX11511;
wire WX7017;
wire WX8696;
wire II18876;
wire WX9448;
wire II26559;
wire II6069;
wire II10974;
wire II18976;
wire WX488;
wire II19216;
wire WX421;
wire II26583;
wire II6970;
wire WX9857;
wire WX946;
wire II2367;
wire WX2399;
wire II22058;
wire II7279;
wire WX11309;
wire WX1025;
wire II34205;
wire WX5617;
wire WX353;
wire WX318;
wire WX6184;
wire WX10296;
wire II22121;
wire II22340;
wire WX4571;
wire WX8871;
wire II6032;
wire WX3633;
wire II35667;
wire WX4096;
wire WX3400;
wire WX784;
wire II34626;
wire WX5120;
wire WX5606;
wire WX2385;
wire WX1288;
wire WX3380;
wire II26621;
wire WX3671;
wire WX7507;
wire WX4346;
wire WX9811;
wire WX4555;
wire WX1653;
wire II2513;
wire II2482;
wire WX8727;
wire WX8640;
wire WX8440;
wire WX2615;
wire II3351;
wire WX6580;
wire WX3100;
wire WX11269;
wire II7584;
wire WX7901;
wire WX6525;
wire WX9471;
wire WX6638;
wire WX359;
wire II34664;
wire WX6879;
wire II10077;
wire WX6913;
wire II2204;
wire WX3284;
wire II18645;
wire WX4413;
wire WX9299;
wire II26342;
wire WX273;
wire WX9176;
wire II10735;
wire II23117;
wire WX9198;
wire WX3454;
wire WX11429;
wire WX8709;
wire WX9291;
wire WX3808;
wire II10322;
wire II2327;
wire II19584;
wire II2103;
wire II23611;
wire WX9993;
wire II18520;
wire WX11499;
wire WX2983;
wire WX11644;
wire WX5793;
wire II14553;
wire WX4471;
wire WX8502;
wire II7423;
wire II27507;
wire WX7494;
wire WX7077;
wire WX340;
wire II18815;
wire WX6144;
wire II6008;
wire II10355;
wire WX5918;
wire II27522;
wire WX8111;
wire II2669;
wire WX4131;
wire II35197;
wire II22960;
wire WX8847;
wire II27637;
wire WX6117;
wire WX1056;
wire II6792;
wire II30511;
wire WX3224;
wire WX983;
wire WX1574;
wire II6574;
wire WX10709;
wire WX8077;
wire WX65;
wire II34788;
wire WX9671;
wire WX5637;
wire II26388;
wire WX3611;
wire II2267;
wire II22042;
wire II6584;
wire II26032;
wire WX84;
wire II18162;
wire WX7052;
wire WX3020;
wire WX10725;
wire WX1953;
wire WX6411;
wire WX8031;
wire II6427;
wire WX2087;
wire II18940;
wire WX8650;
wire WX1451;
wire WX746;
wire WX7355;
wire WX6714;
wire II22400;
wire II10121;
wire WX5094;
wire WX6610;
wire II23646;
wire II3403;
wire WX9310;
wire WX5373;
wire II22438;
wire II30698;
wire WX1164;
wire WX10503;
wire WX8733;
wire WX3199;
wire II10099;
wire II10309;
wire II7626;
wire WX3663;
wire II23624;
wire II7476;
wire WX479;
wire WX1119;
wire WX1815;
wire II10866;
wire II26972;
wire WX10955;
wire WX10397;
wire II11657;
wire WX3252;
wire II35328;
wire WX5426;
wire WX207;
wire II7483;
wire WX6687;
wire II34927;
wire WX8205;
wire WX4635;
wire II14539;
wire WX2946;
wire WX10158;
wire WX5376;
wire II2389;
wire WX2664;
wire II30510;
wire WX2672;
wire II2832;
wire WX6206;
wire II6041;
wire WX139;
wire WX6874;
wire WX5231;
wire II18326;
wire WX7436;
wire WX2255;
wire WX5234;
wire WX6895;
wire WX9569;
wire WX10600;
wire II22480;
wire II15712;
wire WX5145;
wire II15158;
wire WX2658;
wire II2896;
wire WX7676;
wire WX2931;
wire WX10541;
wire II34571;
wire WX264;
wire WX6843;
wire WX1668;
wire WX7462;
wire WX660;
wire WX2681;
wire WX11226;
wire II14468;
wire WX2876;
wire WX10619;
wire WX11252;
wire WX3029;
wire WX1876;
wire WX6892;
wire WX3128;
wire WX637;
wire WX7699;
wire II11089;
wire II22308;
wire WX7450;
wire WX4316;
wire WX10302;
wire II19450;
wire WX8176;
wire II22587;
wire WX8215;
wire WX4609;
wire WX6772;
wire WX2211;
wire WX6621;
wire WX7998;
wire II2692;
wire WX4846;
wire WX109;
wire WX2115;
wire WX9972;
wire WX3826;
wire II18487;
wire WX5592;
wire II7661;
wire WX9660;
wire II18892;
wire WX9390;
wire WX6997;
wire WX8864;
wire II14320;
wire WX6464;
wire WX3701;
wire WX9182;
wire WX9507;
wire WX10039;
wire WX8152;
wire WX5073;
wire WX5008;
wire WX2804;
wire II22301;
wire II34285;
wire WX75;
wire WX4331;
wire WX6303;
wire WX2759;
wire WX115;
wire II35366;
wire II18800;
wire WX10081;
wire II7519;
wire WX1414;
wire WX1255;
wire WX292;
wire WX2992;
wire WX3968;
wire II14513;
wire WX1147;
wire II10524;
wire WX3396;
wire II35555;
wire WX9255;
wire II30597;
wire WX2409;
wire WX8831;
wire WX3733;
wire WX2017;
wire II26047;
wire WX1881;
wire II26026;
wire WX4369;
wire II14389;
wire WX8159;
wire II23700;
wire II6705;
wire WX432;
wire II18495;
wire II22982;
wire WX4138;
wire WX3562;
wire II2592;
wire WX5723;
wire WX6293;
wire II15159;
wire II23104;
wire WX10390;
wire WX3963;
wire II10573;
wire WX2628;
wire WX5328;
wire II34213;
wire WX9212;
wire WX5296;
wire II6146;
wire II30620;
wire II30970;
wire II30456;
wire WX8059;
wire WX11387;
wire II23610;
wire WX5518;
wire WX3278;
wire II14842;
wire II26995;
wire WX1011;
wire WX7072;
wire WX9953;
wire II2594;
wire II35509;
wire II30347;
wire WX808;
wire II6196;
wire II18550;
wire WX5004;
wire II15690;
wire WX1825;
wire WX7480;
wire WX10461;
wire WX4342;
wire II14981;
wire II10508;
wire WX8284;
wire WX2692;
wire II31514;
wire II22114;
wire WX5012;
wire WX944;
wire WX7487;
wire WX11255;
wire WX8903;
wire II6226;
wire II27588;
wire WX11544;
wire WX3176;
wire WX7335;
wire WX6423;
wire WX5684;
wire WX5820;
wire WX8823;
wire WX9445;
wire II6413;
wire WX7425;
wire II22135;
wire WX7127;
wire WX1245;
wire WX2231;
wire WX240;
wire II11439;
wire WX6667;
wire WX5319;
wire WX1399;
wire II34097;
wire WX7879;
wire II22802;
wire WX4966;
wire WX9369;
wire WX6914;
wire WX10765;
wire WX6649;
wire II26760;
wire WX2075;
wire II10873;
wire II10092;
wire II10155;
wire WX1470;
wire WX7495;
wire II18652;
wire WX7874;
wire WX8392;
wire WX8693;
wire WX904;
wire II34462;
wire WX4284;
wire WX3194;
wire WX11276;
wire WX6060;
wire WX2695;
wire II34553;
wire WX11334;
wire II2160;
wire WX6660;
wire II26019;
wire WX10194;
wire II18165;
wire WX9121;
wire WX4302;
wire WX1364;
wire II2966;
wire II30210;
wire II30589;
wire WX6397;
wire WX11313;
wire WX4713;
wire WX7686;
wire WX3949;
wire WX6762;
wire WX3512;
wire WX8187;
wire II35379;
wire WX4806;
wire WX5970;
wire II30046;
wire II26221;
wire WX11564;
wire WX274;
wire WX4296;
wire WX7652;
wire WX3807;
wire II15458;
wire II34300;
wire II7304;
wire WX6615;
wire II30496;
wire II27530;
wire II34742;
wire WX1700;
wire WX7062;
wire WX2302;
wire WX4881;
wire WX8558;
wire WX732;
wire WX2581;
wire WX7317;
wire II26220;
wire II31746;
wire WX650;
wire WX5406;
wire WX9103;
wire WX7731;
wire II26251;
wire WX6807;
wire WX2577;
wire WX2889;
wire WX9646;
wire II3313;
wire WX2488;
wire II19681;
wire WX238;
wire WX389;
wire WX9682;
wire II30242;
wire II18838;
wire II18559;
wire WX3220;
wire II34440;
wire WX5272;
wire WX2193;
wire WX7668;
wire WX11507;
wire WX6334;
wire II34974;
wire WX7469;
wire WX9941;
wire WX6056;
wire WX1308;
wire II30418;
wire WX1791;
wire WX2826;
wire II2098;
wire WX7347;
wire II11504;
wire II2655;
wire II6673;
wire WX7457;
wire II11701;
wire II15420;
wire II35011;
wire WX3426;
wire II7563;
wire II2780;
wire II6900;
wire II10555;
wire WX630;
wire II1997;
wire WX964;
wire WX9042;
wire WX11403;
wire II15289;
wire II34314;
wire WX7871;
wire WX7906;
wire WX626;
wire WX4529;
wire WX37;
wire II2290;
wire WX5650;
wire WX1731;
wire WX917;
wire WX2880;
wire WX6738;
wire WX9723;
wire WX2728;
wire II3689;
wire II22323;
wire WX4375;
wire WX179;
wire II2143;
wire II10191;
wire WX8929;
wire WX8668;
wire II23248;
wire II14702;
wire II2135;
wire WX6569;
wire WX5800;
wire WX4853;
wire WX1543;
wire WX7305;
wire II6472;
wire WX176;
wire II10511;
wire WX1479;
wire WX6112;
wire II30861;
wire II30162;
wire WX2209;
wire II27529;
wire WX7597;
wire WX295;
wire II18032;
wire WX6606;
wire II22270;
wire II35526;
wire II26368;
wire WX11376;
wire WX4751;
wire WX1682;
wire WX7417;
wire WX8312;
wire II18185;
wire WX11040;
wire WX9925;
wire II15487;
wire WX7540;
wire WX2915;
wire WX8914;
wire II27303;
wire WX6642;
wire WX170;
wire WX7622;
wire II35696;
wire WX603;
wire II23568;
wire WX3054;
wire WX8349;
wire II6860;
wire WX1538;
wire WX6405;
wire WX10553;
wire II14730;
wire WX11601;
wire II10959;
wire II22424;
wire II14748;
wire WX6560;
wire WX6274;
wire II6379;
wire II3158;
wire WX10210;
wire II15315;
wire WX10552;
wire II6358;
wire WX190;
wire WX2774;
wire II15586;
wire WX10688;
wire WX698;
wire II30410;
wire WX6756;
wire II22347;
wire WX7818;
wire WX11296;
wire WX10559;
wire WX4987;
wire II10136;
wire WX10223;
wire WX9903;
wire II3443;
wire II26714;
wire WX6083;
wire II18767;
wire II2653;
wire II11324;
wire II27693;
wire II34183;
wire II22865;
wire WX4114;
wire WX7472;
wire II26492;
wire WX5846;
wire WX10241;
wire II18340;
wire WX10880;
wire II6513;
wire WX9500;
wire WX9497;
wire WX2153;
wire WX500;
wire WX2934;
wire WX10181;
wire II6652;
wire WX1005;
wire WX7261;
wire WX4421;
wire II22464;
wire WX7724;
wire WX3969;
wire WX1530;
wire WX10952;
wire WX1505;
wire WX3978;
wire II10167;
wire WX3499;
wire II26746;
wire WX1733;
wire II30116;
wire WX9284;
wire II2012;
wire WX3336;
wire II19613;
wire WX9147;
wire WX2949;
wire II26823;
wire WX8149;
wire II18907;
wire II10611;
wire WX10432;
wire WX11126;
wire II10718;
wire WX1310;
wire WX2911;
wire II30707;
wire WX6528;
wire WX1449;
wire WX1711;
wire WX6364;
wire WX11140;
wire WX5037;
wire WX704;
wire II18140;
wire WX3206;
wire WX9406;
wire II30837;
wire WX3492;
wire WX9095;
wire WX6242;
wire WX10122;
wire II23539;
wire II31663;
wire II22656;
wire II18389;
wire WX927;
wire II35469;
wire WX935;
wire WX7939;
wire WX7524;
wire WX4325;
wire WX2341;
wire WX6433;
wire WX5562;
wire WX2529;
wire WX756;
wire II26855;
wire WX6813;
wire II30425;
wire II34981;
wire II15529;
wire WX9737;
wire II6264;
wire II3130;
wire WX5337;
wire WX4457;
wire WX9651;
wire WX7086;
wire WX8891;
wire WX3918;
wire WX7570;
wire II27251;
wire WX490;
wire WX8738;
wire II30610;
wire II11525;
wire WX5229;
wire II26156;
wire WX3716;
wire WX6050;
wire II7709;
wire II35562;
wire WX4060;
wire WX3820;
wire WX2520;
wire WX4782;
wire WX1465;
wire II31712;
wire II18155;
wire WX370;
wire II27253;
wire II35367;
wire II3565;
wire WX4075;
wire WX8206;
wire II26233;
wire II22748;
wire II10486;
wire II15557;
wire WX10531;
wire II31192;
wire WX5551;
wire WX11409;
wire II22261;
wire II18720;
wire WX9674;
wire WX5706;
wire II2516;
wire II7526;
wire WX10102;
wire II22021;
wire II26079;
wire WX8771;
wire WX6799;
wire II11652;
wire II18094;
wire WX415;
wire WX6196;
wire WX2984;
wire WX9654;
wire II31593;
wire WX9775;
wire WX7414;
wire II14694;
wire II30744;
wire WX4233;
wire II15249;
wire II2253;
wire II11141;
wire II31257;
wire II18071;
wire II23687;
wire WX4043;
wire II15656;
wire WX7831;
wire WX9411;
wire WX8012;
wire WX4034;
wire II6086;
wire WX1681;
wire II2049;
wire WX1842;
wire II23680;
wire WX11624;
wire WX1410;
wire WX10739;
wire II30117;
wire WX8630;
wire II30729;
wire WX4595;
wire WX5643;
wire WX4266;
wire WX8510;
wire II22569;
wire WX8118;
wire II18729;
wire WX3597;
wire WX1548;
wire II18589;
wire II30784;
wire WX1499;
wire WX5587;
wire II2331;
wire II10704;
wire II23602;
wire II35547;
wire WX7023;
wire WX1510;
wire WX10912;
wire WX1605;
wire II22549;
wire WX9861;
wire II27514;
wire WX2879;
wire WX694;
wire WX7822;
wire WX1566;
wire WX11481;
wire WX8532;
wire II30396;
wire WX6354;
wire II26963;
wire WX7988;
wire WX10216;
wire II6599;
wire WX5854;
wire WX9128;
wire WX5798;
wire WX7745;
wire II22547;
wire II6078;
wire II18580;
wire II18931;
wire WX7502;
wire WX5858;
wire WX4358;
wire II26419;
wire II18668;
wire II31284;
wire II18349;
wire WX10337;
wire WX10273;
wire II31592;
wire II14095;
wire II6699;
wire II10765;
wire II34345;
wire WX10793;
wire WX2788;
wire WX3474;
wire WX4147;
wire WX6626;
wire WX10445;
wire II14640;
wire WX5569;
wire WX1072;
wire II14932;
wire WX5074;
wire WX868;
wire WX6518;
wire II7239;
wire WX5809;
wire WX2264;
wire WX9093;
wire WX6788;
wire WX10042;
wire WX5647;
wire II27628;
wire WX1596;
wire II30324;
wire WX5103;
wire II14035;
wire II10291;
wire II19504;
wire WX9288;
wire WX10770;
wire WX3384;
wire WX6680;
wire WX8412;
wire II27671;
wire WX6360;
wire WX5654;
wire WX7209;
wire WX7066;
wire II7293;
wire WX8065;
wire WX2465;
wire WX1076;
wire II15514;
wire II6063;
wire WX7912;
wire WX1963;
wire II2066;
wire WX6759;
wire WX6671;
wire II19674;
wire WX7038;
wire II30200;
wire II22872;
wire II22154;
wire WX7815;
wire II22184;
wire WX4868;
wire WX4629;
wire II27266;
wire WX2069;
wire WX10470;
wire II34090;
wire II27344;
wire II6256;
wire II30293;
wire WX11352;
wire WX1328;
wire II14584;
wire WX6869;
wire WX2274;
wire WX8238;
wire WX3880;
wire WX5042;
wire WX2792;
wire WX1688;
wire WX11272;
wire II30853;
wire II31347;
wire WX1702;
wire II26296;
wire WX69;
wire II26609;
wire II18867;
wire WX11423;
wire II15355;
wire WX1274;
wire WX2081;
wire WX9835;
wire WX8720;
wire II19254;
wire II22354;
wire WX9465;
wire WX8754;
wire WX9248;
wire WX2107;
wire WX7201;
wire WX11536;
wire WX1585;
wire II18813;
wire WX9713;
wire WX8810;
wire WX3360;
wire WX10848;
wire WX9222;
wire II10844;
wire II14871;
wire II10880;
wire WX1374;
wire II10278;
wire II2887;
wire WX362;
wire II2360;
wire WX6496;
wire WX6949;
wire II35263;
wire WX8853;
wire WX9341;
wire II22477;
wire II11076;
wire WX10202;
wire WX1622;
wire II31440;
wire WX8710;
wire WX8957;
wire WX11142;
wire II6853;
wire WX1642;
wire WX52;
wire WX2674;
wire WX6931;
wire WX10586;
wire WX3912;
wire WX7617;
wire WX10452;
wire II2855;
wire II23630;
wire WX10410;
wire WX4517;
wire WX7922;
wire WX8673;
wire WX326;
wire WX5276;
wire II14777;
wire WX1759;
wire II2119;
wire WX9851;
wire WX2956;
wire WX3310;
wire WX1231;
wire II14817;
wire WX6402;
wire WX9783;
wire II26481;
wire WX8878;
wire II14273;
wire WX7842;
wire WX7719;
wire WX9200;
wire II27713;
wire WX5411;
wire II2212;
wire II26329;
wire II3327;
wire WX3753;
wire II34192;
wire WX5263;
wire WX237;
wire WX7990;
wire II18952;
wire II6465;
wire WX3750;
wire II3273;
wire II26143;
wire II7638;
wire WX8676;
wire II14656;
wire WX1855;
wire II31102;
wire II22510;
wire WX2444;
wire II10821;
wire II6177;
wire II15544;
wire II23518;
wire WX9436;
wire II26862;
wire II19230;
wire II31427;
wire WX8606;
wire WX2417;
wire WX5688;
wire WX10114;
wire II3431;
wire II34856;
wire WX3856;
wire WX9155;
wire II31634;
wire WX8396;
wire II2917;
wire II35133;
wire WX7767;
wire WX7098;
wire II30022;
wire II1986;
wire WX10623;
wire II34595;
wire II2779;
wire WX5252;
wire WX11190;
wire WX2387;
wire WX4673;
wire WX7671;
wire II14869;
wire WX7339;
wire WX80;
wire WX1932;
wire II6558;
wire II18233;
wire WX7663;
wire WX10424;
wire WX10593;
wire WX8353;
wire WX4823;
wire II10634;
wire WX2245;
wire WX243;
wire II10836;
wire WX1205;
wire II31478;
wire WX2897;
wire WX11416;
wire II35302;
wire WX11528;
wire WX9187;
wire II26257;
wire II31491;
wire WX10057;
wire II34081;
wire WX578;
wire WX7795;
wire II19228;
wire WX5744;
wire WX4193;
wire WX6006;
wire WX4121;
wire II34261;
wire WX1258;
wire II18056;
wire WX10633;
wire II10982;
wire WX377;
wire II30536;
wire WX1394;
wire WX5135;
wire II2050;
wire WX7585;
wire WX6150;
wire WX1890;
wire WX11501;
wire II15329;
wire WX10816;
wire II10014;
wire II15108;
wire WX4954;
wire II35275;
wire II26297;
wire WX10825;
wire II10742;
wire WX1770;
wire WX9519;
wire II2823;
wire II6939;
wire II34834;
wire WX5734;
wire II2641;
wire WX5224;
wire WX2767;
wire WX8943;
wire II2755;
wire WX11259;
wire WX6102;
wire WX4833;
wire WX7538;
wire WX3642;
wire WX5766;
wire WX3704;
wire II2972;
wire WX8131;
wire II14948;
wire II14808;
wire II18194;
wire WX2228;
wire WX9709;
wire WX10408;
wire WX1829;
wire WX6690;
wire WX1747;
wire WX7783;
wire WX6245;
wire WX6268;
wire II10464;
wire WX1639;
wire WX10052;
wire WX4016;
wire WX5347;
wire WX3862;
wire WX7697;
wire II30264;
wire II35185;
wire WX1522;
wire WX3146;
wire WX3155;
wire II14012;
wire WX6940;
wire II15601;
wire II2888;
wire II2802;
wire WX2551;
wire WX9343;
wire II11722;
wire II6125;
wire WX9000;
wire WX4925;
wire WX4013;
wire WX8967;
wire WX8661;
wire II11180;
wire WX5281;
wire II31586;
wire WX10987;
wire WX1847;
wire WX10742;
wire II7506;
wire II30714;
wire II34424;
wire WX6646;
wire WX4611;
wire WX6299;
wire II35288;
wire WX7600;
wire WX4816;
wire WX6961;
wire WX4923;
wire WX10986;
wire WX4255;
wire II34646;
wire II19332;
wire II14088;
wire II34764;
wire WX10367;
wire WX7835;
wire WX8097;
wire II35661;
wire WX5027;
wire II15622;
wire WX10329;
wire WX2410;
wire WX2854;
wire WX9891;
wire II23337;
wire WX464;
wire WX728;
wire II15719;
wire II26785;
wire II14211;
wire WX2121;
wire WX9086;
wire WX6338;
wire WX7323;
wire II27096;
wire II30092;
wire WX7544;
wire II26063;
wire II18069;
wire WX1900;
wire WX10777;
wire II35539;
wire WX7714;
wire II22951;
wire WX6231;
wire WX1981;
wire WX3616;
wire WX10151;
wire WX1106;
wire II2021;
wire II3591;
wire WX8018;
wire WX9263;
wire WX6227;
wire II14699;
wire WX5974;
wire WX11492;
wire WX9981;
wire II14048;
wire WX7395;
wire II14041;
wire II14662;
wire WX2336;
wire WX3582;
wire WX10937;
wire WX7035;
wire WX2502;
wire II2637;
wire WX4891;
wire II30892;
wire WX8863;
wire WX1430;
wire II26164;
wire WX2737;
wire WX1921;
wire WX7227;
wire II34491;
wire II14545;
wire WX428;
wire WX10784;
wire II2051;
wire II34670;
wire II14420;
wire WX4270;
wire II2352;
wire WX3169;
wire II26554;
wire WX3545;
wire WX8258;
wire WX3004;
wire WX8432;
wire WX7271;
wire WX1408;
wire WX6905;
wire WX11303;
wire WX3763;
wire WX2233;
wire WX9533;
wire WX7962;
wire II6053;
wire II6829;
wire II34695;
wire II2616;
wire II34609;
wire WX1137;
wire II2074;
wire WX2290;
wire II30156;
wire WX4601;
wire WX10657;
wire WX5908;
wire II26468;
wire II6553;
wire WX11329;
wire WX1897;
wire WX1345;
wire II35612;
wire II7383;
wire II10943;
wire II30691;
wire WX10805;
wire II14966;
wire WX5470;
wire II26776;
wire II6529;
wire WX2622;
wire II2260;
wire WX4461;
wire WX4112;
wire WX10437;
wire II30673;
wire WX2688;
wire II19492;
wire WX7159;
wire WX3041;
wire II26869;
wire WX1707;
wire II26406;
wire II23389;
wire WX7930;
wire II10208;
wire WX7111;
wire II6311;
wire WX10882;
wire WX474;
wire WX3569;
wire WX4731;
wire WX6175;
wire WX5577;
wire II34867;
wire II30836;
wire WX6531;
wire II35404;
wire WX502;
wire WX6346;
wire II30735;
wire II14925;
wire WX10274;
wire WX10172;
wire WX2972;
wire WX5912;
wire WX5866;
wire II22883;
wire WX1484;
wire II26816;
wire WX9015;
wire WX10641;
wire WX3038;
wire II27726;
wire II23502;
wire II6496;
wire WX599;
wire II15444;
wire II22818;
wire II10394;
wire II35745;
wire WX4053;
wire WX7483;
wire II18132;
wire II23496;
wire WX6036;
wire WX6938;
wire WX7102;
wire WX6172;
wire WX9234;
wire II14916;
wire II14435;
wire WX11585;
wire WX11014;
wire WX7960;
wire WX4309;
wire II35314;
wire WX10707;
wire WX6409;
wire II14019;
wire II18147;
wire II18131;
wire II18674;
wire II34401;
wire II7213;
wire WX4701;
wire WX6851;
wire WX8309;
wire II34578;
wire WX1224;
wire WX8638;
wire WX10495;
wire WX2595;
wire WX2494;
wire II35106;
wire II6070;
wire II30450;
wire II10719;
wire WX256;
wire II30907;
wire WX444;
wire II35701;
wire WX2328;
wire WX4201;
wire WX8107;
wire II14141;
wire II23090;
wire II26979;
wire II7492;
wire II2391;
wire II30130;
wire WX2373;
wire WX3306;
wire WX7628;
wire II30061;
wire WX921;
wire WX3724;
wire II22842;
wire II7058;
wire II2452;
wire WX8932;
wire II34252;
wire WX2951;
wire WX11230;
wire WX1121;
wire WX9012;
wire WX8937;
wire WX8962;
wire WX2175;
wire WX8548;
wire II6666;
wire II14104;
wire WX9054;
wire II15706;
wire II26903;
wire WX7605;
wire II10727;
wire II34557;
wire II2127;
wire WX6817;
wire WX2181;
wire WX2814;
wire II15171;
wire WX468;
wire WX4063;
wire II2625;
wire WX563;
wire WX2648;
wire II22292;
wire II26097;
wire II3222;
wire WX10064;
wire WX6327;
wire WX4174;
wire II22015;
wire WX9024;
wire II26946;
wire II30582;
wire WX3228;
wire WX3656;
wire WX986;
wire WX4212;
wire II26538;
wire II27291;
wire II27649;
wire WX6906;
wire WX6653;
wire WX3422;
wire WX9907;
wire II2599;
wire WX102;
wire II6534;
wire II10084;
wire WX6703;
wire II27566;
wire WX6106;
wire WX8359;
wire WX2797;
wire WX7389;
wire WX8210;
wire WX8270;
wire WX6718;
wire II30644;
wire WX966;
wire WX8219;
wire WX4799;
wire WX5815;
wire WX4001;
wire II27409;
wire WX5141;
wire II30574;
wire WX2929;
wire WX3555;
wire II15508;
wire WX5463;
wire II30884;
wire WX2718;
wire WX11595;
wire WX10722;
wire WX414;
wire II35688;
wire II11538;
wire II26708;
wire WX3834;
wire II2810;
wire WX7596;
wire WX8526;
wire WX6711;
wire II2243;
wire WX11194;
wire WX2752;
wire WX5601;
wire WX3067;
wire II19384;
wire II35006;
wire WX5187;
wire II6801;
wire II30936;
wire WX1140;
wire WX5623;
wire WX1335;
wire II11532;
wire II14594;
wire II18512;
wire WX5704;
wire WX9600;
wire II18914;
wire WX566;
wire WX6596;
wire WX4275;
wire II22138;
wire WX10896;
wire II14490;
wire WX6163;
wire WX2251;
wire II34383;
wire WX592;
wire II2796;
wire II18657;
wire II26459;
wire WX9692;
wire II2809;
wire WX828;
wire WX7579;
wire WX5785;
wire II11559;
wire WX2637;
wire WX1382;
wire WX10903;
wire WX9451;
wire WX2436;
wire WX7105;
wire WX3798;
wire II26227;
wire WX8026;
wire II2531;
wire WX2360;
wire II6544;
wire II23143;
wire WX874;
wire II30921;
wire II26181;
wire WX7554;
wire WX5308;
wire WX11104;
wire WX331;
wire WX8365;
wire WX393;
wire II31283;
wire WX9030;
wire WX8129;
wire WX4990;
wire WX10046;
wire WX9258;
wire WX7886;
wire II14763;
wire WX8978;
wire II34541;
wire WX1044;
wire II26616;
wire II30566;
wire WX3955;
wire WX6018;
wire II2221;
wire II30055;
wire WX3124;
wire II2453;
wire WX9414;
wire II6363;
wire II35496;
wire II26670;
wire WX6697;
wire WX544;
wire WX5521;
wire WX8300;
wire WX10698;
wire II18831;
wire WX7422;
wire II3522;
wire WX8993;
wire WX9805;
wire WX10763;
wire II11387;
wire II22524;
wire WX3213;
wire WX1779;
wire WX11559;
wire II2950;
wire WX6305;
wire WX8328;
wire II19571;
wire WX7632;
wire WX372;
wire WX2900;
wire II30488;
wire II26667;
wire II11518;
wire WX1084;
wire WX1458;
wire II19731;
wire II2684;
wire WX10996;
wire II11375;
wire II22082;
wire WX11573;
wire WX2369;
wire II34393;
wire II34454;
wire II2716;
wire WX2013;
wire WX6415;
wire WX4173;
wire WX9612;
wire WX618;
wire WX5495;
wire II23666;
wire WX8061;
wire WX11509;
wire II19688;
wire WX11060;
wire WX8985;
wire II34756;
wire WX3572;
wire WX3992;
wire WX1028;
wire II26072;
wire II14220;
wire WX3986;
wire WX3872;
wire WX6507;
wire WX2698;
wire II30249;
wire II30520;
wire WX5396;
wire WX6727;
wire WX6837;
wire II30521;
wire II19203;
wire WX4446;
wire WX3540;
wire II1989;
wire II31492;
wire WX5450;
wire WX2456;
wire II2284;
wire II22445;
wire II3209;
wire WX4999;
wire II15543;
wire WX5342;
wire WX5958;
wire II9999;
wire WX3534;
wire II3182;
wire WX4972;
wire WX2998;
wire WX4661;
wire II3641;
wire WX288;
wire WX11172;
wire WX11281;
wire II35540;
wire II14577;
wire WX9841;
wire WX4403;
wire WX3776;
wire II19241;
wire II30627;
wire II10914;
wire II22642;
wire II10151;
wire II26357;
wire WX6092;
wire WX688;
wire II2476;
wire II10494;
wire II14268;
wire II6180;
wire WX6576;
wire II30427;
wire WX10013;
wire II14978;
wire WX8019;
wire WX9006;
wire WX2536;
wire WX6790;
wire II11510;
wire WX7648;
wire WX9373;
wire WX9348;
wire WX888;
wire II14206;
wire II6659;
wire II31297;
wire II34377;
wire WX1529;
wire WX7388;
wire WX4312;
wire WX8741;
wire WX5439;
wire II30393;
wire WX2746;
wire II26676;
wire II10852;
wire WX1318;
wire WX2355;
wire II22921;
wire WX10333;
wire II27174;
wire WX300;
wire II2033;
wire II11142;
wire II6923;
wire WX644;
wire II26888;
wire II3390;
wire WX3594;
wire WX3929;
wire WX1922;
wire II26500;
wire WX10758;
wire WX812;
wire WX8765;
wire WX10661;
wire WX11263;
wire II2421;
wire II6489;
wire WX6802;
wire WX3791;
wire WX977;
wire WX3682;
wire WX6632;
wire WX910;
wire WX1248;
wire WX3460;
wire WX10751;
wire II26545;
wire WX5992;
wire WX2923;
wire WX8806;
wire WX1379;
wire II26576;
wire WX8190;
wire WX634;
wire WX2760;
wire II3619;
wire II10200;
wire II6977;
wire WX2801;
wire WX10096;
wire II11413;
wire II30829;
wire II26915;
wire WX7363;
wire II19557;
wire II18380;
wire WX10681;
wire WX6731;
wire II30503;
wire II26523;
wire WX213;
wire WX10079;
wire II22733;
wire WX2215;
wire II26042;
wire WX3446;
wire WX10747;
wire II34278;
wire WX6748;
wire II14467;
wire II31647;
wire WX8749;
wire II14723;
wire WX5876;
wire II23208;
wire WX214;
wire WX11290;
wire WX6594;
wire WX3999;
wire WX1261;
wire WX11612;
wire WX5087;
wire WX3200;
wire WX2307;
wire II23325;
wire WX3248;
wire II18108;
wire II18450;
wire WX11038;
wire II10833;
wire WX6922;
wire WX5322;
wire WX3378;
wire WX8222;
wire II34774;
wire II30185;
wire II3418;
wire II14050;
wire WX9795;
wire WX4593;
wire WX9441;
wire II7319;
wire WX6072;
wire WX8895;
wire WX9112;
wire WX8718;
wire II11350;
wire II2150;
wire II30319;
wire WX6135;
wire WX3172;
wire WX3915;
wire II11531;
wire WX1387;
wire WX1421;
wire II15081;
wire II3486;
wire II34174;
wire WX4934;
wire WX10025;
wire WX220;
wire II15531;
wire II11127;
wire II30753;
wire WX9513;
wire WX1918;
wire WX4224;
wire WX9325;
wire WX7972;
wire WX9317;
wire WX3620;
wire II6117;
wire WX4156;
wire WX11345;
wire WX10691;
wire II22702;
wire II26320;
wire WX8141;
wire WX4236;
wire II19321;
wire WX91;
wire WX4655;
wire II10757;
wire WX8777;
wire WX5112;
wire WX3011;
wire WX7802;
wire II2157;
wire II23588;
wire WX4217;
wire WX629;
wire WX11319;
wire WX1407;
wire II6103;
wire WX5364;
wire II14312;
wire II10052;
wire WX8290;
wire WX6044;
wire II30945;
wire II10635;
wire II26134;
wire WX5727;
wire II14599;
wire II22277;
wire WX3531;
wire II27187;
wire II19399;
wire II26693;
wire WX2834;
wire WX8368;
wire II27002;
wire WX152;
wire WX4952;
wire WX2719;
wire II30822;
wire II22712;
wire WX8045;
wire II19697;
wire II10601;
wire II19295;
wire WX4107;
wire WX11534;
wire WX7958;
wire WX10383;
wire WX4745;
wire WX6619;
wire WX4024;
wire WX44;
wire WX6099;
wire II23737;
wire II14810;
wire II18085;
wire WX6314;
wire II19268;
wire WX5756;
wire WX1977;
wire II10353;
wire II3052;
wire WX10448;
wire WX7095;
wire II2763;
wire II2297;
wire II30703;
wire II6212;
wire II6791;
wire WX5065;
wire WX1882;
wire II22060;
wire WX7943;
wire WX4321;
wire WX7259;
wire WX10716;
wire II14259;
wire II31739;
wire WX10961;
wire WX11668;
wire WX5777;
wire WX1769;
wire WX742;
wire WX5960;
wire WX9958;
wire II14770;
wire WX5596;
wire II27240;
wire WX2742;
wire WX10639;
wire II6838;
wire WX8038;
wire II30991;
wire WX1813;
wire WX7528;
wire II6279;
wire WX3037;
wire WX9278;
wire WX9300;
wire WX7749;
wire II34942;
wire WX2243;
wire WX6054;
wire WX9733;
wire WX11406;
wire II31007;
wire II7461;
wire WX11355;
wire II19475;
wire WX3667;
wire WX8700;
wire II10139;
wire WX7936;
wire WX8682;
wire II34913;
wire II30163;
wire WX6555;
wire II6770;
wire WX1885;
wire WX7041;
wire WX2119;
wire II30085;
wire II22046;
wire II22230;
wire WX10575;
wire II3066;
wire WX9351;
wire II6961;
wire II22260;
wire II14888;
wire II7254;
wire WX9845;
wire WX10728;
wire WX8156;
wire WX5230;
wire II27734;
wire II2089;
wire II14212;
wire WX9490;
wire WX232;
wire WX5487;
wire II27630;
wire WX10075;
wire II31527;
wire II18861;
wire WX3274;
wire WX8664;
wire WX1803;
wire WX9280;
wire WX5914;
wire WX3496;
wire WX1570;
wire WX3024;
wire II27448;
wire WX9755;
wire II10616;
wire WX5634;
wire WX9358;
wire II30107;
wire II26244;
wire WX10319;
wire WX8843;
wire WX229;
wire WX5418;
wire II2577;
wire WX5880;
wire II6677;
wire WX2942;
wire WX10729;
wire WX3914;
wire WX6570;
wire WX3589;
wire WX9565;
wire II10401;
wire II22493;
wire II30192;
wire WX2611;
wire II26476;
wire WX2135;
wire WX1064;
wire WX10483;
wire II18629;
wire WX10035;
wire WX1872;
wire II3288;
wire WX7475;
wire WX9161;
wire WX9623;
wire WX1342;
wire II2648;
wire WX4481;
wire II18475;
wire WX8121;
wire WX10615;
wire WX120;
wire WX8444;
wire WX9402;
wire WX941;
wire WX3839;
wire II18628;
wire WX1613;
wire WX3092;
wire WX7285;
wire WX4164;
wire II11643;
wire WX5504;
wire II22130;
wire WX9385;
wire WX5208;
wire WX6460;
wire WX9429;
wire II11231;
wire WX1213;
wire II2678;
wire II18217;
wire WX778;
wire WX11488;
wire WX3614;
wire WX8776;
wire WX10215;
wire WX296;
wire II18776;
wire WX4262;
wire WX4527;
wire WX11467;
wire II22557;
wire WX5117;
wire II10527;
wire II10764;
wire II26638;
wire WX6993;
wire II22882;
wire WX2736;
wire WX8070;
wire WX10678;
wire WX5024;
wire WX3151;
wire II7534;
wire II2236;
wire II6456;
wire II10627;
wire II34718;
wire II6357;
wire II3550;
wire II34672;
wire WX8001;
wire WX3525;
wire WX3436;
wire WX4237;
wire WX3288;
wire II11283;
wire II10379;
wire WX664;
wire WX4339;
wire II22904;
wire II22092;
wire WX1879;
wire WX3588;
wire II22943;
wire II7124;
wire WX5751;
wire WX3254;
wire II19625;
wire II18062;
wire WX5001;
wire WX3868;
wire WX7441;
wire WX1495;
wire II19267;
wire WX2668;
wire WX4863;
wire II6590;
wire WX2848;
wire WX1723;
wire WX111;
wire WX9628;
wire II7589;
wire WX622;
wire WX5630;
wire WX2548;
wire II3649;
wire WX1091;
wire II22485;
wire WX9875;
wire II18366;
wire II26521;
wire WX1163;
wire WX4941;
wire II27487;
wire WX6248;
wire II2948;
wire WX2841;
wire II26103;
wire II10897;
wire WX4030;
wire II6272;
wire WX2624;
wire WX4134;
wire WX2405;
wire WX10960;
wire II7541;
wire WX6643;
wire WX10277;
wire II2740;
wire WX2506;
wire WX1691;
wire II15493;
wire WX4511;
wire WX4769;
wire WX2976;
wire II23637;
wire WX1391;
wire WX1766;
wire II34230;
wire WX5243;
wire II10733;
wire II6441;
wire WX1134;
wire II31451;
wire WX8514;
wire II18611;
wire WX7394;
wire II10532;
wire WX1418;
wire WX3195;
wire WX8820;
wire WX4365;
wire WX6113;
wire WX9889;
wire WX5435;
wire WX2206;
wire WX1544;
wire WX11542;
wire WX8169;
wire WX930;
wire II2126;
wire II23260;
wire II6171;
wire II19437;
wire WX4779;
wire WX1725;
wire WX7814;
wire II18442;
wire WX11502;
wire II18519;
wire II26795;
wire WX7245;
wire II10423;
wire WX3694;
wire II7357;
wire WX8829;
wire II19100;
wire WX2873;
wire II22912;
wire WX8797;
wire WX5714;
wire WX6917;
wire II18781;
wire WX3737;
wire WX10250;
wire II6434;
wire WX9821;
wire WX1753;
wire WX2603;
wire WX8322;
wire II35730;
wire WX449;
wire WX1192;
wire II14065;
wire WX1232;
wire WX10583;
wire II14686;
wire WX9013;
wire WX11132;
wire WX4643;
wire II6723;
wire II19520;
wire WX5430;
wire WX7925;
wire WX2380;
wire WX11440;
wire II10060;
wire WX2257;
wire WX344;
wire WX3730;
wire WX3219;
wire WX4834;
wire WX2317;
wire WX7368;
wire WX2476;
wire WX2471;
wire II10408;
wire II7598;
wire WX9251;
wire II19709;
wire WX8135;
wire II7136;
wire WX5446;
wire WX11162;
wire WX11445;
wire WX10377;
wire WX5139;
wire II23625;
wire WX3188;
wire WX11279;
wire WX425;
wire WX7429;
wire WX5181;
wire II22650;
wire II7597;
wire WX4440;
wire WX5124;
wire II27123;
wire WX2968;
wire WX11476;
wire WX3710;
wire WX3003;
wire WX10369;
wire II6505;
wire II31522;
wire WX11236;
wire WX6217;
wire WX10548;
wire WX4468;
wire WX6306;
wire WX10088;
wire II6931;
wire WX1433;
wire WX183;
wire WX1156;
wire WX7359;
wire WX9482;
wire II7369;
wire WX2227;
wire WX145;
wire II6808;
wire II10433;
wire II34850;
wire WX4651;
wire II22766;
wire WX5301;
wire II26724;
wire WX2822;
wire WX8166;
wire II22772;
wire WX10759;
wire WX6323;
wire II22052;
wire II22833;
wire WX686;
wire WX1375;
wire WX985;
wire II30294;
wire II2902;
wire II2703;
wire WX3272;
wire WX5513;
wire WX7408;
wire WX314;
wire WX6126;
wire II6342;
wire II6372;
wire WX357;
wire II14654;
wire WX3508;
wire WX3190;
wire WX3819;
wire WX3638;
wire II35708;
wire WX3578;
wire II3326;
wire II27214;
wire II18862;
wire II30858;
wire WX3942;
wire WX8990;
wire WX2724;
wire II2857;
wire WX383;
wire II18039;
wire WX9997;
wire II35157;
wire II7603;
wire WX6684;
wire WX8997;
wire WX7710;
wire WX9609;
wire II14003;
wire II2095;
wire WX4900;
wire WX3842;
wire II2375;
wire WX3886;
wire WX8748;
wire WX9315;
wire II2486;
wire WX10004;
wire II31464;
wire II27651;
wire WX10144;
wire II2181;
wire WX4501;
wire WX1749;
wire WX11305;
wire WX10305;
wire WX7580;
wire II19534;
wire II6480;
wire WX10259;
wire WX6753;
wire WX8644;
wire II14870;
wire WX10224;
wire WX4230;
wire WX3930;
wire II30583;
wire II35512;
wire WX4506;
wire WX2817;
wire II15677;
wire WX9331;
wire II35619;
wire II30443;
wire WX5546;
wire WX5225;
wire WX4429;
wire II31507;
wire II22672;
wire II2517;
wire WX248;
wire II14935;
wire II31556;
wire WX10917;
wire WX11380;
wire WX277;
wire WX11648;
wire II31323;
wire II18296;
wire II34416;
wire WX6404;
wire II22958;
wire II18054;
wire II14343;
wire II6491;
wire WX8232;
wire II34166;
wire WX7073;
wire WX142;
wire WX780;
wire WX1657;
wire WX2987;
wire II11219;
wire II23481;
wire WX7707;
wire II22967;
wire II23681;
wire II22201;
wire WX4181;
wire WX336;
wire WX5468;
wire II18844;
wire WX8705;
wire WX3603;
wire WX11346;
wire WX6833;
wire II18971;
wire II6335;
wire WX10436;
wire WX10811;
wire WX6388;
wire WX3974;
wire WX9090;
wire WX6191;
wire WX528;
wire II3599;
wire WX61;
wire WX4347;
wire WX9678;
wire WX9493;
wire WX10008;
wire WX1867;
wire WX482;
wire WX10909;
wire WX3711;
wire II31691;
wire WX4071;
wire WX6488;
wire II6389;
wire WX5062;
wire WX606;
wire II19139;
wire WX2217;
wire II15565;
wire II22788;
wire WX7550;
wire WX1676;
wire WX155;
wire WX301;
wire WX11316;
wire II10124;
wire WX96;
wire II14677;
wire WX7861;
wire II14824;
wire WX2945;
wire WX8280;
wire WX10245;
wire WX6317;
wire WX2220;
wire II30634;
wire II18706;
wire II26306;
wire WX10983;
wire WX2031;
wire WX10105;
wire II22246;
wire WX8761;
wire WX2345;
wire WX10963;
wire II14156;
wire II14252;
wire II10820;
wire II6418;
wire WX5038;
wire II2400;
wire WX5033;
wire WX10282;
wire WX9099;
wire II14112;
wire II18264;
wire II30812;
wire WX88;
wire II18761;
wire WX9347;
wire II22371;
wire WX5034;
wire WX2260;
wire II18984;
wire II10449;
wire II18474;
wire II2145;
wire WX4409;
wire WX10441;
wire II10788;
wire WX4533;
wire WX3655;
wire WX476;
wire II14128;
wire WX1101;
wire II26893;
wire WX6981;
wire WX7476;
wire WX7728;
wire WX1441;
wire WX8648;
wire WX4329;
wire II14497;
wire WX7082;
wire WX9399;
wire II6396;
wire II23404;
wire II30479;
wire WX3013;
wire WX2095;
wire WX6255;
wire II14423;
wire WX1114;
wire WX8383;
wire WX10684;
wire II30614;
wire WX10699;
wire WX2486;
wire WX1888;
wire II3627;
wire WX4885;
wire II18249;
wire WX1864;
wire WX3775;
wire II34650;
wire WX5400;
wire II7187;
wire II18103;
wire WX9510;
wire WX8572;
wire WX5292;
wire II30797;
wire WX11247;
wire WX3675;
wire II26389;
wire II14669;
wire II35633;
wire WX6512;
wire II30465;
wire WX6734;
wire WX586;
wire WX5256;
wire WX11417;
wire II7652;
wire WX3202;
wire WX11064;
wire WX5850;
wire WX10533;
wire WX6149;
wire WX3112;
wire II31549;
wire WX8726;
wire WX11260;
wire WX10797;
wire II35659;
wire WX5773;
wire WX9973;
wire II18542;
wire WX1601;
wire WX10521;
wire II14973;
wire WX6899;
wire II31438;
wire WX4717;
wire II34478;
wire WX8264;
wire II2036;
wire II18017;
wire WX6784;
wire WX8456;
wire WX9457;
wire II14857;
wire WX9140;
wire WX9659;
wire II15663;
wire WX4755;
wire WX9664;
wire WX10756;
wire II6320;
wire WX10738;
wire WX1251;
wire WX10749;
wire WX939;
wire WX5862;
wire WX9779;
wire II3682;
wire II10231;
wire II18265;
wire II18241;
wire WX3669;
wire WX8907;
wire WX1266;
wire WX10735;
wire WX10373;
wire II27083;
wire WX8724;
wire WX1221;
wire II22416;
wire II18661;
wire WX3983;
wire WX8331;
wire II19507;
wire II15132;
wire II14903;
wire WX218;
wire WX4227;
wire WX8536;
wire II18063;
wire WX1228;
wire WX4243;
wire II34841;
wire II6304;
wire WX4047;
wire II15263;
wire II2407;
wire WX11371;
wire II22719;
wire II34679;
wire II6968;
wire WX11122;
wire WX3154;
wire II18025;
wire II2764;
wire WX3164;
wire WX9107;
wire WX1002;
wire WX3404;
wire WX10416;
wire WX970;
wire WX7934;
wire II18768;
wire WX9124;
wire WX1009;
wire WX7373;
wire WX796;
wire II26336;
wire WX5565;
wire WX5718;
wire II34882;
wire II30526;
wire WX9378;
wire WX5616;
wire II6946;
wire II18744;
wire II22542;
wire WX8922;
wire WX676;
wire II22151;
wire WX708;
wire WX9879;
wire WX11022;
wire WX4040;
wire II11207;
wire WX3344;
wire WX2348;
wire II22108;
wire II3300;
wire WX2199;
wire WX3059;
wire WX11044;
wire WX8183;
wire II26934;
wire WX530;
wire II18970;
wire WX720;
wire WX10349;
wire II34029;
wire II11567;
wire II31088;
wire II22237;
wire II31245;
wire WX5680;
wire WX1474;
wire WX3130;
wire II23430;
wire II6767;
wire II22693;
wire WX3945;
wire WX9649;
wire II34997;
wire WX8886;
wire II19662;
wire WX8580;
wire WX1718;
wire II6783;
wire WX554;
wire II10255;
wire II3494;
wire WX6359;
wire WX9642;
wire WX6020;
wire II10935;
wire WX11338;
wire WX7275;
wire WX512;
wire WX10506;
wire WX11485;
wire WX5335;
wire WX135;
wire II6040;
wire WX5016;
wire WX7175;
wire WX7638;
wire II31542;
wire WX1563;
wire II18203;
wire II30133;
wire WX9486;
wire WX5393;
wire II30766;
wire II14032;
wire II10549;
wire WX452;
wire II14345;
wire WX6664;
wire WX6564;
wire WX7564;
wire WX2918;
wire II6744;
wire WX1358;
wire II11155;
wire WX5299;
wire WX4306;
wire II6007;
wire II14451;
wire WX611;
wire WX461;
wire WX7309;
wire II11694;
wire WX6611;
wire II31747;
wire WX3034;
wire II14160;
wire II14297;
wire WX4787;
wire II2941;
wire WX8554;
wire II19632;
wire WX2696;
wire II7708;
wire II34354;
wire WX8925;
wire WX1086;
wire II34789;
wire WX10084;
wire WX9207;
wire WX6945;
wire II2545;
wire WX7491;
wire II19598;
wire WX1453;
wire II34338;
wire II3471;
wire WX3516;
wire WX3746;
wire II11546;
wire WX8992;
wire II3612;
wire WX2632;
wire II2175;
wire II35750;
wire WX5527;
wire II18125;
wire WX5696;
wire WX2885;
wire II22843;
wire WX2051;
wire WX8999;
wire II6450;
wire II14366;
wire WX1462;
wire WX10518;
wire WX7656;
wire II34246;
wire II15615;
wire WX9365;
wire II6518;
wire WX4982;
wire WX7682;
wire II26484;
wire II18334;
wire II15290;
wire WX8867;
wire WX8315;
wire II26382;
wire WX4587;
wire WX10221;
wire WX8362;
wire WX10673;
wire WX1436;
wire WX4092;
wire WX2439;
wire II22097;
wire WX9921;
wire WX8816;
wire WX11330;
wire II22564;
wire WX8751;
wire WX5600;
wire WX5357;
wire WX202;
wire WX11451;
wire II30371;
wire II26073;
wire WX1469;
wire WX9686;
wire II34533;
wire WX6689;
wire II10578;
wire WX1365;
wire II11638;
wire II30495;
wire WX8628;
wire WX2714;
wire WX6330;
wire WX106;
wire II30557;
wire WX10190;
wire WX9225;
wire WX2733;
wire II6319;
wire WX900;
wire WX4847;
wire WX736;
wire WX7123;
wire WX1908;
wire WX9046;
wire WX7503;
wire II18962;
wire WX10186;
wire WX1534;
wire WX7343;
wire II10215;
wire II23170;
wire WX10890;
wire II14621;
wire WX3466;
wire II22440;
wire WX4430;
wire WX8333;
wire WX3558;
wire WX6155;
wire II6636;
wire WX3223;
wire WX2793;
wire WX6602;
wire WX4196;
wire II7397;
wire II26831;
wire WX400;
wire WX7878;
wire II7449;
wire II19463;
wire II15394;
wire II22805;
wire WX1738;
wire WX10893;
wire II14189;
wire WX2519;
wire II6088;
wire WX7909;
wire WX1280;
wire II26764;
wire WX1302;
wire II10495;
wire WX5352;
wire II30938;
wire II14484;
wire II26454;
wire WX5543;
wire II2315;
wire II23561;
wire WX7875;
wire WX8317;
wire II2724;
wire WX11547;
wire WX4860;
wire II11678;
wire WX8783;
wire WX10924;
wire II27684;
wire WX4360;
wire WX7777;
wire II30875;
wire II15685;
wire WX6590;
wire WX10403;
wire II2017;
wire II23209;
wire WX4259;
wire II26599;
wire WX4017;
wire WX10746;
wire WX8566;
wire WX9985;
wire WX7513;
wire WX7091;
wire II10416;
wire WX5628;
wire II7583;
wire II2671;
wire WX8200;
wire II6444;
wire II23441;
wire II22470;
wire II2244;
wire II7226;
wire WX7401;
wire WX10420;
wire II10193;
wire WX10147;
wire WX10838;
wire WX4379;
wire WX11589;
wire WX1760;
wire II31565;
wire II10130;
wire II34104;
wire WX3142;
wire WX1904;
wire WX440;
wire WX2512;
wire II27318;
wire WX10363;
wire II26686;
wire WX10780;
wire WX9082;
wire WX3965;
wire WX2463;
wire II34429;
wire WX7453;
wire WX1038;
wire II15551;
wire II26213;
wire WX304;
wire II34587;
wire WX10886;
wire WX284;
wire II6094;
wire II22945;
wire WX10526;
wire WX10947;
wire II22570;
wire WX7053;
wire WX506;
wire II19647;
wire WX9393;
wire WX3850;
wire WX8436;
wire WX5374;
wire WX8889;
wire II14516;
wire WX2547;
wire WX5237;
wire WX9456;
wire WX10568;
wire II7632;
wire II10905;
wire WX6586;
wire WX10155;
wire II35583;
wire II11589;
wire WX2493;
wire II14625;
wire WX4088;
wire II19113;
wire II18599;
wire WX5247;
wire WX7560;
wire WX6123;
wire II22074;
wire WX1853;
wire WX1183;
wire WX2127;
wire WX5213;
wire WX10646;
wire II30923;
wire WX7399;
wire II27728;
wire WX4319;
wire WX1577;
wire WX8787;
wire II3247;
wire II34634;
wire WX967;
wire II30783;
wire WX638;
wire WX1925;
wire II2957;
wire WX1635;
wire WX2295;
wire WX437;
wire II10067;
wire WX4249;
wire II31374;
wire II6404;
wire WX8216;
wire WX6951;
wire WX9307;
wire II10045;
wire WX3392;
wire II10803;
wire WX9130;
wire II30123;
wire WX6884;
wire WX1951;
wire II18784;
wire WX11108;
wire II10867;
wire II30257;
wire II34956;
wire II30967;
wire WX1513;
wire II22755;
wire WX11325;
wire WX7525;
wire II6057;
wire II3515;
wire II3703;
wire WX7694;
wire II22208;
wire II30038;
wire WX2237;
wire WX1349;
wire WX6823;
wire WX2278;
wire II26871;
wire II19163;
wire WX9801;
wire WX10854;
wire II34229;
wire WX2753;
wire II15500;
wire II26878;
wire WX6934;
wire II22027;
wire WX10844;
wire II10300;
wire WX6545;
wire WX9963;
wire II14570;
wire II15484;
wire WX6068;
wire WX7847;
wire WX7378;
wire II31570;
wire WX1665;
wire WX11572;
wire II10455;
wire II31349;
wire WX7379;
wire WX10427;
wire WX8054;
wire II11595;
wire WX7966;
wire II30752;
wire WX9230;
wire WX3348;
wire WX10704;
wire WX2655;
wire WX8194;
wire II26206;
wire WX3971;
wire WX4465;
wire II26956;
wire II3620;
wire WX6536;
wire II18551;
wire WX1783;
wire II6621;
wire WX10592;
wire WX1632;
wire II14590;
wire WX410;
wire WX3045;
wire WX6432;
wire WX8090;
wire WX10967;
wire WX6909;
wire II34138;
wire WX8598;
wire WX7602;
wire WX10801;
wire WX11034;
wire WX2927;
wire II18681;
wire II34298;
wire WX4842;
wire II19306;
wire WX2858;
wire II14637;
wire II18428;
wire II6611;
wire II3377;
wire WX4010;
wire II19098;
wire WX2677;
wire II34439;
wire WX5788;
wire II34649;
wire WX5269;
wire II6876;
wire II30101;
wire WX6787;
wire II2834;
wire II2733;
wire II3677;
wire II35144;
wire WX5106;
wire WX6298;
wire WX8209;
wire WX9268;
wire WX1083;
wire WX5203;
wire II34897;
wire WX11010;
wire WX5573;
wire WX5368;
wire II3091;
wire WX1098;
wire WX6965;
wire II26089;
wire WX3676;
wire II19497;
wire WX6264;
wire WX8103;
wire II18590;
wire II23596;
wire II35327;
wire WX8402;
wire II22756;
wire II30573;
wire II6883;
wire WX4535;
wire II11246;
wire WX1329;
wire WX9591;
wire WX4928;
wire II26467;
wire WX3660;
wire WX1671;
wire WX10208;
wire WX2868;
wire WX5429;
wire II10542;
wire II27238;
wire WX2306;
wire II6565;
wire II14560;
wire WX2784;
wire II11465;
wire WX2861;
wire WX760;
wire WX4170;
wire II35723;
wire WX11498;
wire WX5672;
wire II34863;
wire WX8714;
wire WX4875;
wire WX9638;
wire WX10268;
wire II22664;
wire WX524;
wire WX5324;
wire II6257;
wire II27175;
wire II2687;
wire WX4220;
wire WX6189;
wire WX319;
wire II26577;
wire WX10030;
wire II14004;
wire II22972;
wire II6294;
wire WX6324;
wire WX5658;
wire WX10165;
wire WX9831;
wire WX10070;
wire II14911;
wire II6015;
wire II23468;
wire II14180;
wire WX4486;
wire WX6286;
wire WX2103;
wire II15699;
wire II22386;
wire WX1626;
wire WX6743;
wire WX5066;
wire II15537;
wire WX11518;
wire WX4168;
wire WX4056;
wire II23707;
wire WX9190;
wire WX5884;
wire WX2662;
wire WX7145;
wire II18357;
wire WX8399;
wire WX10261;
wire II14165;
wire II26530;
wire WX3230;
wire II26326;
wire WX8757;
wire WX10413;
wire WX8274;
wire WX10246;
wire WX406;
wire WX2372;
wire II19527;
wire WX3788;
wire WX4128;
wire WX5584;
wire WX9717;
wire II2299;
wire WX9449;
wire WX4179;
wire II27502;
wire WX9516;
wire II2190;
wire WX5720;
wire II26569;
wire WX1608;
wire WX6865;
wire WX4437;
wire WX365;
wire II26562;
wire WX3374;
wire II35248;
wire WX9469;
wire II11309;
wire II30844;
wire II27622;
wire II34727;
wire II6109;
wire WX7109;
wire II35430;
wire WX3757;
wire WX1024;
wire II30056;
wire II3197;
wire WX3102;
wire WX7613;
wire WX2432;
wire WX5458;
wire WX11523;
wire II31703;
wire WX3210;
wire WX2827;
wire WX10562;
wire II7646;
wire WX3779;
wire WX92;
wire II19541;
wire WX7763;
wire WX2499;
wire II22269;
wire WX3651;
wire II22618;
wire II22611;
wire WX1949;
wire WX3923;
wire WX4496;
wire II34640;
wire WX6836;
wire II6466;
wire II10774;
wire WX7589;
wire WX5789;
wire II27226;
wire WX10944;
wire WX2440;
wire II22858;
wire WX2468;
wire II18828;
wire WX5386;
wire WX9203;
wire WX582;
wire WX9977;
wire II23527;
wire WX4125;
wire II2632;
wire WX11437;
wire WX5220;
wire II10663;
wire WX7432;
wire WX1200;
wire WX194;
wire WX5415;
wire WX7534;
wire II6172;
wire WX10582;
wire WX5177;
wire WX10823;
wire WX10607;
wire II34322;
wire WX11341;
wire II22414;
wire WX10933;
wire WX3517;
wire WX960;
wire WX7094;
wire WX5131;
wire WX573;
wire II22167;
wire II22456;
wire II6759;
wire WX6180;
wire II31413;
wire WX10717;
wire WX8874;
wire WX5532;
wire II35235;
wire WX6278;
wire WX3709;
wire II6100;
wire WX1742;
wire II22997;
wire II31656;
wire WX55;
wire WX299;
wire WX10024;
wire II7591;
wire WX6220;
wire WX2065;
wire WX9247;
wire II34277;
wire WX5730;
wire WX9151;
wire II23416;
wire WX2047;
wire WX3698;
wire WX8125;
wire WX11602;
wire WX3766;
wire WX72;
wire WX6501;
wire WX4163;
wire WX4083;
wire WX8959;
wire WX5539;
wire WX494;
wire WX9244;
wire WX3898;
wire WX1292;
wire WX5221;
wire II22409;
wire WX6548;
wire WX8173;
wire WX8492;
wire WX10626;
wire WX1937;
wire II22779;
wire WX2396;
wire WX7644;
wire WX4958;
wire II23391;
wire WX6458;
wire WX7916;
wire WX10353;
wire II15366;
wire WX151;
wire WX4790;
wire II3210;
wire WX5762;
wire WX269;
wire WX7297;
wire WX3646;
wire II7645;
wire II3536;
wire WX10768;
wire WX7426;
wire WX3168;
wire WX7049;
wire WX9787;
wire WX6676;
wire WX1127;
wire II26661;
wire II6239;
wire WX1356;
wire II22035;
wire WX8857;
wire WX9749;
wire II22603;
wire WX7557;
wire II31231;
wire II26514;
wire II26095;
wire II34702;
wire WX10694;
wire II34657;
wire II11192;
wire II2568;
wire WX11530;
wire WX6171;
wire WX5218;
wire II6024;
wire II11374;
wire II11310;
wire WX11082;
wire WX1926;
wire WX9295;
wire WX3118;
wire II15594;
wire WX6556;
wire WX8989;
wire WX10664;
wire WX6372;
wire WX5936;
wire WX4699;
wire II26414;
wire WX2554;
wire WX217;
wire WX9275;
wire WX11466;
wire II35646;
wire II26949;
wire WX11363;
wire II26652;
wire WX11537;
wire WX2789;
wire II18466;
wire WX9767;
wire II26188;
wire WX9318;
wire WX10712;
wire WX2532;
wire WX10982;
wire WX8947;
wire II14218;
wire WX9551;
wire WX11368;
wire WX6283;
wire II11062;
wire WX4353;
wire II18899;
wire WX6806;
wire WX2313;
wire II3429;
wire II34910;
wire WX11393;
wire II26730;
wire II14056;
wire II34361;
wire II3079;
wire II18991;
wire WX4020;
wire II31361;
wire II18985;
wire WX6794;
wire II22425;
wire II10688;
wire WX4615;
wire WX5490;
wire II15068;
wire WX5051;
wire II15121;
wire WX7860;
wire WX3590;
wire WX1660;
wire WX2351;
wire WX4931;
wire WX4520;
wire II26846;
wire WX2763;
wire II10641;
wire WX1552;
wire II14718;
wire II14205;
wire II27474;
wire II26919;
wire II15649;
wire II14191;
wire II27658;
wire II18210;
wire WX7410;
wire II11680;
wire WX8115;
wire WX10017;
wire II30366;
wire WX7385;
wire WX3794;
wire WX4119;
wire II10260;
wire WX5023;
wire II7202;
wire II2445;
wire WX2009;
wire II30224;
wire WX8329;
wire II15515;
wire WX7953;
wire II6150;
wire WX4559;
wire II23287;
wire II14477;
wire WX682;
wire WX609;
wire WX9002;
wire WX10236;
wire WX5748;
wire WX10174;
wire WX6572;
wire II18434;
wire WX9380;
wire II26515;
wire WX10900;
wire WX7793;
wire II2506;
wire WX3501;
wire II3171;
wire WX6898;
wire II34315;
wire WX8972;
wire WX3933;
wire II7694;
wire II15210;
wire WX5666;
wire WX1595;
wire WX8343;
wire II10378;
wire II6847;
wire WX4320;
wire WX10630;
wire II7343;
wire II10837;
wire WX4027;
wire WX8802;
wire II30195;
wire WX7058;
wire II2172;
wire WX457;
wire WX8416;
wire II31621;
wire WX7384;
wire WX2684;
wire WX127;
wire WX79;
wire WX376;
wire II15093;
wire II26202;
wire WX2481;
wire II19711;
wire WX7471;
wire WX5128;
wire WX1181;
wire WX9619;
wire II3654;
wire WX8689;
wire WX2890;
wire WX2838;
wire WX5611;
wire WX7977;
wire WX10653;
wire WX3244;
wire II2491;
wire II34903;
wire II34432;
wire WX8254;
wire WX3686;
wire WX3624;
wire WX167;
wire II3053;
wire II14358;
wire WX3926;
wire WX5767;
wire WX10971;
wire II18573;
wire WX4458;
wire WX2323;
wire WX9663;
wire WX1079;
wire II10043;
wire II34445;
wire WX4490;
wire II23674;
wire II31335;
wire II30303;
wire II14399;
wire WX8088;
wire WX6861;
wire II15080;
wire II18286;
wire WX6178;
wire II2121;
wire II6813;
wire II30448;
wire WX6139;
wire II35605;
wire WX7807;
wire WX7205;
wire WX9329;
wire WX8478;
wire WX6382;
wire WX47;
wire II30683;
wire WX4100;
wire WX3523;
wire WX6435;
wire WX9417;
wire WX10579;
wire II34517;
wire WX4916;
wire II10006;
wire II31270;
wire II27422;
wire WX10474;
wire WX6076;
wire II30651;
wire WX8040;
wire WX6259;
wire WX4741;
wire WX2749;
wire II34564;
wire WX10029;
wire WX11058;
wire WX253;
wire WX8750;
wire WX9111;
wire WX4248;
wire WX9116;
wire II35744;
wire WX118;
wire II23653;
wire II6000;
wire II26376;
wire WX2634;
wire WX11198;
wire WX6070;
wire WX2167;
wire II23554;
wire WX5046;
wire WX3137;
wire II31375;
wire WX9815;
wire WX1589;
wire WX1914;
wire II18418;
wire WX11402;
wire WX10150;
wire WX4037;
wire II2041;
wire II22433;
wire II11167;
wire WX7541;
wire II10928;
wire WX4064;
wire II30487;
wire WX1706;
wire WX5363;
wire II35519;
wire WX907;
wire II10588;
wire WX5115;
wire II14483;
wire II30480;
wire WX8081;
wire II22632;
wire WX2332;
wire II11103;
wire II26110;
wire II15238;
wire II31400;
wire II26802;
wire II10564;
wire WX5700;
wire WX9487;
wire WX8699;
wire WX6657;
wire II3697;
wire WX4271;
wire II15224;
wire II6775;
wire II23562;
wire II26491;
wire WX6707;
wire WX2818;
wire II10105;
wire II18751;
wire WX2955;
wire II27147;
wire WX2777;
wire WX3551;
wire WX10012;
wire WX4995;
wire II34967;
wire WX4151;
wire II18272;
wire WX3544;
wire WX8544;
wire WX9933;
wire II26809;
wire II10185;
wire II2322;
wire II34610;
wire WX2994;
wire WX7947;
wire II34074;
wire II22812;
wire WX6392;
wire WX5344;
wire II6348;
wire WX3830;
wire WX40;
wire WX1858;
wire WX2027;
wire II31534;
wire II3578;
wire WX3813;
wire WX5314;
wire WX3565;
wire WX2701;
wire II10038;
wire II14671;
wire WX2770;
wire II6906;
wire II30140;
wire II34848;
wire II18037;
wire II23299;
wire II14406;
wire II19204;
wire WX1559;
wire WX7983;
wire WX6551;
wire WX1339;
wire WX6329;
wire II6909;
wire II22332;
wire WX5467;
wire WX567;
wire WX9050;
wire II11554;
wire WX7715;
wire WX8917;
wire WX1617;
wire WX7067;
wire WX4252;
wire WX594;
wire WX1775;
wire II2569;
wire WX11462;
wire WX4067;
wire II26275;
wire II35456;
wire II22665;
wire II2935;
wire II30372;
wire WX9604;
wire II6684;
wire WX1402;
wire II27581;
wire II27594;
wire II34495;
wire WX8522;
wire WX2730;
wire II27517;
wire II10819;
wire WX548;
wire WX4808;
wire II10248;
wire WX824;
wire WX9525;
wire II18301;
wire II30952;
wire II15184;
wire WX11112;
wire WX9072;
wire II11687;
wire II18503;
wire WX7486;
wire WX8324;
wire WX5441;
wire WX8358;
wire II6157;
wire II34880;
wire WX10238;
wire II2438;
wire WX10118;
wire WX1647;
wire WX4208;
wire WX6650;
wire II19548;
wire WX258;
wire II14523;
wire II23364;
wire WX201;
wire WX3488;
wire II22146;
wire WX187;
wire WX5383;
wire WX7147;
wire WX6918;
wire II26080;
wire WX3063;
wire II6164;
wire II7533;
wire WX1709;
wire WX10479;
wire WX3549;
wire WX5175;
wire II30031;
wire II3456;
wire WX973;
wire II26126;
wire WX11579;
wire WX5812;
wire WX4837;
wire WX9226;
wire II2771;
wire WX1332;
wire WX6342;
wire WX8304;
wire II14986;
wire WX2907;
wire II14738;
wire II7410;
wire WX3084;
wire II14614;
wire II18224;
wire WX1508;
wire II26399;
wire II14445;
wire WX8824;
wire II34802;
wire WX7616;
wire WX4977;
wire II34244;
wire II26755;
wire WX193;
wire II6583;
wire WX6166;
wire WX11555;
wire II6133;
wire WX10256;
wire II11573;
wire WX4005;
wire WX10936;
wire WX2298;
wire II15552;
wire II18318;
wire WX8769;
wire II22011;
wire WX4286;
wire WX7827;
wire WX9697;
wire II31579;
wire WX7531;
wire WX2587;
wire WX11166;
wire II14942;
wire II23157;
wire II11624;
wire WX3959;
wire II14864;
wire WX3576;
wire WX7185;
wire II18311;
wire WX724;
wire II2739;
wire WX1035;
wire WX2359;
wire WX10068;
wire II31717;
wire WX8981;
wire WX161;
wire WX10341;
wire WX7680;
wire II15198;
wire WX10516;
wire WX6723;
wire WX5082;
wire WX7882;
wire II3571;
wire WX3700;
wire WX5477;
wire II26900;
wire WX4978;
wire WX10773;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX485 <= 0;
  else
    WX485 <= WX484;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX487 <= 0;
  else
    WX487 <= WX486;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX489 <= 0;
  else
    WX489 <= WX488;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX491 <= 0;
  else
    WX491 <= WX490;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX493 <= 0;
  else
    WX493 <= WX492;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX495 <= 0;
  else
    WX495 <= WX494;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX497 <= 0;
  else
    WX497 <= WX496;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX499 <= 0;
  else
    WX499 <= WX498;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX501 <= 0;
  else
    WX501 <= WX500;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX503 <= 0;
  else
    WX503 <= WX502;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX505 <= 0;
  else
    WX505 <= WX504;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX507 <= 0;
  else
    WX507 <= WX506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX509 <= 0;
  else
    WX509 <= WX508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX511 <= 0;
  else
    WX511 <= WX510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX513 <= 0;
  else
    WX513 <= WX512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX515 <= 0;
  else
    WX515 <= WX514;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX517 <= 0;
  else
    WX517 <= WX516;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX519 <= 0;
  else
    WX519 <= WX518;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX521 <= 0;
  else
    WX521 <= WX520;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX523 <= 0;
  else
    WX523 <= WX522;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX525 <= 0;
  else
    WX525 <= WX524;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX527 <= 0;
  else
    WX527 <= WX526;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX529 <= 0;
  else
    WX529 <= WX528;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX531 <= 0;
  else
    WX531 <= WX530;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX533 <= 0;
  else
    WX533 <= WX532;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX535 <= 0;
  else
    WX535 <= WX534;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX537 <= 0;
  else
    WX537 <= WX536;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX539 <= 0;
  else
    WX539 <= WX538;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX541 <= 0;
  else
    WX541 <= WX540;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX543 <= 0;
  else
    WX543 <= WX542;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX545 <= 0;
  else
    WX545 <= WX544;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX547 <= 0;
  else
    WX547 <= WX546;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX645 <= 0;
  else
    WX645 <= WX644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX647 <= 0;
  else
    WX647 <= WX646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX649 <= 0;
  else
    WX649 <= WX648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX651 <= 0;
  else
    WX651 <= WX650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX653 <= 0;
  else
    WX653 <= WX652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX655 <= 0;
  else
    WX655 <= WX654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX657 <= 0;
  else
    WX657 <= WX656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX659 <= 0;
  else
    WX659 <= WX658;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX661 <= 0;
  else
    WX661 <= WX660;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX663 <= 0;
  else
    WX663 <= WX662;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX665 <= 0;
  else
    WX665 <= WX664;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX667 <= 0;
  else
    WX667 <= WX666;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX669 <= 0;
  else
    WX669 <= WX668;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX671 <= 0;
  else
    WX671 <= WX670;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX673 <= 0;
  else
    WX673 <= WX672;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX675 <= 0;
  else
    WX675 <= WX674;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX677 <= 0;
  else
    WX677 <= WX676;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX679 <= 0;
  else
    WX679 <= WX678;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX681 <= 0;
  else
    WX681 <= WX680;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX683 <= 0;
  else
    WX683 <= WX682;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX685 <= 0;
  else
    WX685 <= WX684;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX687 <= 0;
  else
    WX687 <= WX686;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX689 <= 0;
  else
    WX689 <= WX688;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX691 <= 0;
  else
    WX691 <= WX690;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX693 <= 0;
  else
    WX693 <= WX692;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX695 <= 0;
  else
    WX695 <= WX694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX697 <= 0;
  else
    WX697 <= WX696;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX699 <= 0;
  else
    WX699 <= WX698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX701 <= 0;
  else
    WX701 <= WX700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX703 <= 0;
  else
    WX703 <= WX702;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX705 <= 0;
  else
    WX705 <= WX704;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX707 <= 0;
  else
    WX707 <= WX706;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX709 <= 0;
  else
    WX709 <= WX708;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX711 <= 0;
  else
    WX711 <= WX710;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX713 <= 0;
  else
    WX713 <= WX712;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX715 <= 0;
  else
    WX715 <= WX714;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX717 <= 0;
  else
    WX717 <= WX716;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX719 <= 0;
  else
    WX719 <= WX718;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX721 <= 0;
  else
    WX721 <= WX720;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX723 <= 0;
  else
    WX723 <= WX722;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX725 <= 0;
  else
    WX725 <= WX724;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX727 <= 0;
  else
    WX727 <= WX726;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX729 <= 0;
  else
    WX729 <= WX728;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX731 <= 0;
  else
    WX731 <= WX730;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX733 <= 0;
  else
    WX733 <= WX732;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX735 <= 0;
  else
    WX735 <= WX734;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX737 <= 0;
  else
    WX737 <= WX736;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX739 <= 0;
  else
    WX739 <= WX738;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX741 <= 0;
  else
    WX741 <= WX740;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX743 <= 0;
  else
    WX743 <= WX742;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX745 <= 0;
  else
    WX745 <= WX744;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX747 <= 0;
  else
    WX747 <= WX746;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX749 <= 0;
  else
    WX749 <= WX748;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX751 <= 0;
  else
    WX751 <= WX750;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX753 <= 0;
  else
    WX753 <= WX752;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX755 <= 0;
  else
    WX755 <= WX754;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX757 <= 0;
  else
    WX757 <= WX756;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX759 <= 0;
  else
    WX759 <= WX758;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX761 <= 0;
  else
    WX761 <= WX760;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX763 <= 0;
  else
    WX763 <= WX762;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX765 <= 0;
  else
    WX765 <= WX764;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX767 <= 0;
  else
    WX767 <= WX766;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX769 <= 0;
  else
    WX769 <= WX768;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX771 <= 0;
  else
    WX771 <= WX770;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX773 <= 0;
  else
    WX773 <= WX772;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX775 <= 0;
  else
    WX775 <= WX774;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX777 <= 0;
  else
    WX777 <= WX776;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX779 <= 0;
  else
    WX779 <= WX778;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX781 <= 0;
  else
    WX781 <= WX780;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX783 <= 0;
  else
    WX783 <= WX782;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX785 <= 0;
  else
    WX785 <= WX784;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX787 <= 0;
  else
    WX787 <= WX786;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX789 <= 0;
  else
    WX789 <= WX788;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX791 <= 0;
  else
    WX791 <= WX790;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX793 <= 0;
  else
    WX793 <= WX792;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX795 <= 0;
  else
    WX795 <= WX794;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX797 <= 0;
  else
    WX797 <= WX796;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX799 <= 0;
  else
    WX799 <= WX798;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX801 <= 0;
  else
    WX801 <= WX800;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX803 <= 0;
  else
    WX803 <= WX802;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX805 <= 0;
  else
    WX805 <= WX804;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX807 <= 0;
  else
    WX807 <= WX806;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX809 <= 0;
  else
    WX809 <= WX808;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX811 <= 0;
  else
    WX811 <= WX810;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX813 <= 0;
  else
    WX813 <= WX812;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX815 <= 0;
  else
    WX815 <= WX814;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX817 <= 0;
  else
    WX817 <= WX816;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX819 <= 0;
  else
    WX819 <= WX818;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX821 <= 0;
  else
    WX821 <= WX820;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX823 <= 0;
  else
    WX823 <= WX822;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX825 <= 0;
  else
    WX825 <= WX824;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX827 <= 0;
  else
    WX827 <= WX826;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX829 <= 0;
  else
    WX829 <= WX828;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX831 <= 0;
  else
    WX831 <= WX830;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX833 <= 0;
  else
    WX833 <= WX832;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX835 <= 0;
  else
    WX835 <= WX834;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX837 <= 0;
  else
    WX837 <= WX836;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX839 <= 0;
  else
    WX839 <= WX838;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX841 <= 0;
  else
    WX841 <= WX840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX843 <= 0;
  else
    WX843 <= WX842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX845 <= 0;
  else
    WX845 <= WX844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX847 <= 0;
  else
    WX847 <= WX846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX849 <= 0;
  else
    WX849 <= WX848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX851 <= 0;
  else
    WX851 <= WX850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX853 <= 0;
  else
    WX853 <= WX852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX855 <= 0;
  else
    WX855 <= WX854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX857 <= 0;
  else
    WX857 <= WX856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX859 <= 0;
  else
    WX859 <= WX858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX861 <= 0;
  else
    WX861 <= WX860;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX863 <= 0;
  else
    WX863 <= WX862;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX865 <= 0;
  else
    WX865 <= WX864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX867 <= 0;
  else
    WX867 <= WX866;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX869 <= 0;
  else
    WX869 <= WX868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX871 <= 0;
  else
    WX871 <= WX870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX873 <= 0;
  else
    WX873 <= WX872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX875 <= 0;
  else
    WX875 <= WX874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX877 <= 0;
  else
    WX877 <= WX876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX879 <= 0;
  else
    WX879 <= WX878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX881 <= 0;
  else
    WX881 <= WX880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX883 <= 0;
  else
    WX883 <= WX882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX885 <= 0;
  else
    WX885 <= WX884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX887 <= 0;
  else
    WX887 <= WX886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX889 <= 0;
  else
    WX889 <= WX888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX891 <= 0;
  else
    WX891 <= WX890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX893 <= 0;
  else
    WX893 <= WX892;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX895 <= 0;
  else
    WX895 <= WX894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX897 <= 0;
  else
    WX897 <= WX896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX899 <= 0;
  else
    WX899 <= WX898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2077_ <= 0;
  else
    _2077_ <= WX1264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2078_ <= 0;
  else
    _2078_ <= WX1266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2079_ <= 0;
  else
    _2079_ <= WX1268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2080_ <= 0;
  else
    _2080_ <= WX1270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2081_ <= 0;
  else
    _2081_ <= WX1272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2082_ <= 0;
  else
    _2082_ <= WX1274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2083_ <= 0;
  else
    _2083_ <= WX1276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2084_ <= 0;
  else
    _2084_ <= WX1278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2085_ <= 0;
  else
    _2085_ <= WX1280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2086_ <= 0;
  else
    _2086_ <= WX1282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2087_ <= 0;
  else
    _2087_ <= WX1284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2088_ <= 0;
  else
    _2088_ <= WX1286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2089_ <= 0;
  else
    _2089_ <= WX1288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2090_ <= 0;
  else
    _2090_ <= WX1290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2091_ <= 0;
  else
    _2091_ <= WX1292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2092_ <= 0;
  else
    _2092_ <= WX1294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2093_ <= 0;
  else
    _2093_ <= WX1296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2094_ <= 0;
  else
    _2094_ <= WX1298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2095_ <= 0;
  else
    _2095_ <= WX1300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2096_ <= 0;
  else
    _2096_ <= WX1302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2097_ <= 0;
  else
    _2097_ <= WX1304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2098_ <= 0;
  else
    _2098_ <= WX1306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2099_ <= 0;
  else
    _2099_ <= WX1308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2100_ <= 0;
  else
    _2100_ <= WX1310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2101_ <= 0;
  else
    _2101_ <= WX1312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2102_ <= 0;
  else
    _2102_ <= WX1314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2103_ <= 0;
  else
    _2103_ <= WX1316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2104_ <= 0;
  else
    _2104_ <= WX1318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2105_ <= 0;
  else
    _2105_ <= WX1320;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2106_ <= 0;
  else
    _2106_ <= WX1322;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2107_ <= 0;
  else
    _2107_ <= WX1324;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2108_ <= 0;
  else
    _2108_ <= WX1326;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1778 <= 0;
  else
    WX1778 <= WX1777;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1780 <= 0;
  else
    WX1780 <= WX1779;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1782 <= 0;
  else
    WX1782 <= WX1781;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1784 <= 0;
  else
    WX1784 <= WX1783;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1786 <= 0;
  else
    WX1786 <= WX1785;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1788 <= 0;
  else
    WX1788 <= WX1787;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1790 <= 0;
  else
    WX1790 <= WX1789;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1792 <= 0;
  else
    WX1792 <= WX1791;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1794 <= 0;
  else
    WX1794 <= WX1793;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1796 <= 0;
  else
    WX1796 <= WX1795;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1798 <= 0;
  else
    WX1798 <= WX1797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1800 <= 0;
  else
    WX1800 <= WX1799;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1802 <= 0;
  else
    WX1802 <= WX1801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1804 <= 0;
  else
    WX1804 <= WX1803;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1806 <= 0;
  else
    WX1806 <= WX1805;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1808 <= 0;
  else
    WX1808 <= WX1807;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1810 <= 0;
  else
    WX1810 <= WX1809;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1812 <= 0;
  else
    WX1812 <= WX1811;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1814 <= 0;
  else
    WX1814 <= WX1813;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1816 <= 0;
  else
    WX1816 <= WX1815;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1818 <= 0;
  else
    WX1818 <= WX1817;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1820 <= 0;
  else
    WX1820 <= WX1819;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1822 <= 0;
  else
    WX1822 <= WX1821;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1824 <= 0;
  else
    WX1824 <= WX1823;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1826 <= 0;
  else
    WX1826 <= WX1825;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1828 <= 0;
  else
    WX1828 <= WX1827;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1830 <= 0;
  else
    WX1830 <= WX1829;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1832 <= 0;
  else
    WX1832 <= WX1831;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1834 <= 0;
  else
    WX1834 <= WX1833;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1836 <= 0;
  else
    WX1836 <= WX1835;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1838 <= 0;
  else
    WX1838 <= WX1837;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1840 <= 0;
  else
    WX1840 <= WX1839;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1938 <= 0;
  else
    WX1938 <= WX1937;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1940 <= 0;
  else
    WX1940 <= WX1939;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1942 <= 0;
  else
    WX1942 <= WX1941;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1944 <= 0;
  else
    WX1944 <= WX1943;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1946 <= 0;
  else
    WX1946 <= WX1945;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1948 <= 0;
  else
    WX1948 <= WX1947;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1950 <= 0;
  else
    WX1950 <= WX1949;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1952 <= 0;
  else
    WX1952 <= WX1951;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1954 <= 0;
  else
    WX1954 <= WX1953;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1956 <= 0;
  else
    WX1956 <= WX1955;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1958 <= 0;
  else
    WX1958 <= WX1957;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1960 <= 0;
  else
    WX1960 <= WX1959;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1962 <= 0;
  else
    WX1962 <= WX1961;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1964 <= 0;
  else
    WX1964 <= WX1963;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1966 <= 0;
  else
    WX1966 <= WX1965;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1968 <= 0;
  else
    WX1968 <= WX1967;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1970 <= 0;
  else
    WX1970 <= WX1969;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1972 <= 0;
  else
    WX1972 <= WX1971;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1974 <= 0;
  else
    WX1974 <= WX1973;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1976 <= 0;
  else
    WX1976 <= WX1975;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1978 <= 0;
  else
    WX1978 <= WX1977;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1980 <= 0;
  else
    WX1980 <= WX1979;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1982 <= 0;
  else
    WX1982 <= WX1981;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1984 <= 0;
  else
    WX1984 <= WX1983;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1986 <= 0;
  else
    WX1986 <= WX1985;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1988 <= 0;
  else
    WX1988 <= WX1987;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1990 <= 0;
  else
    WX1990 <= WX1989;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1992 <= 0;
  else
    WX1992 <= WX1991;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1994 <= 0;
  else
    WX1994 <= WX1993;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1996 <= 0;
  else
    WX1996 <= WX1995;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX1998 <= 0;
  else
    WX1998 <= WX1997;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2000 <= 0;
  else
    WX2000 <= WX1999;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2002 <= 0;
  else
    WX2002 <= WX2001;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2004 <= 0;
  else
    WX2004 <= WX2003;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2006 <= 0;
  else
    WX2006 <= WX2005;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2008 <= 0;
  else
    WX2008 <= WX2007;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2010 <= 0;
  else
    WX2010 <= WX2009;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2012 <= 0;
  else
    WX2012 <= WX2011;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2014 <= 0;
  else
    WX2014 <= WX2013;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2016 <= 0;
  else
    WX2016 <= WX2015;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2018 <= 0;
  else
    WX2018 <= WX2017;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2020 <= 0;
  else
    WX2020 <= WX2019;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2022 <= 0;
  else
    WX2022 <= WX2021;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2024 <= 0;
  else
    WX2024 <= WX2023;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2026 <= 0;
  else
    WX2026 <= WX2025;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2028 <= 0;
  else
    WX2028 <= WX2027;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2030 <= 0;
  else
    WX2030 <= WX2029;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2032 <= 0;
  else
    WX2032 <= WX2031;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2034 <= 0;
  else
    WX2034 <= WX2033;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2036 <= 0;
  else
    WX2036 <= WX2035;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2038 <= 0;
  else
    WX2038 <= WX2037;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2040 <= 0;
  else
    WX2040 <= WX2039;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2042 <= 0;
  else
    WX2042 <= WX2041;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2044 <= 0;
  else
    WX2044 <= WX2043;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2046 <= 0;
  else
    WX2046 <= WX2045;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2048 <= 0;
  else
    WX2048 <= WX2047;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2050 <= 0;
  else
    WX2050 <= WX2049;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2052 <= 0;
  else
    WX2052 <= WX2051;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2054 <= 0;
  else
    WX2054 <= WX2053;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2056 <= 0;
  else
    WX2056 <= WX2055;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2058 <= 0;
  else
    WX2058 <= WX2057;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2060 <= 0;
  else
    WX2060 <= WX2059;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2062 <= 0;
  else
    WX2062 <= WX2061;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2064 <= 0;
  else
    WX2064 <= WX2063;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2066 <= 0;
  else
    WX2066 <= WX2065;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2068 <= 0;
  else
    WX2068 <= WX2067;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2070 <= 0;
  else
    WX2070 <= WX2069;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2072 <= 0;
  else
    WX2072 <= WX2071;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2074 <= 0;
  else
    WX2074 <= WX2073;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2076 <= 0;
  else
    WX2076 <= WX2075;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2078 <= 0;
  else
    WX2078 <= WX2077;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2080 <= 0;
  else
    WX2080 <= WX2079;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2082 <= 0;
  else
    WX2082 <= WX2081;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2084 <= 0;
  else
    WX2084 <= WX2083;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2086 <= 0;
  else
    WX2086 <= WX2085;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2088 <= 0;
  else
    WX2088 <= WX2087;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2090 <= 0;
  else
    WX2090 <= WX2089;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2092 <= 0;
  else
    WX2092 <= WX2091;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2094 <= 0;
  else
    WX2094 <= WX2093;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2096 <= 0;
  else
    WX2096 <= WX2095;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2098 <= 0;
  else
    WX2098 <= WX2097;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2100 <= 0;
  else
    WX2100 <= WX2099;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2102 <= 0;
  else
    WX2102 <= WX2101;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2104 <= 0;
  else
    WX2104 <= WX2103;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2106 <= 0;
  else
    WX2106 <= WX2105;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2108 <= 0;
  else
    WX2108 <= WX2107;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2110 <= 0;
  else
    WX2110 <= WX2109;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2112 <= 0;
  else
    WX2112 <= WX2111;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2114 <= 0;
  else
    WX2114 <= WX2113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2116 <= 0;
  else
    WX2116 <= WX2115;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2118 <= 0;
  else
    WX2118 <= WX2117;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2120 <= 0;
  else
    WX2120 <= WX2119;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2122 <= 0;
  else
    WX2122 <= WX2121;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2124 <= 0;
  else
    WX2124 <= WX2123;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2126 <= 0;
  else
    WX2126 <= WX2125;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2128 <= 0;
  else
    WX2128 <= WX2127;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2130 <= 0;
  else
    WX2130 <= WX2129;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2132 <= 0;
  else
    WX2132 <= WX2131;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2134 <= 0;
  else
    WX2134 <= WX2133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2136 <= 0;
  else
    WX2136 <= WX2135;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2138 <= 0;
  else
    WX2138 <= WX2137;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2140 <= 0;
  else
    WX2140 <= WX2139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2142 <= 0;
  else
    WX2142 <= WX2141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2144 <= 0;
  else
    WX2144 <= WX2143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2146 <= 0;
  else
    WX2146 <= WX2145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2148 <= 0;
  else
    WX2148 <= WX2147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2150 <= 0;
  else
    WX2150 <= WX2149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2152 <= 0;
  else
    WX2152 <= WX2151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2154 <= 0;
  else
    WX2154 <= WX2153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2156 <= 0;
  else
    WX2156 <= WX2155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2158 <= 0;
  else
    WX2158 <= WX2157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2160 <= 0;
  else
    WX2160 <= WX2159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2162 <= 0;
  else
    WX2162 <= WX2161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2164 <= 0;
  else
    WX2164 <= WX2163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2166 <= 0;
  else
    WX2166 <= WX2165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2168 <= 0;
  else
    WX2168 <= WX2167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2170 <= 0;
  else
    WX2170 <= WX2169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2172 <= 0;
  else
    WX2172 <= WX2171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2174 <= 0;
  else
    WX2174 <= WX2173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2176 <= 0;
  else
    WX2176 <= WX2175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2178 <= 0;
  else
    WX2178 <= WX2177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2180 <= 0;
  else
    WX2180 <= WX2179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2182 <= 0;
  else
    WX2182 <= WX2181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2184 <= 0;
  else
    WX2184 <= WX2183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2186 <= 0;
  else
    WX2186 <= WX2185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2188 <= 0;
  else
    WX2188 <= WX2187;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2190 <= 0;
  else
    WX2190 <= WX2189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX2192 <= 0;
  else
    WX2192 <= WX2191;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2109_ <= 0;
  else
    _2109_ <= WX2557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2110_ <= 0;
  else
    _2110_ <= WX2559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2111_ <= 0;
  else
    _2111_ <= WX2561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2112_ <= 0;
  else
    _2112_ <= WX2563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2113_ <= 0;
  else
    _2113_ <= WX2565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2114_ <= 0;
  else
    _2114_ <= WX2567;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2115_ <= 0;
  else
    _2115_ <= WX2569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2116_ <= 0;
  else
    _2116_ <= WX2571;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2117_ <= 0;
  else
    _2117_ <= WX2573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2118_ <= 0;
  else
    _2118_ <= WX2575;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2119_ <= 0;
  else
    _2119_ <= WX2577;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2120_ <= 0;
  else
    _2120_ <= WX2579;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2121_ <= 0;
  else
    _2121_ <= WX2581;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2122_ <= 0;
  else
    _2122_ <= WX2583;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2123_ <= 0;
  else
    _2123_ <= WX2585;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2124_ <= 0;
  else
    _2124_ <= WX2587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2125_ <= 0;
  else
    _2125_ <= WX2589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2126_ <= 0;
  else
    _2126_ <= WX2591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2127_ <= 0;
  else
    _2127_ <= WX2593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2128_ <= 0;
  else
    _2128_ <= WX2595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2129_ <= 0;
  else
    _2129_ <= WX2597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2130_ <= 0;
  else
    _2130_ <= WX2599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2131_ <= 0;
  else
    _2131_ <= WX2601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2132_ <= 0;
  else
    _2132_ <= WX2603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2133_ <= 0;
  else
    _2133_ <= WX2605;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2134_ <= 0;
  else
    _2134_ <= WX2607;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2135_ <= 0;
  else
    _2135_ <= WX2609;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2136_ <= 0;
  else
    _2136_ <= WX2611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2137_ <= 0;
  else
    _2137_ <= WX2613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2138_ <= 0;
  else
    _2138_ <= WX2615;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2139_ <= 0;
  else
    _2139_ <= WX2617;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2140_ <= 0;
  else
    _2140_ <= WX2619;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3071 <= 0;
  else
    WX3071 <= WX3070;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3073 <= 0;
  else
    WX3073 <= WX3072;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3075 <= 0;
  else
    WX3075 <= WX3074;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3077 <= 0;
  else
    WX3077 <= WX3076;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3079 <= 0;
  else
    WX3079 <= WX3078;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3081 <= 0;
  else
    WX3081 <= WX3080;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3083 <= 0;
  else
    WX3083 <= WX3082;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3085 <= 0;
  else
    WX3085 <= WX3084;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3087 <= 0;
  else
    WX3087 <= WX3086;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3089 <= 0;
  else
    WX3089 <= WX3088;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3091 <= 0;
  else
    WX3091 <= WX3090;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3093 <= 0;
  else
    WX3093 <= WX3092;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3095 <= 0;
  else
    WX3095 <= WX3094;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3097 <= 0;
  else
    WX3097 <= WX3096;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3099 <= 0;
  else
    WX3099 <= WX3098;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3101 <= 0;
  else
    WX3101 <= WX3100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3103 <= 0;
  else
    WX3103 <= WX3102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3105 <= 0;
  else
    WX3105 <= WX3104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3107 <= 0;
  else
    WX3107 <= WX3106;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3109 <= 0;
  else
    WX3109 <= WX3108;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3111 <= 0;
  else
    WX3111 <= WX3110;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3113 <= 0;
  else
    WX3113 <= WX3112;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3115 <= 0;
  else
    WX3115 <= WX3114;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3117 <= 0;
  else
    WX3117 <= WX3116;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3119 <= 0;
  else
    WX3119 <= WX3118;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3121 <= 0;
  else
    WX3121 <= WX3120;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3123 <= 0;
  else
    WX3123 <= WX3122;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3125 <= 0;
  else
    WX3125 <= WX3124;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3127 <= 0;
  else
    WX3127 <= WX3126;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3129 <= 0;
  else
    WX3129 <= WX3128;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3131 <= 0;
  else
    WX3131 <= WX3130;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3133 <= 0;
  else
    WX3133 <= WX3132;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3231 <= 0;
  else
    WX3231 <= WX3230;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3233 <= 0;
  else
    WX3233 <= WX3232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3235 <= 0;
  else
    WX3235 <= WX3234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3237 <= 0;
  else
    WX3237 <= WX3236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3239 <= 0;
  else
    WX3239 <= WX3238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3241 <= 0;
  else
    WX3241 <= WX3240;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3243 <= 0;
  else
    WX3243 <= WX3242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3245 <= 0;
  else
    WX3245 <= WX3244;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3247 <= 0;
  else
    WX3247 <= WX3246;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3249 <= 0;
  else
    WX3249 <= WX3248;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3251 <= 0;
  else
    WX3251 <= WX3250;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3253 <= 0;
  else
    WX3253 <= WX3252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3255 <= 0;
  else
    WX3255 <= WX3254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3257 <= 0;
  else
    WX3257 <= WX3256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3259 <= 0;
  else
    WX3259 <= WX3258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3261 <= 0;
  else
    WX3261 <= WX3260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3263 <= 0;
  else
    WX3263 <= WX3262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3265 <= 0;
  else
    WX3265 <= WX3264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3267 <= 0;
  else
    WX3267 <= WX3266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3269 <= 0;
  else
    WX3269 <= WX3268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3271 <= 0;
  else
    WX3271 <= WX3270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3273 <= 0;
  else
    WX3273 <= WX3272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3275 <= 0;
  else
    WX3275 <= WX3274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3277 <= 0;
  else
    WX3277 <= WX3276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3279 <= 0;
  else
    WX3279 <= WX3278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3281 <= 0;
  else
    WX3281 <= WX3280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3283 <= 0;
  else
    WX3283 <= WX3282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3285 <= 0;
  else
    WX3285 <= WX3284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3287 <= 0;
  else
    WX3287 <= WX3286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3289 <= 0;
  else
    WX3289 <= WX3288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3291 <= 0;
  else
    WX3291 <= WX3290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3293 <= 0;
  else
    WX3293 <= WX3292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3295 <= 0;
  else
    WX3295 <= WX3294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3297 <= 0;
  else
    WX3297 <= WX3296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3299 <= 0;
  else
    WX3299 <= WX3298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3301 <= 0;
  else
    WX3301 <= WX3300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3303 <= 0;
  else
    WX3303 <= WX3302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3305 <= 0;
  else
    WX3305 <= WX3304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3307 <= 0;
  else
    WX3307 <= WX3306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3309 <= 0;
  else
    WX3309 <= WX3308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3311 <= 0;
  else
    WX3311 <= WX3310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3313 <= 0;
  else
    WX3313 <= WX3312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3315 <= 0;
  else
    WX3315 <= WX3314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3317 <= 0;
  else
    WX3317 <= WX3316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3319 <= 0;
  else
    WX3319 <= WX3318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3321 <= 0;
  else
    WX3321 <= WX3320;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3323 <= 0;
  else
    WX3323 <= WX3322;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3325 <= 0;
  else
    WX3325 <= WX3324;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3327 <= 0;
  else
    WX3327 <= WX3326;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3329 <= 0;
  else
    WX3329 <= WX3328;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3331 <= 0;
  else
    WX3331 <= WX3330;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3333 <= 0;
  else
    WX3333 <= WX3332;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3335 <= 0;
  else
    WX3335 <= WX3334;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3337 <= 0;
  else
    WX3337 <= WX3336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3339 <= 0;
  else
    WX3339 <= WX3338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3341 <= 0;
  else
    WX3341 <= WX3340;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3343 <= 0;
  else
    WX3343 <= WX3342;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3345 <= 0;
  else
    WX3345 <= WX3344;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3347 <= 0;
  else
    WX3347 <= WX3346;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3349 <= 0;
  else
    WX3349 <= WX3348;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3351 <= 0;
  else
    WX3351 <= WX3350;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3353 <= 0;
  else
    WX3353 <= WX3352;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3355 <= 0;
  else
    WX3355 <= WX3354;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3357 <= 0;
  else
    WX3357 <= WX3356;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3359 <= 0;
  else
    WX3359 <= WX3358;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3361 <= 0;
  else
    WX3361 <= WX3360;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3363 <= 0;
  else
    WX3363 <= WX3362;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3365 <= 0;
  else
    WX3365 <= WX3364;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3367 <= 0;
  else
    WX3367 <= WX3366;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3369 <= 0;
  else
    WX3369 <= WX3368;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3371 <= 0;
  else
    WX3371 <= WX3370;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3373 <= 0;
  else
    WX3373 <= WX3372;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3375 <= 0;
  else
    WX3375 <= WX3374;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3377 <= 0;
  else
    WX3377 <= WX3376;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3379 <= 0;
  else
    WX3379 <= WX3378;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3381 <= 0;
  else
    WX3381 <= WX3380;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3383 <= 0;
  else
    WX3383 <= WX3382;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3385 <= 0;
  else
    WX3385 <= WX3384;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3387 <= 0;
  else
    WX3387 <= WX3386;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3389 <= 0;
  else
    WX3389 <= WX3388;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3391 <= 0;
  else
    WX3391 <= WX3390;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3393 <= 0;
  else
    WX3393 <= WX3392;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3395 <= 0;
  else
    WX3395 <= WX3394;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3397 <= 0;
  else
    WX3397 <= WX3396;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3399 <= 0;
  else
    WX3399 <= WX3398;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3401 <= 0;
  else
    WX3401 <= WX3400;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3403 <= 0;
  else
    WX3403 <= WX3402;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3405 <= 0;
  else
    WX3405 <= WX3404;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3407 <= 0;
  else
    WX3407 <= WX3406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3409 <= 0;
  else
    WX3409 <= WX3408;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3411 <= 0;
  else
    WX3411 <= WX3410;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3413 <= 0;
  else
    WX3413 <= WX3412;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3415 <= 0;
  else
    WX3415 <= WX3414;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3417 <= 0;
  else
    WX3417 <= WX3416;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3419 <= 0;
  else
    WX3419 <= WX3418;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3421 <= 0;
  else
    WX3421 <= WX3420;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3423 <= 0;
  else
    WX3423 <= WX3422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3425 <= 0;
  else
    WX3425 <= WX3424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3427 <= 0;
  else
    WX3427 <= WX3426;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3429 <= 0;
  else
    WX3429 <= WX3428;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3431 <= 0;
  else
    WX3431 <= WX3430;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3433 <= 0;
  else
    WX3433 <= WX3432;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3435 <= 0;
  else
    WX3435 <= WX3434;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3437 <= 0;
  else
    WX3437 <= WX3436;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3439 <= 0;
  else
    WX3439 <= WX3438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3441 <= 0;
  else
    WX3441 <= WX3440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3443 <= 0;
  else
    WX3443 <= WX3442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3445 <= 0;
  else
    WX3445 <= WX3444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3447 <= 0;
  else
    WX3447 <= WX3446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3449 <= 0;
  else
    WX3449 <= WX3448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3451 <= 0;
  else
    WX3451 <= WX3450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3453 <= 0;
  else
    WX3453 <= WX3452;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3455 <= 0;
  else
    WX3455 <= WX3454;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3457 <= 0;
  else
    WX3457 <= WX3456;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3459 <= 0;
  else
    WX3459 <= WX3458;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3461 <= 0;
  else
    WX3461 <= WX3460;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3463 <= 0;
  else
    WX3463 <= WX3462;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3465 <= 0;
  else
    WX3465 <= WX3464;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3467 <= 0;
  else
    WX3467 <= WX3466;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3469 <= 0;
  else
    WX3469 <= WX3468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3471 <= 0;
  else
    WX3471 <= WX3470;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3473 <= 0;
  else
    WX3473 <= WX3472;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3475 <= 0;
  else
    WX3475 <= WX3474;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3477 <= 0;
  else
    WX3477 <= WX3476;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3479 <= 0;
  else
    WX3479 <= WX3478;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3481 <= 0;
  else
    WX3481 <= WX3480;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3483 <= 0;
  else
    WX3483 <= WX3482;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX3485 <= 0;
  else
    WX3485 <= WX3484;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2141_ <= 0;
  else
    _2141_ <= WX3850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2142_ <= 0;
  else
    _2142_ <= WX3852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2143_ <= 0;
  else
    _2143_ <= WX3854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2144_ <= 0;
  else
    _2144_ <= WX3856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2145_ <= 0;
  else
    _2145_ <= WX3858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2146_ <= 0;
  else
    _2146_ <= WX3860;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2147_ <= 0;
  else
    _2147_ <= WX3862;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2148_ <= 0;
  else
    _2148_ <= WX3864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2149_ <= 0;
  else
    _2149_ <= WX3866;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2150_ <= 0;
  else
    _2150_ <= WX3868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2151_ <= 0;
  else
    _2151_ <= WX3870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2152_ <= 0;
  else
    _2152_ <= WX3872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2153_ <= 0;
  else
    _2153_ <= WX3874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2154_ <= 0;
  else
    _2154_ <= WX3876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2155_ <= 0;
  else
    _2155_ <= WX3878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2156_ <= 0;
  else
    _2156_ <= WX3880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2157_ <= 0;
  else
    _2157_ <= WX3882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2158_ <= 0;
  else
    _2158_ <= WX3884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2159_ <= 0;
  else
    _2159_ <= WX3886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2160_ <= 0;
  else
    _2160_ <= WX3888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2161_ <= 0;
  else
    _2161_ <= WX3890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2162_ <= 0;
  else
    _2162_ <= WX3892;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2163_ <= 0;
  else
    _2163_ <= WX3894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2164_ <= 0;
  else
    _2164_ <= WX3896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2165_ <= 0;
  else
    _2165_ <= WX3898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2166_ <= 0;
  else
    _2166_ <= WX3900;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2167_ <= 0;
  else
    _2167_ <= WX3902;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2168_ <= 0;
  else
    _2168_ <= WX3904;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2169_ <= 0;
  else
    _2169_ <= WX3906;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2170_ <= 0;
  else
    _2170_ <= WX3908;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2171_ <= 0;
  else
    _2171_ <= WX3910;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2172_ <= 0;
  else
    _2172_ <= WX3912;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4364 <= 0;
  else
    WX4364 <= WX4363;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4366 <= 0;
  else
    WX4366 <= WX4365;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4368 <= 0;
  else
    WX4368 <= WX4367;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4370 <= 0;
  else
    WX4370 <= WX4369;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4372 <= 0;
  else
    WX4372 <= WX4371;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4374 <= 0;
  else
    WX4374 <= WX4373;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4376 <= 0;
  else
    WX4376 <= WX4375;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4378 <= 0;
  else
    WX4378 <= WX4377;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4380 <= 0;
  else
    WX4380 <= WX4379;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4382 <= 0;
  else
    WX4382 <= WX4381;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4384 <= 0;
  else
    WX4384 <= WX4383;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4386 <= 0;
  else
    WX4386 <= WX4385;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4388 <= 0;
  else
    WX4388 <= WX4387;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4390 <= 0;
  else
    WX4390 <= WX4389;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4392 <= 0;
  else
    WX4392 <= WX4391;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4394 <= 0;
  else
    WX4394 <= WX4393;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4396 <= 0;
  else
    WX4396 <= WX4395;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4398 <= 0;
  else
    WX4398 <= WX4397;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4400 <= 0;
  else
    WX4400 <= WX4399;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4402 <= 0;
  else
    WX4402 <= WX4401;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4404 <= 0;
  else
    WX4404 <= WX4403;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4406 <= 0;
  else
    WX4406 <= WX4405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4408 <= 0;
  else
    WX4408 <= WX4407;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4410 <= 0;
  else
    WX4410 <= WX4409;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4412 <= 0;
  else
    WX4412 <= WX4411;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4414 <= 0;
  else
    WX4414 <= WX4413;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4416 <= 0;
  else
    WX4416 <= WX4415;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4418 <= 0;
  else
    WX4418 <= WX4417;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4420 <= 0;
  else
    WX4420 <= WX4419;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4422 <= 0;
  else
    WX4422 <= WX4421;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4424 <= 0;
  else
    WX4424 <= WX4423;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4426 <= 0;
  else
    WX4426 <= WX4425;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4524 <= 0;
  else
    WX4524 <= WX4523;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4526 <= 0;
  else
    WX4526 <= WX4525;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4528 <= 0;
  else
    WX4528 <= WX4527;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4530 <= 0;
  else
    WX4530 <= WX4529;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4532 <= 0;
  else
    WX4532 <= WX4531;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4534 <= 0;
  else
    WX4534 <= WX4533;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4536 <= 0;
  else
    WX4536 <= WX4535;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4538 <= 0;
  else
    WX4538 <= WX4537;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4540 <= 0;
  else
    WX4540 <= WX4539;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4542 <= 0;
  else
    WX4542 <= WX4541;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4544 <= 0;
  else
    WX4544 <= WX4543;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4546 <= 0;
  else
    WX4546 <= WX4545;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4548 <= 0;
  else
    WX4548 <= WX4547;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4550 <= 0;
  else
    WX4550 <= WX4549;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4552 <= 0;
  else
    WX4552 <= WX4551;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4554 <= 0;
  else
    WX4554 <= WX4553;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4556 <= 0;
  else
    WX4556 <= WX4555;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4558 <= 0;
  else
    WX4558 <= WX4557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4560 <= 0;
  else
    WX4560 <= WX4559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4562 <= 0;
  else
    WX4562 <= WX4561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4564 <= 0;
  else
    WX4564 <= WX4563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4566 <= 0;
  else
    WX4566 <= WX4565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4568 <= 0;
  else
    WX4568 <= WX4567;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4570 <= 0;
  else
    WX4570 <= WX4569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4572 <= 0;
  else
    WX4572 <= WX4571;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4574 <= 0;
  else
    WX4574 <= WX4573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4576 <= 0;
  else
    WX4576 <= WX4575;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4578 <= 0;
  else
    WX4578 <= WX4577;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4580 <= 0;
  else
    WX4580 <= WX4579;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4582 <= 0;
  else
    WX4582 <= WX4581;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4584 <= 0;
  else
    WX4584 <= WX4583;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4586 <= 0;
  else
    WX4586 <= WX4585;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4588 <= 0;
  else
    WX4588 <= WX4587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4590 <= 0;
  else
    WX4590 <= WX4589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4592 <= 0;
  else
    WX4592 <= WX4591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4594 <= 0;
  else
    WX4594 <= WX4593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4596 <= 0;
  else
    WX4596 <= WX4595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4598 <= 0;
  else
    WX4598 <= WX4597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4600 <= 0;
  else
    WX4600 <= WX4599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4602 <= 0;
  else
    WX4602 <= WX4601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4604 <= 0;
  else
    WX4604 <= WX4603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4606 <= 0;
  else
    WX4606 <= WX4605;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4608 <= 0;
  else
    WX4608 <= WX4607;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4610 <= 0;
  else
    WX4610 <= WX4609;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4612 <= 0;
  else
    WX4612 <= WX4611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4614 <= 0;
  else
    WX4614 <= WX4613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4616 <= 0;
  else
    WX4616 <= WX4615;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4618 <= 0;
  else
    WX4618 <= WX4617;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4620 <= 0;
  else
    WX4620 <= WX4619;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4622 <= 0;
  else
    WX4622 <= WX4621;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4624 <= 0;
  else
    WX4624 <= WX4623;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4626 <= 0;
  else
    WX4626 <= WX4625;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4628 <= 0;
  else
    WX4628 <= WX4627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4630 <= 0;
  else
    WX4630 <= WX4629;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4632 <= 0;
  else
    WX4632 <= WX4631;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4634 <= 0;
  else
    WX4634 <= WX4633;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4636 <= 0;
  else
    WX4636 <= WX4635;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4638 <= 0;
  else
    WX4638 <= WX4637;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4640 <= 0;
  else
    WX4640 <= WX4639;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4642 <= 0;
  else
    WX4642 <= WX4641;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4644 <= 0;
  else
    WX4644 <= WX4643;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4646 <= 0;
  else
    WX4646 <= WX4645;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4648 <= 0;
  else
    WX4648 <= WX4647;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4650 <= 0;
  else
    WX4650 <= WX4649;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4652 <= 0;
  else
    WX4652 <= WX4651;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4654 <= 0;
  else
    WX4654 <= WX4653;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4656 <= 0;
  else
    WX4656 <= WX4655;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4658 <= 0;
  else
    WX4658 <= WX4657;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4660 <= 0;
  else
    WX4660 <= WX4659;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4662 <= 0;
  else
    WX4662 <= WX4661;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4664 <= 0;
  else
    WX4664 <= WX4663;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4666 <= 0;
  else
    WX4666 <= WX4665;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4668 <= 0;
  else
    WX4668 <= WX4667;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4670 <= 0;
  else
    WX4670 <= WX4669;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4672 <= 0;
  else
    WX4672 <= WX4671;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4674 <= 0;
  else
    WX4674 <= WX4673;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4676 <= 0;
  else
    WX4676 <= WX4675;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4678 <= 0;
  else
    WX4678 <= WX4677;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4680 <= 0;
  else
    WX4680 <= WX4679;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4682 <= 0;
  else
    WX4682 <= WX4681;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4684 <= 0;
  else
    WX4684 <= WX4683;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4686 <= 0;
  else
    WX4686 <= WX4685;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4688 <= 0;
  else
    WX4688 <= WX4687;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4690 <= 0;
  else
    WX4690 <= WX4689;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4692 <= 0;
  else
    WX4692 <= WX4691;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4694 <= 0;
  else
    WX4694 <= WX4693;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4696 <= 0;
  else
    WX4696 <= WX4695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4698 <= 0;
  else
    WX4698 <= WX4697;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4700 <= 0;
  else
    WX4700 <= WX4699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4702 <= 0;
  else
    WX4702 <= WX4701;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4704 <= 0;
  else
    WX4704 <= WX4703;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4706 <= 0;
  else
    WX4706 <= WX4705;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4708 <= 0;
  else
    WX4708 <= WX4707;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4710 <= 0;
  else
    WX4710 <= WX4709;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4712 <= 0;
  else
    WX4712 <= WX4711;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4714 <= 0;
  else
    WX4714 <= WX4713;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4716 <= 0;
  else
    WX4716 <= WX4715;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4718 <= 0;
  else
    WX4718 <= WX4717;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4720 <= 0;
  else
    WX4720 <= WX4719;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4722 <= 0;
  else
    WX4722 <= WX4721;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4724 <= 0;
  else
    WX4724 <= WX4723;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4726 <= 0;
  else
    WX4726 <= WX4725;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4728 <= 0;
  else
    WX4728 <= WX4727;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4730 <= 0;
  else
    WX4730 <= WX4729;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4732 <= 0;
  else
    WX4732 <= WX4731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4734 <= 0;
  else
    WX4734 <= WX4733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4736 <= 0;
  else
    WX4736 <= WX4735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4738 <= 0;
  else
    WX4738 <= WX4737;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4740 <= 0;
  else
    WX4740 <= WX4739;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4742 <= 0;
  else
    WX4742 <= WX4741;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4744 <= 0;
  else
    WX4744 <= WX4743;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4746 <= 0;
  else
    WX4746 <= WX4745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4748 <= 0;
  else
    WX4748 <= WX4747;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4750 <= 0;
  else
    WX4750 <= WX4749;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4752 <= 0;
  else
    WX4752 <= WX4751;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4754 <= 0;
  else
    WX4754 <= WX4753;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4756 <= 0;
  else
    WX4756 <= WX4755;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4758 <= 0;
  else
    WX4758 <= WX4757;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4760 <= 0;
  else
    WX4760 <= WX4759;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4762 <= 0;
  else
    WX4762 <= WX4761;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4764 <= 0;
  else
    WX4764 <= WX4763;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4766 <= 0;
  else
    WX4766 <= WX4765;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4768 <= 0;
  else
    WX4768 <= WX4767;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4770 <= 0;
  else
    WX4770 <= WX4769;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4772 <= 0;
  else
    WX4772 <= WX4771;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4774 <= 0;
  else
    WX4774 <= WX4773;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4776 <= 0;
  else
    WX4776 <= WX4775;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX4778 <= 0;
  else
    WX4778 <= WX4777;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2173_ <= 0;
  else
    _2173_ <= WX5143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2174_ <= 0;
  else
    _2174_ <= WX5145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2175_ <= 0;
  else
    _2175_ <= WX5147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2176_ <= 0;
  else
    _2176_ <= WX5149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2177_ <= 0;
  else
    _2177_ <= WX5151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2178_ <= 0;
  else
    _2178_ <= WX5153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2179_ <= 0;
  else
    _2179_ <= WX5155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2180_ <= 0;
  else
    _2180_ <= WX5157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2181_ <= 0;
  else
    _2181_ <= WX5159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2182_ <= 0;
  else
    _2182_ <= WX5161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2183_ <= 0;
  else
    _2183_ <= WX5163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2184_ <= 0;
  else
    _2184_ <= WX5165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2185_ <= 0;
  else
    _2185_ <= WX5167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2186_ <= 0;
  else
    _2186_ <= WX5169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2187_ <= 0;
  else
    _2187_ <= WX5171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2188_ <= 0;
  else
    _2188_ <= WX5173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2189_ <= 0;
  else
    _2189_ <= WX5175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2190_ <= 0;
  else
    _2190_ <= WX5177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2191_ <= 0;
  else
    _2191_ <= WX5179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2192_ <= 0;
  else
    _2192_ <= WX5181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2193_ <= 0;
  else
    _2193_ <= WX5183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2194_ <= 0;
  else
    _2194_ <= WX5185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2195_ <= 0;
  else
    _2195_ <= WX5187;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2196_ <= 0;
  else
    _2196_ <= WX5189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2197_ <= 0;
  else
    _2197_ <= WX5191;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2198_ <= 0;
  else
    _2198_ <= WX5193;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2199_ <= 0;
  else
    _2199_ <= WX5195;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2200_ <= 0;
  else
    _2200_ <= WX5197;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2201_ <= 0;
  else
    _2201_ <= WX5199;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2202_ <= 0;
  else
    _2202_ <= WX5201;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2203_ <= 0;
  else
    _2203_ <= WX5203;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2204_ <= 0;
  else
    _2204_ <= WX5205;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5657 <= 0;
  else
    WX5657 <= WX5656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5659 <= 0;
  else
    WX5659 <= WX5658;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5661 <= 0;
  else
    WX5661 <= WX5660;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5663 <= 0;
  else
    WX5663 <= WX5662;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5665 <= 0;
  else
    WX5665 <= WX5664;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5667 <= 0;
  else
    WX5667 <= WX5666;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5669 <= 0;
  else
    WX5669 <= WX5668;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5671 <= 0;
  else
    WX5671 <= WX5670;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5673 <= 0;
  else
    WX5673 <= WX5672;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5675 <= 0;
  else
    WX5675 <= WX5674;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5677 <= 0;
  else
    WX5677 <= WX5676;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5679 <= 0;
  else
    WX5679 <= WX5678;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5681 <= 0;
  else
    WX5681 <= WX5680;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5683 <= 0;
  else
    WX5683 <= WX5682;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5685 <= 0;
  else
    WX5685 <= WX5684;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5687 <= 0;
  else
    WX5687 <= WX5686;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5689 <= 0;
  else
    WX5689 <= WX5688;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5691 <= 0;
  else
    WX5691 <= WX5690;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5693 <= 0;
  else
    WX5693 <= WX5692;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5695 <= 0;
  else
    WX5695 <= WX5694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5697 <= 0;
  else
    WX5697 <= WX5696;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5699 <= 0;
  else
    WX5699 <= WX5698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5701 <= 0;
  else
    WX5701 <= WX5700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5703 <= 0;
  else
    WX5703 <= WX5702;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5705 <= 0;
  else
    WX5705 <= WX5704;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5707 <= 0;
  else
    WX5707 <= WX5706;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5709 <= 0;
  else
    WX5709 <= WX5708;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5711 <= 0;
  else
    WX5711 <= WX5710;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5713 <= 0;
  else
    WX5713 <= WX5712;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5715 <= 0;
  else
    WX5715 <= WX5714;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5717 <= 0;
  else
    WX5717 <= WX5716;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5719 <= 0;
  else
    WX5719 <= WX5718;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5817 <= 0;
  else
    WX5817 <= WX5816;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5819 <= 0;
  else
    WX5819 <= WX5818;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5821 <= 0;
  else
    WX5821 <= WX5820;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5823 <= 0;
  else
    WX5823 <= WX5822;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5825 <= 0;
  else
    WX5825 <= WX5824;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5827 <= 0;
  else
    WX5827 <= WX5826;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5829 <= 0;
  else
    WX5829 <= WX5828;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5831 <= 0;
  else
    WX5831 <= WX5830;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5833 <= 0;
  else
    WX5833 <= WX5832;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5835 <= 0;
  else
    WX5835 <= WX5834;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5837 <= 0;
  else
    WX5837 <= WX5836;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5839 <= 0;
  else
    WX5839 <= WX5838;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5841 <= 0;
  else
    WX5841 <= WX5840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5843 <= 0;
  else
    WX5843 <= WX5842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5845 <= 0;
  else
    WX5845 <= WX5844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5847 <= 0;
  else
    WX5847 <= WX5846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5849 <= 0;
  else
    WX5849 <= WX5848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5851 <= 0;
  else
    WX5851 <= WX5850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5853 <= 0;
  else
    WX5853 <= WX5852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5855 <= 0;
  else
    WX5855 <= WX5854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5857 <= 0;
  else
    WX5857 <= WX5856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5859 <= 0;
  else
    WX5859 <= WX5858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5861 <= 0;
  else
    WX5861 <= WX5860;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5863 <= 0;
  else
    WX5863 <= WX5862;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5865 <= 0;
  else
    WX5865 <= WX5864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5867 <= 0;
  else
    WX5867 <= WX5866;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5869 <= 0;
  else
    WX5869 <= WX5868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5871 <= 0;
  else
    WX5871 <= WX5870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5873 <= 0;
  else
    WX5873 <= WX5872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5875 <= 0;
  else
    WX5875 <= WX5874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5877 <= 0;
  else
    WX5877 <= WX5876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5879 <= 0;
  else
    WX5879 <= WX5878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5881 <= 0;
  else
    WX5881 <= WX5880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5883 <= 0;
  else
    WX5883 <= WX5882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5885 <= 0;
  else
    WX5885 <= WX5884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5887 <= 0;
  else
    WX5887 <= WX5886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5889 <= 0;
  else
    WX5889 <= WX5888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5891 <= 0;
  else
    WX5891 <= WX5890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5893 <= 0;
  else
    WX5893 <= WX5892;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5895 <= 0;
  else
    WX5895 <= WX5894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5897 <= 0;
  else
    WX5897 <= WX5896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5899 <= 0;
  else
    WX5899 <= WX5898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5901 <= 0;
  else
    WX5901 <= WX5900;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5903 <= 0;
  else
    WX5903 <= WX5902;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5905 <= 0;
  else
    WX5905 <= WX5904;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5907 <= 0;
  else
    WX5907 <= WX5906;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5909 <= 0;
  else
    WX5909 <= WX5908;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5911 <= 0;
  else
    WX5911 <= WX5910;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5913 <= 0;
  else
    WX5913 <= WX5912;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5915 <= 0;
  else
    WX5915 <= WX5914;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5917 <= 0;
  else
    WX5917 <= WX5916;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5919 <= 0;
  else
    WX5919 <= WX5918;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5921 <= 0;
  else
    WX5921 <= WX5920;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5923 <= 0;
  else
    WX5923 <= WX5922;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5925 <= 0;
  else
    WX5925 <= WX5924;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5927 <= 0;
  else
    WX5927 <= WX5926;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5929 <= 0;
  else
    WX5929 <= WX5928;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5931 <= 0;
  else
    WX5931 <= WX5930;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5933 <= 0;
  else
    WX5933 <= WX5932;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5935 <= 0;
  else
    WX5935 <= WX5934;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5937 <= 0;
  else
    WX5937 <= WX5936;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5939 <= 0;
  else
    WX5939 <= WX5938;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5941 <= 0;
  else
    WX5941 <= WX5940;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5943 <= 0;
  else
    WX5943 <= WX5942;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5945 <= 0;
  else
    WX5945 <= WX5944;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5947 <= 0;
  else
    WX5947 <= WX5946;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5949 <= 0;
  else
    WX5949 <= WX5948;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5951 <= 0;
  else
    WX5951 <= WX5950;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5953 <= 0;
  else
    WX5953 <= WX5952;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5955 <= 0;
  else
    WX5955 <= WX5954;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5957 <= 0;
  else
    WX5957 <= WX5956;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5959 <= 0;
  else
    WX5959 <= WX5958;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5961 <= 0;
  else
    WX5961 <= WX5960;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5963 <= 0;
  else
    WX5963 <= WX5962;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5965 <= 0;
  else
    WX5965 <= WX5964;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5967 <= 0;
  else
    WX5967 <= WX5966;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5969 <= 0;
  else
    WX5969 <= WX5968;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5971 <= 0;
  else
    WX5971 <= WX5970;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5973 <= 0;
  else
    WX5973 <= WX5972;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5975 <= 0;
  else
    WX5975 <= WX5974;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5977 <= 0;
  else
    WX5977 <= WX5976;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5979 <= 0;
  else
    WX5979 <= WX5978;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5981 <= 0;
  else
    WX5981 <= WX5980;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5983 <= 0;
  else
    WX5983 <= WX5982;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5985 <= 0;
  else
    WX5985 <= WX5984;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5987 <= 0;
  else
    WX5987 <= WX5986;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5989 <= 0;
  else
    WX5989 <= WX5988;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5991 <= 0;
  else
    WX5991 <= WX5990;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5993 <= 0;
  else
    WX5993 <= WX5992;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5995 <= 0;
  else
    WX5995 <= WX5994;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5997 <= 0;
  else
    WX5997 <= WX5996;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX5999 <= 0;
  else
    WX5999 <= WX5998;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6001 <= 0;
  else
    WX6001 <= WX6000;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6003 <= 0;
  else
    WX6003 <= WX6002;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6005 <= 0;
  else
    WX6005 <= WX6004;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6007 <= 0;
  else
    WX6007 <= WX6006;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6009 <= 0;
  else
    WX6009 <= WX6008;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6011 <= 0;
  else
    WX6011 <= WX6010;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6013 <= 0;
  else
    WX6013 <= WX6012;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6015 <= 0;
  else
    WX6015 <= WX6014;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6017 <= 0;
  else
    WX6017 <= WX6016;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6019 <= 0;
  else
    WX6019 <= WX6018;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6021 <= 0;
  else
    WX6021 <= WX6020;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6023 <= 0;
  else
    WX6023 <= WX6022;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6025 <= 0;
  else
    WX6025 <= WX6024;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6027 <= 0;
  else
    WX6027 <= WX6026;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6029 <= 0;
  else
    WX6029 <= WX6028;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6031 <= 0;
  else
    WX6031 <= WX6030;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6033 <= 0;
  else
    WX6033 <= WX6032;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6035 <= 0;
  else
    WX6035 <= WX6034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6037 <= 0;
  else
    WX6037 <= WX6036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6039 <= 0;
  else
    WX6039 <= WX6038;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6041 <= 0;
  else
    WX6041 <= WX6040;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6043 <= 0;
  else
    WX6043 <= WX6042;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6045 <= 0;
  else
    WX6045 <= WX6044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6047 <= 0;
  else
    WX6047 <= WX6046;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6049 <= 0;
  else
    WX6049 <= WX6048;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6051 <= 0;
  else
    WX6051 <= WX6050;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6053 <= 0;
  else
    WX6053 <= WX6052;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6055 <= 0;
  else
    WX6055 <= WX6054;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6057 <= 0;
  else
    WX6057 <= WX6056;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6059 <= 0;
  else
    WX6059 <= WX6058;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6061 <= 0;
  else
    WX6061 <= WX6060;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6063 <= 0;
  else
    WX6063 <= WX6062;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6065 <= 0;
  else
    WX6065 <= WX6064;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6067 <= 0;
  else
    WX6067 <= WX6066;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6069 <= 0;
  else
    WX6069 <= WX6068;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6071 <= 0;
  else
    WX6071 <= WX6070;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2205_ <= 0;
  else
    _2205_ <= WX6436;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2206_ <= 0;
  else
    _2206_ <= WX6438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2207_ <= 0;
  else
    _2207_ <= WX6440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2208_ <= 0;
  else
    _2208_ <= WX6442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2209_ <= 0;
  else
    _2209_ <= WX6444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2210_ <= 0;
  else
    _2210_ <= WX6446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2211_ <= 0;
  else
    _2211_ <= WX6448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2212_ <= 0;
  else
    _2212_ <= WX6450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2213_ <= 0;
  else
    _2213_ <= WX6452;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2214_ <= 0;
  else
    _2214_ <= WX6454;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2215_ <= 0;
  else
    _2215_ <= WX6456;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2216_ <= 0;
  else
    _2216_ <= WX6458;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2217_ <= 0;
  else
    _2217_ <= WX6460;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2218_ <= 0;
  else
    _2218_ <= WX6462;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2219_ <= 0;
  else
    _2219_ <= WX6464;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2220_ <= 0;
  else
    _2220_ <= WX6466;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2221_ <= 0;
  else
    _2221_ <= WX6468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2222_ <= 0;
  else
    _2222_ <= WX6470;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2223_ <= 0;
  else
    _2223_ <= WX6472;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2224_ <= 0;
  else
    _2224_ <= WX6474;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2225_ <= 0;
  else
    _2225_ <= WX6476;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2226_ <= 0;
  else
    _2226_ <= WX6478;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2227_ <= 0;
  else
    _2227_ <= WX6480;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2228_ <= 0;
  else
    _2228_ <= WX6482;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2229_ <= 0;
  else
    _2229_ <= WX6484;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2230_ <= 0;
  else
    _2230_ <= WX6486;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2231_ <= 0;
  else
    _2231_ <= WX6488;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2232_ <= 0;
  else
    _2232_ <= WX6490;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2233_ <= 0;
  else
    _2233_ <= WX6492;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2234_ <= 0;
  else
    _2234_ <= WX6494;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2235_ <= 0;
  else
    _2235_ <= WX6496;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2236_ <= 0;
  else
    _2236_ <= WX6498;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6950 <= 0;
  else
    WX6950 <= WX6949;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6952 <= 0;
  else
    WX6952 <= WX6951;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6954 <= 0;
  else
    WX6954 <= WX6953;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6956 <= 0;
  else
    WX6956 <= WX6955;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6958 <= 0;
  else
    WX6958 <= WX6957;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6960 <= 0;
  else
    WX6960 <= WX6959;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6962 <= 0;
  else
    WX6962 <= WX6961;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6964 <= 0;
  else
    WX6964 <= WX6963;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6966 <= 0;
  else
    WX6966 <= WX6965;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6968 <= 0;
  else
    WX6968 <= WX6967;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6970 <= 0;
  else
    WX6970 <= WX6969;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6972 <= 0;
  else
    WX6972 <= WX6971;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6974 <= 0;
  else
    WX6974 <= WX6973;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6976 <= 0;
  else
    WX6976 <= WX6975;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6978 <= 0;
  else
    WX6978 <= WX6977;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6980 <= 0;
  else
    WX6980 <= WX6979;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6982 <= 0;
  else
    WX6982 <= WX6981;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6984 <= 0;
  else
    WX6984 <= WX6983;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6986 <= 0;
  else
    WX6986 <= WX6985;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6988 <= 0;
  else
    WX6988 <= WX6987;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6990 <= 0;
  else
    WX6990 <= WX6989;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6992 <= 0;
  else
    WX6992 <= WX6991;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6994 <= 0;
  else
    WX6994 <= WX6993;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6996 <= 0;
  else
    WX6996 <= WX6995;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX6998 <= 0;
  else
    WX6998 <= WX6997;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7000 <= 0;
  else
    WX7000 <= WX6999;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7002 <= 0;
  else
    WX7002 <= WX7001;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7004 <= 0;
  else
    WX7004 <= WX7003;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7006 <= 0;
  else
    WX7006 <= WX7005;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7008 <= 0;
  else
    WX7008 <= WX7007;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7010 <= 0;
  else
    WX7010 <= WX7009;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7012 <= 0;
  else
    WX7012 <= WX7011;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7110 <= 0;
  else
    WX7110 <= WX7109;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7112 <= 0;
  else
    WX7112 <= WX7111;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7114 <= 0;
  else
    WX7114 <= WX7113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7116 <= 0;
  else
    WX7116 <= WX7115;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7118 <= 0;
  else
    WX7118 <= WX7117;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7120 <= 0;
  else
    WX7120 <= WX7119;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7122 <= 0;
  else
    WX7122 <= WX7121;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7124 <= 0;
  else
    WX7124 <= WX7123;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7126 <= 0;
  else
    WX7126 <= WX7125;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7128 <= 0;
  else
    WX7128 <= WX7127;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7130 <= 0;
  else
    WX7130 <= WX7129;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7132 <= 0;
  else
    WX7132 <= WX7131;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7134 <= 0;
  else
    WX7134 <= WX7133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7136 <= 0;
  else
    WX7136 <= WX7135;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7138 <= 0;
  else
    WX7138 <= WX7137;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7140 <= 0;
  else
    WX7140 <= WX7139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7142 <= 0;
  else
    WX7142 <= WX7141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7144 <= 0;
  else
    WX7144 <= WX7143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7146 <= 0;
  else
    WX7146 <= WX7145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7148 <= 0;
  else
    WX7148 <= WX7147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7150 <= 0;
  else
    WX7150 <= WX7149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7152 <= 0;
  else
    WX7152 <= WX7151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7154 <= 0;
  else
    WX7154 <= WX7153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7156 <= 0;
  else
    WX7156 <= WX7155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7158 <= 0;
  else
    WX7158 <= WX7157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7160 <= 0;
  else
    WX7160 <= WX7159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7162 <= 0;
  else
    WX7162 <= WX7161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7164 <= 0;
  else
    WX7164 <= WX7163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7166 <= 0;
  else
    WX7166 <= WX7165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7168 <= 0;
  else
    WX7168 <= WX7167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7170 <= 0;
  else
    WX7170 <= WX7169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7172 <= 0;
  else
    WX7172 <= WX7171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7174 <= 0;
  else
    WX7174 <= WX7173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7176 <= 0;
  else
    WX7176 <= WX7175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7178 <= 0;
  else
    WX7178 <= WX7177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7180 <= 0;
  else
    WX7180 <= WX7179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7182 <= 0;
  else
    WX7182 <= WX7181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7184 <= 0;
  else
    WX7184 <= WX7183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7186 <= 0;
  else
    WX7186 <= WX7185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7188 <= 0;
  else
    WX7188 <= WX7187;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7190 <= 0;
  else
    WX7190 <= WX7189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7192 <= 0;
  else
    WX7192 <= WX7191;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7194 <= 0;
  else
    WX7194 <= WX7193;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7196 <= 0;
  else
    WX7196 <= WX7195;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7198 <= 0;
  else
    WX7198 <= WX7197;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7200 <= 0;
  else
    WX7200 <= WX7199;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7202 <= 0;
  else
    WX7202 <= WX7201;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7204 <= 0;
  else
    WX7204 <= WX7203;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7206 <= 0;
  else
    WX7206 <= WX7205;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7208 <= 0;
  else
    WX7208 <= WX7207;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7210 <= 0;
  else
    WX7210 <= WX7209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7212 <= 0;
  else
    WX7212 <= WX7211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7214 <= 0;
  else
    WX7214 <= WX7213;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7216 <= 0;
  else
    WX7216 <= WX7215;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7218 <= 0;
  else
    WX7218 <= WX7217;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7220 <= 0;
  else
    WX7220 <= WX7219;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7222 <= 0;
  else
    WX7222 <= WX7221;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7224 <= 0;
  else
    WX7224 <= WX7223;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7226 <= 0;
  else
    WX7226 <= WX7225;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7228 <= 0;
  else
    WX7228 <= WX7227;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7230 <= 0;
  else
    WX7230 <= WX7229;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7232 <= 0;
  else
    WX7232 <= WX7231;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7234 <= 0;
  else
    WX7234 <= WX7233;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7236 <= 0;
  else
    WX7236 <= WX7235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7238 <= 0;
  else
    WX7238 <= WX7237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7240 <= 0;
  else
    WX7240 <= WX7239;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7242 <= 0;
  else
    WX7242 <= WX7241;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7244 <= 0;
  else
    WX7244 <= WX7243;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7246 <= 0;
  else
    WX7246 <= WX7245;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7248 <= 0;
  else
    WX7248 <= WX7247;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7250 <= 0;
  else
    WX7250 <= WX7249;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7252 <= 0;
  else
    WX7252 <= WX7251;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7254 <= 0;
  else
    WX7254 <= WX7253;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7256 <= 0;
  else
    WX7256 <= WX7255;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7258 <= 0;
  else
    WX7258 <= WX7257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7260 <= 0;
  else
    WX7260 <= WX7259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7262 <= 0;
  else
    WX7262 <= WX7261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7264 <= 0;
  else
    WX7264 <= WX7263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7266 <= 0;
  else
    WX7266 <= WX7265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7268 <= 0;
  else
    WX7268 <= WX7267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7270 <= 0;
  else
    WX7270 <= WX7269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7272 <= 0;
  else
    WX7272 <= WX7271;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7274 <= 0;
  else
    WX7274 <= WX7273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7276 <= 0;
  else
    WX7276 <= WX7275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7278 <= 0;
  else
    WX7278 <= WX7277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7280 <= 0;
  else
    WX7280 <= WX7279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7282 <= 0;
  else
    WX7282 <= WX7281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7284 <= 0;
  else
    WX7284 <= WX7283;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7286 <= 0;
  else
    WX7286 <= WX7285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7288 <= 0;
  else
    WX7288 <= WX7287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7290 <= 0;
  else
    WX7290 <= WX7289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7292 <= 0;
  else
    WX7292 <= WX7291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7294 <= 0;
  else
    WX7294 <= WX7293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7296 <= 0;
  else
    WX7296 <= WX7295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7298 <= 0;
  else
    WX7298 <= WX7297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7300 <= 0;
  else
    WX7300 <= WX7299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7302 <= 0;
  else
    WX7302 <= WX7301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7304 <= 0;
  else
    WX7304 <= WX7303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7306 <= 0;
  else
    WX7306 <= WX7305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7308 <= 0;
  else
    WX7308 <= WX7307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7310 <= 0;
  else
    WX7310 <= WX7309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7312 <= 0;
  else
    WX7312 <= WX7311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7314 <= 0;
  else
    WX7314 <= WX7313;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7316 <= 0;
  else
    WX7316 <= WX7315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7318 <= 0;
  else
    WX7318 <= WX7317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7320 <= 0;
  else
    WX7320 <= WX7319;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7322 <= 0;
  else
    WX7322 <= WX7321;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7324 <= 0;
  else
    WX7324 <= WX7323;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7326 <= 0;
  else
    WX7326 <= WX7325;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7328 <= 0;
  else
    WX7328 <= WX7327;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7330 <= 0;
  else
    WX7330 <= WX7329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7332 <= 0;
  else
    WX7332 <= WX7331;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7334 <= 0;
  else
    WX7334 <= WX7333;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7336 <= 0;
  else
    WX7336 <= WX7335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7338 <= 0;
  else
    WX7338 <= WX7337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7340 <= 0;
  else
    WX7340 <= WX7339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7342 <= 0;
  else
    WX7342 <= WX7341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7344 <= 0;
  else
    WX7344 <= WX7343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7346 <= 0;
  else
    WX7346 <= WX7345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7348 <= 0;
  else
    WX7348 <= WX7347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7350 <= 0;
  else
    WX7350 <= WX7349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7352 <= 0;
  else
    WX7352 <= WX7351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7354 <= 0;
  else
    WX7354 <= WX7353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7356 <= 0;
  else
    WX7356 <= WX7355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7358 <= 0;
  else
    WX7358 <= WX7357;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7360 <= 0;
  else
    WX7360 <= WX7359;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7362 <= 0;
  else
    WX7362 <= WX7361;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX7364 <= 0;
  else
    WX7364 <= WX7363;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2237_ <= 0;
  else
    _2237_ <= WX7729;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2238_ <= 0;
  else
    _2238_ <= WX7731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2239_ <= 0;
  else
    _2239_ <= WX7733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2240_ <= 0;
  else
    _2240_ <= WX7735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2241_ <= 0;
  else
    _2241_ <= WX7737;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2242_ <= 0;
  else
    _2242_ <= WX7739;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2243_ <= 0;
  else
    _2243_ <= WX7741;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2244_ <= 0;
  else
    _2244_ <= WX7743;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2245_ <= 0;
  else
    _2245_ <= WX7745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2246_ <= 0;
  else
    _2246_ <= WX7747;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2247_ <= 0;
  else
    _2247_ <= WX7749;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2248_ <= 0;
  else
    _2248_ <= WX7751;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2249_ <= 0;
  else
    _2249_ <= WX7753;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2250_ <= 0;
  else
    _2250_ <= WX7755;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2251_ <= 0;
  else
    _2251_ <= WX7757;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2252_ <= 0;
  else
    _2252_ <= WX7759;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2253_ <= 0;
  else
    _2253_ <= WX7761;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2254_ <= 0;
  else
    _2254_ <= WX7763;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2255_ <= 0;
  else
    _2255_ <= WX7765;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2256_ <= 0;
  else
    _2256_ <= WX7767;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2257_ <= 0;
  else
    _2257_ <= WX7769;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2258_ <= 0;
  else
    _2258_ <= WX7771;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2259_ <= 0;
  else
    _2259_ <= WX7773;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2260_ <= 0;
  else
    _2260_ <= WX7775;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2261_ <= 0;
  else
    _2261_ <= WX7777;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2262_ <= 0;
  else
    _2262_ <= WX7779;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2263_ <= 0;
  else
    _2263_ <= WX7781;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2264_ <= 0;
  else
    _2264_ <= WX7783;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2265_ <= 0;
  else
    _2265_ <= WX7785;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2266_ <= 0;
  else
    _2266_ <= WX7787;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2267_ <= 0;
  else
    _2267_ <= WX7789;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2268_ <= 0;
  else
    _2268_ <= WX7791;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8243 <= 0;
  else
    WX8243 <= WX8242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8245 <= 0;
  else
    WX8245 <= WX8244;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8247 <= 0;
  else
    WX8247 <= WX8246;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8249 <= 0;
  else
    WX8249 <= WX8248;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8251 <= 0;
  else
    WX8251 <= WX8250;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8253 <= 0;
  else
    WX8253 <= WX8252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8255 <= 0;
  else
    WX8255 <= WX8254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8257 <= 0;
  else
    WX8257 <= WX8256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8259 <= 0;
  else
    WX8259 <= WX8258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8261 <= 0;
  else
    WX8261 <= WX8260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8263 <= 0;
  else
    WX8263 <= WX8262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8265 <= 0;
  else
    WX8265 <= WX8264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8267 <= 0;
  else
    WX8267 <= WX8266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8269 <= 0;
  else
    WX8269 <= WX8268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8271 <= 0;
  else
    WX8271 <= WX8270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8273 <= 0;
  else
    WX8273 <= WX8272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8275 <= 0;
  else
    WX8275 <= WX8274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8277 <= 0;
  else
    WX8277 <= WX8276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8279 <= 0;
  else
    WX8279 <= WX8278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8281 <= 0;
  else
    WX8281 <= WX8280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8283 <= 0;
  else
    WX8283 <= WX8282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8285 <= 0;
  else
    WX8285 <= WX8284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8287 <= 0;
  else
    WX8287 <= WX8286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8289 <= 0;
  else
    WX8289 <= WX8288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8291 <= 0;
  else
    WX8291 <= WX8290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8293 <= 0;
  else
    WX8293 <= WX8292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8295 <= 0;
  else
    WX8295 <= WX8294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8297 <= 0;
  else
    WX8297 <= WX8296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8299 <= 0;
  else
    WX8299 <= WX8298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8301 <= 0;
  else
    WX8301 <= WX8300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8303 <= 0;
  else
    WX8303 <= WX8302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8305 <= 0;
  else
    WX8305 <= WX8304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8403 <= 0;
  else
    WX8403 <= WX8402;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8405 <= 0;
  else
    WX8405 <= WX8404;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8407 <= 0;
  else
    WX8407 <= WX8406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8409 <= 0;
  else
    WX8409 <= WX8408;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8411 <= 0;
  else
    WX8411 <= WX8410;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8413 <= 0;
  else
    WX8413 <= WX8412;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8415 <= 0;
  else
    WX8415 <= WX8414;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8417 <= 0;
  else
    WX8417 <= WX8416;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8419 <= 0;
  else
    WX8419 <= WX8418;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8421 <= 0;
  else
    WX8421 <= WX8420;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8423 <= 0;
  else
    WX8423 <= WX8422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8425 <= 0;
  else
    WX8425 <= WX8424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8427 <= 0;
  else
    WX8427 <= WX8426;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8429 <= 0;
  else
    WX8429 <= WX8428;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8431 <= 0;
  else
    WX8431 <= WX8430;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8433 <= 0;
  else
    WX8433 <= WX8432;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8435 <= 0;
  else
    WX8435 <= WX8434;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8437 <= 0;
  else
    WX8437 <= WX8436;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8439 <= 0;
  else
    WX8439 <= WX8438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8441 <= 0;
  else
    WX8441 <= WX8440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8443 <= 0;
  else
    WX8443 <= WX8442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8445 <= 0;
  else
    WX8445 <= WX8444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8447 <= 0;
  else
    WX8447 <= WX8446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8449 <= 0;
  else
    WX8449 <= WX8448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8451 <= 0;
  else
    WX8451 <= WX8450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8453 <= 0;
  else
    WX8453 <= WX8452;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8455 <= 0;
  else
    WX8455 <= WX8454;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8457 <= 0;
  else
    WX8457 <= WX8456;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8459 <= 0;
  else
    WX8459 <= WX8458;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8461 <= 0;
  else
    WX8461 <= WX8460;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8463 <= 0;
  else
    WX8463 <= WX8462;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8465 <= 0;
  else
    WX8465 <= WX8464;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8467 <= 0;
  else
    WX8467 <= WX8466;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8469 <= 0;
  else
    WX8469 <= WX8468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8471 <= 0;
  else
    WX8471 <= WX8470;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8473 <= 0;
  else
    WX8473 <= WX8472;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8475 <= 0;
  else
    WX8475 <= WX8474;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8477 <= 0;
  else
    WX8477 <= WX8476;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8479 <= 0;
  else
    WX8479 <= WX8478;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8481 <= 0;
  else
    WX8481 <= WX8480;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8483 <= 0;
  else
    WX8483 <= WX8482;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8485 <= 0;
  else
    WX8485 <= WX8484;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8487 <= 0;
  else
    WX8487 <= WX8486;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8489 <= 0;
  else
    WX8489 <= WX8488;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8491 <= 0;
  else
    WX8491 <= WX8490;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8493 <= 0;
  else
    WX8493 <= WX8492;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8495 <= 0;
  else
    WX8495 <= WX8494;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8497 <= 0;
  else
    WX8497 <= WX8496;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8499 <= 0;
  else
    WX8499 <= WX8498;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8501 <= 0;
  else
    WX8501 <= WX8500;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8503 <= 0;
  else
    WX8503 <= WX8502;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8505 <= 0;
  else
    WX8505 <= WX8504;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8507 <= 0;
  else
    WX8507 <= WX8506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8509 <= 0;
  else
    WX8509 <= WX8508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8511 <= 0;
  else
    WX8511 <= WX8510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8513 <= 0;
  else
    WX8513 <= WX8512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8515 <= 0;
  else
    WX8515 <= WX8514;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8517 <= 0;
  else
    WX8517 <= WX8516;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8519 <= 0;
  else
    WX8519 <= WX8518;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8521 <= 0;
  else
    WX8521 <= WX8520;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8523 <= 0;
  else
    WX8523 <= WX8522;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8525 <= 0;
  else
    WX8525 <= WX8524;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8527 <= 0;
  else
    WX8527 <= WX8526;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8529 <= 0;
  else
    WX8529 <= WX8528;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8531 <= 0;
  else
    WX8531 <= WX8530;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8533 <= 0;
  else
    WX8533 <= WX8532;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8535 <= 0;
  else
    WX8535 <= WX8534;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8537 <= 0;
  else
    WX8537 <= WX8536;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8539 <= 0;
  else
    WX8539 <= WX8538;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8541 <= 0;
  else
    WX8541 <= WX8540;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8543 <= 0;
  else
    WX8543 <= WX8542;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8545 <= 0;
  else
    WX8545 <= WX8544;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8547 <= 0;
  else
    WX8547 <= WX8546;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8549 <= 0;
  else
    WX8549 <= WX8548;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8551 <= 0;
  else
    WX8551 <= WX8550;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8553 <= 0;
  else
    WX8553 <= WX8552;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8555 <= 0;
  else
    WX8555 <= WX8554;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8557 <= 0;
  else
    WX8557 <= WX8556;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8559 <= 0;
  else
    WX8559 <= WX8558;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8561 <= 0;
  else
    WX8561 <= WX8560;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8563 <= 0;
  else
    WX8563 <= WX8562;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8565 <= 0;
  else
    WX8565 <= WX8564;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8567 <= 0;
  else
    WX8567 <= WX8566;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8569 <= 0;
  else
    WX8569 <= WX8568;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8571 <= 0;
  else
    WX8571 <= WX8570;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8573 <= 0;
  else
    WX8573 <= WX8572;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8575 <= 0;
  else
    WX8575 <= WX8574;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8577 <= 0;
  else
    WX8577 <= WX8576;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8579 <= 0;
  else
    WX8579 <= WX8578;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8581 <= 0;
  else
    WX8581 <= WX8580;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8583 <= 0;
  else
    WX8583 <= WX8582;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8585 <= 0;
  else
    WX8585 <= WX8584;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8587 <= 0;
  else
    WX8587 <= WX8586;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8589 <= 0;
  else
    WX8589 <= WX8588;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8591 <= 0;
  else
    WX8591 <= WX8590;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8593 <= 0;
  else
    WX8593 <= WX8592;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8595 <= 0;
  else
    WX8595 <= WX8594;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8597 <= 0;
  else
    WX8597 <= WX8596;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8599 <= 0;
  else
    WX8599 <= WX8598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8601 <= 0;
  else
    WX8601 <= WX8600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8603 <= 0;
  else
    WX8603 <= WX8602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8605 <= 0;
  else
    WX8605 <= WX8604;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8607 <= 0;
  else
    WX8607 <= WX8606;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8609 <= 0;
  else
    WX8609 <= WX8608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8611 <= 0;
  else
    WX8611 <= WX8610;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8613 <= 0;
  else
    WX8613 <= WX8612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8615 <= 0;
  else
    WX8615 <= WX8614;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8617 <= 0;
  else
    WX8617 <= WX8616;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8619 <= 0;
  else
    WX8619 <= WX8618;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8621 <= 0;
  else
    WX8621 <= WX8620;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8623 <= 0;
  else
    WX8623 <= WX8622;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8625 <= 0;
  else
    WX8625 <= WX8624;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8627 <= 0;
  else
    WX8627 <= WX8626;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8629 <= 0;
  else
    WX8629 <= WX8628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8631 <= 0;
  else
    WX8631 <= WX8630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8633 <= 0;
  else
    WX8633 <= WX8632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8635 <= 0;
  else
    WX8635 <= WX8634;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8637 <= 0;
  else
    WX8637 <= WX8636;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8639 <= 0;
  else
    WX8639 <= WX8638;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8641 <= 0;
  else
    WX8641 <= WX8640;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8643 <= 0;
  else
    WX8643 <= WX8642;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8645 <= 0;
  else
    WX8645 <= WX8644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8647 <= 0;
  else
    WX8647 <= WX8646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8649 <= 0;
  else
    WX8649 <= WX8648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8651 <= 0;
  else
    WX8651 <= WX8650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8653 <= 0;
  else
    WX8653 <= WX8652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8655 <= 0;
  else
    WX8655 <= WX8654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX8657 <= 0;
  else
    WX8657 <= WX8656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2269_ <= 0;
  else
    _2269_ <= WX9022;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2270_ <= 0;
  else
    _2270_ <= WX9024;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2271_ <= 0;
  else
    _2271_ <= WX9026;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2272_ <= 0;
  else
    _2272_ <= WX9028;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2273_ <= 0;
  else
    _2273_ <= WX9030;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2274_ <= 0;
  else
    _2274_ <= WX9032;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2275_ <= 0;
  else
    _2275_ <= WX9034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2276_ <= 0;
  else
    _2276_ <= WX9036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2277_ <= 0;
  else
    _2277_ <= WX9038;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2278_ <= 0;
  else
    _2278_ <= WX9040;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2279_ <= 0;
  else
    _2279_ <= WX9042;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2280_ <= 0;
  else
    _2280_ <= WX9044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2281_ <= 0;
  else
    _2281_ <= WX9046;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2282_ <= 0;
  else
    _2282_ <= WX9048;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2283_ <= 0;
  else
    _2283_ <= WX9050;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2284_ <= 0;
  else
    _2284_ <= WX9052;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2285_ <= 0;
  else
    _2285_ <= WX9054;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2286_ <= 0;
  else
    _2286_ <= WX9056;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2287_ <= 0;
  else
    _2287_ <= WX9058;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2288_ <= 0;
  else
    _2288_ <= WX9060;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2289_ <= 0;
  else
    _2289_ <= WX9062;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2290_ <= 0;
  else
    _2290_ <= WX9064;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2291_ <= 0;
  else
    _2291_ <= WX9066;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2292_ <= 0;
  else
    _2292_ <= WX9068;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2293_ <= 0;
  else
    _2293_ <= WX9070;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2294_ <= 0;
  else
    _2294_ <= WX9072;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2295_ <= 0;
  else
    _2295_ <= WX9074;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2296_ <= 0;
  else
    _2296_ <= WX9076;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2297_ <= 0;
  else
    _2297_ <= WX9078;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2298_ <= 0;
  else
    _2298_ <= WX9080;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2299_ <= 0;
  else
    _2299_ <= WX9082;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2300_ <= 0;
  else
    _2300_ <= WX9084;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9536 <= 0;
  else
    WX9536 <= WX9535;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9538 <= 0;
  else
    WX9538 <= WX9537;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9540 <= 0;
  else
    WX9540 <= WX9539;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9542 <= 0;
  else
    WX9542 <= WX9541;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9544 <= 0;
  else
    WX9544 <= WX9543;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9546 <= 0;
  else
    WX9546 <= WX9545;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9548 <= 0;
  else
    WX9548 <= WX9547;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9550 <= 0;
  else
    WX9550 <= WX9549;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9552 <= 0;
  else
    WX9552 <= WX9551;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9554 <= 0;
  else
    WX9554 <= WX9553;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9556 <= 0;
  else
    WX9556 <= WX9555;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9558 <= 0;
  else
    WX9558 <= WX9557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9560 <= 0;
  else
    WX9560 <= WX9559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9562 <= 0;
  else
    WX9562 <= WX9561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9564 <= 0;
  else
    WX9564 <= WX9563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9566 <= 0;
  else
    WX9566 <= WX9565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9568 <= 0;
  else
    WX9568 <= WX9567;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9570 <= 0;
  else
    WX9570 <= WX9569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9572 <= 0;
  else
    WX9572 <= WX9571;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9574 <= 0;
  else
    WX9574 <= WX9573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9576 <= 0;
  else
    WX9576 <= WX9575;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9578 <= 0;
  else
    WX9578 <= WX9577;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9580 <= 0;
  else
    WX9580 <= WX9579;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9582 <= 0;
  else
    WX9582 <= WX9581;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9584 <= 0;
  else
    WX9584 <= WX9583;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9586 <= 0;
  else
    WX9586 <= WX9585;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9588 <= 0;
  else
    WX9588 <= WX9587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9590 <= 0;
  else
    WX9590 <= WX9589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9592 <= 0;
  else
    WX9592 <= WX9591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9594 <= 0;
  else
    WX9594 <= WX9593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9596 <= 0;
  else
    WX9596 <= WX9595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9598 <= 0;
  else
    WX9598 <= WX9597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9696 <= 0;
  else
    WX9696 <= WX9695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9698 <= 0;
  else
    WX9698 <= WX9697;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9700 <= 0;
  else
    WX9700 <= WX9699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9702 <= 0;
  else
    WX9702 <= WX9701;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9704 <= 0;
  else
    WX9704 <= WX9703;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9706 <= 0;
  else
    WX9706 <= WX9705;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9708 <= 0;
  else
    WX9708 <= WX9707;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9710 <= 0;
  else
    WX9710 <= WX9709;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9712 <= 0;
  else
    WX9712 <= WX9711;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9714 <= 0;
  else
    WX9714 <= WX9713;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9716 <= 0;
  else
    WX9716 <= WX9715;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9718 <= 0;
  else
    WX9718 <= WX9717;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9720 <= 0;
  else
    WX9720 <= WX9719;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9722 <= 0;
  else
    WX9722 <= WX9721;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9724 <= 0;
  else
    WX9724 <= WX9723;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9726 <= 0;
  else
    WX9726 <= WX9725;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9728 <= 0;
  else
    WX9728 <= WX9727;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9730 <= 0;
  else
    WX9730 <= WX9729;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9732 <= 0;
  else
    WX9732 <= WX9731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9734 <= 0;
  else
    WX9734 <= WX9733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9736 <= 0;
  else
    WX9736 <= WX9735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9738 <= 0;
  else
    WX9738 <= WX9737;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9740 <= 0;
  else
    WX9740 <= WX9739;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9742 <= 0;
  else
    WX9742 <= WX9741;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9744 <= 0;
  else
    WX9744 <= WX9743;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9746 <= 0;
  else
    WX9746 <= WX9745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9748 <= 0;
  else
    WX9748 <= WX9747;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9750 <= 0;
  else
    WX9750 <= WX9749;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9752 <= 0;
  else
    WX9752 <= WX9751;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9754 <= 0;
  else
    WX9754 <= WX9753;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9756 <= 0;
  else
    WX9756 <= WX9755;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9758 <= 0;
  else
    WX9758 <= WX9757;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9760 <= 0;
  else
    WX9760 <= WX9759;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9762 <= 0;
  else
    WX9762 <= WX9761;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9764 <= 0;
  else
    WX9764 <= WX9763;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9766 <= 0;
  else
    WX9766 <= WX9765;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9768 <= 0;
  else
    WX9768 <= WX9767;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9770 <= 0;
  else
    WX9770 <= WX9769;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9772 <= 0;
  else
    WX9772 <= WX9771;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9774 <= 0;
  else
    WX9774 <= WX9773;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9776 <= 0;
  else
    WX9776 <= WX9775;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9778 <= 0;
  else
    WX9778 <= WX9777;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9780 <= 0;
  else
    WX9780 <= WX9779;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9782 <= 0;
  else
    WX9782 <= WX9781;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9784 <= 0;
  else
    WX9784 <= WX9783;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9786 <= 0;
  else
    WX9786 <= WX9785;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9788 <= 0;
  else
    WX9788 <= WX9787;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9790 <= 0;
  else
    WX9790 <= WX9789;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9792 <= 0;
  else
    WX9792 <= WX9791;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9794 <= 0;
  else
    WX9794 <= WX9793;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9796 <= 0;
  else
    WX9796 <= WX9795;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9798 <= 0;
  else
    WX9798 <= WX9797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9800 <= 0;
  else
    WX9800 <= WX9799;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9802 <= 0;
  else
    WX9802 <= WX9801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9804 <= 0;
  else
    WX9804 <= WX9803;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9806 <= 0;
  else
    WX9806 <= WX9805;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9808 <= 0;
  else
    WX9808 <= WX9807;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9810 <= 0;
  else
    WX9810 <= WX9809;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9812 <= 0;
  else
    WX9812 <= WX9811;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9814 <= 0;
  else
    WX9814 <= WX9813;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9816 <= 0;
  else
    WX9816 <= WX9815;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9818 <= 0;
  else
    WX9818 <= WX9817;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9820 <= 0;
  else
    WX9820 <= WX9819;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9822 <= 0;
  else
    WX9822 <= WX9821;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9824 <= 0;
  else
    WX9824 <= WX9823;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9826 <= 0;
  else
    WX9826 <= WX9825;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9828 <= 0;
  else
    WX9828 <= WX9827;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9830 <= 0;
  else
    WX9830 <= WX9829;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9832 <= 0;
  else
    WX9832 <= WX9831;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9834 <= 0;
  else
    WX9834 <= WX9833;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9836 <= 0;
  else
    WX9836 <= WX9835;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9838 <= 0;
  else
    WX9838 <= WX9837;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9840 <= 0;
  else
    WX9840 <= WX9839;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9842 <= 0;
  else
    WX9842 <= WX9841;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9844 <= 0;
  else
    WX9844 <= WX9843;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9846 <= 0;
  else
    WX9846 <= WX9845;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9848 <= 0;
  else
    WX9848 <= WX9847;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9850 <= 0;
  else
    WX9850 <= WX9849;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9852 <= 0;
  else
    WX9852 <= WX9851;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9854 <= 0;
  else
    WX9854 <= WX9853;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9856 <= 0;
  else
    WX9856 <= WX9855;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9858 <= 0;
  else
    WX9858 <= WX9857;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9860 <= 0;
  else
    WX9860 <= WX9859;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9862 <= 0;
  else
    WX9862 <= WX9861;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9864 <= 0;
  else
    WX9864 <= WX9863;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9866 <= 0;
  else
    WX9866 <= WX9865;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9868 <= 0;
  else
    WX9868 <= WX9867;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9870 <= 0;
  else
    WX9870 <= WX9869;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9872 <= 0;
  else
    WX9872 <= WX9871;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9874 <= 0;
  else
    WX9874 <= WX9873;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9876 <= 0;
  else
    WX9876 <= WX9875;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9878 <= 0;
  else
    WX9878 <= WX9877;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9880 <= 0;
  else
    WX9880 <= WX9879;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9882 <= 0;
  else
    WX9882 <= WX9881;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9884 <= 0;
  else
    WX9884 <= WX9883;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9886 <= 0;
  else
    WX9886 <= WX9885;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9888 <= 0;
  else
    WX9888 <= WX9887;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9890 <= 0;
  else
    WX9890 <= WX9889;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9892 <= 0;
  else
    WX9892 <= WX9891;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9894 <= 0;
  else
    WX9894 <= WX9893;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9896 <= 0;
  else
    WX9896 <= WX9895;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9898 <= 0;
  else
    WX9898 <= WX9897;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9900 <= 0;
  else
    WX9900 <= WX9899;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9902 <= 0;
  else
    WX9902 <= WX9901;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9904 <= 0;
  else
    WX9904 <= WX9903;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9906 <= 0;
  else
    WX9906 <= WX9905;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9908 <= 0;
  else
    WX9908 <= WX9907;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9910 <= 0;
  else
    WX9910 <= WX9909;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9912 <= 0;
  else
    WX9912 <= WX9911;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9914 <= 0;
  else
    WX9914 <= WX9913;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9916 <= 0;
  else
    WX9916 <= WX9915;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9918 <= 0;
  else
    WX9918 <= WX9917;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9920 <= 0;
  else
    WX9920 <= WX9919;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9922 <= 0;
  else
    WX9922 <= WX9921;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9924 <= 0;
  else
    WX9924 <= WX9923;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9926 <= 0;
  else
    WX9926 <= WX9925;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9928 <= 0;
  else
    WX9928 <= WX9927;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9930 <= 0;
  else
    WX9930 <= WX9929;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9932 <= 0;
  else
    WX9932 <= WX9931;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9934 <= 0;
  else
    WX9934 <= WX9933;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9936 <= 0;
  else
    WX9936 <= WX9935;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9938 <= 0;
  else
    WX9938 <= WX9937;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9940 <= 0;
  else
    WX9940 <= WX9939;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9942 <= 0;
  else
    WX9942 <= WX9941;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9944 <= 0;
  else
    WX9944 <= WX9943;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9946 <= 0;
  else
    WX9946 <= WX9945;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9948 <= 0;
  else
    WX9948 <= WX9947;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX9950 <= 0;
  else
    WX9950 <= WX9949;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2301_ <= 0;
  else
    _2301_ <= WX10315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2302_ <= 0;
  else
    _2302_ <= WX10317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2303_ <= 0;
  else
    _2303_ <= WX10319;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2304_ <= 0;
  else
    _2304_ <= WX10321;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2305_ <= 0;
  else
    _2305_ <= WX10323;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2306_ <= 0;
  else
    _2306_ <= WX10325;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2307_ <= 0;
  else
    _2307_ <= WX10327;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2308_ <= 0;
  else
    _2308_ <= WX10329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2309_ <= 0;
  else
    _2309_ <= WX10331;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2310_ <= 0;
  else
    _2310_ <= WX10333;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2311_ <= 0;
  else
    _2311_ <= WX10335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2312_ <= 0;
  else
    _2312_ <= WX10337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2313_ <= 0;
  else
    _2313_ <= WX10339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2314_ <= 0;
  else
    _2314_ <= WX10341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2315_ <= 0;
  else
    _2315_ <= WX10343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2316_ <= 0;
  else
    _2316_ <= WX10345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2317_ <= 0;
  else
    _2317_ <= WX10347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2318_ <= 0;
  else
    _2318_ <= WX10349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2319_ <= 0;
  else
    _2319_ <= WX10351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2320_ <= 0;
  else
    _2320_ <= WX10353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2321_ <= 0;
  else
    _2321_ <= WX10355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2322_ <= 0;
  else
    _2322_ <= WX10357;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2323_ <= 0;
  else
    _2323_ <= WX10359;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2324_ <= 0;
  else
    _2324_ <= WX10361;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2325_ <= 0;
  else
    _2325_ <= WX10363;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2326_ <= 0;
  else
    _2326_ <= WX10365;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2327_ <= 0;
  else
    _2327_ <= WX10367;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2328_ <= 0;
  else
    _2328_ <= WX10369;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2329_ <= 0;
  else
    _2329_ <= WX10371;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2330_ <= 0;
  else
    _2330_ <= WX10373;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2331_ <= 0;
  else
    _2331_ <= WX10375;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2332_ <= 0;
  else
    _2332_ <= WX10377;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10829 <= 0;
  else
    WX10829 <= WX10828;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10831 <= 0;
  else
    WX10831 <= WX10830;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10833 <= 0;
  else
    WX10833 <= WX10832;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10835 <= 0;
  else
    WX10835 <= WX10834;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10837 <= 0;
  else
    WX10837 <= WX10836;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10839 <= 0;
  else
    WX10839 <= WX10838;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10841 <= 0;
  else
    WX10841 <= WX10840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10843 <= 0;
  else
    WX10843 <= WX10842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10845 <= 0;
  else
    WX10845 <= WX10844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10847 <= 0;
  else
    WX10847 <= WX10846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10849 <= 0;
  else
    WX10849 <= WX10848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10851 <= 0;
  else
    WX10851 <= WX10850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10853 <= 0;
  else
    WX10853 <= WX10852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10855 <= 0;
  else
    WX10855 <= WX10854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10857 <= 0;
  else
    WX10857 <= WX10856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10859 <= 0;
  else
    WX10859 <= WX10858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10861 <= 0;
  else
    WX10861 <= WX10860;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10863 <= 0;
  else
    WX10863 <= WX10862;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10865 <= 0;
  else
    WX10865 <= WX10864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10867 <= 0;
  else
    WX10867 <= WX10866;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10869 <= 0;
  else
    WX10869 <= WX10868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10871 <= 0;
  else
    WX10871 <= WX10870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10873 <= 0;
  else
    WX10873 <= WX10872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10875 <= 0;
  else
    WX10875 <= WX10874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10877 <= 0;
  else
    WX10877 <= WX10876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10879 <= 0;
  else
    WX10879 <= WX10878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10881 <= 0;
  else
    WX10881 <= WX10880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10883 <= 0;
  else
    WX10883 <= WX10882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10885 <= 0;
  else
    WX10885 <= WX10884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10887 <= 0;
  else
    WX10887 <= WX10886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10889 <= 0;
  else
    WX10889 <= WX10888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10891 <= 0;
  else
    WX10891 <= WX10890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10989 <= 0;
  else
    WX10989 <= WX10988;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10991 <= 0;
  else
    WX10991 <= WX10990;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10993 <= 0;
  else
    WX10993 <= WX10992;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10995 <= 0;
  else
    WX10995 <= WX10994;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10997 <= 0;
  else
    WX10997 <= WX10996;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX10999 <= 0;
  else
    WX10999 <= WX10998;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11001 <= 0;
  else
    WX11001 <= WX11000;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11003 <= 0;
  else
    WX11003 <= WX11002;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11005 <= 0;
  else
    WX11005 <= WX11004;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11007 <= 0;
  else
    WX11007 <= WX11006;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11009 <= 0;
  else
    WX11009 <= WX11008;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11011 <= 0;
  else
    WX11011 <= WX11010;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11013 <= 0;
  else
    WX11013 <= WX11012;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11015 <= 0;
  else
    WX11015 <= WX11014;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11017 <= 0;
  else
    WX11017 <= WX11016;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11019 <= 0;
  else
    WX11019 <= WX11018;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11021 <= 0;
  else
    WX11021 <= WX11020;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11023 <= 0;
  else
    WX11023 <= WX11022;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11025 <= 0;
  else
    WX11025 <= WX11024;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11027 <= 0;
  else
    WX11027 <= WX11026;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11029 <= 0;
  else
    WX11029 <= WX11028;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11031 <= 0;
  else
    WX11031 <= WX11030;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11033 <= 0;
  else
    WX11033 <= WX11032;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11035 <= 0;
  else
    WX11035 <= WX11034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11037 <= 0;
  else
    WX11037 <= WX11036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11039 <= 0;
  else
    WX11039 <= WX11038;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11041 <= 0;
  else
    WX11041 <= WX11040;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11043 <= 0;
  else
    WX11043 <= WX11042;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11045 <= 0;
  else
    WX11045 <= WX11044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11047 <= 0;
  else
    WX11047 <= WX11046;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11049 <= 0;
  else
    WX11049 <= WX11048;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11051 <= 0;
  else
    WX11051 <= WX11050;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11053 <= 0;
  else
    WX11053 <= WX11052;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11055 <= 0;
  else
    WX11055 <= WX11054;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11057 <= 0;
  else
    WX11057 <= WX11056;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11059 <= 0;
  else
    WX11059 <= WX11058;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11061 <= 0;
  else
    WX11061 <= WX11060;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11063 <= 0;
  else
    WX11063 <= WX11062;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11065 <= 0;
  else
    WX11065 <= WX11064;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11067 <= 0;
  else
    WX11067 <= WX11066;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11069 <= 0;
  else
    WX11069 <= WX11068;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11071 <= 0;
  else
    WX11071 <= WX11070;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11073 <= 0;
  else
    WX11073 <= WX11072;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11075 <= 0;
  else
    WX11075 <= WX11074;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11077 <= 0;
  else
    WX11077 <= WX11076;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11079 <= 0;
  else
    WX11079 <= WX11078;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11081 <= 0;
  else
    WX11081 <= WX11080;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11083 <= 0;
  else
    WX11083 <= WX11082;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11085 <= 0;
  else
    WX11085 <= WX11084;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11087 <= 0;
  else
    WX11087 <= WX11086;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11089 <= 0;
  else
    WX11089 <= WX11088;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11091 <= 0;
  else
    WX11091 <= WX11090;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11093 <= 0;
  else
    WX11093 <= WX11092;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11095 <= 0;
  else
    WX11095 <= WX11094;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11097 <= 0;
  else
    WX11097 <= WX11096;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11099 <= 0;
  else
    WX11099 <= WX11098;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11101 <= 0;
  else
    WX11101 <= WX11100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11103 <= 0;
  else
    WX11103 <= WX11102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11105 <= 0;
  else
    WX11105 <= WX11104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11107 <= 0;
  else
    WX11107 <= WX11106;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11109 <= 0;
  else
    WX11109 <= WX11108;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11111 <= 0;
  else
    WX11111 <= WX11110;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11113 <= 0;
  else
    WX11113 <= WX11112;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11115 <= 0;
  else
    WX11115 <= WX11114;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11117 <= 0;
  else
    WX11117 <= WX11116;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11119 <= 0;
  else
    WX11119 <= WX11118;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11121 <= 0;
  else
    WX11121 <= WX11120;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11123 <= 0;
  else
    WX11123 <= WX11122;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11125 <= 0;
  else
    WX11125 <= WX11124;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11127 <= 0;
  else
    WX11127 <= WX11126;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11129 <= 0;
  else
    WX11129 <= WX11128;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11131 <= 0;
  else
    WX11131 <= WX11130;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11133 <= 0;
  else
    WX11133 <= WX11132;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11135 <= 0;
  else
    WX11135 <= WX11134;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11137 <= 0;
  else
    WX11137 <= WX11136;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11139 <= 0;
  else
    WX11139 <= WX11138;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11141 <= 0;
  else
    WX11141 <= WX11140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11143 <= 0;
  else
    WX11143 <= WX11142;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11145 <= 0;
  else
    WX11145 <= WX11144;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11147 <= 0;
  else
    WX11147 <= WX11146;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11149 <= 0;
  else
    WX11149 <= WX11148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11151 <= 0;
  else
    WX11151 <= WX11150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11153 <= 0;
  else
    WX11153 <= WX11152;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11155 <= 0;
  else
    WX11155 <= WX11154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11157 <= 0;
  else
    WX11157 <= WX11156;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11159 <= 0;
  else
    WX11159 <= WX11158;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11161 <= 0;
  else
    WX11161 <= WX11160;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11163 <= 0;
  else
    WX11163 <= WX11162;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11165 <= 0;
  else
    WX11165 <= WX11164;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11167 <= 0;
  else
    WX11167 <= WX11166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11169 <= 0;
  else
    WX11169 <= WX11168;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11171 <= 0;
  else
    WX11171 <= WX11170;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11173 <= 0;
  else
    WX11173 <= WX11172;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11175 <= 0;
  else
    WX11175 <= WX11174;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11177 <= 0;
  else
    WX11177 <= WX11176;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11179 <= 0;
  else
    WX11179 <= WX11178;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11181 <= 0;
  else
    WX11181 <= WX11180;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11183 <= 0;
  else
    WX11183 <= WX11182;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11185 <= 0;
  else
    WX11185 <= WX11184;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11187 <= 0;
  else
    WX11187 <= WX11186;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11189 <= 0;
  else
    WX11189 <= WX11188;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11191 <= 0;
  else
    WX11191 <= WX11190;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11193 <= 0;
  else
    WX11193 <= WX11192;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11195 <= 0;
  else
    WX11195 <= WX11194;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11197 <= 0;
  else
    WX11197 <= WX11196;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11199 <= 0;
  else
    WX11199 <= WX11198;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11201 <= 0;
  else
    WX11201 <= WX11200;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11203 <= 0;
  else
    WX11203 <= WX11202;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11205 <= 0;
  else
    WX11205 <= WX11204;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11207 <= 0;
  else
    WX11207 <= WX11206;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11209 <= 0;
  else
    WX11209 <= WX11208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11211 <= 0;
  else
    WX11211 <= WX11210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11213 <= 0;
  else
    WX11213 <= WX11212;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11215 <= 0;
  else
    WX11215 <= WX11214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11217 <= 0;
  else
    WX11217 <= WX11216;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11219 <= 0;
  else
    WX11219 <= WX11218;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11221 <= 0;
  else
    WX11221 <= WX11220;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11223 <= 0;
  else
    WX11223 <= WX11222;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11225 <= 0;
  else
    WX11225 <= WX11224;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11227 <= 0;
  else
    WX11227 <= WX11226;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11229 <= 0;
  else
    WX11229 <= WX11228;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11231 <= 0;
  else
    WX11231 <= WX11230;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11233 <= 0;
  else
    WX11233 <= WX11232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11235 <= 0;
  else
    WX11235 <= WX11234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11237 <= 0;
  else
    WX11237 <= WX11236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11239 <= 0;
  else
    WX11239 <= WX11238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11241 <= 0;
  else
    WX11241 <= WX11240;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    WX11243 <= 0;
  else
    WX11243 <= WX11242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2333_ <= 0;
  else
    _2333_ <= WX11608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2334_ <= 0;
  else
    _2334_ <= WX11610;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2335_ <= 0;
  else
    _2335_ <= WX11612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2336_ <= 0;
  else
    _2336_ <= WX11614;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2337_ <= 0;
  else
    _2337_ <= WX11616;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2338_ <= 0;
  else
    _2338_ <= WX11618;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2339_ <= 0;
  else
    _2339_ <= WX11620;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2340_ <= 0;
  else
    _2340_ <= WX11622;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2341_ <= 0;
  else
    _2341_ <= WX11624;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2342_ <= 0;
  else
    _2342_ <= WX11626;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2343_ <= 0;
  else
    _2343_ <= WX11628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2344_ <= 0;
  else
    _2344_ <= WX11630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2345_ <= 0;
  else
    _2345_ <= WX11632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2346_ <= 0;
  else
    _2346_ <= WX11634;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2347_ <= 0;
  else
    _2347_ <= WX11636;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2348_ <= 0;
  else
    _2348_ <= WX11638;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2349_ <= 0;
  else
    _2349_ <= WX11640;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2350_ <= 0;
  else
    _2350_ <= WX11642;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2351_ <= 0;
  else
    _2351_ <= WX11644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2352_ <= 0;
  else
    _2352_ <= WX11646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2353_ <= 0;
  else
    _2353_ <= WX11648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2354_ <= 0;
  else
    _2354_ <= WX11650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2355_ <= 0;
  else
    _2355_ <= WX11652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2356_ <= 0;
  else
    _2356_ <= WX11654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2357_ <= 0;
  else
    _2357_ <= WX11656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2358_ <= 0;
  else
    _2358_ <= WX11658;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2359_ <= 0;
  else
    _2359_ <= WX11660;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2360_ <= 0;
  else
    _2360_ <= WX11662;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2361_ <= 0;
  else
    _2361_ <= WX11664;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2362_ <= 0;
  else
    _2362_ <= WX11666;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2363_ <= 0;
  else
    _2363_ <= WX11668;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _2364_ <= 0;
  else
    _2364_ <= WX11670;
assign II22507 = ((~II22517))|((~II22518));
assign II26071 = ((~II26047))|((~II26063));
assign WX6414 = ((~II19591))|((~II19592));
assign II22128 = ((~II22104))|((~II22120));
assign II6147 = ((~II6149))|((~II6150));
assign WX9613 = ((~WX10044));
assign WX7987 = ((~WX7978));
assign II26918 = ((~WX8760))|((~II26917));
assign WX2450 = (WX2448)|(WX2447);
assign II2229 = ((~II2219))|((~II2227));
assign II30149 = ((~WX9704))|((~II30147));
assign II2963 = ((~II2965))|((~II2966));
assign WX8188 = (WX8186)|(WX8185);
assign II30497 = ((~II30487))|((~II30495));
assign WX3931 = (WX3929)|(WX3928);
assign WX7670 = ((~WX7470));
assign WX6302 = ((~WX6301));
assign II15655 = ((~WX4509))|((~_2185_));
assign WX2888 = (WX2894&WX2889);
assign II19689 = ((~WX5807))|((~II19688));
assign II22743 = ((~WX7348))|((~II22741));
assign WX4303 = (WX4301)|(WX4300);
assign WX10189 = ((~WX10188));
assign II22919 = ((~WX7232))|((~II22911));
assign WX3340 = (WX3277&RESET);
assign WX6164 = ((~WX6086));
assign WX239 = (WX513&WX1004);
assign WX2459 = ((~WX2458));
assign WX330 = (WX336&WX331);
assign WX5710 = (WX5713&RESET);
assign II2018 = ((~II2020))|((~II2021));
assign II3642 = ((~_2089_))|((~II3640));
assign II26018 = ((~WX8759))|((~WX8403));
assign II15405 = ((~WX4485))|((~WX4416));
assign II15147 = ((~WX4376))|((~II15145));
assign WX9021 = ((~WX8988));
assign WX9060 = (WX9005&WX9021);
assign II2144 = ((~WX1001))|((~II2143));
assign WX615 = ((~WX843));
assign WX2904 = (WX2902)|(WX2901);
assign II34120 = ((~II34122))|((~II34123));
assign WX8882 = ((~WX8881));
assign WX1732 = ((~WX1723));
assign WX5365 = (_2225_&WX6176);
assign WX8975 = (WX8974&WX8763);
assign WX5343 = ((~WX6176));
assign II2492 = ((~WX741))|((~II2491));
assign II14615 = ((~II14590))|((~II14614));
assign WX516 = (WX519&RESET);
assign WX11312 = ((~WX11246));
assign WX1466 = ((~WX1457));
assign WX3563 = ((~WX3562));
assign WX8062 = (WX8060)|(WX8059);
assign WX4905 = ((~WX4904));
assign WX2751 = (_2163_&WX3590);
assign WX7523 = ((~WX7470));
assign WX1607 = ((~WX1606));
assign II14260 = ((~II14250))|((~II14258));
assign II34743 = ((~WX11035))|((~II34741));
assign WX1525 = (WX1531&WX1526);
assign WX9603 = ((~WX10024));
assign II19294 = ((~WX5769))|((~II19293));
assign II19696 = ((~WX5808))|((~II19695));
assign II30287 = ((~WX9840))|((~II30286));
assign II30045 = ((~II30021))|((~II30037));
assign WX3734 = (WX3186&WX3735);
assign WX1406 = (WX1788&WX2297);
assign WX8364 = ((~WX8332));
assign II10585 = ((~II10595))|((~II10596));
assign WX11054 = (WX10991&RESET);
assign II34796 = ((~II34786))|((~II34794));
assign II14826 = ((~WX4768))|((~II14824));
assign WX4953 = ((~WX4952));
assign II14222 = ((~WX4538))|((~II14220));
assign II10239 = ((~II10229))|((~II10237));
assign II2499 = ((~WX805))|((~WX869));
assign II1988 = ((~WX1001))|((~WX645));
assign WX628 = ((~WX869));
assign II26172 = ((~II26174))|((~II26175));
assign II26856 = ((~WX8760))|((~II26855));
assign II19682 = ((~WX5806))|((~II19681));
assign WX268 = (DATA_9_15&WX269);
assign WX8837 = ((~WX8763));
assign II10315 = ((~WX3315))|((~II10307));
assign II30248 = ((~WX9774))|((~II30247));
assign II26252 = ((~WX8609))|((~II26250));
assign II7562 = ((~WX1910))|((~II7561));
assign WX8313 = ((~WX8737));
assign WX8793 = (WX8792&WX8763);
assign II30929 = ((~WX9818))|((~II30921));
assign WX2627 = ((~WX3590));
assign WX4973 = (WX4971)|(WX4970);
assign II34098 = ((~WX11057))|((~II34097));
assign WX388 = (WX386)|(WX385);
assign WX11574 = ((~RESET));
assign WX11360 = ((~WX11349));
assign WX2993 = (WX3123&WX3590);
assign WX11558 = ((~WX11557));
assign II26791 = ((~II26801))|((~II26802));
assign II27699 = ((~WX8393))|((~II27698));
assign II15587 = ((~_2196_))|((~II15585));
assign WX10544 = (WX10542)|(WX10541);
assign WX7501 = (WX7049&WX7502);
assign WX9283 = (WX9289&WX9284);
assign WX10599 = ((~WX11348));
assign WX10618 = (WX10624&WX10619);
assign WX4974 = ((~WX4973));
assign WX153 = ((~WX1004));
assign II2436 = ((~II2438))|((~II2439));
assign WX7151 = (WX6807&RESET);
assign II34975 = ((~WX11241))|((~II34973));
assign II30419 = ((~II30409))|((~II30417));
assign WX5271 = (WX5665&WX6176);
assign II18597 = ((~WX6174))|((~WX5855));
assign WX5460 = (WX5466&WX5461);
assign II18093 = ((~II18068))|((~II18092));
assign WX4967 = ((~WX4966));
assign WX8768 = (WX8766)|(WX8765);
assign II34167 = ((~WX11125))|((~WX11189));
assign WX11251 = ((~II34268))|((~II34269));
assign WX3030 = (WX3028)|(WX3027);
assign II2685 = ((~WX817))|((~WX881));
assign WX5407 = (_2222_&WX6176);
assign II34214 = ((~WX11345))|((~WX11001));
assign II11517 = ((~_2144_))|((~II11509));
assign II35012 = ((~II34987))|((~II35011));
assign WX3659 = (WX3657)|(WX3656);
assign II30280 = ((~II30270))|((~II30278));
assign WX5451 = ((~WX6176));
assign II2214 = ((~II2204))|((~II2212));
assign WX3416 = (WX3353&RESET);
assign WX1581 = (WX1587&WX1582);
assign II18658 = ((~II18660))|((~II18661));
assign II34750 = ((~II34740))|((~II34748));
assign WX6728 = (_2252_&WX7469);
assign WX10418 = (WX10416)|(WX10415);
assign WX929 = ((~II2910))|((~II2911));
assign WX4489 = ((~WX4457));
assign WX10790 = (DATA_0_2&WX10791);
assign WX5064 = (WX5062)|(WX5061);
assign II26259 = ((~II26249))|((~II26257));
assign II18100 = ((~II18102))|((~II18103));
assign WX5449 = (_2219_&WX6176);
assign WX11506 = (WX10946&WX11507);
assign WX5280 = (WX5278)|(WX5277);
assign WX9273 = (WX11447&WX9274);
assign WX6424 = ((~II19661))|((~II19662));
assign WX8596 = (WX8533&RESET);
assign II3509 = ((~II3499))|((~II3507));
assign WX3714 = ((~WX3591));
assign WX5285 = (WX5667&WX6176);
assign II23455 = ((~WX7074))|((~II23454));
assign WX2773 = ((~WX2764));
assign WX5524 = (WX6338&WX5525);
assign WX555 = ((~WX979));
assign II10587 = ((~WX3588))|((~WX3269));
assign WX1457 = (WX1455)|(WX1454);
assign II30288 = ((~WX9904))|((~II30286));
assign WX3489 = ((~II10114))|((~II10115));
assign WX2358 = ((~WX2298));
assign DATA_9_0 = ((~WX1228));
assign II11440 = ((~WX3195))|((~II11439));
assign II2801 = ((~WX761))|((~II2793));
assign II2624 = ((~WX813))|((~II2623));
assign WX4831 = ((~WX4805));
assign WX11256 = ((~II34423))|((~II34424));
assign II18830 = ((~WX5997))|((~II18829));
assign WX11342 = ((~TM0));
assign WX6651 = (WX6649)|(WX6648);
assign WX6356 = ((~WX6177));
assign WX10762 = (DATA_0_4&WX10763);
assign WX7488 = ((~WX7470));
assign WX3825 = ((~II11560))|((~II11561));
assign WX7677 = ((~WX7470));
assign WX8391 = ((~WX8637));
assign WX3548 = ((~WX3517));
assign WX2361 = ((~WX2360));
assign II30954 = ((~WX10053))|((~II30953));
assign WX2055 = (WX1992&RESET);
assign II18743 = ((~II18719))|((~II18735));
assign II35702 = ((~WX10978))|((~II35701));
assign II34818 = ((~WX11167))|((~WX11231));
assign WX11012 = (WX10560&RESET);
assign II19099 = ((~WX5754))|((~II19098));
assign WX6816 = (WX6994&WX7469);
assign II34780 = ((~WX11101))|((~II34779));
assign WX1560 = (WX1810&WX2297);
assign WX6698 = ((~WX7468));
assign II22850 = ((~WX7467))|((~WX7164));
assign WX9931 = (WX9868&RESET);
assign II10936 = ((~WX3355))|((~II10935));
assign WX9078 = (WX8996&WX9021);
assign WX7864 = (WX7870&WX7865);
assign WX10766 = (WX11545&WX10767);
assign WX101 = ((~WX1004));
assign II7109 = ((~WX1877))|((~WX1786));
assign II2276 = ((~II2266))|((~II2274));
assign WX7129 = (WX6653&RESET);
assign WX3962 = ((~WX4883));
assign WX7279 = (WX7216&RESET);
assign WX11600 = ((~II35709))|((~II35710));
assign WX11294 = ((~WX11269));
assign II34928 = ((~WX11346))|((~II34927));
assign II30781 = ((~II30783))|((~II30784));
assign WX6662 = (WX6972&WX7469);
assign WX6396 = (WX6395&WX6177);
assign WX5348 = (WX5354&WX5349);
assign WX241 = ((~WX1004));
assign WX2693 = ((~WX3589));
assign WX10168 = ((~WX10167));
assign II10883 = ((~WX3479))|((~II10881));
assign WX1604 = ((~WX2297));
assign II18254 = ((~II18264))|((~II18265));
assign WX456 = (WX462&WX457);
assign WX1539 = (WX1545&WX1540);
assign II11545 = ((~WX3200))|((~_2169_));
assign II22176 = ((~WX7184))|((~II22175));
assign WX5651 = ((~WX6176));
assign WX7424 = ((~WX7423));
assign II1990 = ((~WX645))|((~II1988));
assign WX5338 = (WX7540&WX5339);
assign WX10934 = ((~WX10902));
assign WX800 = (WX737&RESET);
assign WX6335 = ((~WX6177));
assign II30489 = ((~WX10052))|((~II30488));
assign WX10138 = (WX10136)|(WX10135);
assign WX7873 = ((~WX8762));
assign WX5072 = ((~WX5071));
assign WX5013 = (WX4477&WX5014);
assign II26700 = ((~WX8760))|((~WX8447));
assign II30379 = ((~WX9846))|((~WX9910));
assign WX5212 = (WX7477&WX5213);
assign WX10080 = (WX9634&WX10081);
assign WX9691 = ((~WX9944));
assign WX3662 = ((~II11193))|((~II11194));
assign II15720 = ((~_2174_))|((~II15718));
assign WX4838 = ((~WX4837));
assign II6735 = ((~II6745))|((~II6746));
assign II26668 = ((~II26670))|((~II26671));
assign WX8488 = (WX8425&RESET);
assign WX1714 = (WX1832&WX2297);
assign II22314 = ((~II22290))|((~II22306));
assign II3119 = ((~WX495))|((~II3117));
assign WX8904 = ((~II27343))|((~II27344));
assign WX989 = ((~WX988));
assign II34308 = ((~WX11345))|((~II34307));
assign II6543 = ((~II6518))|((~II6542));
assign II18171 = ((~WX5891))|((~II18170));
assign WX3742 = ((~WX3591));
assign II30170 = ((~II30145))|((~II30169));
assign WX3511 = ((~II10796))|((~II10797));
assign II19570 = ((~WX5788))|((~II19569));
assign WX1567 = (WX1573&WX1568);
assign II18651 = ((~II18626))|((~II18650));
assign WX991 = ((~WX990));
assign II30831 = ((~WX9748))|((~II30829));
assign WX11377 = ((~WX11376));
assign II6615 = ((~WX1978))|((~II6613));
assign II18208 = ((~II18210))|((~II18211));
assign II10029 = ((~WX3587))|((~WX3233));
assign WX4872 = ((~WX4871));
assign WX11118 = (WX11055&RESET);
assign WX8250 = (WX8253&RESET);
assign II11427 = ((~WX3194))|((~II11426));
assign WX2565 = (WX2526&WX2556);
assign WX8089 = ((~WX8761));
assign II30759 = ((~II30734))|((~II30758));
assign II23701 = ((~WX7101))|((~II23700));
assign II23667 = ((~_2249_))|((~II23665));
assign WX404 = (WX2487&WX405);
assign II7475 = ((~WX1920))|((~_2140_));
assign II22541 = ((~WX7467))|((~II22540));
assign II2011 = ((~II1986))|((~II2010));
assign WX7621 = ((~WX7470));
assign II27623 = ((~_2289_))|((~II27621));
assign II23645 = ((~WX7091))|((~II23644));
assign WX6095 = ((~II18744))|((~II18745));
assign WX2796 = (WX2794)|(WX2793);
assign II19577 = ((~WX5789))|((~II19576));
assign WX5622 = (WX6387&WX5623);
assign II30411 = ((~WX9848))|((~II30410));
assign II34238 = ((~II34228))|((~II34236));
assign WX4242 = ((~WX4883));
assign WX10193 = ((~WX10056));
assign WX1428 = ((~WX2296));
assign WX6026 = (WX5963&RESET);
assign WX1941 = (WX1369&RESET);
assign II2064 = ((~II2066))|((~II2067));
assign WX10670 = (WX10668)|(WX10667);
assign WX2715 = ((~WX3590));
assign WX2230 = ((~WX2229));
assign WX10644 = ((~WX10643));
assign WX11335 = ((~WX11334));
assign WX6599 = (WX6605&WX6600);
assign WX550 = ((~WX969));
assign WX8582 = (WX8519&RESET);
assign WX4739 = (WX4676&RESET);
assign WX2922 = (WX2920)|(WX2919);
assign WX9897 = (WX9834&RESET);
assign WX1284 = (WX1254&WX1263);
assign WX3450 = (WX3387&RESET);
assign WX10152 = (WX10150)|(WX10149);
assign WX5826 = (WX5290&RESET);
assign II23569 = ((~_2264_))|((~II23567));
assign WX4873 = ((~WX4794));
assign WX2914 = ((~WX2913));
assign II18915 = ((~WX5939))|((~II18914));
assign WX2543 = ((~II7632))|((~II7633));
assign II18533 = ((~II18543))|((~II18544));
assign WX7809 = ((~WX8761));
assign II35563 = ((~_2363_))|((~II35561));
assign WX4172 = ((~WX4883));
assign WX7625 = ((~II23364))|((~II23365));
assign WX8268 = (WX8271&RESET);
assign II30118 = ((~WX9702))|((~II30116));
assign WX591 = ((~WX559));
assign WX9102 = ((~WX10054));
assign WX901 = ((~II2042))|((~II2043));
assign WX7295 = (WX7232&RESET);
assign II7072 = ((~WX1780))|((~II7070));
assign WX918 = ((~II2569))|((~II2570));
assign WX10014 = ((~WX10013));
assign II30490 = ((~WX9726))|((~II30488));
assign WX3991 = (WX3989)|(WX3988);
assign II18186 = ((~II18161))|((~II18185));
assign II35687 = ((~WX10975))|((~_2344_));
assign WX4986 = ((~WX4884));
assign II15314 = ((~WX4478))|((~WX4402));
assign II30643 = ((~WX10053))|((~WX9736));
assign II15288 = ((~WX4476))|((~WX4398));
assign WX6696 = (WX6707&WX7468);
assign WX5604 = (WX7673&WX5605);
assign WX3810 = (WX3809&WX3591);
assign II23583 = ((~_2262_))|((~II23581));
assign WX7061 = ((~WX7029));
assign WX1708 = ((~WX2296));
assign II35005 = ((~WX11179))|((~II35004));
assign WX10213 = (WX9653&WX10214);
assign WX971 = ((~WX970));
assign WX10687 = (WX10698&WX11347);
assign WX11282 = ((~WX11263));
assign WX565 = ((~WX935));
assign II23207 = ((~WX7055))|((~WX6970));
assign II19489 = ((~II19491))|((~II19492));
assign WX5086 = ((~WX5085));
assign WX8756 = ((~TM0));
assign II22461 = ((~II22463))|((~II22464));
assign WX3064 = (WX3815&WX3065);
assign WX954 = ((~WX927));
assign WX3080 = (WX3083&RESET);
assign WX1739 = (WX3801&WX1740);
assign WX7445 = ((~WX7373));
assign II15486 = ((~WX4506))|((~II15485));
assign WX7007 = (WX7010&RESET);
assign WX6561 = (WX8798&WX6562);
assign II30505 = ((~WX9918))|((~II30503));
assign WX11092 = (WX11029&RESET);
assign WX10051 = ((~TM1));
assign WX7723 = ((~II23708))|((~II23709));
assign II2895 = ((~WX767))|((~II2894));
assign WX8614 = (WX8551&RESET);
assign WX536 = (WX539&RESET);
assign WX10888 = (WX10891&RESET);
assign WX9361 = (WX10196&WX9362);
assign WX171 = ((~WX1004));
assign II22431 = ((~WX7264))|((~WX7328));
assign WX10237 = ((~WX10236));
assign WX1383 = ((~WX1382));
assign II14051 = ((~WX4718))|((~II14049));
assign II6009 = ((~WX2066))|((~II6008));
assign WX10558 = (WX10556)|(WX10555);
assign II2808 = ((~II2810))|((~II2811));
assign WX6607 = (WX7526&WX6608);
assign II10951 = ((~II10926))|((~II10950));
assign WX7887 = ((~WX8762));
assign II15711 = ((~WX4519))|((~_2175_));
assign WX522 = (WX525&RESET);
assign WX6136 = ((~WX6072));
assign WX4341 = (WX4339)|(WX4338);
assign II3691 = ((~_2081_))|((~II3689));
assign WX10173 = (WX10171)|(WX10170);
assign II3444 = ((~WX545))|((~II3442));
assign WX1354 = ((~WX1345));
assign II19669 = ((~_2216_))|((~II19667));
assign WX7817 = ((~WX8762));
assign WX9949 = (WX9886&RESET);
assign WX1050 = (WX586&WX1051);
assign WX9695 = (WX9099&RESET);
assign II18581 = ((~WX5981))|((~WX6045));
assign WX10524 = (DATA_0_21&WX10525);
assign WX6757 = (WX8896&WX6758);
assign II34991 = ((~WX11051))|((~II34989));
assign II30435 = ((~II30425))|((~II30433));
assign DATA_9_18 = ((~WX1102));
assign WX2521 = ((~WX2520));
assign II27368 = ((~WX8360))|((~WX8287));
assign WX3440 = (WX3377&RESET);
assign WX5171 = (WX5130&WX5142);
assign WX3848 = ((~II11721))|((~II11722));
assign II23736 = ((~WX7107))|((~II23735));
assign II14284 = ((~WX4542))|((~II14282));
assign WX8963 = ((~WX8763));
assign II18797 = ((~II18799))|((~II18800));
assign WX3178 = ((~WX3146));
assign II6901 = ((~II6891))|((~II6899));
assign II26451 = ((~II26453))|((~II26454));
assign WX3175 = ((~WX3143));
assign WX2187 = (WX2124&RESET);
assign WX2125 = (WX2062&RESET);
assign II19542 = ((~WX5784))|((~II19541));
assign WX3502 = ((~II10517))|((~II10518));
assign II2166 = ((~II2141))|((~II2165));
assign WX2703 = ((~WX2694));
assign II18883 = ((~WX5937))|((~II18875));
assign WX3722 = (WX3720)|(WX3719);
assign II14965 = ((~WX4881))|((~II14964));
assign WX3567 = ((~WX3566));
assign II30340 = ((~WX9780))|((~II30332));
assign WX6838 = ((~WX7468));
assign WX10860 = (WX10863&RESET);
assign II14893 = ((~II14869))|((~II14885));
assign WX2709 = (_2166_&WX3590);
assign WX7022 = ((~WX7448));
assign WX8899 = (WX8357&WX8900);
assign WX9751 = (WX9491&RESET);
assign II22796 = ((~WX7224))|((~II22795));
assign WX8286 = (WX8289&RESET);
assign II34741 = ((~WX11346))|((~WX11035));
assign WX11300 = ((~WX11272));
assign WX10551 = (_2352_&WX11348);
assign II14762 = ((~WX4700))|((~WX4764));
assign II7695 = ((~WX1931))|((~II7694));
assign II6643 = ((~II6645))|((~II6646));
assign II10175 = ((~II10151))|((~II10167));
assign II6219 = ((~II6209))|((~II6217));
assign WX8025 = (WX8275&WX8762);
assign WX3366 = (WX3303&RESET);
assign II27252 = ((~WX8351))|((~II27251));
assign WX838 = (WX775&RESET);
assign WX5473 = (WX5484&WX6175);
assign WX10200 = ((~WX10056));
assign WX10951 = ((~WX10919));
assign II10217 = ((~WX3245))|((~II10215));
assign WX1638 = ((~WX2296));
assign WX5116 = ((~II15551))|((~II15552));
assign WX627 = ((~WX867));
assign WX4993 = ((~WX4884));
assign WX3227 = ((~WX3481));
assign II18273 = ((~WX6025))|((~II18271));
assign II15211 = ((~WX4470))|((~II15210));
assign II2451 = ((~II2461))|((~II2462));
assign WX10100 = (WX10099&WX10056);
assign WX4278 = (WX4289&WX4882);
assign II30565 = ((~WX9858))|((~WX9922));
assign WX10981 = ((~WX11231));
assign WX6720 = ((~WX7469));
assign II19111 = ((~WX5755))|((~WX5663));
assign II30145 = ((~II30155))|((~II30156));
assign WX1663 = ((~WX1662));
assign II27515 = ((~WX8390))|((~_2300_));
assign WX11596 = ((~II35681))|((~II35682));
assign WX10063 = ((~WX10062));
assign WX1478 = ((~WX2297));
assign WX11543 = (WX11541)|(WX11540);
assign WX7880 = (WX7878)|(WX7877);
assign II19730 = ((~WX5814))|((~_2205_));
assign WX1553 = (WX1559&WX1554);
assign WX4297 = (WX6373&WX4298);
assign WX177 = ((~WX1003));
assign II18232 = ((~WX5895))|((~II18224));
assign II27304 = ((~WX8355))|((~II27303));
assign II6922 = ((~II6924))|((~II6925));
assign WX2687 = ((~WX3590));
assign WX4575 = (WX4291&RESET);
assign II11270 = ((~WX3182))|((~WX3103));
assign II2615 = ((~WX749))|((~II2607));
assign WX8692 = ((~WX8675));
assign II30706 = ((~WX10053))|((~II30705));
assign WX4004 = ((~WX4883));
assign II34540 = ((~WX11149))|((~II34539));
assign II14351 = ((~WX4610))|((~II14343));
assign WX2910 = (WX3738&WX2911);
assign WX6739 = (WX6745&WX6740);
assign WX1631 = (WX2452&WX1632);
assign WX631 = ((~WX875));
assign II30474 = ((~WX9916))|((~II30472));
assign WX7598 = (WX7597&WX7470);
assign II11495 = ((~WX3218))|((~_2172_));
assign WX6654 = (WX6665&WX7468);
assign WX9579 = (WX9582&RESET);
assign WX2825 = (WX3099&WX3590);
assign II30805 = ((~WX9810))|((~II30797));
assign II30394 = ((~II30396))|((~II30397));
assign WX10697 = ((~WX11348));
assign II26490 = ((~WX8497))|((~II26482));
assign II27290 = ((~WX8354))|((~WX8275));
assign WX2426 = (WX2425&WX2298);
assign II15067 = ((~WX4459))|((~WX4364));
assign II6682 = ((~WX2046))|((~II6674));
assign WX5316 = (WX5314)|(WX5313);
assign WX4350 = ((~WX4882));
assign II2136 = ((~II2126))|((~II2134));
assign WX2645 = ((~WX3590));
assign II2811 = ((~WX889))|((~II2809));
assign II14506 = ((~WX4620))|((~II14498));
assign WX5179 = (WX5127&WX5142);
assign WX922 = ((~II2693))|((~II2694));
assign II31563 = ((~WX9664))|((~_2330_));
assign WX7713 = ((~II23638))|((~II23639));
assign WX3777 = ((~WX3591));
assign WX6741 = (WX6739)|(WX6738);
assign WX6365 = ((~WX6364));
assign WX1776 = ((~WX1778));
assign II11388 = ((~WX3191))|((~II11387));
assign II10244 = ((~II10254))|((~II10255));
assign WX5816 = (WX5220&RESET);
assign WX1640 = (_2118_&WX2297);
assign WX10101 = (WX9637&WX10102);
assign WX8728 = ((~WX8661));
assign II35577 = ((~_2361_))|((~II35575));
assign WX8380 = ((~WX8615));
assign II14855 = ((~WX4706))|((~WX4770));
assign II6861 = ((~WX2295))|((~WX1994));
assign II27001 = ((~II26977))|((~II26993));
assign WX4919 = ((~WX4918));
assign WX3537 = ((~WX3536));
assign WX9849 = (WX9786&RESET);
assign II3487 = ((~_2108_))|((~II3485));
assign II34980 = ((~II34956))|((~II34972));
assign II34771 = ((~II34773))|((~II34774));
assign II30424 = ((~II30434))|((~II30435));
assign WX3681 = ((~WX3680));
assign WX10840 = (WX10843&RESET);
assign II14057 = ((~II14032))|((~II14056));
assign WX10690 = (WX10688)|(WX10687);
assign WX1835 = (WX1838&RESET);
assign WX10000 = ((~WX9999));
assign WX3530 = ((~WX3508));
assign WX508 = (WX511&RESET);
assign II34510 = ((~WX11211))|((~II34508));
assign WX9650 = ((~WX9618));
assign WX11359 = (WX10925&WX11360);
assign WX4216 = (WX4406&WX4883);
assign II3605 = ((~WX624))|((~_2095_));
assign II23510 = ((~WX7097))|((~_2268_));
assign WX6378 = (WX6376)|(WX6375);
assign WX10019 = ((~WX9953));
assign II34801 = ((~II34811))|((~II34812));
assign WX8056 = (WX8054)|(WX8053);
assign WX4589 = (WX4526&RESET);
assign WX10499 = (WX10845&WX11348);
assign WX1680 = ((~WX2296));
assign WX339 = ((~WX1004));
assign II7577 = ((~_2132_))|((~II7575));
assign WX5589 = (_2209_&WX6176);
assign II31642 = ((~_2319_))|((~II31640));
assign II19512 = ((~_2215_))|((~II19504));
assign II11414 = ((~WX3193))|((~II11413));
assign II31614 = ((~_2323_))|((~II31612));
assign WX8294 = (WX8297&RESET);
assign WX5030 = ((~WX5029));
assign II34453 = ((~II34429))|((~II34445));
assign WX2941 = ((~WX2932));
assign WX3715 = (WX3713)|(WX3712);
assign WX936 = ((~WX918));
assign II2034 = ((~WX775))|((~WX839));
assign II26754 = ((~II26729))|((~II26753));
assign WX6313 = (WX5771&WX6314);
assign WX8342 = ((~WX8310));
assign WX6042 = (WX5979&RESET);
assign WX399 = (WX410&WX1003);
assign WX6814 = ((~WX7469));
assign II3477 = ((~_2092_))|((~II3469));
assign WX1359 = (WX1357)|(WX1356);
assign WX36 = (WX42&WX37);
assign II14359 = ((~WX4674))|((~WX4738));
assign II11524 = ((~WX3229))|((~_2172_));
assign WX8670 = ((~II26413))|((~II26414));
assign WX10471 = (WX10841&WX11348);
assign WX2497 = (WX1901&WX2498);
assign II22508 = ((~II22510))|((~II22511));
assign WX8735 = ((~WX8734));
assign WX570 = ((~WX945));
assign II14854 = ((~II14856))|((~II14857));
assign WX4328 = (WX4422&WX4883);
assign WX10669 = ((~WX11348));
assign WX10537 = (_2353_&WX11348);
assign WX8207 = (WX8301&WX8762);
assign II22804 = ((~WX7288))|((~II22803));
assign WX4074 = ((~WX4883));
assign WX9036 = (WX9015&WX9021);
assign WX4613 = (WX4550&RESET);
assign II31689 = ((~WX9684))|((~_2310_));
assign WX8772 = (WX8771&WX8763);
assign WX5910 = (WX5847&RESET);
assign WX896 = (WX833&RESET);
assign II18759 = ((~WX5929))|((~II18751));
assign WX378 = (WX376)|(WX375);
assign WX8474 = (WX8411&RESET);
assign WX10447 = ((~WX10438));
assign WX4456 = ((~WX4838));
assign II6225 = ((~WX2080))|((~WX2144));
assign II11714 = ((~WX3227))|((~II11713));
assign II3564 = ((~WX618))|((~II3563));
assign II22749 = ((~II22724))|((~II22748));
assign II10470 = ((~WX3325))|((~II10462));
assign II14315 = ((~WX4544))|((~II14313));
assign II10485 = ((~II10461))|((~II10477));
assign II34950 = ((~II34925))|((~II34949));
assign WX4887 = (WX4459&WX4888);
assign WX1042 = (WX1041&WX1005);
assign WX10925 = ((~WX10893));
assign WX10240 = (WX10239&WX10056);
assign WX5264 = (WX5270&WX5265);
assign WX4561 = (WX4193&RESET);
assign WX9129 = (WX9135&WX9130);
assign WX5760 = ((~WX5728));
assign WX4438 = ((~WX4866));
assign WX2909 = (WX3111&WX3590);
assign II14931 = ((~II14941))|((~II14942));
assign II26157 = ((~WX8539))|((~WX8603));
assign II10341 = ((~WX3253))|((~II10339));
assign II10053 = ((~II10043))|((~II10051));
assign II22476 = ((~II22486))|((~II22487));
assign WX9355 = (WX9353)|(WX9352);
assign II31232 = ((~WX9558))|((~II31230));
assign II22192 = ((~II22182))|((~II22190));
assign WX5542 = ((~WX5541));
assign WX1334 = ((~WX2297));
assign II31193 = ((~WX9552))|((~II31191));
assign II10834 = ((~II10836))|((~II10837));
assign WX6510 = ((~WX7469));
assign II2762 = ((~II2764))|((~II2765));
assign II18750 = ((~II18760))|((~II18761));
assign WX621 = ((~WX855));
assign WX9547 = (WX9550&RESET);
assign WX6749 = (WX6747)|(WX6746);
assign WX6434 = ((~II19731))|((~II19732));
assign WX9675 = ((~WX9912));
assign WX5559 = ((~WX6175));
assign WX1861 = ((~WX2234));
assign II34291 = ((~WX11133))|((~WX11197));
assign II34696 = ((~WX11223))|((~II34694));
assign II27109 = ((~WX8340))|((~II27108));
assign WX10549 = ((~WX11347));
assign WX7415 = ((~WX7390));
assign WX5199 = (WX5117&WX5142);
assign II14034 = ((~WX4880))|((~WX4526));
assign WX7896 = (WX10112&WX7897);
assign II14745 = ((~II14755))|((~II14756));
assign WX8223 = ((~WX8762));
assign II18721 = ((~WX6174))|((~WX5863));
assign WX10492 = (WX10498&WX10493);
assign II2493 = ((~II2483))|((~II2491));
assign WX8011 = (WX8273&WX8762);
assign II34346 = ((~WX11073))|((~II34345));
assign II31670 = ((~_2314_))|((~II31668));
assign II18008 = ((~WX6173))|((~WX5817));
assign II35313 = ((~WX10941))|((~WX10863));
assign II27692 = ((~WX8392))|((~II27691));
assign II22216 = ((~WX7314))|((~II22214));
assign II18285 = ((~II18295))|((~II18296));
assign II18766 = ((~II18768))|((~II18769));
assign WX8892 = (WX8356&WX8893);
assign WX1237 = ((~II3536))|((~II3537));
assign WX4899 = ((~II15094))|((~II15095));
assign II2654 = ((~WX815))|((~WX879));
assign WX6868 = (_2242_&WX7469);
assign II2250 = ((~II2252))|((~II2253));
assign WX1734 = (WX1745&WX2296);
assign WX6527 = ((~WX6526));
assign II22680 = ((~WX7280))|((~II22679));
assign II2461 = ((~WX739))|((~II2460));
assign II6156 = ((~WX2012))|((~II6155));
assign WX10464 = (WX10470&WX10465);
assign WX10286 = ((~II31557))|((~II31558));
assign WX3719 = (WX3718&WX3591);
assign II14532 = ((~WX4558))|((~II14530));
assign WX1917 = ((~WX2154));
assign II18783 = ((~WX6174))|((~WX5867));
assign WX10093 = (WX10092&WX10056);
assign WX8387 = ((~WX8629));
assign WX7837 = ((~WX8761));
assign II31256 = ((~WX9644))|((~WX9562));
assign II23532 = ((~_2240_))|((~II23524));
assign WX225 = (WX511&WX1004);
assign WX8376 = ((~WX8607));
assign WX7195 = (WX7132&RESET);
assign WX9498 = ((~WX10055));
assign WX9413 = (WX11517&WX9414);
assign WX7800 = (WX7798)|(WX7797);
assign WX3017 = (_2144_&WX3590);
assign II3485 = ((~WX632))|((~_2108_));
assign WX9126 = ((~WX9117));
assign WX8337 = ((~WX8721));
assign WX6086 = ((~II18465))|((~II18466));
assign II18211 = ((~WX6021))|((~II18209));
assign WX8973 = ((~WX8972));
assign WX4537 = (WX4025&RESET);
assign WX8855 = ((~II27252))|((~II27253));
assign WX4693 = (WX4630&RESET);
assign II10958 = ((~II10960))|((~II10961));
assign WX1531 = (WX1529)|(WX1528);
assign WX10272 = ((~WX10271));
assign II34386 = ((~WX11203))|((~II34384));
assign WX4603 = (WX4540&RESET);
assign II22423 = ((~WX7200))|((~II22415));
assign II30316 = ((~II30318))|((~II30319));
assign II26430 = ((~II26420))|((~II26428));
assign WX3207 = ((~WX3441));
assign WX6977 = (WX6980&RESET);
assign WX6926 = ((~WX7469));
assign II22655 = ((~II22631))|((~II22647));
assign WX2093 = (WX2030&RESET);
assign II6031 = ((~WX2004))|((~II6023));
assign WX5121 = ((~II15586))|((~II15587));
assign WX1177 = ((~WX1005));
assign WX4781 = ((~II14088))|((~II14089));
assign WX8744 = ((~WX8669));
assign II18567 = ((~WX6174))|((~II18566));
assign WX9913 = (WX9850&RESET);
assign WX1620 = ((~WX1611));
assign WX2248 = ((~WX2247));
assign II11337 = ((~WX3113))|((~II11335));
assign WX9227 = (WX9233&WX9228);
assign WX10574 = ((~WX10573));
assign II34686 = ((~WX11095))|((~II34678));
assign II26692 = ((~II26667))|((~II26691));
assign II10206 = ((~II10182))|((~II10198));
assign WX2732 = ((~WX2731));
assign WX1006 = ((~II3053))|((~II3054));
assign WX6243 = (WX5761&WX6244);
assign II19412 = ((~WX5709))|((~II19410));
assign WX7015 = ((~WX7434));
assign WX9146 = (_2328_&WX10055);
assign II10168 = ((~WX3369))|((~WX3433));
assign WX10978 = ((~WX11225));
assign WX6078 = ((~II18217))|((~II18218));
assign II27553 = ((~_2299_))|((~II27551));
assign WX11130 = (WX11067&RESET);
assign WX4894 = (WX4460&WX4895);
assign WX1807 = (WX1810&RESET);
assign WX605 = ((~WX573));
assign WX9514 = (WX9596&WX10055);
assign II19126 = ((~WX5665))|((~II19124));
assign WX10386 = (WX10384)|(WX10383);
assign WX8576 = (WX8513&RESET);
assign WX4854 = ((~WX4853));
assign WX3033 = ((~WX3590));
assign WX597 = ((~WX565));
assign II10184 = ((~WX3587))|((~WX3243));
assign WX7810 = (WX7808)|(WX7807);
assign II14174 = ((~WX4662))|((~II14173));
assign II10446 = ((~II10448))|((~II10449));
assign WX1540 = ((~WX2296));
assign WX8508 = (WX8445&RESET);
assign II26733 = ((~WX8449))|((~II26731));
assign WX10123 = ((~WX10056));
assign WX164 = (WX162)|(WX161);
assign II18481 = ((~WX5911))|((~II18480));
assign WX7801 = (WX8243&WX8762);
assign WX9171 = (WX9177&WX9172);
assign WX2935 = ((~WX3590));
assign II26822 = ((~II26832))|((~II26833));
assign WX10431 = ((~WX11348));
assign II14159 = ((~WX4880))|((~II14158));
assign II34182 = ((~II34184))|((~II34185));
assign II30815 = ((~WX9938))|((~II30813));
assign II19660 = ((~WX5802))|((~_2217_));
assign WX5906 = (WX5843&RESET);
assign WX6252 = (WX6250)|(WX6249);
assign WX1448 = (WX1794&WX2297);
assign WX6780 = (WX6791&WX7468);
assign II10647 = ((~II10657))|((~II10658));
assign WX10662 = (WX10660)|(WX10659);
assign WX6153 = ((~WX6152));
assign II27601 = ((~WX8377))|((~II27600));
assign II3131 = ((~WX586))|((~II3130));
assign II18636 = ((~WX5921))|((~II18635));
assign WX10295 = ((~II31620))|((~II31621));
assign II18192 = ((~II18202))|((~II18203));
assign WX6519 = (WX8777&WX6520);
assign WX11482 = ((~WX11481));
assign WX9581 = (WX9584&RESET);
assign WX6730 = ((~WX7469));
assign II18698 = ((~WX5925))|((~II18697));
assign II18373 = ((~II18363))|((~II18371));
assign WX2722 = (WX2720)|(WX2719);
assign WX11026 = (WX10658&RESET);
assign II30721 = ((~WX9868))|((~II30720));
assign WX7980 = (WX10154&WX7981);
assign WX9962 = ((~II30387))|((~II30388));
assign WX3876 = (WX3838&WX3849);
assign WX8805 = ((~WX8804));
assign II22957 = ((~II22959))|((~II22960));
assign WX7591 = (WX7590&WX7470);
assign WX4106 = ((~WX4883));
assign WX8703 = ((~WX8702));
assign WX83 = ((~WX1004));
assign WX11582 = ((~II35583))|((~II35584));
assign WX1007 = (WX1006&WX1005);
assign WX792 = (WX729&RESET);
assign II27186 = ((~WX8346))|((~WX8259));
assign WX1862 = ((~WX2236));
assign II27316 = ((~WX8356))|((~WX8279));
assign WX5572 = (WX5578&WX5573);
assign II31360 = ((~WX9652))|((~WX9578));
assign WX4317 = (WX4315)|(WX4314);
assign WX11271 = ((~II34888))|((~II34889));
assign II6349 = ((~WX2088))|((~WX2152));
assign WX5932 = (WX5869&RESET);
assign II22278 = ((~WX7318))|((~II22276));
assign WX3797 = (WX3195&WX3798);
assign II26546 = ((~WX8760))|((~II26545));
assign WX413 = (WX424&WX1003);
assign II35094 = ((~WX10829))|((~II35092));
assign II6598 = ((~WX2104))|((~II6597));
assign WX8007 = (_2285_&WX8762);
assign WX998 = ((~TM0));
assign II18502 = ((~II18512))|((~II18513));
assign II2142 = ((~II2144))|((~II2145));
assign WX5020 = (WX4478&WX5021);
assign WX8246 = (WX8249&RESET);
assign II34825 = ((~II34801))|((~II34817));
assign II30891 = ((~WX10053))|((~WX9752));
assign WX2212 = ((~II6605))|((~II6606));
assign II6241 = ((~WX2294))|((~WX1954));
assign WX3998 = (WX4009&WX4882);
assign II2793 = ((~II2795))|((~II2796));
assign WX11531 = ((~WX11530));
assign II10292 = ((~WX3377))|((~WX3441));
assign WX7669 = (WX7073&WX7670);
assign II11622 = ((~WX3211))|((~_2158_));
assign WX4944 = ((~WX4884));
assign II22247 = ((~WX7316))|((~II22245));
assign II10269 = ((~II10244))|((~II10268));
assign WX210 = (WX208)|(WX207);
assign WX11529 = (WX11527)|(WX11526);
assign WX3482 = (WX3419&RESET);
assign II22531 = ((~II22507))|((~II22523));
assign II18348 = ((~II18350))|((~II18351));
assign II2422 = ((~WX1001))|((~WX673));
assign II18953 = ((~WX6005))|((~WX6069));
assign II30898 = ((~WX9816))|((~II30890));
assign II27714 = ((~_2274_))|((~II27712));
assign WX11326 = ((~WX11253));
assign WX11369 = ((~WX11368));
assign WX5982 = (WX5919&RESET);
assign WX9741 = (WX9421&RESET);
assign WX10680 = (WX10678)|(WX10677);
assign WX6625 = ((~WX6624));
assign WX10532 = ((~WX10531));
assign WX5757 = ((~WX5725));
assign WX5560 = (WX5558)|(WX5557);
assign WX1695 = (WX1693)|(WX1692);
assign WX3074 = (WX3077&RESET);
assign II7520 = ((~WX1936))|((~II7519));
assign II10090 = ((~II10092))|((~II10093));
assign II22045 = ((~WX7466))|((~II22044));
assign WX9909 = (WX9846&RESET);
assign II19556 = ((~WX5786))|((~II19555));
assign II6139 = ((~II6115))|((~II6131));
assign WX9412 = (_2309_&WX10055);
assign WX2844 = ((~WX2843));
assign WX9382 = ((~WX10054));
assign WX4523 = (WX3927&RESET);
assign WX5808 = ((~WX6057));
assign WX2729 = ((~WX3590));
assign WX844 = (WX781&RESET);
assign II19074 = ((~WX5657))|((~II19072));
assign WX1597 = (WX1595)|(WX1594);
assign II22113 = ((~WX7180))|((~II22105));
assign WX7931 = ((~WX7922));
assign WX5648 = (WX5646)|(WX5645);
assign WX5355 = (WX5677&WX6176);
assign WX2787 = ((~WX2778));
assign WX8954 = (WX8953&WX8763);
assign WX5104 = (WX4490&WX5105);
assign WX10041 = ((~WX9964));
assign WX4117 = (WX4115)|(WX4114);
assign WX10799 = (WX10810&WX11347);
assign II14747 = ((~WX4881))|((~WX4572));
assign WX10907 = ((~WX11339));
assign WX7942 = (WX8840&WX7943);
assign WX10752 = (WX11538&WX10753);
assign WX6486 = (WX6413&WX6435);
assign II14094 = ((~II14104))|((~II14105));
assign WX10748 = (DATA_0_5&WX10749);
assign WX10446 = (WX10444)|(WX10443);
assign WX9372 = ((~WX10055));
assign WX9131 = (WX9129)|(WX9128);
assign WX2267 = ((~WX2198));
assign II22697 = ((~WX7154))|((~II22695));
assign II3634 = ((~WX629))|((~II3633));
assign WX9871 = (WX9808&RESET);
assign WX10146 = ((~WX10145));
assign WX5832 = (WX5332&RESET);
assign WX9115 = (WX9121&WX9116);
assign II10709 = ((~II10719))|((~II10720));
assign WX7269 = (WX7206&RESET);
assign WX7971 = ((~WX8762));
assign II14228 = ((~WX4602))|((~II14227));
assign WX1923 = ((~WX2166));
assign WX4579 = (WX4319&RESET);
assign WX4479 = ((~WX4447));
assign WX7830 = (WX8784&WX7831);
assign WX6789 = (WX7617&WX6790);
assign WX6197 = ((~WX6196));
assign II30209 = ((~WX10052))|((~WX9708));
assign WX7575 = ((~WX7574));
assign II30985 = ((~WX10053))|((~II30984));
assign WX1549 = (WX1547)|(WX1546);
assign II22866 = ((~WX7292))|((~II22865));
assign II10604 = ((~WX3461))|((~II10602));
assign II26235 = ((~WX8759))|((~WX8417));
assign WX416 = (WX414)|(WX413);
assign WX397 = ((~WX388));
assign WX1118 = ((~II3261))|((~II3262));
assign WX4994 = (WX4992)|(WX4991);
assign WX6791 = (WX6789)|(WX6788);
assign WX5552 = (WX6352&WX5553);
assign WX10239 = ((~II31426))|((~II31427));
assign II35548 = ((~_2336_))|((~II35547));
assign II34136 = ((~WX11123))|((~WX11187));
assign II18908 = ((~WX6174))|((~II18907));
assign II10363 = ((~II10353))|((~II10361));
assign WX4476 = ((~WX4444));
assign WX6798 = (_2247_&WX7469);
assign WX7080 = ((~WX7308));
assign WX3664 = (WX3176&WX3665);
assign WX2867 = (WX3105&WX3590);
assign II10913 = ((~WX3417))|((~II10912));
assign WX4044 = (_2195_&WX4883);
assign WX10515 = ((~WX11348));
assign WX4109 = ((~WX4108));
assign II14522 = ((~II14497))|((~II14521));
assign WX7662 = (WX7072&WX7663);
assign WX9501 = (WX10266&WX9502);
assign II35666 = ((~WX10972))|((~_2347_));
assign II7554 = ((~WX1909))|((~_2135_));
assign II27587 = ((~WX8375))|((~II27586));
assign II34989 = ((~WX11346))|((~WX11051));
assign WX8130 = (WX8136&WX8131);
assign WX4933 = ((~WX4932));
assign WX4033 = (WX4031)|(WX4030);
assign II22538 = ((~II22548))|((~II22549));
assign WX10734 = (DATA_0_6&WX10735);
assign WX6384 = ((~WX6177));
assign WX4543 = (WX4067&RESET);
assign WX5737 = ((~WX6107));
assign WX1910 = ((~WX2140));
assign WX9797 = (WX9734&RESET);
assign WX90 = ((~WX89));
assign II6085 = ((~II6087))|((~II6088));
assign WX2005 = (WX1942&RESET);
assign WX5644 = (WX5642)|(WX5641);
assign II6263 = ((~II6239))|((~II6255));
assign WX1000 = ((~TM1));
assign WX6577 = (WX6575)|(WX6574);
assign WX6326 = (WX6325&WX6177);
assign II26537 = ((~II26512))|((~II26536));
assign II10703 = ((~II10678))|((~II10702));
assign II35432 = ((~WX10881))|((~II35430));
assign II6325 = ((~II6301))|((~II6317));
assign WX328 = ((~WX327));
assign II26350 = ((~II26326))|((~II26342));
assign WX2391 = (WX2390&WX2298);
assign WX7251 = (WX7188&RESET);
assign II31738 = ((~WX9692))|((~_2302_));
assign WX7645 = ((~WX7644));
assign WX1843 = ((~WX2262));
assign WX244 = ((~WX243));
assign WX10620 = (WX10618)|(WX10617);
assign WX1689 = (WX1687)|(WX1686);
assign II30611 = ((~II30613))|((~II30614));
assign WX1395 = (WX1393)|(WX1392);
assign WX1498 = ((~WX2296));
assign WX6886 = (WX7004&WX7469);
assign WX10911 = ((~WX11283));
assign WX672 = (WX244&RESET);
assign WX5978 = (WX5915&RESET);
assign WX9260 = ((~WX10055));
assign II7701 = ((~WX1933))|((~_2111_));
assign WX1411 = ((~WX1410));
assign II6488 = ((~II6490))|((~II6491));
assign WX5582 = (WX5580)|(WX5579);
assign WX10990 = (WX10406&RESET);
assign II22548 = ((~WX7208))|((~II22547));
assign II19449 = ((~WX5781))|((~WX5715));
assign WX8988 = ((~RESET));
assign WX8372 = ((~WX8599));
assign WX11287 = ((~WX11286));
assign WX4223 = (WX4229&WX4224);
assign WX860 = (WX797&RESET);
assign II15629 = ((~_2190_))|((~II15627));
assign II3521 = ((~WX612))|((~_2107_));
assign WX10821 = (WX10891&WX11348);
assign WX5946 = (WX5883&RESET);
assign II10702 = ((~II10678))|((~II10694));
assign WX10486 = (WX11405&WX10487);
assign WX4385 = (WX4388&RESET);
assign WX2511 = (WX1903&WX2512);
assign WX6371 = (WX6369)|(WX6368);
assign WX9653 = ((~WX9621));
assign WX5938 = (WX5875&RESET);
assign WX7704 = ((~II23575))|((~II23576));
assign WX4663 = (WX4600&RESET);
assign II18921 = ((~II18923))|((~II18924));
assign WX4122 = ((~WX4113));
assign II18195 = ((~WX6173))|((~II18194));
assign WX8086 = ((~WX8085));
assign II18325 = ((~WX5901))|((~II18317));
assign WX7293 = (WX7230&RESET);
assign II22686 = ((~II22662))|((~II22678));
assign WX1148 = (WX600&WX1149);
assign II35654 = ((~_2350_))|((~II35652));
assign II15524 = ((~II15514))|((~II15522));
assign WX10608 = (DATA_0_15&WX10609);
assign WX6422 = ((~II19647))|((~II19648));
assign WX6348 = (WX5776&WX6349);
assign WX1697 = (WX3780&WX1698);
assign WX3258 = (WX2830&RESET);
assign II18309 = ((~II18285))|((~II18301));
assign WX4082 = (WX4093&WX4882);
assign WX6355 = (WX5777&WX6356);
assign WX1278 = (WX1257&WX1263);
assign WX5185 = (WX5124&WX5142);
assign WX266 = (WX264)|(WX263);
assign WX9313 = (WX9311)|(WX9310);
assign WX9994 = ((~WX9993));
assign II31519 = ((~II31521))|((~II31522));
assign II26219 = ((~WX8543))|((~WX8607));
assign WX9007 = ((~II27650))|((~II27651));
assign WX4957 = (WX4469&WX4958);
assign WX10148 = ((~II31257))|((~II31258));
assign WX7852 = (WX7850)|(WX7849);
assign II23118 = ((~WX6956))|((~II23116));
assign WX8028 = (WX8026)|(WX8025);
assign WX5797 = ((~WX6035));
assign WX5157 = (WX5136&WX5142);
assign II26218 = ((~II26220))|((~II26221));
assign II2971 = ((~II2947))|((~II2963));
assign WX850 = (WX787&RESET);
assign II7633 = ((~_2123_))|((~II7631));
assign WX3754 = (WX3753&WX3591);
assign WX10257 = (WX10255)|(WX10254);
assign II22616 = ((~II22618))|((~II22619));
assign WX6508 = (WX6950&WX7469);
assign WX2447 = (WX2446&WX2298);
assign II3556 = ((~WX617))|((~_2102_));
assign II30533 = ((~II30535))|((~II30536));
assign II34175 = ((~II34150))|((~II34174));
assign WX8852 = (WX8850)|(WX8849);
assign WX10264 = (WX10262)|(WX10261);
assign II14769 = ((~II14745))|((~II14761));
assign WX5425 = (WX5687&WX6176);
assign II10666 = ((~WX3465))|((~II10664));
assign II26174 = ((~WX8759))|((~II26173));
assign WX10815 = ((~WX11347));
assign WX10065 = (WX10064&WX10056);
assign WX234 = (WX232)|(WX231);
assign WX3691 = (WX3690&WX3591);
assign II23378 = ((~WX6996))|((~II23376));
assign WX6101 = ((~II18930))|((~II18931));
assign II2413 = ((~II2389))|((~II2405));
assign WX11408 = (WX10932&WX11409);
assign WX8414 = (WX7890&RESET);
assign WX5794 = ((~WX6029));
assign WX8163 = ((~WX8762));
assign WX5588 = (WX5586)|(WX5585);
assign II35681 = ((~WX10974))|((~II35680));
assign WX9026 = (WX9019&WX9021);
assign WX10116 = ((~WX10056));
assign WX3940 = ((~WX3931));
assign WX8494 = (WX8431&RESET);
assign WX5262 = ((~WX5261));
assign WX2364 = (WX1882&WX2365);
assign II35132 = ((~WX10927))|((~II35131));
assign WX10136 = (WX9642&WX10137);
assign WX10585 = ((~WX11348));
assign WX5302 = (WX5300)|(WX5299);
assign WX4451 = ((~WX4828));
assign II14807 = ((~II14817))|((~II14818));
assign WX3996 = ((~WX3987));
assign II31166 = ((~WX9637))|((~II31165));
assign II10695 = ((~WX3403))|((~WX3467));
assign II22190 = ((~II22166))|((~II22182));
assign WX6446 = (WX6431&WX6435);
assign WX11605 = ((~II35744))|((~II35745));
assign II10919 = ((~II10895))|((~II10911));
assign II34275 = ((~II34277))|((~II34278));
assign WX2294 = ((~WX2293));
assign II27615 = ((~WX8379))|((~II27614));
assign II6940 = ((~WX2190))|((~II6938));
assign WX4946 = ((~WX4945));
assign WX418 = (WX2494&WX419);
assign II27712 = ((~WX8395))|((~_2274_));
assign II14816 = ((~WX4640))|((~II14808));
assign II6566 = ((~WX2102))|((~WX2166));
assign WX5412 = (WX6282&WX5413);
assign WX435 = (WX541&WX1004);
assign WX5662 = (WX5665&RESET);
assign II30357 = ((~II30347))|((~II30355));
assign II3704 = ((~WX641))|((~II3703));
assign WX5765 = ((~WX5733));
assign II26204 = ((~WX8759))|((~WX8415));
assign II27343 = ((~WX8358))|((~II27342));
assign WX1204 = (WX608&WX1205);
assign WX74 = (WX72)|(WX71);
assign WX8146 = (WX8144)|(WX8143);
assign II27121 = ((~WX8341))|((~WX8249));
assign WX6260 = ((~WX6259));
assign WX5755 = ((~WX5723));
assign II23517 = ((~_2247_))|((~II23509));
assign II10673 = ((~II10663))|((~II10671));
assign II34739 = ((~II34749))|((~II34750));
assign WX1935 = ((~WX2190));
assign WX6130 = ((~WX6101));
assign II15340 = ((~WX4480))|((~WX4406));
assign II18993 = ((~II18983))|((~II18991));
assign WX2552 = ((~II7695))|((~II7696));
assign II3514 = ((~WX643))|((~_2108_));
assign II22013 = ((~WX7466))|((~WX7110));
assign II2865 = ((~II2855))|((~II2863));
assign WX9214 = ((~WX10054));
assign II14236 = ((~WX4666))|((~II14235));
assign WX5480 = (WX5478)|(WX5477);
assign WX4783 = ((~II14150))|((~II14151));
assign WX4826 = ((~WX4825));
assign WX1496 = (WX1507&WX2296);
assign II22129 = ((~II22104))|((~II22128));
assign WX2208 = ((~II6481))|((~II6482));
assign WX4807 = ((~II14894))|((~II14895));
assign WX10945 = ((~WX10913));
assign WX3598 = ((~WX3597));
assign WX10317 = (WX10313&WX10314);
assign WX7921 = ((~WX8761));
assign II10294 = ((~WX3441))|((~II10292));
assign II26391 = ((~WX8759))|((~II26390));
assign WX1254 = ((~II3655))|((~II3656));
assign WX5044 = ((~WX5043));
assign WX1961 = (WX1509&RESET);
assign II18929 = ((~II18905))|((~II18921));
assign II18619 = ((~II18595))|((~II18611));
assign WX186 = (WX184)|(WX183);
assign WX5924 = (WX5861&RESET);
assign WX6844 = (WX6998&WX7469);
assign WX1346 = (_2139_&WX2297);
assign WX10313 = ((~II31746))|((~II31747));
assign II7682 = ((~_2115_))|((~II7680));
assign WX11658 = (WX11585&WX11607);
assign WX8220 = (WX8218)|(WX8217);
assign WX6456 = (WX6426&WX6435);
assign WX7522 = (WX7052&WX7523);
assign WX2141 = (WX2078&RESET);
assign WX10478 = (WX10484&WX10479);
assign WX6622 = ((~WX7469));
assign WX4647 = (WX4584&RESET);
assign WX9353 = (WX9359&WX9354);
assign WX9979 = ((~II30914))|((~II30915));
assign II11496 = ((~WX3218))|((~II11495));
assign II19217 = ((~WX5679))|((~II19215));
assign WX3900 = (WX3827&WX3849);
assign WX5554 = (WX5552)|(WX5551);
assign WX6876 = ((~WX6867));
assign II31115 = ((~WX9540))|((~II31113));
assign II26421 = ((~WX8759))|((~WX8429));
assign II22022 = ((~II22012))|((~II22020));
assign II14129 = ((~WX4532))|((~II14127));
assign WX1388 = (_2136_&WX2297);
assign WX11242 = (WX11179&RESET);
assign WX9298 = ((~WX10054));
assign II31550 = ((~WX9694))|((~II31549));
assign II18046 = ((~WX5883))|((~II18038));
assign II10115 = ((~II10105))|((~II10113));
assign WX3157 = ((~WX3533));
assign WX3787 = ((~WX3786));
assign WX1931 = ((~WX2182));
assign WX7231 = (WX7168&RESET);
assign II11713 = ((~WX3227))|((~_2142_));
assign II6730 = ((~II6720))|((~II6728));
assign WX6294 = (WX6292)|(WX6291);
assign WX2452 = ((~WX2451));
assign II22965 = ((~II22941))|((~II22957));
assign WX4811 = ((~WX4795));
assign WX5173 = (WX5129&WX5142);
assign II10430 = ((~II10440))|((~II10441));
assign WX3613 = ((~II11102))|((~II11103));
assign II26330 = ((~WX8423))|((~II26328));
assign WX6213 = ((~II19138))|((~II19139));
assign WX10830 = (WX10833&RESET);
assign WX7040 = ((~WX7420));
assign II27395 = ((~WX8362))|((~II27394));
assign WX1629 = (WX1627)|(WX1626);
assign WX7451 = ((~WX7376));
assign WX5750 = ((~WX6133));
assign WX5002 = ((~WX5001));
assign II23688 = ((~_2245_))|((~II23686));
assign WX9249 = (WX10140&WX9250);
assign WX996 = ((~TM0));
assign II23168 = ((~WX7052))|((~WX6964));
assign WX2370 = (WX2369&WX2298);
assign II10772 = ((~II10774))|((~II10775));
assign II22145 = ((~WX7182))|((~II22144));
assign II31506 = ((~WX9678))|((~II31505));
assign WX5227 = ((~WX6176));
assign WX1506 = ((~WX2297));
assign II34918 = ((~II34894))|((~II34910));
assign WX9334 = ((~WX10055));
assign WX3184 = ((~WX3152));
assign II31719 = ((~_2306_))|((~II31717));
assign WX2810 = (WX2808)|(WX2807);
assign WX9460 = ((~WX10055));
assign II10223 = ((~WX3309))|((~II10222));
assign WX10968 = ((~WX11205));
assign II26698 = ((~II26708))|((~II26709));
assign II14940 = ((~WX4648))|((~II14932));
assign WX226 = (DATA_9_18&WX227);
assign WX10828 = (WX10831&RESET);
assign II6178 = ((~II6180))|((~II6181));
assign WX643 = ((~WX899));
assign WX7187 = (WX7124&RESET);
assign WX4499 = ((~WX4732));
assign WX3864 = (WX3843&WX3849);
assign WX6442 = (WX6432&WX6435);
assign II6706 = ((~WX2295))|((~WX1984));
assign II3430 = ((~WX609))|((~II3429));
assign WX287 = (WX298&WX1003);
assign WX9336 = ((~WX9327));
assign II22874 = ((~II22864))|((~II22872));
assign WX2896 = (WX3731&WX2897);
assign II10154 = ((~WX3587))|((~II10153));
assign II31466 = ((~WX9594))|((~II31464));
assign II30736 = ((~WX10053))|((~WX9742));
assign II15367 = ((~WX4482))|((~II15366));
assign II34594 = ((~WX11089))|((~II34593));
assign II22821 = ((~WX7162))|((~II22819));
assign WX10731 = ((~WX11347));
assign WX3214 = ((~WX3455));
assign WX1893 = ((~WX1861));
assign WX2422 = (WX2420)|(WX2419);
assign WX579 = ((~WX963));
assign II30350 = ((~WX9908))|((~II30348));
assign WX5136 = ((~II15691))|((~II15692));
assign II18010 = ((~WX5817))|((~II18008));
assign WX4055 = (WX4061&WX4056);
assign WX7439 = ((~WX7370));
assign II34911 = ((~WX11173))|((~WX11237));
assign II14328 = ((~WX4672))|((~WX4736));
assign WX7433 = ((~WX7367));
assign WX8996 = ((~II27573))|((~II27574));
assign II7200 = ((~WX1884))|((~WX1800));
assign WX4336 = ((~WX4882));
assign WX7253 = (WX7190&RESET);
assign WX5163 = (WX5133&WX5142);
assign WX4417 = (WX4420&RESET);
assign II6528 = ((~WX2036))|((~II6527));
assign WX3532 = ((~WX3509));
assign II26195 = ((~II26171))|((~II26187));
assign II10633 = ((~WX3399))|((~WX3463));
assign WX8193 = (WX8299&WX8762);
assign II7703 = ((~_2111_))|((~II7701));
assign WX7559 = (WX7557)|(WX7556);
assign WX3751 = ((~WX3750));
assign II10207 = ((~II10182))|((~II10206));
assign WX11086 = (WX11023&RESET);
assign II22036 = ((~II22011))|((~II22035));
assign WX4505 = ((~WX4744));
assign WX2378 = (WX1884&WX2379);
assign II11574 = ((~WX3204))|((~II11573));
assign WX9262 = (WX9560&WX10055);
assign WX2546 = ((~II7653))|((~II7654));
assign WX9470 = ((~WX10055));
assign II22600 = ((~II22610))|((~II22611));
assign II6589 = ((~WX2040))|((~II6581));
assign II18814 = ((~WX6174))|((~WX5869));
assign II18752 = ((~WX6174))|((~WX5865));
assign II18258 = ((~WX5833))|((~II18256));
assign WX6376 = (WX5780&WX6377);
assign II14631 = ((~WX4628))|((~II14630));
assign WX2435 = ((~WX2298));
assign II18513 = ((~II18503))|((~II18511));
assign II2205 = ((~WX1001))|((~WX659));
assign II35392 = ((~WX10947))|((~II35391));
assign WX1756 = (WX1838&WX2297);
assign WX2514 = ((~WX2513));
assign II31178 = ((~WX9638))|((~WX9550));
assign WX11459 = (WX11457)|(WX11456);
assign WX5149 = (WX5139&WX5142);
assign WX7584 = (WX7583&WX7470);
assign WX10567 = ((~WX11348));
assign WX6677 = (WX7561&WX6678);
assign WX10808 = (WX11566&WX10809);
assign WX7794 = (WX7800&WX7795);
assign II34221 = ((~WX11065))|((~II34213));
assign II18172 = ((~II18162))|((~II18170));
assign WX4508 = ((~WX4750));
assign II7332 = ((~WX1820))|((~II7330));
assign WX5729 = ((~WX6155));
assign II14583 = ((~II14559))|((~II14575));
assign II30187 = ((~II30177))|((~II30185));
assign WX7618 = ((~II23351))|((~II23352));
assign WX1021 = (WX1020&WX1005);
assign WX206 = (WX204)|(WX203);
assign II3535 = ((~WX614))|((~_2105_));
assign WX7299 = (WX7236&RESET);
assign II10563 = ((~WX3331))|((~II10555));
assign II2043 = ((~II2033))|((~II2041));
assign WX51 = ((~WX1003));
assign II22316 = ((~II22306))|((~II22314));
assign WX4775 = (WX4712&RESET);
assign WX1727 = (WX1725)|(WX1724);
assign II26352 = ((~II26342))|((~II26350));
assign II10076 = ((~WX3363))|((~II10075));
assign WX2765 = (_2162_&WX3590);
assign II26412 = ((~II26388))|((~II26404));
assign WX11426 = ((~WX11425));
assign II2886 = ((~II2888))|((~II2889));
assign WX2957 = (WX2968&WX3589);
assign WX9229 = (WX9227)|(WX9226);
assign II18444 = ((~WX5845))|((~II18442));
assign WX11642 = (WX11593&WX11607);
assign WX6490 = (WX6411&WX6435);
assign WX1431 = (WX3647&WX1432);
assign WX386 = (WX392&WX387);
assign WX9473 = (WX10252&WX9474);
assign II26702 = ((~WX8447))|((~II26700));
assign WX8813 = ((~II27174))|((~II27175));
assign WX3977 = (WX3975)|(WX3974);
assign WX4519 = ((~WX4772));
assign WX1720 = (WX1731&WX2296);
assign WX8448 = (WX8128&RESET);
assign WX5505 = (_2215_&WX6176);
assign WX2286 = ((~WX2285));
assign II34082 = ((~II34057))|((~II34081));
assign WX7039 = ((~WX7418));
assign WX7032 = ((~WX7404));
assign II26574 = ((~II26584))|((~II26585));
assign II14962 = ((~II14972))|((~II14973));
assign II6651 = ((~WX2044))|((~II6643));
assign WX10778 = (WX10776)|(WX10775);
assign II19514 = ((~II19504))|((~II19512));
assign II19333 = ((~WX5772))|((~II19332));
assign WX1573 = (WX1571)|(WX1570);
assign WX3236 = (WX2676&RESET);
assign II18099 = ((~II18109))|((~II18110));
assign II2343 = ((~II2345))|((~II2346));
assign WX10197 = ((~II31348))|((~II31349));
assign II2104 = ((~II2079))|((~II2103));
assign WX6339 = ((~II19372))|((~II19373));
assign WX6234 = ((~II19177))|((~II19178));
assign II2328 = ((~II2330))|((~II2331));
assign WX8774 = ((~WX8763));
assign WX9627 = ((~WX10008));
assign II2631 = ((~II2606))|((~II2630));
assign II22307 = ((~WX7256))|((~WX7320));
assign II2873 = ((~WX893))|((~II2871));
assign WX315 = (WX326&WX1003);
assign II7460 = ((~WX1904))|((~WX1840));
assign WX4516 = ((~WX4766));
assign WX10658 = ((~WX10657));
assign WX2847 = ((~WX3589));
assign WX4866 = ((~WX4865));
assign WX3388 = (WX3325&RESET);
assign II19282 = ((~WX5689))|((~II19280));
assign II30580 = ((~II30582))|((~II30583));
assign WX10651 = ((~WX11348));
assign II7542 = ((~_2137_))|((~II7540));
assign WX11146 = (WX11083&RESET);
assign II11323 = ((~WX3186))|((~II11322));
assign WX10219 = (WX10218&WX10056);
assign WX4729 = (WX4666&RESET);
assign II26144 = ((~WX8411))|((~II26142));
assign WX10323 = (WX10284&WX10314);
assign II34293 = ((~WX11197))|((~II34291));
assign II11244 = ((~WX3180))|((~WX3099));
assign II14949 = ((~WX4712))|((~II14948));
assign WX8697 = ((~WX8696));
assign II35223 = ((~WX10934))|((~II35222));
assign WX9464 = (WX9475&WX10054);
assign WX5492 = (WX7617&WX5493);
assign WX11636 = (WX11595&WX11607);
assign II34057 = ((~II34067))|((~II34068));
assign II10658 = ((~II10648))|((~II10656));
assign WX3670 = (WX3669&WX3591);
assign WX10923 = ((~WX11307));
assign WX1485 = (WX1483)|(WX1482);
assign II23313 = ((~WX6986))|((~II23311));
assign II30658 = ((~WX9864))|((~WX9928));
assign WX8956 = ((~WX8763));
assign WX9208 = ((~WX10055));
assign II2213 = ((~WX723))|((~II2212));
assign WX1071 = (WX589&WX1072);
assign II34267 = ((~II34243))|((~II34259));
assign II14439 = ((~WX4552))|((~II14437));
assign WX945 = ((~WX944));
assign II34463 = ((~WX11345))|((~II34462));
assign II26629 = ((~II26605))|((~II26621));
assign II15419 = ((~WX4486))|((~II15418));
assign II26081 = ((~WX8759))|((~II26080));
assign II18425 = ((~II18427))|((~II18428));
assign II6894 = ((~WX1996))|((~II6892));
assign WX8715 = ((~WX8714));
assign II2368 = ((~WX733))|((~II2367));
assign WX7391 = ((~II22842))|((~II22843));
assign WX4761 = (WX4698&RESET);
assign WX8272 = (WX8275&RESET);
assign II6234 = ((~II6224))|((~II6232));
assign WX1214 = ((~WX1213));
assign II18939 = ((~WX6174))|((~II18938));
assign II10973 = ((~II10975))|((~II10976));
assign II7717 = ((~_2109_))|((~II7715));
assign II22810 = ((~II22786))|((~II22802));
assign II18877 = ((~WX6174))|((~II18876));
assign WX64 = (WX70&WX65);
assign WX1227 = (WX1225)|(WX1224);
assign II26313 = ((~WX8549))|((~II26312));
assign WX9184 = (WX9195&WX10054);
assign II18713 = ((~II18688))|((~II18712));
assign II10308 = ((~WX3587))|((~WX3251));
assign II2266 = ((~II2268))|((~II2269));
assign WX8422 = (WX7946&RESET);
assign II26289 = ((~II26264))|((~II26288));
assign WX4204 = ((~WX4883));
assign WX5331 = ((~WX5322));
assign II18006 = ((~II18016))|((~II18017));
assign WX9181 = (WX9179)|(WX9178);
assign II15251 = ((~WX4392))|((~II15249));
assign WX2466 = ((~WX2465));
assign II15275 = ((~WX4475))|((~WX4396));
assign II6366 = ((~WX2294))|((~II6365));
assign II6064 = ((~II6054))|((~II6062));
assign WX11351 = (WX11350&WX11349);
assign WX11308 = ((~WX11244));
assign II31682 = ((~WX9682))|((~_2312_));
assign II30542 = ((~II30517))|((~II30541));
assign WX11006 = (WX10518&RESET);
assign DATA_9_28 = ((~WX1032));
assign WX6672 = (_2256_&WX7469);
assign II6971 = ((~WX2192))|((~II6969));
assign WX8915 = (WX8913)|(WX8912);
assign WX3648 = ((~II11167))|((~II11168));
assign WX8832 = ((~WX8831));
assign II26531 = ((~WX8627))|((~II26529));
assign II27265 = ((~WX8352))|((~II27264));
assign II14392 = ((~WX4740))|((~II14390));
assign II3470 = ((~WX627))|((~_2108_));
assign II14087 = ((~II14063))|((~II14079));
assign WX6183 = ((~WX6182));
assign WX1053 = ((~WX1052));
assign II3365 = ((~WX604))|((~II3364));
assign II14144 = ((~WX4724))|((~II14142));
assign II2090 = ((~II2080))|((~II2088));
assign WX2246 = ((~WX2245));
assign II26265 = ((~II26267))|((~II26268));
assign II18388 = ((~WX5905))|((~II18387));
assign WX138 = (WX2354&WX139);
assign WX11512 = (WX11511&WX11349);
assign WX6848 = ((~WX6839));
assign II26205 = ((~WX8759))|((~II26204));
assign II18457 = ((~WX5973))|((~WX6037));
assign WX420 = (WX418)|(WX417);
assign WX4870 = ((~WX4869));
assign II31585 = ((~WX9667))|((~II31584));
assign II35715 = ((~WX10980))|((~_2339_));
assign II34631 = ((~II34633))|((~II34634));
assign WX8139 = ((~WX8762));
assign WX10425 = (_2361_&WX11348);
assign II19690 = ((~_2212_))|((~II19688));
assign WX7839 = (_2297_&WX8762);
assign WX518 = (WX521&RESET);
assign WX9405 = (WX9403)|(WX9402);
assign WX9524 = (_2301_&WX10055);
assign WX4152 = (WX4163&WX4882);
assign II6124 = ((~WX2010))|((~II6116));
assign WX1905 = ((~WX2130));
assign II27551 = ((~WX8370))|((~_2299_));
assign WX2899 = ((~WX2890));
assign II26622 = ((~WX8569))|((~WX8633));
assign WX7018 = ((~WX7440));
assign WX1712 = ((~WX2297));
assign WX11614 = (WX11604&WX11607);
assign WX1216 = ((~II3443))|((~II3444));
assign WX10899 = ((~WX11323));
assign WX4683 = (WX4620&RESET);
assign WX2650 = (WX2656&WX2651);
assign II26848 = ((~II26838))|((~II26846));
assign WX7867 = (_2295_&WX8762);
assign WX2782 = (WX2780)|(WX2779);
assign WX7603 = ((~WX7602));
assign II6118 = ((~WX2294))|((~II6117));
assign WX3280 = (WX2984&RESET);
assign WX6887 = (WX7666&WX6888);
assign II14149 = ((~II14125))|((~II14141));
assign II10725 = ((~II10727))|((~II10728));
assign II2949 = ((~WX1002))|((~WX707));
assign WX6686 = (_2255_&WX7469);
assign WX2745 = ((~WX2736));
assign WX8604 = (WX8541&RESET);
assign II34724 = ((~II34726))|((~II34727));
assign II34616 = ((~II34618))|((~II34619));
assign WX9191 = (WX9189)|(WX9188);
assign WX10453 = (_2359_&WX11348);
assign WX10297 = ((~II31634))|((~II31635));
assign II14538 = ((~WX4622))|((~II14537));
assign II2647 = ((~WX751))|((~II2646));
assign WX9100 = (WX9111&WX10054);
assign WX8034 = (WX8032)|(WX8031);
assign WX2273 = ((~WX2201));
assign WX9370 = (_2312_&WX10055);
assign II22819 = ((~WX7467))|((~WX7162));
assign II15509 = ((~II15499))|((~II15507));
assign WX148 = (WX154&WX149);
assign II35554 = ((~WX10987))|((~_2364_));
assign II26980 = ((~WX8760))|((~II26979));
assign II10439 = ((~WX3323))|((~II10431));
assign II2909 = ((~II2885))|((~II2901));
assign II34284 = ((~WX11069))|((~II34283));
assign II30628 = ((~WX9862))|((~II30627));
assign II18087 = ((~WX6013))|((~II18085));
assign WX5605 = ((~WX6176));
assign WX2678 = (WX2684&WX2679);
assign II30598 = ((~WX9924))|((~II30596));
assign WX6408 = ((~II19549))|((~II19550));
assign WX8789 = (WX8787)|(WX8786);
assign II19491 = ((~WX5799))|((~II19490));
assign WX1483 = (WX1489&WX1484);
assign WX9165 = (WX10098&WX9166);
assign WX4129 = (WX6289&WX4130);
assign WX6224 = (WX6222)|(WX6221);
assign WX4545 = (WX4081&RESET);
assign WX133 = (WX144&WX1003);
assign WX6547 = (WX8791&WX6548);
assign WX1069 = ((~II3170))|((~II3171));
assign WX1111 = ((~II3248))|((~II3249));
assign II22941 = ((~II22951))|((~II22952));
assign WX7090 = ((~WX7328));
assign II34926 = ((~II34928))|((~II34929));
assign II10021 = ((~II9996))|((~II10020));
assign WX8204 = (WX10266&WX8205);
assign WX11156 = (WX11093&RESET);
assign WX7846 = (WX7844)|(WX7843);
assign WX8618 = (WX8555&RESET);
assign WX4361 = ((~WX4360));
assign WX3801 = ((~WX3800));
assign II34197 = ((~II34199))|((~II34200));
assign WX9290 = (WX9564&WX10055);
assign WX10642 = (WX10640)|(WX10639);
assign WX10956 = ((~WX11181));
assign II10301 = ((~II10291))|((~II10299));
assign WX5599 = (WX5610&WX6175);
assign WX2930 = (WX2936&WX2931);
assign WX305 = (_2089_&WX1004);
assign WX602 = ((~WX570));
assign WX6097 = ((~II18806))|((~II18807));
assign II31334 = ((~WX9650))|((~WX9574));
assign II22935 = ((~II22910))|((~II22934));
assign WX6700 = (_2254_&WX7469);
assign WX3554 = ((~WX3488));
assign II35315 = ((~WX10863))|((~II35313));
assign II6025 = ((~WX2294))|((~II6024));
assign II15381 = ((~WX4412))|((~II15379));
assign II11453 = ((~WX3196))|((~II11452));
assign WX668 = (WX216&RESET);
assign WX534 = (WX537&RESET);
assign II34872 = ((~WX11107))|((~II34864));
assign WX2482 = (WX2481&WX2298);
assign WX8153 = ((~WX8762));
assign WX7430 = ((~WX7429));
assign II18403 = ((~II18378))|((~II18402));
assign II3416 = ((~WX608))|((~WX541));
assign WX11277 = ((~WX11276));
assign WX7479 = (WX7478&WX7470);
assign II11596 = ((~_2162_))|((~II11594));
assign II6628 = ((~WX2106))|((~WX2170));
assign WX9237 = (WX9235)|(WX9234);
assign II2787 = ((~II2777))|((~II2785));
assign WX11328 = ((~WX11254));
assign WX5591 = ((~WX6176));
assign II10678 = ((~II10688))|((~II10689));
assign WX10467 = (_2358_&WX11348);
assign WX8838 = (WX8836)|(WX8835);
assign II22711 = ((~WX7282))|((~II22710));
assign II19498 = ((~_2220_))|((~II19497));
assign WX1445 = (WX3654&WX1446);
assign WX2663 = (WX2674&WX3589);
assign WX2925 = ((~WX3590));
assign WX774 = (WX711&RESET);
assign WX5510 = (WX6331&WX5511);
assign II34399 = ((~II34401))|((~II34402));
assign II26994 = ((~WX8593))|((~WX8657));
assign II18409 = ((~II18419))|((~II18420));
assign II7660 = ((~WX1926))|((~II7659));
assign WX9823 = (WX9760&RESET);
assign WX11068 = (WX11005&RESET);
assign II18402 = ((~II18378))|((~II18394));
assign II6281 = ((~II6271))|((~II6279));
assign WX7025 = ((~WX7454));
assign II22059 = ((~WX7240))|((~WX7304));
assign WX7481 = ((~WX7470));
assign WX6246 = ((~WX6245));
assign WX11389 = (WX11387)|(WX11386);
assign WX4843 = ((~WX4779));
assign II35276 = ((~WX10857))|((~II35274));
assign II14785 = ((~WX4638))|((~II14777));
assign II7484 = ((~II7474))|((~II7482));
assign WX10285 = ((~II31550))|((~II31551));
assign WX2495 = ((~II7422))|((~II7423));
assign WX451 = ((~WX1004));
assign II26615 = ((~WX8505))|((~II26614));
assign WX10404 = (WX10402)|(WX10401);
assign WX3524 = ((~WX3505));
assign WX1514 = (_2127_&WX2297);
assign WX9561 = (WX9564&RESET);
assign II26553 = ((~WX8501))|((~II26552));
assign WX2469 = (WX1897&WX2470);
assign WX429 = ((~WX1003));
assign II27558 = ((~WX8371))|((~_2298_));
assign WX4393 = (WX4396&RESET);
assign WX2326 = ((~WX2325));
assign WX5193 = (WX5120&WX5142);
assign WX5900 = (WX5837&RESET);
assign II10015 = ((~WX3423))|((~II10013));
assign II14304 = ((~II14280))|((~II14296));
assign II7647 = ((~_2121_))|((~II7645));
assign WX7775 = (WX7708&WX7728);
assign WX11090 = (WX11027&RESET);
assign WX6955 = (WX6958&RESET);
assign WX6540 = ((~WX6531));
assign WX445 = (_2079_&WX1004);
assign II6467 = ((~II6457))|((~II6465));
assign II31386 = ((~WX9654))|((~WX9582));
assign II22602 = ((~WX7467))|((~WX7148));
assign WX10706 = (DATA_0_8&WX10707);
assign WX6310 = ((~WX6309));
assign WX9425 = (WX9423)|(WX9422);
assign WX2657 = (WX3075&WX3590);
assign II23442 = ((~WX7073))|((~II23441));
assign II14647 = ((~II14637))|((~II14645));
assign II11349 = ((~WX3188))|((~II11348));
assign WX8119 = (_2277_&WX8762);
assign WX6896 = (_2240_&WX7469);
assign WX1894 = ((~WX1862));
assign II3663 = ((~_2085_))|((~II3661));
assign II34811 = ((~WX11103))|((~II34810));
assign II30301 = ((~II30303))|((~II30304));
assign WX3096 = (WX3099&RESET);
assign WX2978 = (WX2976)|(WX2975);
assign WX10594 = (DATA_0_16&WX10595);
assign WX10788 = (WX10786)|(WX10785);
assign II10120 = ((~II10130))|((~II10131));
assign WX8106 = (WX10217&WX8107);
assign II22322 = ((~II22324))|((~II22325));
assign WX2971 = (WX2982&WX3589);
assign WX8944 = ((~WX8943));
assign II19085 = ((~WX5753))|((~WX5659));
assign WX146 = ((~WX145));
assign II34400 = ((~WX11345))|((~WX11013));
assign WX2413 = (WX1889&WX2414);
assign WX6145 = ((~WX6144));
assign WX656 = (WX132&RESET);
assign II7163 = ((~WX1794))|((~II7161));
assign WX10616 = ((~WX10615));
assign WX583 = ((~WX551));
assign WX5475 = ((~WX6175));
assign WX2224 = ((~II6977))|((~II6978));
assign WX458 = (WX456)|(WX455);
assign WX10502 = (WX10500)|(WX10499);
assign WX9432 = ((~WX10055));
assign WX8466 = (WX8403&RESET);
assign WX6904 = ((~WX6895));
assign II31477 = ((~WX9661))|((~WX9596));
assign II31740 = ((~_2302_))|((~II31738));
assign II30908 = ((~WX9944))|((~II30906));
assign WX2428 = ((~WX2298));
assign II35419 = ((~WX10879))|((~II35417));
assign WX712 = (WX649&RESET);
assign II26288 = ((~II26264))|((~II26280));
assign WX9670 = ((~WX9902));
assign II18047 = ((~WX5883))|((~II18046));
assign WX5069 = (WX4485&WX5070);
assign WX880 = (WX817&RESET);
assign II34959 = ((~WX11346))|((~II34958));
assign WX5325 = ((~WX6176));
assign II26779 = ((~WX8643))|((~II26777));
assign WX8177 = ((~WX8762));
assign WX3009 = ((~WX3590));
assign II22625 = ((~II22600))|((~II22624));
assign WX3908 = (WX3823&WX3849);
assign II26877 = ((~II26853))|((~II26869));
assign WX7375 = ((~II22346))|((~II22347));
assign II34305 = ((~II34315))|((~II34316));
assign WX836 = (WX773&RESET);
assign WX9661 = ((~WX9629));
assign II22043 = ((~II22045))|((~II22046));
assign WX9389 = (WX10210&WX9390);
assign WX7241 = (WX7178&RESET);
assign II22983 = ((~II22973))|((~II22981));
assign II18575 = ((~II18565))|((~II18573));
assign WX4470 = ((~WX4438));
assign WX191 = ((~WX1003));
assign WX10494 = (WX10492)|(WX10491);
assign II27560 = ((~_2298_))|((~II27558));
assign II35575 = ((~WX10958))|((~_2361_));
assign WX9342 = (_2314_&WX10055);
assign II19112 = ((~WX5755))|((~II19111));
assign WX6291 = (WX6290&WX6177);
assign WX8252 = (WX8255&RESET);
assign WX3542 = ((~WX3514));
assign WX6715 = (WX8875&WX6716);
assign II22213 = ((~II22215))|((~II22216));
assign II30457 = ((~WX10052))|((~WX9724));
assign WX7519 = ((~WX7518));
assign WX8158 = (WX8164&WX8159);
assign II6148 = ((~WX2294))|((~WX1948));
assign WX1165 = ((~WX1164));
assign WX1031 = (WX1029)|(WX1028);
assign WX982 = ((~WX909));
assign II7278 = ((~WX1890))|((~WX1812));
assign WX5743 = ((~WX6119));
assign II31724 = ((~WX9689))|((~_2305_));
assign WX8846 = ((~WX8845));
assign WX1450 = ((~WX2297));
assign WX740 = (WX677&RESET);
assign WX10787 = ((~WX11347));
assign WX5500 = ((~WX5499));
assign II30590 = ((~II30580))|((~II30588));
assign II27546 = ((~_2300_))|((~II27544));
assign II6522 = ((~WX1972))|((~II6520));
assign WX2271 = ((~WX2200));
assign II26469 = ((~WX8623))|((~II26467));
assign II18068 = ((~II18078))|((~II18079));
assign WX1324 = (WX1236&WX1263);
assign II18535 = ((~WX6174))|((~WX5851));
assign II11700 = ((~WX3224))|((~II11699));
assign II6209 = ((~II6211))|((~II6212));
assign WX5095 = ((~II15458))|((~II15459));
assign WX3702 = ((~WX3701));
assign WX9421 = ((~WX9420));
assign WX10703 = ((~WX11347));
assign WX251 = ((~WX1004));
assign WX4332 = ((~WX4323));
assign II6575 = ((~II6565))|((~II6573));
assign WX9960 = ((~II30325))|((~II30326));
assign II23339 = ((~WX6990))|((~II23337));
assign WX2283 = ((~WX2206));
assign WX4199 = (WX6324&WX4200);
assign WX1085 = (WX591&WX1086);
assign WX9545 = (WX9548&RESET);
assign II34608 = ((~II34584))|((~II34600));
assign II7505 = ((~WX1932))|((~_2140_));
assign WX10636 = (DATA_0_13&WX10637);
assign WX882 = (WX819&RESET);
assign II3655 = ((~WX633))|((~II3654));
assign WX465 = ((~WX1004));
assign II10279 = ((~WX3249))|((~II10277));
assign WX9633 = ((~WX9601));
assign II31426 = ((~WX9657))|((~II31425));
assign WX7854 = (WX10091&WX7855);
assign WX471 = ((~WX1003));
assign WX3320 = (WX3257&RESET);
assign WX6946 = ((~WX6937));
assign II27707 = ((~_2275_))|((~II27705));
assign II11503 = ((~_2151_))|((~II11502));
assign WX6820 = ((~WX6811));
assign WX3318 = (WX3255&RESET);
assign II6095 = ((~II6085))|((~II6093));
assign WX7568 = ((~WX7567));
assign WX7097 = ((~WX7342));
assign WX6526 = ((~WX6517));
assign II7241 = ((~WX1806))|((~II7239));
assign WX8919 = (WX8918&WX8763);
assign WX7193 = (WX7130&RESET);
assign II18496 = ((~II18471))|((~II18495));
assign II2661 = ((~II2637))|((~II2653));
assign WX10561 = (WX10572&WX11347);
assign WX1936 = ((~WX2192));
assign II10129 = ((~WX3303))|((~II10121));
assign II10525 = ((~WX3588))|((~WX3265));
assign WX9453 = (WX9451)|(WX9450);
assign II26027 = ((~II26017))|((~II26025));
assign WX10078 = ((~II31127))|((~II31128));
assign WX9150 = (WX9544&WX10055);
assign WX7398 = ((~WX7397));
assign II26841 = ((~WX8647))|((~II26839));
assign WX10769 = ((~WX10760));
assign II26064 = ((~WX8533))|((~WX8597));
assign II6425 = ((~II6435))|((~II6436));
assign WX8438 = (WX8058&RESET);
assign WX10627 = ((~WX11348));
assign II2227 = ((~II2203))|((~II2219));
assign WX7561 = ((~WX7560));
assign WX6796 = ((~WX7468));
assign WX7995 = ((~WX8762));
assign II10384 = ((~II10386))|((~II10387));
assign WX7545 = (WX7543)|(WX7542);
assign WX1633 = (WX1631)|(WX1630);
assign WX11473 = (WX11471)|(WX11470);
assign WX1501 = (WX3682&WX1502);
assign WX10874 = (WX10877&RESET);
assign WX3266 = (WX2886&RESET);
assign WX8229 = ((~WX8761));
assign WX5676 = (WX5679&RESET);
assign WX9218 = ((~WX10055));
assign WX9515 = (WX10273&WX9516);
assign WX9087 = (WX9093&WX9088);
assign II15160 = ((~WX4378))|((~II15158));
assign WX2501 = ((~WX2500));
assign WX1880 = ((~WX1848));
assign WX8667 = ((~II26320))|((~II26321));
assign II22563 = ((~II22538))|((~II22562));
assign II14074 = ((~II14064))|((~II14072));
assign WX10157 = (WX9645&WX10158);
assign WX3014 = (WX3020&WX3015);
assign WX366 = (DATA_9_8&WX367);
assign WX4879 = ((~TM1));
assign II22571 = ((~WX7467))|((~WX7146));
assign WX85 = (WX491&WX1004);
assign II2593 = ((~WX811))|((~II2592));
assign WX7370 = ((~II22191))|((~II22192));
assign WX7696 = ((~II23503))|((~II23504));
assign II19529 = ((~II19519))|((~II19527));
assign WX6333 = (WX6332&WX6177);
assign WX6583 = ((~WX6582));
assign WX5377 = ((~WX6175));
assign WX3604 = ((~WX3603));
assign II19424 = ((~WX5779))|((~II19423));
assign WX3509 = ((~II10734))|((~II10735));
assign WX8564 = (WX8501&RESET);
assign WX2254 = ((~WX2253));
assign WX8214 = (WX8220&WX8215);
assign WX7137 = (WX6709&RESET);
assign II22430 = ((~II22432))|((~II22433));
assign WX5590 = (WX7666&WX5591);
assign WX6492 = (WX6410&WX6435);
assign II19398 = ((~WX5777))|((~II19397));
assign WX9320 = ((~WX10055));
assign WX9668 = ((~WX9898));
assign WX6173 = ((~WX6172));
assign II18595 = ((~II18605))|((~II18606));
assign II10572 = ((~WX3395))|((~II10571));
assign WX337 = (WX527&WX1004);
assign II18078 = ((~WX5885))|((~II18077));
assign WX7904 = ((~WX7903));
assign WX6558 = ((~WX7468));
assign WX325 = ((~WX1004));
assign WX6930 = ((~WX7469));
assign II30211 = ((~WX9708))|((~II30209));
assign WX3610 = (WX3608)|(WX3607);
assign II26931 = ((~II26933))|((~II26934));
assign II26048 = ((~II26050))|((~II26051));
assign WX5005 = (WX5004&WX4884);
assign WX3847 = ((~II11714))|((~II11715));
assign WX9681 = ((~WX9924));
assign WX4014 = ((~WX4882));
assign II30621 = ((~II30611))|((~II30619));
assign WX9304 = (WX9566&WX10055);
assign WX3964 = (WX4370&WX4883);
assign WX5457 = ((~WX5448));
assign WX7548 = ((~II23221))|((~II23222));
assign WX7915 = ((~WX8762));
assign WX341 = ((~WX332));
assign II18688 = ((~II18698))|((~II18699));
assign WX9489 = (WX9487)|(WX9486);
assign WX7179 = (WX7116&RESET);
assign WX11386 = (WX11385&WX11349);
assign WX5295 = (_2230_&WX6176);
assign WX3852 = (WX3848&WX3849);
assign WX11584 = ((~II35597))|((~II35598));
assign WX6205 = ((~WX6204));
assign WX1750 = ((~WX2296));
assign II3223 = ((~WX511))|((~II3221));
assign WX6575 = (WX8805&WX6576);
assign II30512 = ((~II30502))|((~II30510));
assign WX1584 = (_2122_&WX2297);
assign WX9553 = (WX9556&RESET);
assign WX5878 = (WX5654&RESET);
assign II14841 = ((~WX4881))|((~II14840));
assign WX442 = (WX448&WX443);
assign WX4401 = (WX4404&RESET);
assign WX8074 = (WX8080&WX8075);
assign WX11297 = ((~WX11296));
assign WX4256 = ((~WX4883));
assign II34585 = ((~II34587))|((~II34588));
assign WX7653 = ((~II23416))|((~II23417));
assign WX6265 = ((~WX6177));
assign WX4512 = ((~WX4758));
assign WX11030 = (WX10686&RESET);
assign II14794 = ((~WX4702))|((~II14793));
assign II10198 = ((~II10200))|((~II10201));
assign WX11182 = (WX11119&RESET);
assign WX10235 = ((~WX10056));
assign II14330 = ((~WX4736))|((~II14328));
assign WX2460 = ((~II7357))|((~II7358));
assign WX10053 = ((~WX10049));
assign WX10542 = (WX11433&WX10543);
assign WX1987 = (WX1691&RESET);
assign II22727 = ((~WX7467))|((~II22726));
assign II14469 = ((~WX4880))|((~II14468));
assign II18413 = ((~WX5843))|((~II18411));
assign II10270 = ((~II10260))|((~II10268));
assign WX5242 = (WX5240)|(WX5239);
assign WX872 = (WX809&RESET);
assign II34701 = ((~II34677))|((~II34693));
assign II5991 = ((~II6001))|((~II6002));
assign WX7675 = (WX7674&WX7470);
assign WX11465 = ((~WX11349));
assign WX3147 = ((~WX3577));
assign WX10988 = (WX10392&RESET);
assign II7110 = ((~WX1877))|((~II7109));
assign WX10572 = (WX10570)|(WX10569);
assign WX7108 = ((~WX7364));
assign WX108 = (WX106)|(WX105);
assign WX4892 = ((~II15081))|((~II15082));
assign WX10111 = ((~WX10110));
assign II30690 = ((~WX9866))|((~II30689));
assign II26444 = ((~II26419))|((~II26443));
assign WX636 = ((~WX885));
assign II10237 = ((~II10213))|((~II10229));
assign II35497 = ((~WX10891))|((~II35495));
assign II6884 = ((~II6859))|((~II6883));
assign II35237 = ((~WX10851))|((~II35235));
assign WX1875 = ((~WX1843));
assign II34160 = ((~WX11061))|((~II34159));
assign WX7606 = (WX7064&WX7607);
assign WX6763 = (WX6761)|(WX6760);
assign WX9534 = ((~WX9536));
assign WX9705 = (WX9169&RESET);
assign WX7755 = (WX7717&WX7728);
assign II18893 = ((~WX6065))|((~II18891));
assign WX2680 = (WX2678)|(WX2677);
assign II22077 = ((~WX7114))|((~II22075));
assign WX7213 = (WX7150&RESET);
assign II22852 = ((~WX7164))|((~II22850));
assign II14382 = ((~WX4612))|((~II14374));
assign WX2805 = ((~WX3589));
assign WX4657 = (WX4594&RESET);
assign II2668 = ((~II2678))|((~II2679));
assign II26988 = ((~II26978))|((~II26986));
assign II22555 = ((~WX7272))|((~WX7336));
assign WX5232 = (WX5230)|(WX5229);
assign WX6281 = ((~WX6280));
assign WX5009 = ((~WX5008));
assign WX8550 = (WX8487&RESET);
assign WX4924 = (WX4922)|(WX4921);
assign II22300 = ((~WX7192))|((~II22299));
assign WX6300 = ((~WX6177));
assign WX114 = (DATA_9_26&WX115);
assign WX6783 = (WX6781)|(WX6780);
assign WX8006 = (WX8004)|(WX8003);
assign II31649 = ((~_2318_))|((~II31647));
assign WX9506 = (WX9517&WX10054);
assign WX6647 = (WX6645)|(WX6644);
assign WX1196 = (WX1195&WX1005);
assign II2374 = ((~II2376))|((~II2377));
assign II18133 = ((~WX6173))|((~II18132));
assign WX2671 = (WX3077&WX3590);
assign WX7711 = ((~II23624))|((~II23625));
assign WX648 = (WX76&RESET);
assign II35340 = ((~WX10943))|((~II35339));
assign WX6694 = ((~WX6685));
assign WX9368 = ((~WX10054));
assign II31348 = ((~WX9651))|((~II31347));
assign II14321 = ((~WX4608))|((~II14320));
assign WX2137 = (WX2074&RESET);
assign II2840 = ((~WX827))|((~WX891));
assign II11181 = ((~WX3089))|((~II11179));
assign WX4190 = ((~WX4883));
assign II18488 = ((~WX5975))|((~WX6039));
assign WX9254 = (WX9265&WX10054);
assign II27135 = ((~WX8342))|((~II27134));
assign II2238 = ((~WX661))|((~II2236));
assign II30674 = ((~WX10053))|((~WX9738));
assign WX6129 = ((~WX6128));
assign WX2593 = (WX2541&WX2556);
assign II18256 = ((~WX6173))|((~WX5833));
assign II22586 = ((~WX7274))|((~WX7338));
assign WX7458 = ((~WX7457));
assign WX1799 = (WX1802&RESET);
assign WX8053 = (WX8279&WX8762);
assign WX3070 = (WX3073&RESET);
assign WX5169 = (WX5131&WX5142);
assign II14924 = ((~II14900))|((~II14916));
assign WX9391 = (WX9389)|(WX9388);
assign WX4130 = ((~WX4883));
assign II35250 = ((~WX10853))|((~II35248));
assign II26475 = ((~II26450))|((~II26474));
assign II6869 = ((~WX2058))|((~II6868));
assign WX265 = ((~WX1004));
assign II22170 = ((~WX7120))|((~II22168));
assign II18527 = ((~II18502))|((~II18526));
assign WX5102 = ((~II15471))|((~II15472));
assign WX7353 = (WX7290&RESET);
assign WX7045 = ((~WX7013));
assign WX5531 = ((~WX6175));
assign WX9595 = (WX9598&RESET);
assign WX8128 = ((~WX8127));
assign WX3021 = (WX3127&WX3590);
assign WX11490 = ((~II35353))|((~II35354));
assign II26109 = ((~II26119))|((~II26120));
assign II14428 = ((~II14404))|((~II14420));
assign II10069 = ((~II10059))|((~II10067));
assign II6832 = ((~WX1992))|((~II6830));
assign WX9573 = (WX9576&RESET);
assign WX1615 = (WX1613)|(WX1612);
assign WX2007 = (WX1944&RESET);
assign II34857 = ((~II34832))|((~II34856));
assign WX3042 = (WX3048&WX3043);
assign WX11340 = ((~TM0));
assign WX2928 = ((~WX2927));
assign WX2855 = ((~WX3590));
assign WX9988 = ((~WX9987));
assign WX261 = ((~WX1003));
assign II26343 = ((~WX8551))|((~WX8615));
assign WX961 = ((~WX960));
assign WX10303 = ((~II31676))|((~II31677));
assign WX4922 = (WX4464&WX4923);
assign WX7063 = ((~WX7031));
assign II14731 = ((~WX4698))|((~WX4762));
assign WX3055 = (WX3066&WX3589);
assign II31154 = ((~WX9546))|((~II31152));
assign II18790 = ((~WX5931))|((~II18782));
assign II3442 = ((~WX610))|((~WX545));
assign WX1027 = ((~II3092))|((~II3093));
assign WX666 = (WX202&RESET);
assign WX10195 = ((~WX10194));
assign II31114 = ((~WX9633))|((~II31113));
assign WX10554 = (WX10552)|(WX10551);
assign II26367 = ((~WX8489))|((~II26366));
assign II2555 = ((~II2545))|((~II2553));
assign WX4984 = (WX4983&WX4884);
assign II18947 = ((~II18937))|((~II18945));
assign WX7181 = (WX7118&RESET);
assign WX9621 = ((~WX9996));
assign II19191 = ((~WX5675))|((~II19189));
assign WX6605 = (WX6603)|(WX6602);
assign II15713 = ((~_2175_))|((~II15711));
assign II30645 = ((~WX9736))|((~II30643));
assign WX4798 = ((~II14615))|((~II14616));
assign WX6024 = (WX5961&RESET);
assign WX402 = (WX400)|(WX399);
assign WX4244 = (WX4410&WX4883);
assign WX8211 = ((~WX8202));
assign WX8235 = (WX8305&WX8762);
assign WX6717 = (WX6715)|(WX6714);
assign WX520 = (WX523&RESET);
assign WX11248 = ((~II34175))|((~II34176));
assign WX11344 = ((~TM1));
assign II34678 = ((~II34680))|((~II34681));
assign WX8348 = ((~WX8316));
assign WX1555 = (WX1553)|(WX1552);
assign WX8690 = ((~WX8674));
assign WX3370 = (WX3307&RESET);
assign II19385 = ((~WX5776))|((~II19384));
assign II31205 = ((~WX9640))|((~II31204));
assign II27565 = ((~WX8372))|((~_2297_));
assign WX5818 = (WX5234&RESET);
assign WX4541 = (WX4053&RESET);
assign II2539 = ((~II2529))|((~II2537));
assign II31698 = ((~_2309_))|((~II31696));
assign WX3835 = ((~II11630))|((~II11631));
assign WX2798 = (WX3682&WX2799);
assign II26709 = ((~II26699))|((~II26707));
assign WX3636 = (WX3172&WX3637);
assign WX5724 = ((~WX6145));
assign II2004 = ((~WX773))|((~II2003));
assign II10323 = ((~WX3379))|((~WX3443));
assign WX2912 = (WX2910)|(WX2909);
assign WX6702 = ((~WX7469));
assign II26422 = ((~WX8759))|((~II26421));
assign II11539 = ((~WX3199))|((~II11538));
assign WX10016 = ((~WX10015));
assign WX5602 = (WX5600)|(WX5599);
assign II30944 = ((~II30920))|((~II30936));
assign WX10721 = ((~WX11348));
assign WX8308 = ((~WX8727));
assign WX10288 = ((~II31571))|((~II31572));
assign WX4880 = ((~WX4879));
assign WX10045 = ((~WX9966));
assign WX7803 = ((~WX8762));
assign II10557 = ((~WX3588))|((~II10556));
assign WX5624 = (WX5622)|(WX5621);
assign WX3066 = (WX3064)|(WX3063);
assign WX856 = (WX793&RESET);
assign WX2705 = (WX2716&WX3589);
assign II14507 = ((~WX4620))|((~II14506));
assign II10013 = ((~WX3359))|((~WX3423));
assign WX593 = ((~WX561));
assign WX10689 = ((~WX11347));
assign WX10211 = ((~II31374))|((~II31375));
assign WX10417 = ((~WX11348));
assign WX9379 = ((~WX9378));
assign WX7944 = (WX7942)|(WX7941);
assign WX2920 = (WX5038&WX2921);
assign WX10897 = ((~WX11319));
assign WX5814 = ((~WX6069));
assign WX4791 = ((~II14398))|((~II14399));
assign WX6367 = ((~II19424))|((~II19425));
assign WX7029 = ((~WX7398));
assign WX3557 = ((~WX3556));
assign WX9693 = ((~WX9948));
assign WX916 = ((~II2507))|((~II2508));
assign WX2916 = (WX2922&WX2917);
assign WX9688 = ((~WX9938));
assign WX4155 = (WX4153)|(WX4152);
assign II26826 = ((~WX8455))|((~II26824));
assign II26807 = ((~II26809))|((~II26810));
assign II27408 = ((~WX8363))|((~II27407));
assign WX2717 = ((~WX2708));
assign WX4276 = ((~WX4267));
assign II26933 = ((~WX8589))|((~II26932));
assign II31543 = ((~_2304_))|((~II31542));
assign WX8389 = ((~WX8633));
assign II7436 = ((~WX1836))|((~II7434));
assign WX6186 = (WX6185&WX6177);
assign WX11268 = ((~II34795))|((~II34796));
assign WX7468 = ((~WX7464));
assign II23665 = ((~WX7095))|((~_2249_));
assign II11533 = ((~_2171_))|((~II11531));
assign II14749 = ((~WX4572))|((~II14747));
assign WX6162 = ((~WX6085));
assign WX9374 = (WX9576&WX10055);
assign WX4279 = (WX4285&WX4280);
assign II34579 = ((~II34569))|((~II34577));
assign II23195 = ((~WX7054))|((~II23194));
assign WX7623 = ((~WX7622));
assign WX8612 = (WX8549&RESET);
assign II14754 = ((~WX4636))|((~II14746));
assign WX2194 = ((~II6047))|((~II6048));
assign II34570 = ((~WX11151))|((~WX11215));
assign II11721 = ((~WX3228))|((~II11720));
assign II10246 = ((~WX3587))|((~WX3247));
assign II18511 = ((~WX5913))|((~II18503));
assign WX2252 = ((~WX2251));
assign WX5019 = (WX5018&WX4884);
assign WX6597 = ((~WX6596));
assign WX2301 = (WX1873&WX2302);
assign WX4062 = (WX4384&WX4883);
assign II26033 = ((~WX8531))|((~WX8595));
assign II18109 = ((~WX5887))|((~II18108));
assign WX5735 = ((~WX6167));
assign WX3484 = (WX3421&RESET);
assign WX8504 = (WX8441&RESET);
assign II10554 = ((~II10564))|((~II10565));
assign WX11164 = (WX11101&RESET);
assign WX4343 = (WX5101&WX4344);
assign II6674 = ((~II6676))|((~II6677));
assign II22291 = ((~II22293))|((~II22294));
assign II2778 = ((~WX823))|((~WX887));
assign II18885 = ((~II18875))|((~II18883));
assign WX6609 = (WX6607)|(WX6606);
assign WX7005 = (WX7008&RESET);
assign II7653 = ((~WX1924))|((~II7652));
assign WX6747 = (WX7596&WX6748);
assign WX9673 = ((~WX9908));
assign WX924 = ((~II2755))|((~II2756));
assign WX5370 = (WX6261&WX5371);
assign WX2523 = ((~RESET));
assign II22061 = ((~WX7304))|((~II22059));
assign WX8961 = (WX8960&WX8763);
assign WX2640 = (WX4898&WX2641);
assign WX6120 = ((~WX6096));
assign WX2959 = ((~WX3589));
assign WX9873 = (WX9810&RESET);
assign WX175 = (WX186&WX1003);
assign II6010 = ((~WX2130))|((~II6008));
assign WX564 = ((~WX933));
assign II14980 = ((~WX4714))|((~II14979));
assign II10942 = ((~II10944))|((~II10945));
assign II6381 = ((~WX2090))|((~II6380));
assign WX3040 = ((~WX3039));
assign II11651 = ((~WX3216))|((~II11650));
assign II11088 = ((~WX3168))|((~WX3075));
assign WX2288 = ((~WX2287));
assign WX625 = ((~WX863));
assign II34765 = ((~II34755))|((~II34763));
assign WX2815 = ((~WX2806));
assign WX1336 = (WX1778&WX2297);
assign WX411 = ((~WX402));
assign WX6073 = ((~II18062))|((~II18063));
assign II10339 = ((~WX3587))|((~WX3253));
assign WX8822 = (WX8346&WX8823);
assign II14593 = ((~WX4881))|((~II14592));
assign II7070 = ((~WX1874))|((~WX1780));
assign II7059 = ((~WX1778))|((~II7057));
assign WX10962 = ((~WX11193));
assign WX5471 = ((~WX5462));
assign WX9011 = ((~II27678))|((~II27679));
assign WX4052 = ((~WX4043));
assign II14676 = ((~II14652))|((~II14668));
assign II14373 = ((~II14383))|((~II14384));
assign WX2524 = ((~II7483))|((~II7484));
assign II26902 = ((~WX8587))|((~II26901));
assign WX2557 = (WX2527&WX2556);
assign WX2647 = ((~WX2638));
assign II35003 = ((~II35005))|((~II35006));
assign WX10522 = (WX10520)|(WX10519);
assign WX2823 = ((~WX3590));
assign WX3229 = ((~WX3485));
assign WX2963 = ((~WX3590));
assign II23456 = ((~WX7008))|((~II23454));
assign II22848 = ((~II22858))|((~II22859));
assign WX9665 = ((~WX9892));
assign WX600 = ((~WX568));
assign II2128 = ((~WX781))|((~II2127));
assign II6784 = ((~WX2116))|((~II6783));
assign WX5660 = (WX5663&RESET);
assign WX10513 = (WX10847&WX11348);
assign WX538 = (WX541&RESET);
assign II15669 = ((~WX4512))|((~_2182_));
assign II30161 = ((~II30163))|((~II30164));
assign II34556 = ((~WX11346))|((~II34555));
assign WX3556 = ((~WX3489));
assign WX8552 = (WX8489&RESET);
assign WX10813 = (WX10824&WX11347);
assign WX6241 = ((~II19190))|((~II19191));
assign WX1476 = (WX1798&WX2297);
assign WX4965 = ((~WX4884));
assign WX8278 = (WX8281&RESET);
assign WX3937 = (WX4898&WX3938);
assign II2134 = ((~II2110))|((~II2126));
assign WX7161 = (WX6877&RESET);
assign II27160 = ((~WX8344))|((~WX8255));
assign II6550 = ((~II6552))|((~II6553));
assign WX4352 = (_2173_&WX4883);
assign II30342 = ((~II30332))|((~II30340));
assign II10222 = ((~WX3309))|((~II10214));
assign WX6568 = ((~WX6559));
assign DATA_9_7 = ((~WX1179));
assign WX3452 = (WX3389&RESET);
assign WX10275 = (WX10274&WX10056);
assign WX5318 = ((~WX5317));
assign II11272 = ((~WX3103))|((~II11270));
assign II14801 = ((~II14776))|((~II14800));
assign WX11450 = (WX10938&WX11451);
assign WX6563 = (WX6561)|(WX6560);
assign WX2689 = ((~WX2680));
assign II34045 = ((~WX11181))|((~II34043));
assign II26761 = ((~II26763))|((~II26764));
assign II6217 = ((~WX2016))|((~II6209));
assign WX8913 = (WX8359&WX8914);
assign II1996 = ((~WX709))|((~II1995));
assign WX4002 = (_2198_&WX4883);
assign II30862 = ((~WX9750))|((~II30860));
assign II18799 = ((~WX5995))|((~II18798));
assign II14500 = ((~WX4881))|((~II14499));
assign II35561 = ((~WX10956))|((~_2363_));
assign WX4175 = (WX5017&WX4176);
assign WX1286 = (WX1232&WX1263);
assign WX7496 = (WX7494)|(WX7493);
assign WX8094 = (WX8092)|(WX8091);
assign WX1116 = ((~WX1115));
assign WX4132 = (WX4394&WX4883);
assign WX3723 = ((~WX3722));
assign II34532 = ((~WX11085))|((~II34531));
assign II26647 = ((~II26637))|((~II26645));
assign II27003 = ((~II26993))|((~II27001));
assign WX7627 = (WX7067&WX7628);
assign II22083 = ((~WX7178))|((~II22082));
assign II10161 = ((~WX3305))|((~II10160));
assign II2399 = ((~WX735))|((~II2398));
assign WX7872 = (WX8805&WX7873);
assign WX2711 = ((~WX3590));
assign WX5894 = (WX5831&RESET);
assign WX6320 = (WX5772&WX6321);
assign II30331 = ((~II30341))|((~II30342));
assign WX6386 = ((~WX6385));
assign II34461 = ((~II34463))|((~II34464));
assign WX5508 = (WX5506)|(WX5505);
assign II34455 = ((~II34445))|((~II34453));
assign II2392 = ((~WX1001))|((~II2391));
assign WX11396 = (WX11394)|(WX11393);
assign WX987 = ((~WX986));
assign II3208 = ((~WX592))|((~WX509));
assign II7305 = ((~WX1892))|((~II7304));
assign WX3841 = ((~II11672))|((~II11673));
assign WX6767 = (WX6773&WX6768);
assign WX5142 = ((~WX5109));
assign WX3185 = ((~WX3153));
assign WX3571 = ((~WX3570));
assign II6512 = ((~II6487))|((~II6511));
assign WX2457 = (WX2455)|(WX2454);
assign II34842 = ((~WX11105))|((~II34841));
assign II34554 = ((~II34556))|((~II34557));
assign II6350 = ((~WX2088))|((~II6349));
assign WX6416 = ((~II19605))|((~II19606));
assign WX6090 = ((~II18589))|((~II18590));
assign WX3683 = ((~II11232))|((~II11233));
assign WX11321 = ((~WX11320));
assign WX4009 = (WX4007)|(WX4006);
assign WX4487 = ((~WX4455));
assign WX3985 = (WX3991&WX3986);
assign II34508 = ((~WX11147))|((~WX11211));
assign II22773 = ((~WX7286))|((~II22772));
assign WX7612 = (WX7611&WX7470);
assign II15572 = ((~WX4496))|((~II15571));
assign WX978 = ((~WX907));
assign WX1811 = (WX1814&RESET);
assign WX5950 = (WX5887&RESET);
assign WX7685 = (WX7683)|(WX7682);
assign II14413 = ((~WX4614))|((~II14405));
assign II11376 = ((~WX3119))|((~II11374));
assign WX7985 = ((~WX8762));
assign WX5367 = ((~WX6176));
assign II34228 = ((~II34230))|((~II34231));
assign II7434 = ((~WX1902))|((~WX1836));
assign WX2368 = ((~WX2367));
assign WX2057 = (WX1994&RESET);
assign WX11116 = (WX11053&RESET);
assign WX11210 = (WX11147&RESET);
assign WX557 = ((~WX983));
assign WX8986 = ((~WX8985));
assign WX9745 = (WX9449&RESET);
assign II6535 = ((~WX2100))|((~WX2164));
assign WX2903 = ((~WX3589));
assign WX2234 = ((~WX2233));
assign WX1537 = ((~WX1536));
assign II14606 = ((~II14608))|((~II14609));
assign WX1105 = (WX1104&WX1005);
assign II35495 = ((~WX10955))|((~WX10891));
assign II26815 = ((~II26791))|((~II26807));
assign WX10932 = ((~WX10900));
assign WX4803 = ((~II14770))|((~II14771));
assign WX6269 = ((~II19242))|((~II19243));
assign II30147 = ((~WX10052))|((~WX9704));
assign WX198 = (DATA_9_20&WX199);
assign WX4951 = ((~WX4884));
assign II34569 = ((~II34571))|((~II34572));
assign WX4583 = (WX4347&RESET);
assign WX1464 = ((~WX2297));
assign II34392 = ((~II34367))|((~II34391));
assign II26916 = ((~II26918))|((~II26919));
assign WX6710 = (WX6721&WX7468);
assign WX5494 = (WX5492)|(WX5491);
assign II26769 = ((~WX8515))|((~II26761));
assign II7448 = ((~WX1903))|((~II7447));
assign WX613 = ((~WX839));
assign II22223 = ((~II22213))|((~II22221));
assign WX4447 = ((~WX4820));
assign II31399 = ((~WX9655))|((~WX9584));
assign II26383 = ((~II26373))|((~II26381));
assign II6667 = ((~II6642))|((~II6666));
assign WX2259 = ((~WX2194));
assign WX9982 = ((~II31007))|((~II31008));
assign WX7169 = (WX6933&RESET);
assign II14221 = ((~WX4880))|((~II14220));
assign WX5522 = (WX5520)|(WX5519);
assign WX2991 = ((~WX3590));
assign WX9038 = (WX9014&WX9021);
assign WX5070 = ((~WX4884));
assign WX4167 = (WX4173&WX4168);
assign WX3546 = ((~WX3516));
assign II22137 = ((~WX7466))|((~WX7118));
assign II6305 = ((~WX1958))|((~II6303));
assign WX1542 = (_2125_&WX2297);
assign II22446 = ((~II22448))|((~II22449));
assign II6800 = ((~WX2295))|((~II6799));
assign WX4467 = ((~WX4435));
assign II2803 = ((~II2793))|((~II2801));
assign WX5341 = (WX5675&WX6176);
assign II14120 = ((~II14110))|((~II14118));
assign II6768 = ((~WX2295))|((~WX1988));
assign WX3657 = (WX3175&WX3658);
assign WX5287 = ((~WX6176));
assign WX11367 = ((~WX11349));
assign WX6818 = ((~WX7469));
assign WX6506 = ((~WX7469));
assign WX5350 = (WX5348)|(WX5347);
assign WX7512 = ((~WX7511));
assign WX6832 = ((~WX7469));
assign WX11638 = (WX11594&WX11607);
assign II22981 = ((~WX7236))|((~II22973));
assign II30069 = ((~WX9826))|((~WX9890));
assign II26715 = ((~WX8575))|((~WX8639));
assign WX10028 = ((~WX10027));
assign II10331 = ((~II10306))|((~II10330));
assign WX2198 = ((~II6171))|((~II6172));
assign WX514 = (WX517&RESET);
assign II15571 = ((~WX4496))|((~_2198_));
assign II3640 = ((~WX630))|((~_2089_));
assign II10881 = ((~WX3415))|((~WX3479));
assign WX5297 = ((~WX6176));
assign WX8766 = (WX8338&WX8767);
assign II2351 = ((~II2327))|((~II2343));
assign WX5453 = (WX5691&WX6176);
assign WX2699 = (WX3081&WX3590);
assign II6227 = ((~WX2144))|((~II6225));
assign II30285 = ((~II30287))|((~II30288));
assign II23482 = ((~WX7012))|((~II23480));
assign WX11310 = ((~WX11245));
assign WX9529 = (WX10280&WX9530);
assign WX9271 = (WX9269)|(WX9268);
assign II26793 = ((~WX8760))|((~WX8453));
assign II11489 = ((~II11479))|((~II11487));
assign II30093 = ((~WX9764))|((~II30092));
assign II10728 = ((~WX3469))|((~II10726));
assign WX5397 = (WX5683&WX6176);
assign WX2999 = (WX3010&WX3589);
assign II10619 = ((~WX3588))|((~II10618));
assign WX10347 = (WX10282&WX10314);
assign II14361 = ((~WX4738))|((~II14359));
assign WX6668 = (WX6679&WX7468);
assign WX3412 = (WX3349&RESET);
assign II3314 = ((~WX525))|((~II3312));
assign WX2694 = (WX2692)|(WX2691);
assign WX4961 = ((~WX4960));
assign II35568 = ((~WX10957))|((~_2362_));
assign WX6304 = ((~II19307))|((~II19308));
assign WX8339 = ((~WX8307));
assign WX4937 = ((~WX4884));
assign WX9647 = ((~WX9615));
assign II22516 = ((~WX7206))|((~II22508));
assign WX3491 = ((~II10176))|((~II10177));
assign WX8994 = ((~II27559))|((~II27560));
assign WX6635 = (WX7540&WX6636);
assign WX903 = ((~II2104))|((~II2105));
assign II26165 = ((~II26140))|((~II26164));
assign WX1523 = ((~WX1522));
assign II3507 = ((~_2080_))|((~II3499));
assign II2274 = ((~WX727))|((~II2266));
assign WX1398 = (WX1409&WX2296);
assign WX7635 = ((~WX7470));
assign WX3300 = (WX3237&RESET);
assign II35262 = ((~WX10937))|((~II35261));
assign WX5048 = (WX4482&WX5049);
assign WX3478 = (WX3415&RESET);
assign WX3056 = (WX3062&WX3057);
assign WX6709 = ((~WX6708));
assign II30241 = ((~WX10052))|((~II30240));
assign WX9512 = ((~WX10055));
assign WX5011 = ((~II15302))|((~II15303));
assign WX4330 = ((~WX4883));
assign WX8366 = ((~WX8334));
assign WX3414 = (WX3351&RESET);
assign WX5282 = (WX7512&WX5283);
assign WX7553 = ((~WX7552));
assign WX7862 = ((~WX7861));
assign II15705 = ((~WX4517))|((~II15704));
assign WX8977 = ((~WX8763));
assign WX7885 = (WX8255&WX8762);
assign II15600 = ((~WX4500))|((~II15599));
assign II6549 = ((~II6559))|((~II6560));
assign WX8662 = ((~II26165))|((~II26166));
assign WX2109 = (WX2046&RESET);
assign WX552 = ((~WX973));
assign II31745 = ((~WX9693))|((~_2301_));
assign II14947 = ((~II14949))|((~II14950));
assign II15277 = ((~WX4396))|((~II15275));
assign II27531 = ((~WX8397))|((~II27530));
assign II11311 = ((~WX3109))|((~II11309));
assign II30920 = ((~II30930))|((~II30931));
assign II22115 = ((~II22105))|((~II22113));
assign WX5346 = ((~WX5345));
assign II14661 = ((~WX4630))|((~II14653));
assign II10317 = ((~II10307))|((~II10315));
assign II26228 = ((~II26218))|((~II26226));
assign II31282 = ((~WX9646))|((~WX9566));
assign WX332 = (WX330)|(WX329);
assign II34998 = ((~II34988))|((~II34996));
assign II3613 = ((~WX625))|((~II3612));
assign WX10764 = (WX10762)|(WX10761);
assign WX9911 = (WX9848&RESET);
assign WX2727 = (WX3085&WX3590);
assign WX7631 = ((~WX7630));
assign WX5029 = (WX5027)|(WX5026);
assign WX11337 = ((~WX11336));
assign WX1565 = ((~WX1564));
assign WX5694 = (WX5697&RESET);
assign II22525 = ((~WX7270))|((~II22524));
assign II2818 = ((~II2808))|((~II2816));
assign II15662 = ((~WX4510))|((~_2184_));
assign WX2589 = (WX2524&WX2556);
assign II22324 = ((~WX7466))|((~II22323));
assign WX10613 = ((~WX11348));
assign II18543 = ((~WX5915))|((~II18542));
assign II34151 = ((~II34153))|((~II34154));
assign WX5408 = (WX7575&WX5409);
assign WX10529 = ((~WX11348));
assign WX103 = ((~WX94));
assign WX6426 = ((~II19675))|((~II19676));
assign WX1459 = (WX3661&WX1460);
assign WX11056 = (WX10993&RESET);
assign II6737 = ((~WX2295))|((~WX1986));
assign WX122 = (WX120)|(WX119);
assign II30054 = ((~WX10052))|((~WX9698));
assign II26784 = ((~II26760))|((~II26776));
assign WX6726 = ((~WX7468));
assign II2454 = ((~WX1001))|((~II2453));
assign WX9076 = (WX8997&WX9021);
assign WX11258 = ((~II34485))|((~II34486));
assign WX8578 = (WX8515&RESET);
assign WX8327 = ((~WX8701));
assign WX3927 = ((~WX3926));
assign II23144 = ((~WX6960))|((~II23142));
assign WX9259 = (WX11440&WX9260);
assign WX820 = (WX757&RESET);
assign WX943 = ((~WX942));
assign II15726 = ((~WX4521))|((~II15725));
assign WX8902 = ((~WX8901));
assign WX7464 = ((~TM1));
assign II10145 = ((~II10120))|((~II10144));
assign II30581 = ((~WX10053))|((~WX9732));
assign II22399 = ((~II22401))|((~II22402));
assign WX1361 = (WX3612&WX1362);
assign WX9721 = (WX9281&RESET);
assign WX3790 = (WX3194&WX3791);
assign II11519 = ((~II11509))|((~II11517));
assign II30769 = ((~WX9744))|((~II30767));
assign WX10399 = ((~WX11348));
assign WX2316 = ((~WX2298));
assign WX9937 = (WX9874&RESET);
assign WX6484 = (WX6414&WX6435);
assign WX10634 = (WX10632)|(WX10631);
assign WX6273 = (WX6271)|(WX6270);
assign WX956 = ((~WX928));
assign II11580 = ((~WX3205))|((~_2164_));
assign II2795 = ((~WX1002))|((~II2794));
assign II14096 = ((~WX4880))|((~WX4530));
assign WX3792 = (WX3790)|(WX3789);
assign WX3406 = (WX3343&RESET);
assign II22478 = ((~WX7466))|((~WX7140));
assign II6473 = ((~WX2096))|((~WX2160));
assign WX2308 = (WX1874&WX2309);
assign WX1602 = (WX1816&WX2297);
assign WX9094 = (WX9536&WX10055);
assign WX11273 = ((~II34950))|((~II34951));
assign WX1590 = ((~WX2297));
assign WX6627 = (WX6633&WX6628);
assign WX10043 = ((~WX9965));
assign WX7508 = (WX7050&WX7509);
assign WX1260 = ((~II3697))|((~II3698));
assign WX8266 = (WX8269&RESET);
assign WX2079 = (WX2016&RESET);
assign II14979 = ((~WX4714))|((~WX4778));
assign II34849 = ((~WX11169))|((~WX11233));
assign WX5860 = (WX5528&RESET);
assign WX6801 = (WX6799)|(WX6798);
assign WX2809 = ((~WX3590));
assign II18381 = ((~WX6173))|((~II18380));
assign WX6517 = (WX6515)|(WX6514);
assign WX6395 = ((~II19476))|((~II19477));
assign II19347 = ((~WX5699))|((~II19345));
assign II6978 = ((~II6968))|((~II6976));
assign WX4144 = ((~WX4883));
assign II2424 = ((~WX673))|((~II2422));
assign WX10682 = (WX11503&WX10683);
assign II14909 = ((~WX4646))|((~II14901));
assign WX4407 = (WX4410&RESET);
assign WX1087 = (WX1085)|(WX1084);
assign WX6775 = (WX7610&WX6776);
assign WX10128 = (WX10127&WX10056);
assign WX11220 = (WX11157&RESET);
assign II30968 = ((~WX9884))|((~WX9948));
assign WX9250 = ((~WX10055));
assign WX7905 = (WX7916&WX8761);
assign WX674 = (WX258&RESET);
assign WX9887 = (WX9824&RESET);
assign II26717 = ((~WX8639))|((~II26715));
assign WX6552 = ((~WX7469));
assign WX8000 = (WX7998)|(WX7997);
assign WX5980 = (WX5917&RESET);
assign II26234 = ((~II26236))|((~II26237));
assign WX10292 = ((~II31599))|((~II31600));
assign WX7578 = (WX7060&WX7579);
assign WX9452 = ((~WX10054));
assign WX7087 = ((~WX7322));
assign WX8244 = (WX8247&RESET);
assign WX10109 = ((~WX10056));
assign WX7586 = ((~WX7470));
assign II15107 = ((~WX4462))|((~II15106));
assign WX6855 = (WX8945&WX6856);
assign II23560 = ((~WX7079))|((~_2265_));
assign WX7529 = (WX7053&WX7530);
assign II19371 = ((~WX5775))|((~WX5703));
assign WX10384 = (DATA_0_31&WX10385);
assign WX3072 = (WX3075&RESET);
assign WX1599 = (WX3731&WX1600);
assign II3080 = ((~WX489))|((~II3078));
assign II2849 = ((~II2839))|((~II2847));
assign WX4253 = (WX4251)|(WX4250);
assign II22401 = ((~WX7262))|((~II22400));
assign II6240 = ((~II6242))|((~II6243));
assign WX2756 = (WX3661&WX2757);
assign II10263 = ((~WX3439))|((~II10261));
assign WX10826 = ((~WX10825));
assign II26041 = ((~II26016))|((~II26040));
assign II22394 = ((~II22384))|((~II22392));
assign II19072 = ((~WX5752))|((~WX5657));
assign II6188 = ((~II6178))|((~II6186));
assign WX10530 = (WX10528)|(WX10527);
assign WX10928 = ((~WX10896));
assign II6459 = ((~WX2294))|((~II6458));
assign WX11533 = (WX11532&WX11349);
assign WX6134 = ((~WX6103));
assign WX11028 = (WX10672&RESET);
assign WX4357 = (WX5108&WX4358);
assign WX2214 = ((~II6667))|((~II6668));
assign II6790 = ((~II6766))|((~II6782));
assign WX794 = (WX731&RESET);
assign II14724 = ((~WX4634))|((~II14723));
assign WX3703 = ((~WX3702));
assign WX4625 = (WX4562&RESET);
assign II6698 = ((~II6673))|((~II6697));
assign WX6151 = ((~WX6150));
assign WX6482 = (WX6415&WX6435);
assign II14466 = ((~II14476))|((~II14477));
assign II26142 = ((~WX8759))|((~WX8411));
assign WX4081 = ((~WX4080));
assign WX212 = (DATA_9_19&WX213);
assign WX8009 = ((~WX8762));
assign WX10407 = (WX10418&WX11347);
assign WX8374 = ((~WX8603));
assign II2429 = ((~WX737))|((~II2421));
assign WX3979 = (WX4919&WX3980);
assign WX7517 = (WX7515)|(WX7514);
assign WX8476 = (WX8413&RESET);
assign II19641 = ((~_2221_))|((~II19639));
assign II6398 = ((~WX1964))|((~II6396));
assign WX11469 = ((~II35314))|((~II35315));
assign WX5646 = (WX7694&WX5647);
assign WX10444 = (WX11384&WX10445);
assign WX1493 = (WX1491)|(WX1490);
assign WX8320 = ((~WX8751));
assign II6211 = ((~WX2294))|((~II6210));
assign WX9504 = ((~WX9495));
assign WX431 = (_2080_&WX1004);
assign II19410 = ((~WX5778))|((~WX5709));
assign II7680 = ((~WX1929))|((~_2115_));
assign II10835 = ((~WX3588))|((~WX3285));
assign WX931 = ((~II2972))|((~II2973));
assign WX2189 = (WX2126&RESET);
assign WX1381 = (WX1379)|(WX1378);
assign II27629 = ((~WX8381))|((~II27628));
assign WX818 = (WX755&RESET);
assign WX10175 = ((~WX10174));
assign WX3221 = ((~WX3469));
assign II34378 = ((~II34368))|((~II34376));
assign WX1416 = (_2134_&WX2297);
assign WX2982 = (WX2980)|(WX2979);
assign II34269 = ((~II34259))|((~II34267));
assign II14080 = ((~WX4656))|((~WX4720));
assign II27279 = ((~WX8273))|((~II27277));
assign II18435 = ((~II18425))|((~II18433));
assign WX4685 = (WX4622&RESET);
assign II18745 = ((~II18735))|((~II18743));
assign WX5776 = ((~WX5744));
assign WX10953 = ((~WX10921));
assign WX9687 = ((~WX9936));
assign WX7571 = (WX7059&WX7572);
assign II30362 = ((~II30372))|((~II30373));
assign II22337 = ((~II22339))|((~II22340));
assign II27082 = ((~WX8338))|((~WX8243));
assign WX4639 = (WX4576&RESET);
assign II34371 = ((~WX11011))|((~II34369));
assign II30626 = ((~II30628))|((~II30629));
assign WX8516 = (WX8453&RESET);
assign II22469 = ((~II22445))|((~II22461));
assign II2475 = ((~II2451))|((~II2467));
assign WX5392 = (WX5390)|(WX5389);
assign II22864 = ((~II22866))|((~II22867));
assign II14265 = ((~II14267))|((~II14268));
assign WX9410 = ((~WX10054));
assign WX4935 = (WX4934&WX4884);
assign WX2869 = ((~WX3590));
assign WX5998 = (WX5935&RESET);
assign WX7044 = ((~WX7428));
assign WX9220 = (WX9554&WX10055);
assign II2114 = ((~WX653))|((~II2112));
assign WX6419 = ((~II19626))|((~II19627));
assign II3183 = ((~WX590))|((~II3182));
assign WX4115 = (WX6282&WX4116);
assign WX11124 = (WX11061&RESET);
assign II30813 = ((~WX9874))|((~WX9938));
assign II34982 = ((~II34972))|((~II34980));
assign II30426 = ((~WX10052))|((~WX9722));
assign II10493 = ((~II10495))|((~II10496));
assign WX8023 = ((~WX8762));
assign II15627 = ((~WX4504))|((~_2190_));
assign WX5055 = (WX4483&WX5056);
assign WX10792 = (WX10790)|(WX10789);
assign WX8807 = (WX8806&WX8763);
assign WX1845 = ((~WX2266));
assign II14414 = ((~WX4614))|((~II14413));
assign WX7647 = (WX7646&WX7470);
assign WX7189 = (WX7126&RESET);
assign WX3982 = ((~WX3973));
assign WX690 = (WX370&RESET);
assign WX4042 = ((~WX4882));
assign WX6579 = (WX7512&WX6580);
assign WX5360 = ((~WX5359));
assign WX11076 = (WX11013&RESET);
assign WX98 = (WX96)|(WX95);
assign II10347 = ((~WX3317))|((~II10346));
assign II35118 = ((~WX10926))|((~WX10833));
assign WX1475 = (WX1473)|(WX1472);
assign II35541 = ((~WX10983))|((~II35540));
assign II7556 = ((~_2135_))|((~II7554));
assign WX9583 = (WX9586&RESET);
assign II31140 = ((~WX9635))|((~II31139));
assign WX3442 = (WX3379&RESET);
assign WX5830 = (WX5318&RESET);
assign II10137 = ((~WX3367))|((~WX3431));
assign II35171 = ((~WX10930))|((~II35170));
assign WX10736 = (WX10734)|(WX10733);
assign WX6880 = ((~WX7468));
assign WX4021 = (WX4940&WX4022);
assign WX11264 = ((~II34671))|((~II34672));
assign II2252 = ((~WX789))|((~II2251));
assign WX4104 = (WX4390&WX4883);
assign WX2320 = ((~II7097))|((~II7098));
assign II11298 = ((~WX3107))|((~II11296));
assign WX2833 = ((~WX3589));
assign II31453 = ((~WX9592))|((~II31451));
assign II10602 = ((~WX3397))|((~WX3461));
assign II10983 = ((~II10973))|((~II10981));
assign WX5805 = ((~WX6051));
assign II26887 = ((~WX8760))|((~II26886));
assign WX5795 = ((~WX6031));
assign WX8406 = (WX7834&RESET);
assign WX10757 = (WX10768&WX11347);
assign WX279 = ((~WX1004));
assign II35737 = ((~WX10984))|((~II35736));
assign WX6353 = ((~II19398))|((~II19399));
assign WX10061 = (WX10059)|(WX10058);
assign WX4221 = ((~WX4220));
assign II18630 = ((~WX5857))|((~II18628));
assign II6002 = ((~II5992))|((~II6000));
assign WX4036 = ((~WX4883));
assign II34618 = ((~WX11346))|((~II34617));
assign WX10713 = ((~WX10704));
assign II30433 = ((~WX9786))|((~II30425));
assign WX10392 = ((~WX10391));
assign II34827 = ((~II34817))|((~II34825));
assign WX3330 = (WX3267&RESET);
assign WX10660 = (WX10666&WX10661);
assign WX10184 = (WX10183&WX10056);
assign II35510 = ((~WX10971))|((~_2364_));
assign WX11404 = ((~WX11403));
assign WX3110 = (WX3113&RESET);
assign II27188 = ((~WX8259))|((~II27186));
assign II11402 = ((~WX3123))|((~II11400));
assign WX10795 = ((~WX11348));
assign WX9005 = ((~II27636))|((~II27637));
assign II35527 = ((~_2364_))|((~II35525));
assign WX2541 = ((~II7618))|((~II7619));
assign II30047 = ((~II30037))|((~II30045));
assign II15657 = ((~_2185_))|((~II15655));
assign WX8817 = (WX8815)|(WX8814);
assign WX2356 = (WX2355&WX2298);
assign WX11489 = ((~WX11488));
assign WX5642 = (WX5648&WX5643);
assign II23272 = ((~WX7060))|((~WX6980));
assign WX1687 = (WX2480&WX1688);
assign WX6195 = ((~WX6177));
assign WX11616 = (WX11577&WX11607);
assign II30386 = ((~II30362))|((~II30378));
assign II22523 = ((~II22525))|((~II22526));
assign II7611 = ((~WX1917))|((~II7610));
assign WX2800 = (WX2798)|(WX2797);
assign II6560 = ((~II6550))|((~II6558));
assign WX5544 = (WX5550&WX5545);
assign WX8542 = (WX8479&RESET);
assign II35210 = ((~WX10933))|((~II35209));
assign II30807 = ((~II30797))|((~II30805));
assign WX8330 = ((~WX8707));
assign II7618 = ((~WX1918))|((~II7617));
assign II18660 = ((~WX6174))|((~II18659));
assign II3549 = ((~WX616))|((~_2103_));
assign WX7664 = (WX7662)|(WX7661);
assign II6924 = ((~WX2295))|((~II6923));
assign WX9324 = (WX9335&WX10054);
assign WX4311 = (WX6380&WX4312);
assign II3492 = ((~_2087_))|((~II3484));
assign WX7387 = ((~II22718))|((~II22719));
assign II34161 = ((~II34151))|((~II34159));
assign WX9144 = ((~WX10054));
assign II6715 = ((~II6705))|((~II6713));
assign II34479 = ((~WX11209))|((~II34477));
assign II19648 = ((~_2219_))|((~II19646));
assign II19176 = ((~WX5760))|((~WX5673));
assign WX7442 = ((~WX7441));
assign II15470 = ((~WX4490))|((~WX4426));
assign WX4295 = (WX4293)|(WX4292);
assign WX7215 = (WX7152&RESET);
assign II35584 = ((~_2360_))|((~II35582));
assign WX8046 = (WX8052&WX8047);
assign II30472 = ((~WX9852))|((~WX9916));
assign WX4326 = ((~WX4883));
assign II22353 = ((~II22355))|((~II22356));
assign II18853 = ((~WX5935))|((~II18852));
assign WX8049 = (_2282_&WX8762);
assign II19124 = ((~WX5756))|((~WX5665));
assign WX7821 = (WX7832&WX8761);
assign WX2710 = (WX4933&WX2711);
assign WX4218 = ((~WX4883));
assign WX5988 = (WX5925&RESET);
assign WX1795 = (WX1798&RESET);
assign WX6631 = (WX8833&WX6632);
assign WX4324 = (_2175_&WX4883);
assign WX635 = ((~WX883));
assign WX8171 = (WX8182&WX8761);
assign WX5561 = (_2211_&WX6176);
assign II10051 = ((~II10027))|((~II10043));
assign II2296 = ((~II2306))|((~II2307));
assign WX4301 = (WX5080&WX4302);
assign WX2504 = (WX1902&WX2505);
assign II10425 = ((~II10415))|((~II10423));
assign WX4245 = (WX5052&WX4246);
assign WX1679 = (WX1685&WX1680);
assign WX6040 = (WX5977&RESET);
assign WX10355 = (WX10297&WX10314);
assign II18240 = ((~WX5959))|((~WX6023));
assign WX11578 = ((~II35555))|((~II35556));
assign WX4759 = (WX4696&RESET);
assign II34757 = ((~WX11163))|((~II34756));
assign II7675 = ((~_2116_))|((~II7673));
assign II26135 = ((~II26125))|((~II26133));
assign II30821 = ((~II30796))|((~II30820));
assign WX4910 = (WX4908)|(WX4907);
assign II18350 = ((~WX6173))|((~II18349));
assign WX8742 = ((~WX8668));
assign WX7920 = (WX7926&WX7921);
assign II23728 = ((~WX7106))|((~_2238_));
assign II34067 = ((~WX11055))|((~II34066));
assign WX8292 = (WX8295&RESET);
assign II30397 = ((~WX9720))|((~II30395));
assign WX934 = ((~WX917));
assign II31640 = ((~WX9675))|((~_2319_));
assign WX1034 = ((~II3105))|((~II3106));
assign WX8340 = ((~WX8308));
assign WX6315 = (WX6313)|(WX6312);
assign WX8620 = (WX8557&RESET);
assign II15069 = ((~WX4364))|((~II15067));
assign II31697 = ((~WX9685))|((~II31696));
assign WX10252 = ((~WX10251));
assign WX4076 = (WX4386&WX4883);
assign WX1357 = (WX1363&WX1358);
assign WX1249 = ((~II3620))|((~II3621));
assign II10354 = ((~WX3381))|((~WX3445));
assign II18637 = ((~II18627))|((~II18635));
assign WX3806 = (WX3804)|(WX3803);
assign II34470 = ((~WX11081))|((~II34469));
assign II2283 = ((~WX791))|((~II2282));
assign WX10906 = ((~WX11337));
assign II30325 = ((~II30300))|((~II30324));
assign WX1240 = ((~II3557))|((~II3558));
assign II30800 = ((~WX9746))|((~II30798));
assign WX572 = ((~WX949));
assign II34803 = ((~WX11346))|((~WX11039));
assign WX9563 = (WX9566&RESET);
assign II31731 = ((~WX9691))|((~_2303_));
assign WX10095 = ((~WX10056));
assign WX8382 = ((~WX8619));
assign DATA_9_16 = ((~WX1116));
assign II31296 = ((~WX9647))|((~II31295));
assign WX9340 = ((~WX10054));
assign WX8198 = ((~WX8197));
assign WX1883 = ((~WX1851));
assign WX8452 = (WX8156&RESET);
assign II6033 = ((~II6023))|((~II6031));
assign II18667 = ((~WX5923))|((~II18666));
assign WX4061 = (WX4059)|(WX4058);
assign WX4563 = (WX4207&RESET);
assign II30186 = ((~WX9770))|((~II30185));
assign WX2636 = (WX2642&WX2637);
assign WX9735 = (WX9379&RESET);
assign II15459 = ((~WX4424))|((~II15457));
assign WX4454 = ((~WX4834));
assign WX3744 = ((~WX3743));
assign II14313 = ((~WX4880))|((~WX4544));
assign WX43 = (WX485&WX1004);
assign II10874 = ((~WX3351))|((~II10873));
assign WX10103 = (WX10101)|(WX10100);
assign II6954 = ((~WX2295))|((~WX2000));
assign WX11514 = ((~WX11349));
assign II2501 = ((~WX869))|((~II2499));
assign WX10536 = (WX10534)|(WX10533);
assign WX9433 = (WX9431)|(WX9430);
assign WX6515 = (WX6521&WX6516);
assign WX1502 = ((~WX2297));
assign WX1612 = (_2120_&WX2297);
assign WX1179 = ((~WX1178));
assign WX2579 = (WX2525&WX2556);
assign WX1372 = ((~WX2296));
assign II19612 = ((~WX5794))|((~II19611));
assign WX7655 = (WX7071&WX7656);
assign II23644 = ((~WX7091))|((~_2253_));
assign WX3539 = ((~WX3538));
assign WX45 = ((~WX1004));
assign II18248 = ((~II18223))|((~II18247));
assign WX2919 = (_2151_&WX3590);
assign II34384 = ((~WX11139))|((~WX11203));
assign II18440 = ((~II18450))|((~II18451));
assign II18156 = ((~II18146))|((~II18154));
assign II14258 = ((~WX4604))|((~II14250));
assign II14933 = ((~WX4881))|((~WX4584));
assign WX1643 = (WX1641)|(WX1640);
assign II7098 = ((~WX1784))|((~II7096));
assign II19732 = ((~_2205_))|((~II19730));
assign II14714 = ((~II14724))|((~II14725));
assign II22841 = ((~II22817))|((~II22833));
assign WX9289 = (WX9287)|(WX9286);
assign II14405 = ((~II14407))|((~II14408));
assign II11630 = ((~WX3212))|((~II11629));
assign WX11576 = ((~II35533))|((~II35534));
assign II26895 = ((~II26885))|((~II26893));
assign WX3717 = ((~WX3716));
assign WX1736 = ((~WX2296));
assign WX5920 = (WX5857&RESET);
assign II14150 = ((~II14125))|((~II14149));
assign II11361 = ((~WX3189))|((~WX3117));
assign WX6925 = (WX8980&WX6926);
assign II22928 = ((~WX7296))|((~II22927));
assign WX1122 = (WX1120)|(WX1119);
assign II26304 = ((~WX8485))|((~II26296));
assign WX5041 = (WX4481&WX5042);
assign WX390 = (WX2480&WX391);
assign II7575 = ((~WX1912))|((~_2132_));
assign WX3527 = ((~WX3526));
assign II26056 = ((~WX8469))|((~II26048));
assign WX1420 = (WX1790&WX2297);
assign II6668 = ((~II6658))|((~II6666));
assign WX1516 = ((~WX2297));
assign WX6595 = (WX6593)|(WX6592);
assign WX9867 = (WX9804&RESET);
assign II22657 = ((~II22647))|((~II22655));
assign WX11413 = ((~II35210))|((~II35211));
assign WX10576 = (WX10582&WX10577);
assign WX894 = (WX831&RESET);
assign WX10121 = (WX10120&WX10056);
assign II11129 = ((~WX3081))|((~II11127));
assign WX9316 = ((~WX10055));
assign II30704 = ((~II30706))|((~II30707));
assign II18154 = ((~II18130))|((~II18146));
assign II2067 = ((~WX841))|((~II2065));
assign WX6084 = ((~II18403))|((~II18404));
assign II14353 = ((~II14343))|((~II14351));
assign WX4983 = ((~II15250))|((~II15251));
assign II34773 = ((~WX11346))|((~II34772));
assign WX5579 = (WX5709&WX6176);
assign II30164 = ((~WX9896))|((~II30162));
assign WX9615 = ((~WX9984));
assign WX230 = ((~WX229));
assign WX9522 = ((~WX10054));
assign WX4235 = ((~WX4234));
assign WX7721 = ((~II23694))|((~II23695));
assign WX5111 = ((~II15508))|((~II15509));
assign WX9173 = (WX9171)|(WX9170);
assign WX8574 = (WX8511&RESET);
assign WX10339 = (WX10304&WX10314);
assign II19619 = ((~WX5795))|((~II19618));
assign II3633 = ((~WX629))|((~_2090_));
assign II10570 = ((~II10572))|((~II10573));
assign II3417 = ((~WX608))|((~II3416));
assign WX10976 = ((~WX11221));
assign WX7197 = (WX7134&RESET);
assign II18177 = ((~II18179))|((~II18180));
assign II19269 = ((~WX5687))|((~II19267));
assign WX7413 = ((~WX7389));
assign II3584 = ((~WX621))|((~_2098_));
assign WX308 = (WX306)|(WX305);
assign II23221 = ((~WX7056))|((~II23220));
assign WX3209 = ((~WX3445));
assign WX3201 = ((~WX3429));
assign WX6081 = ((~II18310))|((~II18311));
assign II10609 = ((~II10585))|((~II10601));
assign II6286 = ((~II6288))|((~II6289));
assign WX11285 = ((~WX11284));
assign II30961 = ((~WX9820))|((~II30960));
assign II26113 = ((~WX8409))|((~II26111));
assign WX7473 = (WX7045&WX7474);
assign WX5595 = ((~WX6176));
assign II22330 = ((~WX7194))|((~II22322));
assign II14020 = ((~WX4716))|((~II14018));
assign WX8942 = ((~WX8763));
assign II10596 = ((~II10586))|((~II10594));
assign WX3520 = ((~WX3503));
assign II2189 = ((~WX785))|((~WX849));
assign II22030 = ((~WX7302))|((~II22028));
assign WX4095 = ((~WX4094));
assign II22463 = ((~WX7266))|((~II22462));
assign II15530 = ((~WX4522))|((~II15529));
assign WX2937 = (WX3115&WX3590);
assign WX3916 = ((~WX4882));
assign WX3626 = ((~WX3625));
assign WX7955 = (WX8265&WX8762);
assign WX10629 = ((~WX10620));
assign WX392 = (WX390)|(WX389);
assign WX1170 = ((~WX1005));
assign II30318 = ((~WX9842))|((~II30317));
assign WX3171 = ((~WX3139));
assign WX9096 = ((~WX10055));
assign WX68 = (WX2319&WX69);
assign WX9446 = ((~WX10055));
assign WX2091 = (WX2028&RESET);
assign WX9895 = (WX9832&RESET);
assign II34748 = ((~WX11099))|((~II34740));
assign II5995 = ((~WX1938))|((~II5993));
assign II35710 = ((~_2340_))|((~II35708));
assign WX9969 = ((~II30604))|((~II30605));
assign WX4186 = ((~WX4883));
assign II2188 = ((~II2190))|((~II2191));
assign II31529 = ((~II31519))|((~II31527));
assign WX6254 = ((~WX6253));
assign WX10692 = (DATA_0_9&WX10693);
assign WX3593 = (WX3592&WX3591);
assign WX2059 = (WX1996&RESET);
assign WX8460 = (WX8212&RESET);
assign WX1004 = ((~WX997));
assign WX4265 = (WX4271&WX4266);
assign WX5321 = ((~WX6175));
assign II26824 = ((~WX8760))|((~WX8455));
assign WX8896 = ((~WX8895));
assign WX4856 = ((~WX4855));
assign WX11455 = ((~II35288))|((~II35289));
assign WX10466 = (WX10464)|(WX10463);
assign WX8084 = (WX8082)|(WX8081);
assign II14787 = ((~II14777))|((~II14785));
assign II14172 = ((~II14174))|((~II14175));
assign WX1995 = (WX1747&RESET);
assign WX1837 = (WX1840&RESET);
assign WX1919 = ((~WX2158));
assign WX3621 = (WX3620&WX3591);
assign WX3010 = (WX3008)|(WX3007);
assign WX5311 = ((~WX6176));
assign WX2673 = ((~WX3590));
assign WX5032 = ((~II15341))|((~II15342));
assign WX6585 = (WX6591&WX6586);
assign II14622 = ((~II14624))|((~II14625));
assign WX1013 = ((~II3066))|((~II3067));
assign II18588 = ((~II18564))|((~II18580));
assign WX6529 = (WX6535&WX6530);
assign WX10672 = ((~WX10671));
assign WX4423 = (WX4426&RESET);
assign WX1716 = ((~WX2297));
assign WX3136 = ((~WX3555));
assign WX1789 = (WX1792&RESET);
assign II6962 = ((~WX2064))|((~II6961));
assign WX8778 = ((~II27109))|((~II27110));
assign WX10281 = ((~RESET));
assign WX4283 = (WX6366&WX4284);
assign WX134 = (WX140&WX135);
assign II26321 = ((~II26311))|((~II26319));
assign WX10667 = (WX10869&WX11348);
assign WX2720 = (WX2726&WX2721);
assign II35092 = ((~WX10924))|((~WX10829));
assign II3592 = ((~WX622))|((~II3591));
assign II10758 = ((~WX3407))|((~II10757));
assign II27420 = ((~WX8364))|((~WX8295));
assign WX1701 = (WX2487&WX1702);
assign WX3920 = ((~WX4883));
assign WX2812 = (WX3689&WX2813);
assign WX1623 = (WX1629&WX1624);
assign WX6679 = (WX6677)|(WX6676);
assign WX10203 = ((~WX10202));
assign II2483 = ((~II2485))|((~II2486));
assign WX6637 = (WX6635)|(WX6634);
assign II30395 = ((~WX10052))|((~WX9720));
assign WX5741 = ((~WX6115));
assign WX4507 = ((~WX4748));
assign II14436 = ((~II14438))|((~II14439));
assign II2203 = ((~II2213))|((~II2214));
assign II2111 = ((~II2113))|((~II2114));
assign WX7796 = (WX7794)|(WX7793);
assign WX1993 = (WX1733&RESET);
assign WX2384 = (WX2383&WX2298);
assign II15691 = ((~WX4515))|((~II15690));
assign WX354 = (WX352)|(WX351);
assign II10741 = ((~II10743))|((~II10744));
assign WX2776 = (WX2782&WX2777);
assign WX11444 = ((~WX11349));
assign II26267 = ((~WX8759))|((~II26266));
assign WX10154 = ((~WX10153));
assign WX9177 = (WX9175)|(WX9174);
assign WX10009 = ((~WX9980));
assign WX6468 = (WX6403&WX6435);
assign II14872 = ((~WX4881))|((~II14871));
assign WX9543 = (WX9546&RESET);
assign II23497 = ((~_2268_))|((~II23495));
assign II3338 = ((~WX602))|((~WX529));
assign WX8870 = (WX8869&WX8763);
assign WX9472 = (WX9590&WX10055);
assign II2514 = ((~II2516))|((~II2517));
assign WX8958 = ((~WX8957));
assign II22229 = ((~II22231))|((~II22232));
assign WX8949 = ((~WX8763));
assign WX11170 = (WX11107&RESET);
assign WX8712 = ((~WX8685));
assign II34089 = ((~II34091))|((~II34092));
assign II23589 = ((~WX7083))|((~II23588));
assign II35158 = ((~WX10929))|((~II35157));
assign II26197 = ((~II26187))|((~II26195));
assign II26295 = ((~II26305))|((~II26306));
assign II31635 = ((~_2320_))|((~II31633));
assign WX9199 = (WX9205&WX9200);
assign WX2849 = (_2156_&WX3590);
assign WX221 = (_2095_&WX1004);
assign WX9194 = ((~WX10055));
assign II34525 = ((~WX11346))|((~II34524));
assign WX8815 = (WX8345&WX8816);
assign WX361 = (_2085_&WX1004);
assign WX11522 = (WX11520)|(WX11519);
assign WX3878 = (WX3837&WX3849);
assign WX834 = (WX771&RESET);
assign II22990 = ((~WX7300))|((~II22989));
assign WX6185 = ((~II19086))|((~II19087));
assign WX4514 = ((~WX4762));
assign WX9971 = ((~II30666))|((~II30667));
assign II30077 = ((~II30052))|((~II30076));
assign WX8178 = (WX8176)|(WX8175);
assign II15599 = ((~WX4500))|((~_2194_));
assign WX11088 = (WX11025&RESET);
assign II7540 = ((~WX1907))|((~_2137_));
assign WX1758 = ((~WX2297));
assign WX11519 = (WX11518&WX11349);
assign WX11148 = (WX11085&RESET);
assign WX1744 = ((~WX2297));
assign II7330 = ((~WX1894))|((~WX1820));
assign II26058 = ((~II26048))|((~II26056));
assign WX8378 = ((~WX8611));
assign WX1771 = (WX2522&WX1772);
assign WX9403 = (WX10217&WX9404);
assign WX53 = (_2107_&WX1004);
assign WX10357 = (WX10296&WX10314);
assign II2384 = ((~II2374))|((~II2382));
assign II11644 = ((~WX3215))|((~II11643));
assign WX10656 = (WX10654)|(WX10653);
assign II35694 = ((~WX10977))|((~_2342_));
assign II2600 = ((~II2575))|((~II2599));
assign WX9475 = (WX9473)|(WX9472);
assign WX1370 = (WX1381&WX2296);
assign WX8680 = ((~II26723))|((~II26724));
assign WX7233 = (WX7170&RESET);
assign II2854 = ((~II2864))|((~II2865));
assign WX7078 = ((~WX7304));
assign II14831 = ((~II14807))|((~II14823));
assign II14368 = ((~II14358))|((~II14366));
assign II30869 = ((~II30859))|((~II30867));
assign WX9223 = (WX9221)|(WX9220);
assign II11258 = ((~WX3181))|((~II11257));
assign WX5555 = ((~WX5546));
assign WX7037 = ((~WX7414));
assign II6899 = ((~WX2060))|((~II6891));
assign WX1645 = (WX2459&WX1646);
assign WX7537 = ((~WX7470));
assign WX8706 = ((~WX8682));
assign II22378 = ((~II22368))|((~II22376));
assign WX8325 = ((~WX8697));
assign WX2143 = (WX2080&RESET);
assign WX3602 = ((~WX3591));
assign II18812 = ((~II18822))|((~II18823));
assign WX9292 = ((~WX10055));
assign WX7030 = ((~WX7400));
assign WX1225 = (WX611&WX1226);
assign II27608 = ((~WX8378))|((~II27607));
assign WX1571 = (WX3717&WX1572);
assign WX5653 = ((~WX5644));
assign WX4472 = ((~WX4440));
assign II3234 = ((~WX594))|((~WX513));
assign WX2864 = (WX5010&WX2865);
assign II10806 = ((~WX3283))|((~II10804));
assign WX10199 = (WX9651&WX10200);
assign WX1582 = ((~WX2296));
assign WX8920 = (WX8360&WX8921);
assign WX2726 = (WX2724)|(WX2723);
assign WX8760 = ((~WX8756));
assign WX5792 = ((~WX6025));
assign II30502 = ((~II30504))|((~II30505));
assign II18521 = ((~WX6041))|((~II18519));
assign II14554 = ((~II14544))|((~II14552));
assign WX11527 = (WX10949&WX11528);
assign WX6236 = (WX5760&WX6237);
assign II30201 = ((~II30176))|((~II30200));
assign WX8132 = (WX8130)|(WX8129);
assign II27225 = ((~WX8349))|((~WX8265));
assign WX5410 = (WX5408)|(WX5407);
assign WX2791 = ((~WX3589));
assign II6506 = ((~WX2162))|((~II6504));
assign II27670 = ((~WX8388))|((~_2281_));
assign WX9466 = ((~WX10054));
assign WX6758 = ((~WX7469));
assign WX4903 = (WX4901)|(WX4900);
assign II22183 = ((~WX7248))|((~WX7312));
assign II10966 = ((~WX3357))|((~II10958));
assign WX4763 = (WX4700&RESET);
assign II35626 = ((~_2354_))|((~II35624));
assign WX1055 = ((~II3144))|((~II3145));
assign WX3234 = (WX2662&RESET);
assign II23595 = ((~WX7084))|((~_2260_));
assign II30743 = ((~WX9806))|((~II30735));
assign WX7843 = (WX8249&WX8762);
assign WX6889 = (WX6887)|(WX6886);
assign II10976 = ((~WX3485))|((~II10974));
assign WX9193 = (WX10112&WX9194);
assign WX6681 = ((~WX6680));
assign II2059 = ((~II2049))|((~II2057));
assign II6497 = ((~WX2034))|((~II6496));
assign WX8717 = ((~WX8716));
assign WX4510 = ((~WX4754));
assign WX6983 = (WX6986&RESET);
assign WX3595 = ((~WX3591));
assign WX1648 = ((~WX1639));
assign WX9186 = ((~WX10054));
assign II30874 = ((~II30876))|((~II30877));
assign II22309 = ((~WX7320))|((~II22307));
assign II23324 = ((~WX7064))|((~WX6988));
assign WX3007 = (WX3125&WX3590);
assign II10410 = ((~II10400))|((~II10408));
assign II2065 = ((~WX777))|((~WX841));
assign WX1077 = (WX1076&WX1005);
assign WX10451 = ((~WX11347));
assign WX8616 = (WX8553&RESET);
assign II26584 = ((~WX8503))|((~II26583));
assign II14397 = ((~II14373))|((~II14389));
assign WX2464 = (WX2462)|(WX2461);
assign WX2877 = (_2154_&WX3590);
assign WX422 = (DATA_9_4&WX423);
assign WX280 = (WX278)|(WX277);
assign WX9959 = ((~II30294))|((~II30295));
assign WX5244 = (WX6198&WX5245);
assign WX66 = (WX64)|(WX63);
assign II18187 = ((~II18177))|((~II18185));
assign II14800 = ((~II14776))|((~II14792));
assign WX8484 = (WX8421&RESET);
assign II26452 = ((~WX8759))|((~WX8431));
assign II14639 = ((~WX4692))|((~II14638));
assign WX7816 = (WX8777&WX7817);
assign II18130 = ((~II18140))|((~II18141));
assign WX7405 = ((~WX7385));
assign II18977 = ((~WX5943))|((~II18976));
assign II10920 = ((~II10895))|((~II10919));
assign WX4258 = (WX4412&WX4883);
assign WX2327 = ((~II7110))|((~II7111));
assign WX6368 = (WX6367&WX6177);
assign II10975 = ((~WX3421))|((~II10974));
assign II34732 = ((~II34708))|((~II34724));
assign II7689 = ((~_2114_))|((~II7687));
assign II22122 = ((~WX7244))|((~II22121));
assign II19255 = ((~WX5766))|((~II19254));
assign II18397 = ((~WX6033))|((~II18395));
assign II10030 = ((~WX3587))|((~II10029));
assign WX7530 = ((~WX7470));
assign WX6337 = ((~WX6336));
assign II22989 = ((~WX7300))|((~WX7364));
assign II30798 = ((~WX10053))|((~WX9746));
assign WX8656 = (WX8593&RESET);
assign WX2544 = ((~II7639))|((~II7640));
assign WX11353 = ((~WX11349));
assign II23525 = ((~WX7104))|((~_2268_));
assign WX2398 = (WX2397&WX2298);
assign DATA_9_26 = ((~WX1046));
assign WX2349 = (WX2348&WX2298);
assign WX2473 = ((~WX2472));
assign II14002 = ((~II14004))|((~II14005));
assign WX10622 = (DATA_0_14&WX10623);
assign II6116 = ((~II6118))|((~II6119));
assign II30070 = ((~WX9826))|((~II30069));
assign WX3696 = ((~WX3695));
assign II34662 = ((~II34664))|((~II34665));
assign II6374 = ((~II6364))|((~II6372));
assign WX8239 = ((~WX8230));
assign WX5043 = (WX5041)|(WX5040);
assign WX7865 = ((~WX8761));
assign WX1487 = (WX3675&WX1488);
assign II22817 = ((~II22827))|((~II22828));
assign WX8066 = (WX8064)|(WX8063);
assign WX7011 = (WX6948&RESET);
assign WX2621 = (WX2632&WX3589);
assign WX1167 = ((~II3352))|((~II3353));
assign WX136 = (WX134)|(WX133);
assign WX3634 = ((~II11141))|((~II11142));
assign WX1906 = ((~WX2132));
assign WX2743 = ((~WX3590));
assign II27331 = ((~WX8281))|((~II27329));
assign II2586 = ((~II2576))|((~II2584));
assign WX4484 = ((~WX4452));
assign WX6674 = ((~WX7469));
assign WX10220 = (WX9654&WX10221);
assign WX8753 = ((~WX8752));
assign II6232 = ((~II6208))|((~II6224));
assign WX3408 = (WX3345&RESET);
assign WX2780 = (WX4968&WX2781);
assign II27461 = ((~WX8301))|((~II27459));
assign WX3191 = ((~WX3159));
assign WX5167 = (WX5132&WX5142);
assign WX9183 = ((~WX9182));
assign WX8354 = ((~WX8322));
assign WX6751 = ((~WX6750));
assign II3529 = ((~WX613))|((~II3528));
assign II31479 = ((~WX9596))|((~II31477));
assign WX11253 = ((~II34330))|((~II34331));
assign II30535 = ((~WX9856))|((~II30534));
assign WX8879 = ((~WX8763));
assign WX9630 = ((~WX10014));
assign WX5733 = ((~WX6163));
assign WX4097 = (WX4103&WX4098);
assign WX7889 = ((~WX7880));
assign II18055 = ((~WX5947))|((~II18054));
assign WX1650 = (WX1661&WX2296);
assign II11077 = ((~WX3073))|((~II11075));
assign WX242 = (WX240)|(WX239);
assign II22518 = ((~II22508))|((~II22516));
assign WX2393 = ((~WX2298));
assign II15354 = ((~WX4481))|((~II15353));
assign WX1202 = ((~II3417))|((~II3418));
assign II30905 = ((~II30907))|((~II30908));
assign WX11415 = (WX10933&WX11416);
assign II2439 = ((~WX865))|((~II2437));
assign WX1821 = (WX1824&RESET);
assign WX7702 = ((~II23561))|((~II23562));
assign WX184 = (DATA_9_21&WX185);
assign II26505 = ((~II26481))|((~II26497));
assign II18923 = ((~WX6003))|((~II18922));
assign II10462 = ((~II10464))|((~II10465));
assign II7356 = ((~WX1896))|((~WX1824));
assign WX2535 = ((~II7576))|((~II7577));
assign WX1188 = ((~II3391))|((~II3392));
assign WX323 = (WX525&WX1004);
assign WX3803 = (WX3802&WX3591);
assign II34835 = ((~WX11346))|((~II34834));
assign II6892 = ((~WX2295))|((~WX1996));
assign WX8144 = (WX8150&WX8145);
assign WX8242 = (WX8245&RESET);
assign II7371 = ((~WX1826))|((~II7369));
assign II35146 = ((~WX10837))|((~II35144));
assign WX5803 = ((~WX6047));
assign II23116 = ((~WX7048))|((~WX6956));
assign II2444 = ((~II2420))|((~II2436));
assign WX1393 = (WX2333&WX1394);
assign II10888 = ((~II10864))|((~II10880));
assign WX8393 = ((~WX8641));
assign WX8602 = (WX8539&RESET);
assign WX9243 = (WX9241)|(WX9240);
assign WX6846 = ((~WX7469));
assign WX2965 = (WX3119&WX3590);
assign WX4955 = ((~II15198))|((~II15199));
assign II14926 = ((~II14916))|((~II14924));
assign WX994 = ((~WX915));
assign II3379 = ((~WX535))|((~II3377));
assign WX8161 = (_2274_&WX8762);
assign WX9435 = ((~WX9434));
assign II30332 = ((~II30334))|((~II30335));
assign WX2768 = (WX2766)|(WX2765);
assign WX8496 = (WX8433&RESET);
assign WX1252 = ((~II3641))|((~II3642));
assign II18117 = ((~WX5951))|((~II18116));
assign II27486 = ((~WX8369))|((~II27485));
assign II2824 = ((~II2826))|((~II2827));
assign WX10134 = ((~II31231))|((~II31232));
assign WX38 = (WX36)|(WX35);
assign II6457 = ((~II6459))|((~II6460));
assign WX7753 = (WX7718&WX7728);
assign II18327 = ((~II18317))|((~II18325));
assign WX5533 = (_2213_&WX6176);
assign WX7850 = (WX7856&WX7851);
assign WX6912 = ((~WX7469));
assign WX2229 = ((~WX2211));
assign WX5882 = (WX5819&RESET);
assign WX6878 = (WX6889&WX7468);
assign II26926 = ((~II26916))|((~II26924));
assign WX10089 = (WX10087)|(WX10086);
assign WX9462 = ((~WX9453));
assign II22976 = ((~WX7172))|((~II22974));
assign WX2975 = (_2147_&WX3590);
assign WX6454 = (WX6427&WX6435);
assign WX5284 = (WX5282)|(WX5281);
assign II26575 = ((~II26577))|((~II26578));
assign II3558 = ((~_2102_))|((~II3556));
assign WX140 = (WX138)|(WX137);
assign WX5161 = (WX5134&WX5142);
assign II18371 = ((~II18347))|((~II18363));
assign II18193 = ((~II18195))|((~II18196));
assign WX236 = (WX2403&WX237);
assign II30738 = ((~WX9742))|((~II30736));
assign II2889 = ((~WX703))|((~II2887));
assign II26298 = ((~WX8759))|((~II26297));
assign WX4120 = ((~WX4883));
assign WX5753 = ((~WX5721));
assign II19229 = ((~WX5764))|((~II19228));
assign WX346 = (WX344)|(WX343);
assign II35274 = ((~WX10938))|((~WX10857));
assign II31558 = ((~_2331_))|((~II31556));
assign WX131 = ((~WX122));
assign II30962 = ((~II30952))|((~II30960));
assign II26398 = ((~WX8491))|((~II26397));
assign II14645 = ((~II14621))|((~II14637));
assign WX4649 = (WX4586&RESET);
assign II7640 = ((~_2122_))|((~II7638));
assign WX4809 = ((~II14956))|((~II14957));
assign II3248 = ((~WX595))|((~II3247));
assign WX10161 = ((~WX10160));
assign WX6157 = ((~WX6156));
assign WX5275 = ((~WX5266));
assign WX3120 = (WX3123&RESET);
assign WX6444 = (WX6405&WX6435);
assign II35675 = ((~_2346_))|((~II35673));
assign II35652 = ((~WX10969))|((~_2350_));
assign II19319 = ((~WX5771))|((~WX5695));
assign II3261 = ((~WX596))|((~II3260));
assign WX5422 = (WX7582&WX5423);
assign II14780 = ((~WX4574))|((~II14778));
assign WX10255 = (WX9659&WX10256);
assign WX9992 = ((~WX9991));
assign WX5536 = (WX5534)|(WX5533);
assign II15445 = ((~WX4488))|((~II15444));
assign II22764 = ((~WX7222))|((~II22756));
assign WX10458 = (WX11391&WX10459);
assign II10371 = ((~WX3587))|((~II10370));
assign WX11299 = ((~WX11298));
assign II34726 = ((~WX11161))|((~II34725));
assign II30233 = ((~II30223))|((~II30231));
assign II14776 = ((~II14786))|((~II14787));
assign WX8168 = (WX8166)|(WX8165);
assign WX11428 = (WX11427&WX11349);
assign WX6777 = (WX6775)|(WX6774);
assign WX8672 = ((~II26475))|((~II26476));
assign II18332 = ((~II18334))|((~II18335));
assign WX7769 = (WX7711&WX7728);
assign II30115 = ((~II30117))|((~II30118));
assign WX9483 = (WX11552&WX9484);
assign WX8885 = (WX8355&WX8886);
assign II27473 = ((~WX8368))|((~II27472));
assign II18613 = ((~WX5983))|((~II18612));
assign II18227 = ((~WX5831))|((~II18225));
assign WX5824 = (WX5276&RESET);
assign II26872 = ((~WX8649))|((~II26870));
assign WX9080 = (WX8995&WX9021);
assign WX7075 = ((~WX7043));
assign WX1386 = ((~WX2296));
assign WX1230 = ((~RESET));
assign WX3752 = ((~WX3751));
assign WX447 = ((~WX1004));
assign WX10311 = ((~II31732))|((~II31733));
assign WX8112 = (WX8110)|(WX8109);
assign WX6429 = ((~II19696))|((~II19697));
assign II10697 = ((~WX3467))|((~II10695));
assign II7228 = ((~WX1804))|((~II7226));
assign WX1933 = ((~WX2186));
assign II11511 = ((~WX3225))|((~II11510));
assign II6708 = ((~WX1984))|((~II6706));
assign WX2550 = ((~II7681))|((~II7682));
assign WX4727 = (WX4664&RESET);
assign II19675 = ((~WX5805))|((~II19674));
assign II11602 = ((~WX3208))|((~II11601));
assign WX2445 = ((~WX2444));
assign WX11435 = (WX11434&WX11349);
assign WX5926 = (WX5863&RESET);
assign WX5251 = ((~WX6175));
assign II2530 = ((~WX807))|((~WX871));
assign WX2035 = (WX1972&RESET);
assign II26328 = ((~WX8759))|((~WX8423));
assign II6938 = ((~WX2126))|((~WX2190));
assign WX1242 = ((~II3571))|((~II3572));
assign II6806 = ((~WX2054))|((~II6798));
assign WX10315 = (WX10285&WX10314);
assign WX5290 = ((~WX5289));
assign II22740 = ((~II22742))|((~II22743));
assign II10851 = ((~WX3413))|((~II10850));
assign WX10411 = (_2362_&WX11348);
assign II27200 = ((~WX8347))|((~II27199));
assign II14563 = ((~WX4560))|((~II14561));
assign II34492 = ((~II34494))|((~II34495));
assign II3221 = ((~WX593))|((~WX511));
assign II23632 = ((~_2255_))|((~II23630));
assign II22511 = ((~WX7142))|((~II22509));
assign II30380 = ((~WX9846))|((~II30379));
assign WX6214 = (WX6213&WX6177);
assign II30180 = ((~WX9706))|((~II30178));
assign WX7141 = (WX6737&RESET);
assign II26282 = ((~WX8547))|((~II26281));
assign WX7369 = ((~II22160))|((~II22161));
assign II22263 = ((~WX7126))|((~II22261));
assign WX197 = (WX507&WX1004);
assign WX205 = ((~WX1003));
assign II30021 = ((~II30031))|((~II30032));
assign II14290 = ((~WX4606))|((~II14289));
assign II2746 = ((~II2748))|((~II2749));
assign II30951 = ((~II30961))|((~II30962));
assign WX1504 = (WX1802&WX2297);
assign WX2418 = ((~II7279))|((~II7280));
assign WX10229 = (WX10227)|(WX10226);
assign WX4801 = ((~II14708))|((~II14709));
assign WX5394 = (WX7568&WX5395);
assign WX5183 = (WX5125&WX5142);
assign WX842 = (WX779&RESET);
assign II10108 = ((~WX3429))|((~II10106));
assign WX7856 = (WX7854)|(WX7853);
assign WX4334 = (WX4345&WX4882);
assign II34336 = ((~II34346))|((~II34347));
assign WX9216 = (_2323_&WX10055);
assign WX9240 = (WX9251&WX10054);
assign WX3641 = ((~II11154))|((~II11155));
assign WX2437 = ((~WX2436));
assign WX9206 = (WX9552&WX10055);
assign II30311 = ((~II30301))|((~II30309));
assign WX7527 = ((~II23182))|((~II23183));
assign WX348 = (WX2459&WX349);
assign WX1352 = ((~WX2297));
assign WX4415 = (WX4418&RESET);
assign II18234 = ((~II18224))|((~II18232));
assign WX9363 = (WX9361)|(WX9360);
assign WX3727 = (WX3185&WX3728);
assign WX5289 = ((~WX5280));
assign WX4824 = ((~WX4823));
assign WX762 = (WX699&RESET);
assign WX8404 = (WX7820&RESET);
assign WX11240 = (WX11177&RESET);
assign WX1891 = ((~WX1859));
assign II27657 = ((~WX8386))|((~II27656));
assign WX9322 = ((~WX9313));
assign WX76 = ((~WX75));
assign WX3386 = (WX3323&RESET);
assign II6956 = ((~WX2000))|((~II6954));
assign II23519 = ((~II23509))|((~II23517));
assign WX1854 = ((~WX2284));
assign II23428 = ((~WX7072))|((~WX7004));
assign WX6219 = ((~WX6218));
assign WX272 = ((~WX271));
assign WX9108 = (WX9538&WX10055);
assign WX1049 = (WX1048&WX1005);
assign WX2342 = (WX2341&WX2298);
assign WX81 = (_2105_&WX1004);
assign II30550 = ((~WX10053))|((~WX9730));
assign WX5586 = (WX5592&WX5587);
assign WX11424 = (WX11422)|(WX11421);
assign II2916 = ((~II2926))|((~II2927));
assign II22206 = ((~WX7186))|((~II22198));
assign WX6440 = (WX6433&WX6435);
assign II22346 = ((~II22321))|((~II22345));
assign II10152 = ((~II10154))|((~II10155));
assign WX9332 = (WX9570&WX10055);
assign WX4671 = (WX4608&RESET);
assign WX1150 = (WX1148)|(WX1147);
assign WX9156 = (WX9167&WX10054);
assign WX11480 = (WX11478)|(WX11477);
assign WX9610 = ((~WX10038));
assign II27097 = ((~WX8245))|((~II27095));
assign II14064 = ((~II14066))|((~II14067));
assign WX8811 = ((~WX8810));
assign II10062 = ((~WX3235))|((~II10060));
assign WX5195 = (WX5119&WX5142);
assign WX289 = ((~WX1003));
assign WX7247 = (WX7184&RESET);
assign WX6347 = (WX6346&WX6177);
assign II10386 = ((~WX3383))|((~II10385));
assign WX7543 = (WX7055&WX7544);
assign WX371 = (WX382&WX1003);
assign II2398 = ((~WX735))|((~II2390));
assign WX2376 = ((~II7201))|((~II7202));
assign WX8212 = ((~WX8211));
assign WX2408 = (WX2406)|(WX2405);
assign WX11561 = (WX11560&WX11349);
assign WX10640 = (WX11482&WX10641);
assign WX10603 = (WX10614&WX11347);
assign II23480 = ((~WX7076))|((~WX7012));
assign II10671 = ((~II10647))|((~II10663));
assign WX7968 = (WX7966)|(WX7965);
assign WX5134 = ((~II15677))|((~II15678));
assign II11629 = ((~WX3212))|((~_2157_));
assign WX9264 = ((~WX10055));
assign WX2503 = (WX2502&WX2298);
assign WX1010 = (WX1008)|(WX1007);
assign WX8669 = ((~II26382))|((~II26383));
assign WX577 = ((~WX959));
assign II6752 = ((~WX2114))|((~WX2178));
assign WX10563 = ((~WX11347));
assign WX4460 = ((~WX4428));
assign WX5007 = ((~WX4884));
assign II35249 = ((~WX10936))|((~II35248));
assign WX3368 = (WX3305&RESET);
assign II15650 = ((~_2186_))|((~II15648));
assign WX1235 = ((~II3522))|((~II3523));
assign WX9137 = (WX10084&WX9138);
assign WX2748 = (WX2754&WX2749);
assign WX4192 = ((~WX4183));
assign WX1094 = (WX1092)|(WX1091);
assign II6854 = ((~II6844))|((~II6852));
assign WX5209 = ((~WX6175));
assign WX1929 = ((~WX2178));
assign WX3108 = (WX3111&RESET);
assign WX6969 = (WX6972&RESET);
assign WX10872 = (WX10875&RESET);
assign II2576 = ((~II2578))|((~II2579));
assign WX11491 = (WX11490&WX11349);
assign WX3161 = ((~WX3541));
assign WX3264 = (WX2872&RESET);
assign WX10806 = (WX10804)|(WX10803);
assign WX3581 = ((~WX3580));
assign II18846 = ((~WX6174))|((~II18845));
assign II22950 = ((~WX7234))|((~II22942));
assign WX1886 = ((~WX1854));
assign WX10754 = (WX10752)|(WX10751);
assign WX4794 = ((~II14491))|((~II14492));
assign II14384 = ((~II14374))|((~II14382));
assign II10432 = ((~WX3587))|((~WX3259));
assign II18673 = ((~II18675))|((~II18676));
assign WX9555 = (WX9558&RESET);
assign II35405 = ((~WX10948))|((~II35404));
assign II7409 = ((~WX1900))|((~II7408));
assign II27508 = ((~_2284_))|((~II27507));
assign II14663 = ((~II14653))|((~II14661));
assign WX3619 = ((~WX3618));
assign WX7913 = (WX8259&WX8762);
assign WX1752 = (_2110_&WX2297);
assign II14421 = ((~WX4678))|((~WX4742));
assign WX6450 = (WX6429&WX6435);
assign WX4469 = ((~WX4437));
assign WX8862 = ((~II27265))|((~II27266));
assign WX6146 = ((~WX6077));
assign WX1765 = (WX1763)|(WX1762);
assign II6420 = ((~II6410))|((~II6418));
assign WX7993 = (_2286_&WX8762);
assign II2591 = ((~II2593))|((~II2594));
assign WX9954 = ((~II30139))|((~II30140));
assign WX7071 = ((~WX7039));
assign WX4399 = (WX4402&RESET);
assign II27663 = ((~WX8387))|((~_2282_));
assign II6689 = ((~II6691))|((~II6692));
assign WX4687 = (WX4624&RESET);
assign II14042 = ((~WX4590))|((~II14041));
assign WX7396 = ((~II22997))|((~II22998));
assign WX2291 = ((~TM0));
assign II26102 = ((~II26078))|((~II26094));
assign II18960 = ((~II18936))|((~II18952));
assign II10618 = ((~WX3588))|((~WX3271));
assign WX5246 = (WX5244)|(WX5243);
assign WX2232 = ((~WX2231));
assign II2640 = ((~WX1002))|((~II2639));
assign WX9028 = (WX9018&WX9021);
assign II30349 = ((~WX9844))|((~II30348));
assign WX9989 = ((~WX9970));
assign WX4877 = ((~TM0));
assign WX4059 = (WX6254&WX4060);
assign WX5678 = (WX5681&RESET);
assign WX8562 = (WX8499&RESET);
assign WX9481 = (WX9479)|(WX9478);
assign WX5631 = (_2206_&WX6176);
assign WX7106 = ((~WX7360));
assign II14950 = ((~WX4776))|((~II14948));
assign WX11586 = ((~II35611))|((~II35612));
assign II23091 = ((~WX7046))|((~II23090));
assign II15301 = ((~WX4477))|((~WX4400));
assign WX1060 = ((~WX1059));
assign WX2131 = (WX2068&RESET);
assign WX3854 = (WX3847&WX3849);
assign II19436 = ((~WX5780))|((~WX5713));
assign II23639 = ((~_2254_))|((~II23637));
assign WX2853 = (WX3103&WX3590);
assign WX2738 = (WX4947&WX2739);
assign WX1212 = ((~WX1005));
assign WX4142 = (_2188_&WX4883);
assign II6054 = ((~II6056))|((~II6057));
assign WX8677 = ((~II26630))|((~II26631));
assign WX6765 = ((~WX6764));
assign WX4991 = (WX4990&WX4884);
assign WX4015 = (WX4013)|(WX4012);
assign WX7691 = ((~WX7470));
assign WX6267 = ((~WX6266));
assign II30254 = ((~II30256))|((~II30257));
assign WX5089 = (WX5088&WX4884);
assign II6403 = ((~WX2028))|((~II6395));
assign WX11184 = (WX11121&RESET);
assign WX7938 = (WX10133&WX7939);
assign WX9302 = ((~WX10055));
assign WX6103 = ((~II18992))|((~II18993));
assign WX10178 = (WX9648&WX10179);
assign WX3954 = ((~WX3945));
assign WX3023 = ((~WX3590));
assign WX963 = ((~WX962));
assign WX7923 = (_2291_&WX8762);
assign II34866 = ((~WX11346))|((~II34865));
assign II14847 = ((~WX4642))|((~II14839));
assign II6828 = ((~II6838))|((~II6839));
assign II2617 = ((~II2607))|((~II2615));
assign WX7698 = ((~II23533))|((~II23534));
assign II26608 = ((~WX8760))|((~II26607));
assign II34059 = ((~WX11345))|((~WX10991));
assign WX9178 = (WX9548&WX10055);
assign II22759 = ((~WX7158))|((~II22757));
assign WX1846 = ((~WX2268));
assign WX7608 = (WX7606)|(WX7605);
assign WX1198 = ((~WX1005));
assign II2052 = ((~WX649))|((~II2050));
assign WX6785 = (WX8910&WX6786);
assign II22609 = ((~WX7212))|((~II22601));
assign WX3936 = (WX4366&WX4883);
assign II18378 = ((~II18388))|((~II18389));
assign WX8660 = ((~II26103))|((~II26104));
assign WX1136 = (WX1134)|(WX1133);
assign WX1989 = (WX1705&RESET);
assign WX1300 = (WX1248&WX1263);
assign WX9571 = (WX9574&RESET);
assign WX8968 = (WX8967&WX8763);
assign WX11549 = ((~WX11349));
assign WX1877 = ((~WX1845));
assign WX10723 = (WX10877&WX11348);
assign II30791 = ((~II30781))|((~II30789));
assign II34212 = ((~II34222))|((~II34223));
assign WX7135 = (WX6695&RESET);
assign II7612 = ((~_2127_))|((~II7610));
assign WX6127 = ((~WX6126));
assign WX11622 = (WX11601&WX11607);
assign WX384 = ((~WX383));
assign II30194 = ((~WX9834))|((~II30193));
assign II34206 = ((~II34181))|((~II34205));
assign II26978 = ((~II26980))|((~II26981));
assign WX1797 = (WX1800&RESET);
assign WX10159 = (WX10157)|(WX10156);
assign WX3156 = ((~WX3531));
assign WX8010 = (WX8008)|(WX8007);
assign WX2886 = ((~WX2885));
assign II35289 = ((~WX10859))|((~II35287));
assign II30239 = ((~II30241))|((~II30242));
assign II26407 = ((~WX8619))|((~II26405));
assign II6141 = ((~II6131))|((~II6139));
assign WX9597 = (WX9534&RESET);
assign WX6230 = ((~WX6177));
assign WX8850 = (WX8350&WX8851);
assign II2880 = ((~II2870))|((~II2878));
assign WX2803 = (WX2814&WX3589);
assign WX6111 = ((~WX6110));
assign WX7456 = ((~WX7455));
assign II30087 = ((~WX9700))|((~II30085));
assign WX1669 = (WX3766&WX1670);
assign II30177 = ((~II30179))|((~II30180));
assign WX3028 = (WX3034&WX3029);
assign WX8060 = (WX8066&WX8061);
assign WX4315 = (WX5087&WX4316);
assign WX4926 = ((~WX4925));
assign II26598 = ((~II26574))|((~II26590));
assign II22898 = ((~WX7358))|((~II22896));
assign II15199 = ((~WX4384))|((~II15197));
assign WX10423 = ((~WX11347));
assign WX433 = ((~WX1004));
assign II34708 = ((~II34718))|((~II34719));
assign WX4345 = (WX4343)|(WX4342);
assign WX3145 = ((~WX3573));
assign WX5507 = ((~WX6176));
assign II22387 = ((~WX7134))|((~II22385));
assign WX5052 = ((~WX5051));
assign WX3833 = ((~II11616))|((~II11617));
assign WX293 = ((~WX1004));
assign WX116 = (WX114)|(WX113);
assign WX4363 = (WX4366&RESET);
assign WX3585 = ((~TM1));
assign WX6645 = (WX8840&WX6646);
assign WX10232 = ((~II31413))|((~II31414));
assign WX2785 = ((~WX3590));
assign WX8420 = (WX7932&RESET);
assign WX1945 = (WX1397&RESET);
assign WX7743 = (WX7722&WX7728);
assign WX11463 = (WX11462&WX11349);
assign WX263 = (_2092_&WX1004);
assign WX10649 = (_2345_&WX11348);
assign WX4619 = (WX4556&RESET);
assign II14089 = ((~II14079))|((~II14087));
assign II35184 = ((~WX10931))|((~II35183));
assign WX6524 = ((~WX7469));
assign II35680 = ((~WX10974))|((~_2345_));
assign WX9917 = (WX9854&RESET);
assign II35752 = ((~_2333_))|((~II35750));
assign II22136 = ((~II22138))|((~II22139));
assign WX9428 = ((~WX10055));
assign WX3342 = (WX3279&RESET);
assign II6312 = ((~II6302))|((~II6310));
assign WX2430 = ((~WX2429));
assign WX776 = (WX713&RESET);
assign II2088 = ((~WX715))|((~II2080));
assign WX6852 = ((~WX7468));
assign II23503 = ((~_2252_))|((~II23502));
assign WX467 = ((~WX458));
assign II14142 = ((~WX4660))|((~WX4724));
assign II7174 = ((~WX1882))|((~WX1796));
assign WX9256 = ((~WX10054));
assign WX5419 = ((~WX6175));
assign WX11275 = ((~II35012))|((~II35013));
assign WX4813 = ((~WX4796));
assign WX5489 = ((~WX6175));
assign II15507 = ((~_2183_))|((~II15499));
assign WX9016 = ((~II27713))|((~II27714));
assign WX11062 = (WX10999&RESET);
assign II22090 = ((~WX7242))|((~WX7306));
assign WX4669 = (WX4606&RESET);
assign WX1787 = (WX1790&RESET);
assign II11233 = ((~WX3097))|((~II11231));
assign II14514 = ((~WX4684))|((~WX4748));
assign WX4209 = (WX4215&WX4210);
assign WX6688 = ((~WX7469));
assign WX3298 = (WX3235&RESET);
assign WX9062 = (WX9004&WX9021);
assign WX3039 = ((~WX3030));
assign WX7333 = (WX7270&RESET);
assign II18490 = ((~WX6039))|((~II18488));
assign II7482 = ((~_2124_))|((~II7474));
assign WX4857 = ((~WX4786));
assign II34874 = ((~II34864))|((~II34872));
assign II30518 = ((~II30520))|((~II30521));
assign II10277 = ((~WX3587))|((~WX3249));
assign WX10965 = ((~WX11199));
assign WX980 = ((~WX908));
assign WX9239 = ((~WX9238));
assign WX5763 = ((~WX5731));
assign WX7773 = (WX7709&WX7728);
assign II18945 = ((~WX5941))|((~II18937));
assign WX10596 = (WX10594)|(WX10593);
assign WX4202 = (WX4404&WX4883);
assign WX8202 = (WX8200)|(WX8199);
assign WX6022 = (WX5959&RESET);
assign II2415 = ((~II2405))|((~II2413));
assign WX1762 = (WX1773&WX2296);
assign WX3522 = ((~WX3504));
assign WX9357 = (WX11489&WX9358);
assign WX7727 = ((~II23736))|((~II23737));
assign WX6939 = (WX8987&WX6940);
assign WX5123 = ((~II15600))|((~II15601));
assign WX4084 = ((~WX4882));
assign WX598 = ((~WX566));
assign WX6549 = (WX6547)|(WX6546);
assign WX2947 = (_2149_&WX3590);
assign WX3732 = ((~II11323))|((~II11324));
assign WX4029 = (WX4027)|(WX4026);
assign WX3494 = ((~II10269))|((~II10270));
assign II10325 = ((~WX3443))|((~II10323));
assign II2785 = ((~II2761))|((~II2777));
assign II34402 = ((~WX11013))|((~II34400));
assign II26684 = ((~WX8573))|((~WX8637));
assign II7491 = ((~WX1925))|((~II7490));
assign WX2484 = ((~WX2298));
assign WX9235 = (WX10133&WX9236);
assign WX8032 = (WX8038&WX8033);
assign II7149 = ((~WX1880))|((~II7148));
assign WX1067 = ((~WX1066));
assign II14011 = ((~WX4588))|((~II14010));
assign WX3098 = (WX3101&RESET);
assign II35107 = ((~WX10831))|((~II35105));
assign WX11246 = ((~II34113))|((~II34114));
assign WX4149 = (WX4147)|(WX4146);
assign WX5517 = ((~WX6175));
assign WX5902 = (WX5839&RESET);
assign WX5109 = ((~RESET));
assign II22959 = ((~WX7298))|((~II22958));
assign II26996 = ((~WX8657))|((~II26994));
assign WX5462 = (WX5460)|(WX5459);
assign II23693 = ((~WX7100))|((~_2244_));
assign II23540 = ((~WX7108))|((~II23539));
assign II6428 = ((~WX2294))|((~II6427));
assign WX10708 = (WX10706)|(WX10705);
assign WX2932 = (WX2930)|(WX2929);
assign II34577 = ((~II34553))|((~II34569));
assign WX2821 = (_2158_&WX3590);
assign II14018 = ((~WX4652))|((~WX4716));
assign WX5333 = (WX5344&WX6175);
assign WX2629 = (WX3071&WX3590);
assign WX5265 = ((~WX6175));
assign WX10074 = ((~WX10056));
assign II30993 = ((~II30983))|((~II30991));
assign II10899 = ((~WX3289))|((~II10897));
assign WX10127 = ((~II31218))|((~II31219));
assign WX6827 = (WX8931&WX6828);
assign WX2659 = ((~WX3590));
assign WX11302 = ((~WX11273));
assign II18683 = ((~II18673))|((~II18681));
assign WX9667 = ((~WX9896));
assign II30906 = ((~WX9880))|((~WX9944));
assign WX7709 = ((~II23610))|((~II23611));
assign WX5638 = (WX5636)|(WX5635);
assign WX4695 = (WX4632&RESET);
assign WX257 = ((~WX248));
assign II7161 = ((~WX1881))|((~WX1794));
assign II3661 = ((~WX634))|((~_2085_));
assign II34688 = ((~II34678))|((~II34686));
assign WX718 = (WX655&RESET);
assign WX10298 = ((~II31641))|((~II31642));
assign WX9967 = ((~II30542))|((~II30543));
assign II14544 = ((~II14546))|((~II14547));
assign II34973 = ((~WX11177))|((~WX11241));
assign II30417 = ((~II30393))|((~II30409));
assign WX8073 = (WX8084&WX8761);
assign WX5300 = (WX6226&WX5301);
assign WX10469 = ((~WX11348));
assign WX6202 = ((~WX6177));
assign II30099 = ((~II30101))|((~II30102));
assign WX4845 = ((~WX4780));
assign WX3529 = ((~WX3528));
assign II30272 = ((~WX10052))|((~II30271));
assign WX5635 = (WX5717&WX6176);
assign WX6226 = ((~WX6225));
assign II11218 = ((~WX3178))|((~WX3095));
assign WX8108 = (WX8106)|(WX8105);
assign WX7103 = ((~WX7354));
assign WX6893 = (WX6899&WX6894);
assign WX5093 = ((~WX5092));
assign WX4294 = ((~WX4882));
assign WX10321 = (WX10311&WX10314);
assign WX1896 = ((~WX1864));
assign WX1415 = (WX1413)|(WX1412);
assign II14740 = ((~II14730))|((~II14738));
assign WX5502 = (WX5508&WX5503);
assign WX7437 = ((~WX7369));
assign WX8844 = ((~WX8763));
assign II2313 = ((~WX793))|((~WX857));
assign WX5327 = (WX5673&WX6176);
assign WX4050 = ((~WX4883));
assign II2268 = ((~WX1001))|((~II2267));
assign WX584 = ((~WX552));
assign II23660 = ((~_2250_))|((~II23658));
assign II7382 = ((~WX1898))|((~WX1828));
assign WX5952 = (WX5889&RESET);
assign WX8191 = ((~WX8762));
assign WX5210 = (WX5208)|(WX5207);
assign WX5512 = (WX5510)|(WX5509);
assign WX2335 = (WX2334&WX2298);
assign II31513 = ((~_2316_))|((~II31512));
assign WX6244 = ((~WX6177));
assign WX1692 = (WX1703&WX2296);
assign WX8058 = ((~WX8057));
assign II26838 = ((~II26840))|((~II26841));
assign II22624 = ((~II22600))|((~II22616));
assign WX7961 = (WX7972&WX8761);
assign WX2216 = ((~II6729))|((~II6730));
assign II3712 = ((~_2077_))|((~II3710));
assign WX3679 = ((~WX3591));
assign II31219 = ((~WX9556))|((~II31217));
assign II10463 = ((~WX3587))|((~WX3261));
assign II35196 = ((~WX10932))|((~WX10845));
assign WX2222 = ((~II6915))|((~II6916));
assign WX2665 = ((~WX3589));
assign II35353 = ((~WX10944))|((~II35352));
assign WX6624 = ((~WX6615));
assign II22215 = ((~WX7250))|((~II22214));
assign WX6941 = (WX6939)|(WX6938);
assign WX6542 = (WX6553&WX7468);
assign WX6538 = ((~WX7469));
assign WX9635 = ((~WX9603));
assign WX11204 = (WX11141&RESET);
assign WX3784 = ((~WX3591));
assign WX2831 = (WX2842&WX3589);
assign II27110 = ((~WX8247))|((~II27108));
assign WX2159 = (WX2096&RESET);
assign WX2411 = ((~II7266))|((~II7267));
assign WX6736 = ((~WX6727));
assign II2547 = ((~WX1002))|((~II2546));
assign WX8096 = (WX8917&WX8097);
assign WX4308 = ((~WX4882));
assign WX11449 = (WX11448&WX11349);
assign WX2401 = (WX2399)|(WX2398);
assign WX3764 = (WX3762)|(WX3761);
assign WX8418 = (WX7918&RESET);
assign WX5593 = (WX5711&WX6176);
assign WX6616 = (_2260_&WX7469);
assign II34026 = ((~II34036))|((~II34037));
assign II14049 = ((~WX4654))|((~WX4718));
assign WX1320 = (WX1238&WX1263);
assign WX10031 = ((~WX9959));
assign WX3322 = (WX3259&RESET);
assign II35611 = ((~WX10963))|((~II35610));
assign WX8351 = ((~WX8319));
assign II30937 = ((~WX9882))|((~WX9946));
assign WX10958 = ((~WX11185));
assign WX1424 = ((~WX1415));
assign II30519 = ((~WX10053))|((~WX9728));
assign II2610 = ((~WX685))|((~II2608));
assign WX10785 = (WX10796&WX11347);
assign WX6975 = (WX6978&RESET);
assign WX6822 = (WX6833&WX7468);
assign WX2275 = ((~WX2202));
assign II26460 = ((~WX8495))|((~II26459));
assign WX6948 = ((~WX6950));
assign WX2973 = ((~WX3589));
assign WX4539 = (WX4039&RESET);
assign WX1348 = ((~WX2297));
assign WX6174 = ((~WX6170));
assign WX3580 = ((~WX3501));
assign WX7428 = ((~WX7427));
assign WX8900 = ((~WX8763));
assign II10286 = ((~II10276))|((~II10284));
assign WX10398 = (DATA_0_30&WX10399);
assign WX6539 = (WX6537)|(WX6536);
assign II18969 = ((~WX6174))|((~WX5879));
assign II18163 = ((~WX6173))|((~WX5827));
assign WX5578 = (WX5576)|(WX5575);
assign II18737 = ((~WX5991))|((~II18736));
assign II7507 = ((~_2140_))|((~II7505));
assign WX2894 = (WX2892)|(WX2891);
assign WX11375 = (WX11373)|(WX11372);
assign WX10504 = ((~WX10503));
assign WX6521 = (WX6519)|(WX6518);
assign II6552 = ((~WX2295))|((~II6551));
assign WX11399 = ((~II35184))|((~II35185));
assign WX5239 = (_2234_&WX6176);
assign II18558 = ((~II18533))|((~II18557));
assign II11509 = ((~II11511))|((~II11512));
assign WX4890 = ((~WX4889));
assign WX4867 = ((~WX4791));
assign WX658 = (WX146&RESET);
assign II34763 = ((~II34739))|((~II34755));
assign II15328 = ((~WX4479))|((~II15327));
assign WX10856 = (WX10859&RESET);
assign WX6280 = (WX6278)|(WX6277);
assign II26777 = ((~WX8579))|((~WX8643));
assign WX3316 = (WX3253&RESET);
assign II26817 = ((~II26807))|((~II26815));
assign II34941 = ((~II34943))|((~II34944));
assign II2073 = ((~II2048))|((~II2072));
assign II6605 = ((~II6580))|((~II6604));
assign II35556 = ((~_2364_))|((~II35554));
assign II30459 = ((~WX9724))|((~II30457));
assign II34433 = ((~WX11015))|((~II34431));
assign WX8151 = (WX8293&WX8762);
assign WX3866 = (WX3842&WX3849);
assign WX1427 = (WX1433&WX1428);
assign WX3623 = ((~WX3591));
assign WX1519 = (WX2396&WX1520);
assign DATA_9_14 = ((~WX1130));
assign WX1509 = ((~WX1508));
assign II14151 = ((~II14141))|((~II14149));
assign WX9122 = (WX9540&WX10055);
assign WX473 = (_2077_&WX1004);
assign WX9532 = ((~WX9523));
assign WX8941 = (WX8363&WX8942);
assign II14127 = ((~WX4880))|((~WX4532));
assign WX4886 = (WX4885&WX4884);
assign WX1016 = ((~WX1005));
assign WX6270 = (WX6269&WX6177);
assign WX6735 = (WX6733)|(WX6732);
assign WX4697 = (WX4634&RESET);
assign WX4267 = (WX4265)|(WX4264);
assign WX5545 = ((~WX6175));
assign II14337 = ((~II14327))|((~II14335));
assign WX9032 = (WX9017&WX9021);
assign WX4180 = (WX4191&WX4882);
assign II2507 = ((~II2482))|((~II2506));
assign WX10073 = (WX9633&WX10074);
assign WX8298 = (WX8301&RESET);
assign WX2642 = (WX2640)|(WX2639);
assign II22728 = ((~WX7156))|((~II22726));
assign WX7163 = (WX6891&RESET);
assign II14685 = ((~WX4881))|((~WX4568));
assign WX587 = ((~WX555));
assign WX10244 = ((~WX10243));
assign WX3458 = (WX3395&RESET);
assign WX4281 = (WX4279)|(WX4278);
assign II3668 = ((~WX635))|((~_2084_));
assign WX4915 = (WX4463&WX4916);
assign WX5868 = (WX5584&RESET);
assign WX3550 = ((~WX3486));
assign WX3654 = ((~WX3653));
assign II31669 = ((~WX9680))|((~II31668));
assign II34407 = ((~WX11077))|((~II34399));
assign II7096 = ((~WX1876))|((~WX1784));
assign WX10730 = (WX10736&WX10731);
assign WX5575 = (_2210_&WX6176);
assign WX4250 = (WX4261&WX4882);
assign WX10974 = ((~WX11217));
assign II22449 = ((~WX7138))|((~II22447));
assign WX574 = ((~WX953));
assign II23553 = ((~WX7078))|((~_2266_));
assign II30652 = ((~II30642))|((~II30650));
assign II6807 = ((~WX2054))|((~II6806));
assign II35209 = ((~WX10933))|((~WX10847));
assign II22718 = ((~II22693))|((~II22717));
assign WX10475 = ((~WX10466));
assign WX2638 = (WX2636)|(WX2635);
assign WX4425 = (WX4362&RESET);
assign WX8398 = ((~WX8651));
assign WX1889 = ((~WX1857));
assign WX8276 = (WX8279&RESET);
assign II14253 = ((~WX4540))|((~II14251));
assign II34099 = ((~II34089))|((~II34097));
assign II23652 = ((~WX7093))|((~II23651));
assign WX1686 = (WX1828&WX2297);
assign WX8622 = (WX8559&RESET);
assign WX3012 = ((~WX3011));
assign WX5640 = ((~WX5639));
assign II34755 = ((~II34757))|((~II34758));
assign WX39 = (_2108_&WX1004);
assign WX6336 = (WX6334)|(WX6333);
assign WX3628 = (WX3627&WX3591);
assign II30868 = ((~WX9814))|((~II30867));
assign WX4786 = ((~II14243))|((~II14244));
assign WX10737 = (WX10879&WX11348);
assign II18179 = ((~WX5955))|((~II18178));
assign WX6573 = (WX6571)|(WX6570);
assign WX8654 = (WX8591&RESET);
assign WX6513 = ((~WX6512));
assign WX5401 = ((~WX5392));
assign WX8759 = ((~WX8758));
assign WX8869 = ((~II27278))|((~II27279));
assign WX1440 = (WX1451&WX2296);
assign WX10901 = ((~WX11327));
assign WX10489 = ((~WX10480));
assign II14668 = ((~II14670))|((~II14671));
assign II14190 = ((~WX4880))|((~II14189));
assign WX8082 = (WX8910&WX8083);
assign II22028 = ((~WX7238))|((~WX7302));
assign II2500 = ((~WX805))|((~II2499));
assign WX11470 = (WX11469&WX11349);
assign WX5842 = (WX5402&RESET);
assign II27330 = ((~WX8357))|((~II27329));
assign WX10496 = (DATA_0_23&WX10497);
assign WX6256 = (WX6255&WX6177);
assign WX4068 = (WX4079&WX4882);
assign II26770 = ((~WX8515))|((~II26769));
assign WX2832 = (WX2838&WX2833);
assign II14105 = ((~II14095))|((~II14103));
assign WX2321 = (WX2320&WX2298);
assign II2934 = ((~WX833))|((~II2933));
assign WX6614 = ((~WX7468));
assign II22500 = ((~II22476))|((~II22492));
assign II27656 = ((~WX8386))|((~_2283_));
assign WX6258 = ((~WX6177));
assign WX8332 = ((~WX8711));
assign WX5498 = (WX5496)|(WX5495);
assign II18451 = ((~II18441))|((~II18449));
assign WX8085 = ((~WX8076));
assign WX6870 = ((~WX7469));
assign II23429 = ((~WX7072))|((~II23428));
assign WX8044 = ((~WX8043));
assign WX10720 = (DATA_0_7&WX10721);
assign WX7806 = ((~WX7805));
assign WX11202 = (WX11139&RESET);
assign WX6199 = ((~II19112))|((~II19113));
assign WX7974 = ((~WX7973));
assign WX6821 = ((~WX6820));
assign II6606 = ((~II6596))|((~II6604));
assign WX6148 = ((~WX6078));
assign II26066 = ((~WX8597))|((~II26064));
assign WX10578 = (WX10576)|(WX10575);
assign WX9110 = ((~WX10055));
assign II35743 = ((~WX10985))|((~_2334_));
assign WX6750 = ((~WX6741));
assign WX498 = (WX501&RESET);
assign WX11422 = (WX10934&WX11423);
assign WX6853 = (WX6851)|(WX6850);
assign WX1997 = (WX1761&RESET);
assign II23259 = ((~WX7059))|((~WX6978));
assign II15641 = ((~WX4507))|((~_2187_));
assign WX7485 = ((~II23104))|((~II23105));
assign WX6002 = (WX5939&RESET);
assign II14242 = ((~II14218))|((~II14234));
assign WX10534 = (WX10540&WX10535);
assign WX4124 = (WX4135&WX4882);
assign II11232 = ((~WX3179))|((~II11231));
assign II26381 = ((~II26357))|((~II26373));
assign WX6923 = (WX6921)|(WX6920);
assign WX4565 = (WX4221&RESET);
assign II23504 = ((~II23494))|((~II23502));
assign II14367 = ((~II14342))|((~II14366));
assign WX9319 = (WX10175&WX9320);
assign WX8022 = (WX10175&WX8023);
assign WX10040 = ((~WX10039));
assign WX255 = ((~WX1004));
assign II2847 = ((~II2823))|((~II2839));
assign WX10007 = ((~WX9979));
assign WX5039 = ((~II15354))|((~II15355));
assign WX309 = (WX523&WX1004);
assign II7673 = ((~WX1928))|((~_2116_));
assign WX7558 = ((~WX7470));
assign II26497 = ((~II26499))|((~II26500));
assign WX5742 = ((~WX6117));
assign WX2448 = (WX1894&WX2449);
assign WX154 = (WX152)|(WX151);
assign WX6920 = (WX6931&WX7468);
assign II27149 = ((~WX8253))|((~II27147));
assign II23196 = ((~WX6968))|((~II23194));
assign WX8346 = ((~WX8314));
assign II14250 = ((~II14252))|((~II14253));
assign WX466 = (WX464)|(WX463);
assign II3169 = ((~WX589))|((~WX503));
assign WX6839 = (WX6837)|(WX6836);
assign II15327 = ((~WX4479))|((~WX4404));
assign II2561 = ((~WX809))|((~WX873));
assign WX6192 = ((~II19099))|((~II19100));
assign WX4913 = ((~II15120))|((~II15121));
assign II3528 = ((~WX613))|((~_2106_));
assign WX1677 = ((~WX1676));
assign WX4493 = ((~WX4720));
assign II30039 = ((~WX9824))|((~II30038));
assign WX8686 = ((~II26909))|((~II26910));
assign II14934 = ((~WX4881))|((~II14933));
assign WX5035 = ((~WX4884));
assign WX7907 = ((~WX8761));
assign II9996 = ((~II10006))|((~II10007));
assign WX10718 = (WX10716)|(WX10715);
assign WX7093 = ((~WX7334));
assign II35300 = ((~WX10940))|((~WX10861));
assign WX4026 = (WX4037&WX4882);
assign WX4113 = (WX4111)|(WX4110);
assign WX10631 = (WX10642&WX11347);
assign WX10460 = (WX10458)|(WX10457);
assign WX6389 = (WX6388&WX6177);
assign WX2850 = (WX5003&WX2851);
assign WX7381 = ((~II22532))|((~II22533));
assign II31165 = ((~WX9637))|((~WX9548));
assign II26723 = ((~II26698))|((~II26722));
assign WX5609 = ((~WX6176));
assign WX4093 = (WX4091)|(WX4090);
assign WX9494 = ((~WX10054));
assign II3586 = ((~_2098_))|((~II3584));
assign II18936 = ((~II18946))|((~II18947));
assign WX7380 = ((~II22501))|((~II22502));
assign WX302 = (WX308&WX303);
assign WX1793 = (WX1796&RESET);
assign WX3973 = (WX3971)|(WX3970);
assign II27574 = ((~_2296_))|((~II27572));
assign II14476 = ((~WX4618))|((~II14475));
assign WX10994 = (WX10434&RESET);
assign WX10126 = ((~WX10125));
assign WX7466 = ((~WX7465));
assign II22245 = ((~WX7252))|((~WX7316));
assign II18792 = ((~II18782))|((~II18790));
assign II14010 = ((~WX4588))|((~II14002));
assign WX7976 = (WX7982&WX7977);
assign WX6318 = ((~II19333))|((~II19334));
assign II30032 = ((~II30022))|((~II30030));
assign WX3925 = (WX3923)|(WX3922);
assign II30304 = ((~WX9714))|((~II30302));
assign WX2725 = ((~WX3590));
assign WX11317 = ((~WX11316));
assign II30271 = ((~WX10052))|((~WX9712));
assign WX5566 = (WX6359&WX5567);
assign WX6082 = ((~II18341))|((~II18342));
assign WX7423 = ((~WX7394));
assign WX957 = ((~WX956));
assign WX10104 = ((~WX10103));
assign II18473 = ((~WX6173))|((~WX5847));
assign II34779 = ((~WX11101))|((~II34771));
assign WX9346 = (WX9572&WX10055);
assign WX10964 = ((~WX11197));
assign II3301 = ((~WX523))|((~II3299));
assign WX8931 = ((~WX8930));
assign II18707 = ((~WX6053))|((~II18705));
assign II6845 = ((~WX2120))|((~WX2184));
assign II2151 = ((~WX719))|((~II2150));
assign II34832 = ((~II34842))|((~II34843));
assign II22787 = ((~II22789))|((~II22790));
assign WX6089 = ((~II18558))|((~II18559));
assign WX6973 = (WX6976&RESET);
assign WX5610 = (WX5608)|(WX5607);
assign WX10283 = ((~II31528))|((~II31529));
assign WX5063 = ((~WX4884));
assign II19320 = ((~WX5771))|((~II19319));
assign WX10023 = ((~WX9955));
assign WX2263 = ((~WX2196));
assign II10232 = ((~WX3437))|((~II10230));
assign WX2073 = (WX2010&RESET);
assign WX1080 = (WX1078)|(WX1077);
assign WX1831 = (WX1834&RESET);
assign II6419 = ((~II6394))|((~II6418));
assign II31690 = ((~WX9684))|((~II31689));
assign WX10442 = (WX10440)|(WX10439);
assign WX6176 = ((~WX6169));
assign WX7859 = ((~WX8762));
assign WX10755 = ((~WX10746));
assign WX11160 = (WX11097&RESET);
assign II15643 = ((~_2187_))|((~II15641));
assign WX6744 = ((~WX7469));
assign II18760 = ((~WX5929))|((~II18759));
assign WX311 = ((~WX1004));
assign WX10003 = ((~WX9977));
assign II6714 = ((~WX2048))|((~II6713));
assign WX1172 = ((~WX1171));
assign WX8938 = ((~WX8937));
assign WX4269 = (WX6359&WX4270);
assign WX2839 = (WX3101&WX3590);
assign WX7371 = ((~II22222))|((~II22223));
assign II22377 = ((~II22352))|((~II22376));
assign WX10389 = ((~WX11348));
assign WX4850 = ((~WX4849));
assign WX6156 = ((~WX6082));
assign WX7834 = ((~WX7833));
assign WX7595 = ((~WX7594));
assign WX2268 = ((~WX2267));
assign WX7924 = (WX10126&WX7925);
assign WX5779 = ((~WX5747));
assign WX9865 = (WX9802&RESET);
assign WX5077 = ((~WX4884));
assign II10759 = ((~WX3471))|((~II10757));
assign II34276 = ((~WX11345))|((~WX11005));
assign WX8860 = ((~WX8859));
assign WX8384 = ((~WX8623));
assign II14027 = ((~II14017))|((~II14025));
assign II6692 = ((~WX2174))|((~II6690));
assign WX11494 = (WX11492)|(WX11491);
assign II34671 = ((~II34646))|((~II34670));
assign II22415 = ((~II22417))|((~II22418));
assign WX670 = (WX230&RESET);
assign WX3203 = ((~WX3433));
assign II22786 = ((~II22796))|((~II22797));
assign DATA_9_5 = ((~WX1193));
assign WX7418 = ((~WX7417));
assign WX848 = (WX785&RESET);
assign II26763 = ((~WX8760))|((~II26762));
assign II26552 = ((~WX8501))|((~II26544));
assign WX4143 = (WX6296&WX4144);
assign WX10306 = ((~II31697))|((~II31698));
assign WX9119 = (WX11370&WX9120);
assign II30333 = ((~WX10052))|((~WX9716));
assign WX10401 = (WX10831&WX11348);
assign II6969 = ((~WX2128))|((~WX2192));
assign WX4547 = (WX4095&RESET);
assign WX619 = ((~WX851));
assign WX1368 = ((~WX1359));
assign WX9966 = ((~II30511))|((~II30512));
assign WX4228 = ((~WX4883));
assign WX6987 = (WX6990&RESET);
assign WX3153 = ((~WX3525));
assign WX1262 = ((~II3711))|((~II3712));
assign WX2001 = (WX1938&RESET);
assign II35287 = ((~WX10939))|((~WX10859));
assign WX5100 = ((~WX5099));
assign II30883 = ((~II30858))|((~II30882));
assign II26847 = ((~II26822))|((~II26846));
assign WX3002 = (WX3000)|(WX2999);
assign WX4793 = ((~II14460))|((~II14461));
assign WX11370 = ((~WX11369));
assign DATA_9_30 = ((~WX1018));
assign II22811 = ((~II22786))|((~II22810));
assign WX11158 = (WX11095&RESET);
assign WX5431 = (WX5442&WX6175);
assign WX4381 = (WX4384&RESET);
assign II14311 = ((~II14321))|((~II14322));
assign WX3946 = (_2202_&WX4883);
assign WX4260 = ((~WX4883));
assign WX5749 = ((~WX6131));
assign II14422 = ((~WX4678))|((~II14421));
assign II7396 = ((~WX1899))|((~II7395));
assign WX11477 = (WX11476&WX11349);
assign WX1113 = (WX595&WX1114);
assign II31271 = ((~WX9564))|((~II31269));
assign II18116 = ((~WX5951))|((~WX6015));
assign II14902 = ((~WX4881))|((~WX4582));
assign WX8965 = ((~WX8964));
assign WX9398 = (_2310_&WX10055);
assign WX2161 = (WX2098&RESET);
assign WX8047 = ((~WX8761));
assign II31675 = ((~WX9681))|((~_2313_));
assign II6248 = ((~WX2018))|((~II6240));
assign II11063 = ((~WX3166))|((~II11062));
assign WX8017 = (WX8028&WX8761);
assign WX2764 = (WX2762)|(WX2761);
assign II10952 = ((~II10942))|((~II10950));
assign WX706 = (WX482&RESET);
assign WX1685 = (WX1683)|(WX1682);
assign II6504 = ((~WX2098))|((~WX2162));
assign II6233 = ((~II6208))|((~II6232));
assign WX3559 = ((~WX3558));
assign WX9125 = (WX9123)|(WX9122);
assign II2560 = ((~II2562))|((~II2563));
assign WX6640 = (WX6651&WX7468);
assign WX1473 = (WX3668&WX1474);
assign WX10415 = (WX10833&WX11348);
assign WX2631 = ((~WX3590));
assign WX1100 = ((~WX1005));
assign WX369 = ((~WX360));
assign WX3774 = ((~II11401))|((~II11402));
assign WX790 = (WX727&RESET);
assign WX6593 = (WX7519&WX6594);
assign WX1210 = (WX1209&WX1005);
assign WX9134 = ((~WX10055));
assign WX9003 = ((~II27622))|((~II27623));
assign II2336 = ((~WX731))|((~II2328));
assign II6947 = ((~II6937))|((~II6945));
assign WX10018 = ((~WX10017));
assign WX2573 = (WX2549&WX2556);
assign WX5219 = ((~WX5210));
assign II14460 = ((~II14435))|((~II14459));
assign II3157 = ((~WX588))|((~II3156));
assign II2174 = ((~WX1001))|((~WX657));
assign WX7506 = ((~II23143))|((~II23144));
assign WX9976 = ((~II30821))|((~II30822));
assign II14521 = ((~II14497))|((~II14513));
assign II10261 = ((~WX3375))|((~WX3439));
assign WX4599 = (WX4536&RESET);
assign WX3950 = (WX4368&WX4883);
assign WX9679 = ((~WX9920));
assign II30596 = ((~WX9860))|((~WX9924));
assign II26373 = ((~II26375))|((~II26376));
assign II11582 = ((~_2164_))|((~II11580));
assign WX4553 = (WX4137&RESET);
assign WX6309 = ((~WX6308));
assign WX4703 = (WX4640&RESET);
assign WX7641 = (WX7069&WX7642);
assign WX3163 = ((~WX3545));
assign II30527 = ((~WX9792))|((~II30526));
assign WX1920 = ((~WX2160));
assign WX9685 = ((~WX9932));
assign WX4930 = ((~WX4884));
assign WX9143 = (WX9149&WX9144);
assign WX7665 = ((~WX7664));
assign WX6480 = (WX6416&WX6435);
assign II14204 = ((~WX4664))|((~WX4728));
assign II18754 = ((~WX5865))|((~II18752));
assign II14653 = ((~II14655))|((~II14656));
assign II10859 = ((~II10849))|((~II10857));
assign WX5986 = (WX5923&RESET);
assign II34092 = ((~WX10993))|((~II34090));
assign WX5059 = ((~WX5058));
assign II22152 = ((~WX7246))|((~WX7310));
assign II26335 = ((~WX8487))|((~II26327));
assign II34477 = ((~WX11145))|((~WX11209));
assign WX9458 = (WX9588&WX10055);
assign WX2538 = ((~II7597))|((~II7598));
assign WX9503 = (WX9501)|(WX9500);
assign WX4103 = (WX4101)|(WX4100);
assign II3143 = ((~WX587))|((~WX499));
assign WX8801 = (WX8343&WX8802);
assign WX10693 = ((~WX11348));
assign WX3668 = ((~WX3667));
assign II23673 = ((~WX7096))|((~II23672));
assign WX2375 = ((~WX2374));
assign WX1316 = (WX1240&WX1263);
assign WX9557 = (WX9560&RESET);
assign II23695 = ((~_2244_))|((~II23693));
assign II6527 = ((~WX2036))|((~II6519));
assign WX7870 = (WX7868)|(WX7867);
assign II22641 = ((~WX7214))|((~II22640));
assign WX10794 = (WX11559&WX10795);
assign II7265 = ((~WX1889))|((~WX1810));
assign WX7657 = (WX7655)|(WX7654);
assign WX2043 = (WX1980&RESET);
assign WX2517 = (WX2516&WX2298);
assign WX1866 = ((~WX2244));
assign WX5836 = (WX5360&RESET);
assign WX9883 = (WX9820&RESET);
assign WX3793 = ((~WX3792));
assign II35645 = ((~WX10968))|((~_2351_));
assign II2554 = ((~WX745))|((~II2553));
assign WX6344 = ((~WX6343));
assign WX6795 = (WX6801&WX6796);
assign II18382 = ((~WX5841))|((~II18380));
assign WX3906 = (WX3824&WX3849);
assign II7659 = ((~WX1926))|((~_2118_));
assign WX1020 = ((~II3079))|((~II3080));
assign WX8195 = ((~WX8762));
assign WX1583 = (WX1581)|(WX1580);
assign WX1927 = ((~WX2174));
assign II15671 = ((~_2182_))|((~II15669));
assign WX3533 = ((~WX3532));
assign WX6075 = ((~II18124))|((~II18125));
assign WX2619 = (WX2528&WX2556);
assign II6079 = ((~II6069))|((~II6077));
assign II14678 = ((~II14668))|((~II14676));
assign WX4247 = (WX4245)|(WX4244);
assign II34367 = ((~II34377))|((~II34378));
assign WX7869 = ((~WX8762));
assign II22734 = ((~WX7220))|((~II22733));
assign II3683 = ((~WX637))|((~II3682));
assign II23546 = ((~WX7077))|((~_2267_));
assign WX2559 = (WX2555&WX2556);
assign WX5942 = (WX5879&RESET);
assign WX11538 = ((~WX11537));
assign WX7265 = (WX7202&RESET);
assign II11480 = ((~WX3213))|((~_2172_));
assign II31388 = ((~WX9582))|((~II31386));
assign II6766 = ((~II6776))|((~II6777));
assign WX6030 = (WX5967&RESET);
assign WX4817 = ((~WX4798));
assign WX5772 = ((~WX5740));
assign WX6028 = (WX5965&RESET);
assign WX4861 = ((~WX4788));
assign II34904 = ((~WX11109))|((~II34903));
assign WX3078 = (WX3081&RESET);
assign WX5390 = (WX5396&WX5391);
assign WX816 = (WX753&RESET);
assign WX7331 = (WX7268&RESET);
assign WX9276 = (WX9562&WX10055);
assign WX3114 = (WX3117&RESET);
assign WX7823 = ((~WX8761));
assign WX8540 = (WX8477&RESET);
assign WX10665 = ((~WX11348));
assign WX1097 = ((~II3222))|((~II3223));
assign II14717 = ((~WX4881))|((~II14716));
assign WX11554 = (WX11553&WX11349);
assign WX4211 = (WX4209)|(WX4208);
assign II2035 = ((~WX775))|((~II2034));
assign WX9386 = ((~WX10055));
assign WX8796 = (WX8794)|(WX8793);
assign WX9658 = ((~WX9626));
assign II15678 = ((~_2181_))|((~II15676));
assign WX6375 = (WX6374&WX6177);
assign WX4371 = (WX4374&RESET);
assign WX700 = (WX440&RESET);
assign WX4313 = (WX4311)|(WX4310);
assign WX4354 = ((~WX4883));
assign WX3685 = (WX3179&WX3686);
assign WX3993 = (WX4926&WX3994);
assign WX4859 = ((~WX4787));
assign WX5362 = (WX5368&WX5363);
assign II14119 = ((~II14094))|((~II14118));
assign WX3783 = (WX3193&WX3784);
assign II35445 = ((~WX10883))|((~II35443));
assign II27382 = ((~WX8361))|((~II27381));
assign WX10291 = ((~II31592))|((~II31593));
assign WX10741 = ((~WX10732));
assign II6410 = ((~II6412))|((~II6413));
assign WX6776 = ((~WX7469));
assign II10944 = ((~WX3419))|((~II10943));
assign II27148 = ((~WX8343))|((~II27147));
assign WX8819 = ((~WX8818));
assign WX11080 = (WX11017&RESET);
assign II18242 = ((~WX6023))|((~II18240));
assign II11193 = ((~WX3176))|((~II11192));
assign II3542 = ((~WX615))|((~_2104_));
assign II14098 = ((~WX4530))|((~II14096));
assign WX10482 = (DATA_0_24&WX10483);
assign II6814 = ((~WX2118))|((~WX2182));
assign II18024 = ((~WX5945))|((~II18023));
assign WX8470 = (WX8407&RESET);
assign WX10185 = (WX9649&WX10186);
assign II27532 = ((~_2300_))|((~II27530));
assign WX610 = ((~WX578));
assign WX4307 = (WX4313&WX4308);
assign II6303 = ((~WX2294))|((~WX1958));
assign WX5563 = ((~WX6176));
assign II2158 = ((~WX783))|((~WX847));
assign II30760 = ((~II30750))|((~II30758));
assign WX11364 = ((~II35119))|((~II35120));
assign II30728 = ((~II30703))|((~II30727));
assign II14135 = ((~WX4596))|((~II14134));
assign II6519 = ((~II6521))|((~II6522));
assign WX8809 = ((~WX8763));
assign II34538 = ((~II34540))|((~II34541));
assign WX9106 = ((~WX10055));
assign II6745 = ((~WX2050))|((~II6744));
assign II6736 = ((~II6738))|((~II6739));
assign II26485 = ((~WX8433))|((~II26483));
assign WX10904 = ((~WX11333));
assign WX6724 = (WX6735&WX7468);
assign WX976 = ((~WX906));
assign WX7890 = ((~WX7889));
assign WX1521 = (WX1519)|(WX1518);
assign WX4048 = (WX4382&WX4883);
assign WX5966 = (WX5903&RESET);
assign WX9757 = (WX9533&RESET);
assign II10579 = ((~II10554))|((~II10578));
assign WX5558 = (WX5564&WX5559);
assign WX10942 = ((~WX10910));
assign II14761 = ((~II14763))|((~II14764));
assign WX6504 = (_2268_&WX7469);
assign WX7735 = (WX7725&WX7728);
assign II2747 = ((~WX821))|((~WX885));
assign II26939 = ((~II26915))|((~II26931));
assign II14531 = ((~WX4881))|((~II14530));
assign WX8926 = (WX8925&WX8763);
assign WX7683 = (WX7075&WX7684);
assign WX8632 = (WX8569&RESET);
assign II23182 = ((~WX7053))|((~II23181));
assign WX2285 = ((~WX2207));
assign WX6663 = (WX7554&WX6664);
assign II6451 = ((~II6441))|((~II6449));
assign II2942 = ((~II2932))|((~II2940));
assign II19150 = ((~WX5758))|((~WX5669));
assign WX8367 = ((~WX8335));
assign WX3143 = ((~WX3569));
assign WX7349 = (WX7286&RESET);
assign WX633 = ((~WX879));
assign II7547 = ((~WX1908))|((~_2136_));
assign II34143 = ((~II34119))|((~II34135));
assign II34043 = ((~WX11117))|((~WX11181));
assign WX105 = (WX116&WX1003);
assign II11487 = ((~_2156_))|((~II11479));
assign WX2406 = (WX1888&WX2407);
assign II31600 = ((~_2325_))|((~II31598));
assign WX2037 = (WX1974&RESET);
assign WX8594 = (WX8531&RESET);
assign WX8610 = (WX8547&RESET);
assign II14296 = ((~II14298))|((~II14299));
assign II14407 = ((~WX4880))|((~II14406));
assign II6134 = ((~WX2138))|((~II6132));
assign WX9064 = (WX9003&WX9021);
assign II14485 = ((~WX4746))|((~II14483));
assign WX5047 = (WX5046&WX4884);
assign WX7516 = ((~WX7470));
assign II26924 = ((~WX8525))|((~II26916));
assign WX11100 = (WX11037&RESET);
assign WX270 = (WX268)|(WX267);
assign WX11212 = (WX11149&RESET);
assign WX3858 = (WX3819&WX3849);
assign WX2319 = ((~WX2318));
assign WX10715 = (WX10726&WX11347);
assign II11547 = ((~_2169_))|((~II11545));
assign WX8827 = ((~II27200))|((~II27201));
assign WX1030 = ((~WX1005));
assign WX11590 = ((~II35639))|((~II35640));
assign WX10519 = (WX10530&WX11347);
assign II7085 = ((~WX1782))|((~II7083));
assign WX6910 = (_2239_&WX7469);
assign II34337 = ((~II34339))|((~II34340));
assign WX2438 = ((~WX2437));
assign II18310 = ((~II18285))|((~II18309));
assign II34680 = ((~WX11346))|((~II34679));
assign II3236 = ((~WX513))|((~II3234));
assign WX4802 = ((~II14739))|((~II14740));
assign II31101 = ((~WX9632))|((~II31100));
assign II27537 = ((~_2272_))|((~II27529));
assign WX5496 = (WX6324&WX5497);
assign II18317 = ((~II18319))|((~II18320));
assign II34323 = ((~WX11135))|((~II34322));
assign II6537 = ((~WX2164))|((~II6535));
assign II18544 = ((~II18534))|((~II18542));
assign WX11291 = ((~WX11290));
assign WX10935 = ((~WX10903));
assign II31218 = ((~WX9641))|((~II31217));
assign WX569 = ((~WX943));
assign WX5442 = (WX5440)|(WX5439);
assign WX2884 = (WX2882)|(WX2881);
assign II34531 = ((~WX11085))|((~II34523));
assign WX3090 = (WX3093&RESET);
assign WX6064 = (WX6001&RESET);
assign II18335 = ((~WX6029))|((~II18333));
assign WX7520 = ((~II23169))|((~II23170));
assign WX4979 = ((~WX4884));
assign II34353 = ((~WX11137))|((~WX11201));
assign II22448 = ((~WX7466))|((~II22447));
assign WX162 = (WX168&WX163);
assign WX5528 = ((~WX5527));
assign WX3573 = ((~WX3572));
assign WX9070 = (WX9000&WX9021);
assign WX4981 = ((~WX4980));
assign WX9364 = ((~WX9355));
assign II11154 = ((~WX3173))|((~II11153));
assign WX5081 = ((~II15432))|((~II15433));
assign WX7131 = (WX6667&RESET);
assign WX6328 = ((~WX6177));
assign WX5896 = (WX5833&RESET);
assign WX562 = ((~WX993));
assign WX5956 = (WX5893&RESET);
assign WX5380 = (WX7561&WX5381);
assign WX11565 = ((~WX11564));
assign DATA_9_31 = ((~WX1011));
assign II35013 = ((~II35003))|((~II35011));
assign II18506 = ((~WX5849))|((~II18504));
assign WX5476 = (WX5474)|(WX5473);
assign II34037 = ((~II34027))|((~II34035));
assign WX7372 = ((~II22253))|((~II22254));
assign II31269 = ((~WX9645))|((~WX9564));
assign WX3799 = (WX3797)|(WX3796);
assign WX8752 = ((~WX8673));
assign II10927 = ((~II10929))|((~II10930));
assign WX2569 = (WX2551&WX2556);
assign WX9442 = ((~WX10055));
assign II11206 = ((~WX3177))|((~II11205));
assign II10247 = ((~WX3587))|((~II10246));
assign WX9526 = ((~WX10055));
assign II26884 = ((~II26894))|((~II26895));
assign WX1463 = (WX2368&WX1464);
assign II30765 = ((~II30775))|((~II30776));
assign WX3515 = ((~II10920))|((~II10921));
assign WX906 = ((~II2197))|((~II2198));
assign II14900 = ((~II14910))|((~II14911));
assign II34060 = ((~WX11345))|((~II34059));
assign WX2431 = ((~WX2430));
assign WX3804 = (WX3196&WX3805);
assign WX7957 = ((~WX8762));
assign WX5520 = (WX7631&WX5521);
assign II15573 = ((~_2198_))|((~II15571));
assign WX10527 = (WX10849&WX11348);
assign WX2297 = ((~WX2290));
assign II26614 = ((~WX8505))|((~II26606));
assign II14113 = ((~WX4722))|((~II14111));
assign WX3159 = ((~WX3537));
assign II26226 = ((~II26202))|((~II26218));
assign II11566 = ((~WX3203))|((~_2166_));
assign WX9017 = ((~II27720))|((~II27721));
assign II34106 = ((~WX11121))|((~II34105));
assign WX5340 = (WX5338)|(WX5337);
assign WX9648 = ((~WX9616));
assign WX4963 = (WX4962&WX4884);
assign WX7100 = ((~WX7348));
assign WX7303 = (WX7240&RESET);
assign II22283 = ((~II22259))|((~II22275));
assign WX1074 = ((~WX1073));
assign II18869 = ((~II18859))|((~II18867));
assign II10346 = ((~WX3317))|((~II10338));
assign II30052 = ((~II30062))|((~II30063));
assign WX9444 = (WX9586&WX10055);
assign WX9935 = (WX9872&RESET);
assign WX7028 = ((~WX7460));
assign WX4443 = ((~WX4812));
assign WX2794 = (WX4975&WX2795);
assign WX7826 = (WX10077&WX7827);
assign II10338 = ((~II10340))|((~II10341));
assign WX6420 = ((~II19633))|((~II19634));
assign WX2537 = ((~II7590))|((~II7591));
assign WX10512 = (WX10510)|(WX10509);
assign WX8142 = ((~WX8141));
assign II19723 = ((~WX5813))|((~_2206_));
assign II6165 = ((~WX2140))|((~II6163));
assign WX1107 = ((~WX1005));
assign II11686 = ((~WX3222))|((~II11685));
assign WX6919 = ((~WX6918));
assign WX9905 = (WX9842&RESET);
assign II34484 = ((~II34460))|((~II34476));
assign II31244 = ((~WX9643))|((~II31243));
assign II11428 = ((~WX3127))|((~II11426));
assign WX5870 = (WX5598&RESET);
assign II2220 = ((~WX787))|((~WX851));
assign WX5191 = (WX5121&WX5142);
assign WX7633 = (WX7632&WX7470);
assign II6356 = ((~II6332))|((~II6348));
assign WX10979 = ((~WX11227));
assign II3696 = ((~WX640))|((~_2079_));
assign DATA_9_21 = ((~WX1081));
assign II6580 = ((~II6590))|((~II6591));
assign II31139 = ((~WX9635))|((~WX9544));
assign WX10507 = ((~WX11347));
assign WX10060 = ((~WX10056));
assign WX172 = (WX170)|(WX169);
assign WX1751 = (WX1749)|(WX1748);
assign WX5356 = (WX6254&WX5357);
assign II26111 = ((~WX8759))|((~WX8409));
assign WX3591 = ((~WX3582));
assign WX4051 = (WX4049)|(WX4048);
assign WX6666 = ((~WX6657));
assign II30381 = ((~WX9910))|((~II30379));
assign II34625 = ((~WX11091))|((~II34624));
assign II2406 = ((~WX799))|((~WX863));
assign WX10164 = (WX9646&WX10165);
assign WX4239 = (WX4237)|(WX4236);
assign II10106 = ((~WX3365))|((~WX3429));
assign WX453 = ((~WX444));
assign WX9641 = ((~WX9609));
assign II22640 = ((~WX7214))|((~II22632));
assign WX7637 = ((~WX7636));
assign II11666 = ((~_2150_))|((~II11664));
assign WX6091 = ((~II18620))|((~II18621));
assign WX5438 = (WX5436)|(WX5435);
assign WX3984 = (WX3995&WX4882);
assign WX7883 = ((~WX8762));
assign II10201 = ((~WX3435))|((~II10199));
assign WX6704 = (WX6978&WX7469);
assign WX11339 = ((~WX11338));
assign II3570 = ((~WX619))|((~_2100_));
assign WX8784 = ((~WX8783));
assign WX551 = ((~WX971));
assign WX3493 = ((~II10238))|((~II10239));
assign II11348 = ((~WX3188))|((~WX3115));
assign WX11486 = ((~WX11349));
assign II14624 = ((~WX4881))|((~II14623));
assign WX5787 = ((~WX6015));
assign WX11608 = (WX11578&WX11607);
assign WX5345 = ((~WX5336));
assign WX9485 = (WX9483)|(WX9482);
assign WX6169 = ((~TM0));
assign WX10299 = ((~II31648))|((~II31649));
assign WX2340 = ((~WX2339));
assign II30924 = ((~WX9754))|((~II30922));
assign WX8908 = (WX8906)|(WX8905);
assign WX3302 = (WX3239&RESET);
assign II6782 = ((~II6784))|((~II6785));
assign WX2713 = (WX3083&WX3590);
assign WX9771 = (WX9708&RESET);
assign WX7155 = (WX6835&RESET);
assign II22703 = ((~WX7218))|((~II22702));
assign WX2926 = (WX2924)|(WX2923);
assign WX1579 = ((~WX1578));
assign II34260 = ((~WX11131))|((~WX11195));
assign II26050 = ((~WX8759))|((~II26049));
assign II7162 = ((~WX1881))|((~II7161));
assign II19633 = ((~WX5797))|((~II19632));
assign II10254 = ((~WX3311))|((~II10253));
assign WX394 = (DATA_9_6&WX395);
assign II27292 = ((~WX8275))|((~II27290));
assign II26299 = ((~WX8421))|((~II26297));
assign WX9098 = ((~WX9089));
assign WX3134 = ((~WX3551));
assign WX1710 = (_2113_&WX2297);
assign WX5822 = (WX5262&RESET);
assign II30931 = ((~II30921))|((~II30929));
assign II26443 = ((~II26419))|((~II26435));
assign II14709 = ((~II14699))|((~II14707));
assign WX10047 = ((~TM0));
assign II14344 = ((~WX4880))|((~WX4546));
assign WX913 = ((~II2414))|((~II2415));
assign II18564 = ((~II18574))|((~II18575));
assign WX10177 = (WX10176&WX10056);
assign WX2778 = (WX2776)|(WX2775);
assign II15264 = ((~WX4394))|((~II15262));
assign WX6275 = ((~WX6274));
assign WX4848 = ((~WX4847));
assign II6087 = ((~WX2294))|((~II6086));
assign II14733 = ((~WX4762))|((~II14731));
assign WX10580 = (DATA_0_17&WX10581);
assign WX923 = ((~II2724))|((~II2725));
assign II6635 = ((~II6611))|((~II6627));
assign WX2649 = (WX2660&WX3589);
assign WX7291 = (WX7228&RESET);
assign WX11222 = (WX11159&RESET);
assign WX1029 = (WX583&WX1030);
assign WX2177 = (WX2114&RESET);
assign II15664 = ((~_2184_))|((~II15662));
assign WX1556 = (_2124_&WX2297);
assign WX5728 = ((~WX6153));
assign II30946 = ((~II30936))|((~II30944));
assign II15648 = ((~WX4508))|((~_2186_));
assign WX5017 = ((~WX5016));
assign II27162 = ((~WX8255))|((~II27160));
assign WX2683 = ((~WX3590));
assign II23721 = ((~WX7105))|((~_2239_));
assign II27678 = ((~WX8389))|((~II27677));
assign WX7946 = ((~WX7945));
assign WX4000 = ((~WX4882));
assign II27567 = ((~_2297_))|((~II27565));
assign WX6603 = (WX8819&WX6604);
assign II6397 = ((~WX2294))|((~II6396));
assign II26453 = ((~WX8759))|((~II26452));
assign WX7081 = ((~WX7310));
assign WX228 = (WX226)|(WX225);
assign WX6393 = ((~WX6392));
assign WX7003 = (WX7006&RESET);
assign WX9945 = (WX9882&RESET);
assign WX11008 = (WX10532&RESET);
assign II34028 = ((~WX11345))|((~WX10989));
assign WX3747 = (WX3746&WX3591);
assign WX10556 = (WX11440&WX10557);
assign WX8506 = (WX8443&RESET);
assign WX1135 = ((~WX1005));
assign II26645 = ((~WX8507))|((~II26637));
assign WX4257 = (WX4255)|(WX4254);
assign II15095 = ((~WX4368))|((~II15093));
assign II14444 = ((~WX4616))|((~II14436));
assign II6976 = ((~II6952))|((~II6968));
assign WX926 = ((~II2817))|((~II2818));
assign II27595 = ((~_2293_))|((~II27593));
assign II6676 = ((~WX2295))|((~II6675));
assign WX7950 = (WX7948)|(WX7947);
assign WX1535 = (WX1533)|(WX1532);
assign WX4274 = ((~WX4883));
assign WX6658 = (_2257_&WX7469);
assign WX750 = (WX687&RESET);
assign II34703 = ((~II34693))|((~II34701));
assign WX4359 = (WX4357)|(WX4356);
assign WX10683 = ((~WX11348));
assign WX7281 = (WX7218&RESET);
assign WX7549 = (WX7548&WX7470);
assign WX11070 = (WX11007&RESET);
assign II7253 = ((~WX1888))|((~II7252));
assign WX4197 = (WX4195)|(WX4194);
assign WX7607 = ((~WX7470));
assign WX10382 = (WX10380)|(WX10379);
assign II30247 = ((~WX9774))|((~II30239));
assign II34996 = ((~WX11115))|((~II34988));
assign WX2561 = (WX2554&WX2556);
assign WX7937 = (_2290_&WX8762);
assign WX2518 = (WX1904&WX2519);
assign WX2997 = ((~WX2988));
assign WX3060 = (WX5108&WX3061);
assign II14833 = ((~II14823))|((~II14831));
assign II10479 = ((~WX3389))|((~II10478));
assign WX9287 = (WX11454&WX9288);
assign WX2525 = ((~II7498))|((~II7499));
assign WX9622 = ((~WX9998));
assign WX804 = (WX741&RESET);
assign WX1772 = ((~WX2297));
assign WX5996 = (WX5933&RESET);
assign WX7068 = ((~WX7036));
assign WX4008 = ((~WX4883));
assign II23298 = ((~WX7062))|((~WX6984));
assign II2307 = ((~II2297))|((~II2305));
assign II18016 = ((~WX5881))|((~II18015));
assign II7201 = ((~WX1884))|((~II7200));
assign WX3430 = (WX3367&RESET);
assign WX4023 = (WX4021)|(WX4020);
assign WX9056 = (WX9007&WX9021);
assign WX10422 = (WX10428&WX10423);
assign WX10067 = ((~WX10056));
assign WX8334 = ((~WX8715));
assign WX9201 = (WX9199)|(WX9198);
assign II18216 = ((~II18192))|((~II18208));
assign II30939 = ((~WX9946))|((~II30937));
assign WX1197 = (WX607&WX1198);
assign WX4300 = (WX4418&WX4883);
assign WX7555 = ((~II23234))|((~II23235));
assign WX6331 = ((~WX6330));
assign WX4827 = ((~WX4803));
assign II6839 = ((~II6829))|((~II6837));
assign WX4627 = (WX4564&RESET);
assign WX9607 = ((~WX10032));
assign WX8318 = ((~WX8747));
assign II2548 = ((~WX681))|((~II2546));
assign WX11050 = (WX10826&RESET);
assign II14818 = ((~II14808))|((~II14816));
assign II2725 = ((~II2715))|((~II2723));
assign WX8586 = (WX8523&RESET);
assign WX1909 = ((~WX2138));
assign II27733 = ((~WX8399))|((~_2270_));
assign WX10227 = (WX9655&WX10228);
assign II22293 = ((~WX7466))|((~II22292));
assign II10385 = ((~WX3383))|((~WX3447));
assign WX5778 = ((~WX5746));
assign WX1646 = ((~WX2297));
assign WX10233 = (WX10232&WX10056);
assign WX4431 = ((~WX4852));
assign II22107 = ((~WX7466))|((~II22106));
assign II14482 = ((~II14484))|((~II14485));
assign WX10894 = ((~WX11313));
assign WX1454 = (WX1465&WX2296);
assign II26274 = ((~WX8483))|((~II26273));
assign II27642 = ((~WX8383))|((~_2286_));
assign II10216 = ((~WX3587))|((~II10215));
assign WX7059 = ((~WX7027));
assign WX6160 = ((~WX6084));
assign WX542 = (WX545&RESET);
assign II26901 = ((~WX8587))|((~WX8651));
assign II26190 = ((~WX8605))|((~II26188));
assign II3598 = ((~WX623))|((~_2096_));
assign II18692 = ((~WX5861))|((~II18690));
assign WX1401 = (WX1399)|(WX1398);
assign II26839 = ((~WX8583))|((~WX8647));
assign II30504 = ((~WX9854))|((~II30503));
assign WX3838 = ((~II11651))|((~II11652));
assign WX3058 = (WX3056)|(WX3055);
assign WX10810 = (WX10808)|(WX10807);
assign II19618 = ((~WX5795))|((~_2224_));
assign II11168 = ((~WX3087))|((~II11166));
assign WX11452 = (WX11450)|(WX11449);
assign II14360 = ((~WX4674))|((~II14359));
assign WX8184 = ((~WX8183));
assign II22392 = ((~WX7198))|((~II22384));
assign II18302 = ((~WX5963))|((~WX6027));
assign II14578 = ((~WX4752))|((~II14576));
assign II10580 = ((~II10570))|((~II10578));
assign WX483 = ((~WX485));
assign WX9377 = (WX9375)|(WX9374);
assign WX6361 = (WX6360&WX6177);
assign II7422 = ((~WX1901))|((~II7421));
assign WX11354 = (WX11352)|(WX11351);
assign II34245 = ((~WX11345))|((~WX11003));
assign II6661 = ((~WX2172))|((~II6659));
assign WX5655 = ((~WX5657));
assign II2748 = ((~WX821))|((~II2747));
assign II27084 = ((~WX8243))|((~II27082));
assign II31401 = ((~WX9584))|((~II31399));
assign WX10204 = ((~II31361))|((~II31362));
assign WX5464 = (WX7603&WX5465);
assign II22068 = ((~II22058))|((~II22066));
assign II6520 = ((~WX2295))|((~WX1972));
assign WX2149 = (WX2086&RESET);
assign WX8361 = ((~WX8329));
assign II6318 = ((~WX2086))|((~WX2150));
assign WX11567 = ((~II35496))|((~II35497));
assign II26428 = ((~WX8493))|((~II26420));
assign WX2750 = (WX2748)|(WX2747);
assign WX4970 = (WX4969&WX4884);
assign WX802 = (WX739&RESET);
assign II26528 = ((~II26530))|((~II26531));
assign WX1437 = (WX1435)|(WX1434);
assign WX11331 = ((~WX11330));
assign WX7449 = ((~WX7375));
assign II18278 = ((~II18254))|((~II18270));
assign II27435 = ((~WX8297))|((~II27433));
assign WX10779 = (WX10885&WX11348);
assign II31089 = ((~WX9536))|((~II31087));
assign II22633 = ((~WX7467))|((~WX7150));
assign WX5627 = (WX5638&WX6175);
assign WX10345 = (WX10301&WX10314);
assign II18946 = ((~WX5941))|((~II18945));
assign WX10560 = ((~WX10559));
assign WX11461 = ((~WX11460));
assign II14591 = ((~II14593))|((~II14594));
assign WX5313 = (WX5671&WX6176);
assign WX940 = ((~WX920));
assign WX1528 = (_2126_&WX2297);
assign WX7897 = ((~WX8762));
assign II3647 = ((~WX631))|((~_2088_));
assign II10617 = ((~II10619))|((~II10620));
assign WX5153 = (WX5138&WX5142);
assign II30558 = ((~WX9794))|((~II30557));
assign II22867 = ((~WX7356))|((~II22865));
assign II19653 = ((~WX5801))|((~_2218_));
assign II23715 = ((~WX7103))|((~II23714));
assign WX3332 = (WX3269&RESET);
assign II7057 = ((~WX1873))|((~WX1778));
assign WX9853 = (WX9790&RESET);
assign II26057 = ((~WX8469))|((~II26056));
assign II26591 = ((~WX8567))|((~WX8631));
assign WX3892 = (WX3831&WX3849);
assign WX3814 = ((~WX3813));
assign WX3844 = ((~II11693))|((~II11694));
assign II11637 = ((~WX3214))|((~II11636));
assign WX3444 = (WX3381&RESET);
assign WX4280 = ((~WX4882));
assign WX9837 = (WX9774&RESET);
assign II11553 = ((~WX3201))|((~II11552));
assign WX9326 = ((~WX10054));
assign WX3543 = ((~WX3542));
assign WX5813 = ((~WX6067));
assign II23273 = ((~WX7060))|((~II23272));
assign WX2706 = (WX2712&WX2707);
assign WX3910 = (WX3822&WX3849);
assign WX9575 = (WX9578&RESET);
assign WX2799 = ((~WX3590));
assign II19590 = ((~WX5791))|((~_2228_));
assign WX1717 = (WX1715)|(WX1714);
assign II34524 = ((~WX11346))|((~WX11021));
assign II10176 = ((~II10151))|((~II10175));
assign WX4293 = (WX4299&WX4294);
assign WX107 = ((~WX1003));
assign WX1246 = ((~II3599))|((~II3600));
assign II34330 = ((~II34305))|((~II34329));
assign II2110 = ((~II2120))|((~II2121));
assign WX8681 = ((~II26754))|((~II26755));
assign II6646 = ((~WX1980))|((~II6644));
assign II31152 = ((~WX9636))|((~WX9546));
assign II26358 = ((~II26360))|((~II26361));
assign WX9224 = ((~WX9215));
assign WX2454 = (WX2453&WX2298);
assign WX5702 = (WX5705&RESET);
assign WX11630 = (WX11576&WX11607);
assign WX11520 = (WX10948&WX11521);
assign II3391 = ((~WX606))|((~II3390));
assign WX6565 = (WX7505&WX6566);
assign II23541 = ((~_2268_))|((~II23539));
assign WX9761 = (WX9698&RESET);
assign II35339 = ((~WX10943))|((~WX10867));
assign WX3960 = (_2201_&WX4883);
assign II22494 = ((~WX7268))|((~II22493));
assign WX6959 = (WX6962&RESET);
assign WX8462 = (WX8226&RESET);
assign WX7751 = (WX7697&WX7728);
assign WX11383 = ((~WX11382));
assign WX4188 = (WX4402&WX4883);
assign WX1160 = ((~II3339))|((~II3340));
assign WX5633 = ((~WX6176));
assign II18961 = ((~II18936))|((~II18960));
assign II26243 = ((~WX8481))|((~II26242));
assign WX1898 = ((~WX1866));
assign II31626 = ((~WX9673))|((~_2321_));
assign WX3046 = (WX5101&WX3047);
assign WX6343 = (WX6341)|(WX6340);
assign WX7217 = (WX7154&RESET);
assign WX10545 = ((~WX10536));
assign II31528 = ((~_2311_))|((~II31527));
assign WX11456 = (WX11455&WX11349);
assign WX1338 = ((~WX2297));
assign II6629 = ((~WX2106))|((~II6628));
assign II18806 = ((~II18781))|((~II18805));
assign WX7679 = ((~WX7678));
assign WX11152 = (WX11089&RESET);
assign II22724 = ((~II22734))|((~II22735));
assign II6914 = ((~II6890))|((~II6906));
assign II26544 = ((~II26546))|((~II26547));
assign WX1350 = (WX1780&WX2297);
assign WX6116 = ((~WX6094));
assign II10400 = ((~II10402))|((~II10403));
assign WX8732 = ((~WX8663));
assign II22671 = ((~WX7216))|((~II22663));
assign WX8951 = ((~WX8950));
assign WX4238 = ((~WX4882));
assign II22579 = ((~WX7210))|((~II22578));
assign II18086 = ((~WX5949))|((~II18085));
assign WX10858 = (WX10861&RESET);
assign II10843 = ((~WX3349))|((~II10842));
assign II2940 = ((~II2916))|((~II2932));
assign II14374 = ((~II14376))|((~II14377));
assign WX2021 = (WX1958&RESET);
assign II30983 = ((~II30985))|((~II30986));
assign II26264 = ((~II26274))|((~II26275));
assign WX8157 = (WX8168&WX8761);
assign WX9634 = ((~WX9602));
assign WX8357 = ((~WX8325));
assign WX6221 = (WX6220&WX6177);
assign II31180 = ((~WX9550))|((~II31178));
assign WX5486 = ((~WX5485));
assign WX5904 = (WX5841&RESET);
assign WX3528 = ((~WX3507));
assign II18621 = ((~II18611))|((~II18619));
assign WX3198 = ((~WX3423));
assign WX4397 = (WX4400&RESET);
assign WX2023 = (WX1960&RESET);
assign WX3495 = ((~II10300))|((~II10301));
assign II23417 = ((~WX7002))|((~II23415));
assign WX6544 = ((~WX7468));
assign II10031 = ((~WX3233))|((~II10029));
assign II18627 = ((~II18629))|((~II18630));
assign II11389 = ((~WX3121))|((~II11387));
assign II2827 = ((~WX699))|((~II2825));
assign II7514 = ((~II7504))|((~II7512));
assign WX4482 = ((~WX4450));
assign WX11560 = ((~II35483))|((~II35484));
assign WX9409 = (WX9415&WX9410);
assign WX5028 = ((~WX4884));
assign WX4195 = (WX4201&WX4196);
assign II14235 = ((~WX4666))|((~WX4730));
assign II7668 = ((~_2117_))|((~II7666));
assign WX9162 = ((~WX10055));
assign WX1065 = ((~WX1005));
assign II22757 = ((~WX7467))|((~WX7158));
assign WX7899 = (WX8257&WX8762);
assign WX6778 = ((~WX6769));
assign II3577 = ((~WX620))|((~_2099_));
assign WX3350 = (WX3287&RESET);
assign II26786 = ((~II26776))|((~II26784));
assign II26088 = ((~WX8471))|((~II26087));
assign II14561 = ((~WX4881))|((~WX4560));
assign II6877 = ((~WX2122))|((~II6876));
assign II30256 = ((~WX9838))|((~II30255));
assign WX123 = (_2102_&WX1004);
assign II34259 = ((~II34261))|((~II34262));
assign II10620 = ((~WX3271))|((~II10618));
assign II6890 = ((~II6900))|((~II6901));
assign WX5267 = (_2232_&WX6176);
assign II18612 = ((~WX5983))|((~WX6047));
assign WX10612 = (WX11468&WX10613);
assign WX9637 = ((~WX9605));
assign WX9620 = ((~WX9994));
assign II19535 = ((~WX5815))|((~II19534));
assign II14778 = ((~WX4881))|((~WX4574));
assign WX1715 = (WX2494&WX1716);
assign II6287 = ((~WX2084))|((~WX2148));
assign WX6228 = (WX6227&WX6177);
assign WX1610 = ((~WX2296));
assign II30697 = ((~II30672))|((~II30696));
assign WX9384 = (_2311_&WX10055);
assign II34309 = ((~WX11007))|((~II34307));
assign II18139 = ((~WX5889))|((~II18131));
assign II6551 = ((~WX2295))|((~WX1974));
assign WX5125 = ((~II15614))|((~II15615));
assign WX10034 = ((~WX10033));
assign WX8071 = ((~WX8062));
assign WX6882 = (_2241_&WX7469);
assign II2080 = ((~II2082))|((~II2083));
assign WX159 = ((~WX150));
assign WX6522 = (WX6952&WX7469);
assign WX1259 = ((~II3690))|((~II3691));
assign WX8102 = (WX8108&WX8103);
assign II35105 = ((~WX10925))|((~WX10831));
assign II31490 = ((~WX9662))|((~WX9598));
assign II10533 = ((~WX3329))|((~II10532));
assign WX9359 = (WX9357)|(WX9356);
assign II14546 = ((~WX4686))|((~II14545));
assign II30975 = ((~II30951))|((~II30967));
assign WX9233 = (WX9231)|(WX9230);
assign II7498 = ((~_2119_))|((~II7497));
assign II30572 = ((~II30548))|((~II30564));
assign II14249 = ((~II14259))|((~II14260));
assign WX7718 = ((~II23673))|((~II23674));
assign WX8775 = (WX8773)|(WX8772);
assign WX4605 = (WX4542&RESET);
assign II30269 = ((~II30279))|((~II30280));
assign II3669 = ((~WX635))|((~II3668));
assign II19307 = ((~WX5770))|((~II19306));
assign II18642 = ((~II18644))|((~II18645));
assign WX6937 = (WX6935)|(WX6934);
assign WX1461 = (WX1459)|(WX1458);
assign II6614 = ((~WX2295))|((~II6613));
assign WX10036 = ((~WX10035));
assign WX8316 = ((~WX8743));
assign WX8122 = (WX8120)|(WX8119);
assign WX1128 = ((~WX1005));
assign WX9267 = ((~WX9266));
assign WX1672 = (WX1826&WX2297);
assign II34912 = ((~WX11173))|((~II34911));
assign WX195 = ((~WX1004));
assign II18906 = ((~II18908))|((~II18909));
assign WX11397 = ((~WX11396));
assign II6101 = ((~WX2072))|((~WX2136));
assign WX6824 = ((~WX7468));
assign WX9964 = ((~II30449))|((~II30450));
assign WX3260 = (WX2844&RESET);
assign WX788 = (WX725&RESET);
assign WX9827 = (WX9764&RESET);
assign WX5235 = (WX5246&WX6175);
assign II34546 = ((~II34522))|((~II34538));
assign WX10674 = (WX10680&WX10675);
assign II30613 = ((~WX10053))|((~II30612));
assign II14880 = ((~II14870))|((~II14878));
assign WX5613 = (WX5624&WX6175);
assign WX949 = ((~WX948));
assign WX7787 = (WX7702&WX7728);
assign WX2337 = ((~WX2298));
assign WX2425 = ((~II7292))|((~II7293));
assign WX9279 = (WX9277)|(WX9276);
assign WX3505 = ((~II10610))|((~II10611));
assign WX4434 = ((~WX4858));
assign WX10393 = (WX10404&WX11347);
assign WX2667 = (_2169_&WX3590);
assign WX7935 = ((~WX8761));
assign WX770 = (WX707&RESET);
assign II23235 = ((~WX6974))|((~II23233));
assign II14887 = ((~WX4708))|((~II14886));
assign WX8307 = ((~WX8725));
assign WX8842 = (WX8841&WX8763);
assign WX8217 = (_2270_&WX8762);
assign WX9530 = ((~WX10055));
assign WX5944 = (WX5881&RESET);
assign WX128 = (DATA_9_25&WX129);
assign WX1099 = (WX593&WX1100);
assign II26863 = ((~WX8521))|((~II26862));
assign II19476 = ((~WX5783))|((~II19475));
assign WX2242 = ((~WX2241));
assign II19576 = ((~WX5789))|((~_2230_));
assign WX8486 = (WX8423&RESET);
assign II26683 = ((~II26685))|((~II26686));
assign WX7963 = ((~WX8761));
assign II30999 = ((~WX9886))|((~WX9950));
assign WX4889 = (WX4887)|(WX4886);
assign WX8201 = ((~WX8761));
assign II15501 = ((~WX4511))|((~II15500));
assign II14917 = ((~WX4710))|((~WX4774));
assign II22259 = ((~II22269))|((~II22270));
assign II15471 = ((~WX4490))|((~II15470));
assign WX8560 = (WX8497&RESET);
assign WX4950 = (WX4468&WX4951);
assign WX4908 = (WX4462&WX4909);
assign WX4291 = ((~WX4290));
assign WX8037 = ((~WX8762));
assign WX5781 = ((~WX5749));
assign WX3890 = (WX3832&WX3849);
assign II10465 = ((~WX3261))|((~II10463));
assign WX203 = (WX214&WX1003);
assign II6837 = ((~WX2056))|((~II6829));
assign WX5155 = (WX5137&WX5142);
assign II30124 = ((~WX9766))|((~II30123));
assign WX10484 = (WX10482)|(WX10481);
assign II2485 = ((~WX1002))|((~II2484));
assign WX441 = (WX452&WX1003);
assign II30682 = ((~WX9802))|((~II30681));
assign WX419 = ((~WX1004));
assign II30689 = ((~WX9866))|((~WX9930));
assign WX9308 = ((~WX9299));
assign WX6942 = (WX7012&WX7469);
assign WX5888 = (WX5825&RESET);
assign WX3106 = (WX3109&RESET);
assign WX10115 = (WX9639&WX10116);
assign WX10438 = (WX10436)|(WX10435);
assign WX7672 = ((~WX7671));
assign II11336 = ((~WX3187))|((~II11335));
assign WX5099 = (WX5097)|(WX5096);
assign WX764 = (WX701&RESET);
assign WX1884 = ((~WX1852));
assign II18620 = ((~II18595))|((~II18619));
assign II35354 = ((~WX10869))|((~II35352));
assign WX8078 = (WX10203&WX8079);
assign II22905 = ((~II22895))|((~II22903));
assign WX2003 = (WX1940&RESET);
assign II23078 = ((~WX7045))|((~II23077));
assign WX652 = (WX104&RESET);
assign WX2277 = ((~WX2203));
assign WX10598 = (WX11461&WX10599);
assign WX2700 = (WX3633&WX2701);
assign II23603 = ((~WX7085))|((~II23602));
assign WX2513 = (WX2511)|(WX2510);
assign II34717 = ((~WX11097))|((~II34709));
assign WX8834 = ((~II27213))|((~II27214));
assign II10275 = ((~II10285))|((~II10286));
assign WX5298 = (WX5296)|(WX5295);
assign WX5090 = (WX4488&WX5091);
assign WX7133 = (WX6681&RESET);
assign WX1233 = ((~II3508))|((~II3509));
assign WX3726 = (WX3725&WX3591);
assign WX11324 = ((~WX11252));
assign II10012 = ((~II10014))|((~II10015));
assign II31619 = ((~WX9672))|((~_2322_));
assign II30138 = ((~II30114))|((~II30130));
assign II15276 = ((~WX4475))|((~II15275));
assign II18225 = ((~WX6173))|((~WX5831));
assign WX6908 = ((~WX7468));
assign WX8683 = ((~II26816))|((~II26817));
assign WX6532 = (_2266_&WX7469);
assign WX8114 = ((~WX8113));
assign WX9375 = (WX10203&WX9376);
assign WX10289 = ((~II31578))|((~II31579));
assign WX2244 = ((~WX2243));
assign II10756 = ((~II10758))|((~II10759));
assign WX8888 = ((~WX8887));
assign WX169 = (WX503&WX1004);
assign WX4725 = (WX4662&RESET);
assign WX11186 = (WX11123&RESET);
assign II30084 = ((~II30086))|((~II30087));
assign WX3970 = (WX3981&WX4882);
assign WX1636 = (WX1647&WX2296);
assign WX1039 = ((~WX1038));
assign WX6554 = ((~WX6545));
assign WX5358 = (WX5356)|(WX5355);
assign WX11208 = (WX11145&RESET);
assign II26483 = ((~WX8759))|((~WX8433));
assign II6475 = ((~WX2160))|((~II6473));
assign II14118 = ((~II14094))|((~II14110));
assign WX8663 = ((~II26196))|((~II26197));
assign WX9729 = (WX9337&RESET);
assign WX2989 = (_2146_&WX3590);
assign II22486 = ((~WX7204))|((~II22485));
assign WX1157 = (WX1155)|(WX1154);
assign WX11447 = ((~WX11446));
assign WX6587 = (WX6585)|(WX6584);
assign II30877 = ((~WX9942))|((~II30875));
assign II31633 = ((~WX9674))|((~_2320_));
assign II10037 = ((~WX3297))|((~II10036));
assign WX878 = (WX815&RESET);
assign II34648 = ((~WX11346))|((~WX11029));
assign WX9303 = (WX9301)|(WX9300);
assign WX8786 = (WX8785&WX8763);
assign WX6290 = ((~II19281))|((~II19282));
assign II22750 = ((~II22740))|((~II22748));
assign WX3740 = (WX3739&WX3591);
assign WX10020 = ((~WX10019));
assign WX5315 = ((~WX6176));
assign II2578 = ((~WX1002))|((~II2577));
assign WX6571 = (WX6577&WX6572);
assign WX5583 = ((~WX5574));
assign WX11261 = ((~II34578))|((~II34579));
assign II30774 = ((~WX9808))|((~II30766));
assign II7568 = ((~WX1911))|((~_2133_));
assign II30108 = ((~II30083))|((~II30107));
assign WX4087 = (WX6268&WX4088);
assign WX3018 = (WX5087&WX3019);
assign WX10940 = ((~WX10908));
assign WX9401 = (WX9399)|(WX9398);
assign WX2549 = ((~II7674))|((~II7675));
assign WX1724 = (_2112_&WX2297);
assign WX2623 = ((~WX3589));
assign WX10058 = (WX10057&WX10056);
assign WX7900 = (WX8819&WX7901);
assign II34633 = ((~WX11155))|((~II34632));
assign WX6124 = ((~WX6098));
assign WX3179 = ((~WX3147));
assign II26104 = ((~II26094))|((~II26102));
assign II26971 = ((~II26946))|((~II26970));
assign WX6578 = (WX6960&WX7469);
assign WX438 = (WX436)|(WX435);
assign WX2840 = (WX3703&WX2841);
assign II14508 = ((~II14498))|((~II14506));
assign WX11446 = ((~WX11445));
assign II22073 = ((~II22083))|((~II22084));
assign WX7781 = (WX7705&WX7728);
assign WX4305 = ((~WX4304));
assign WX6793 = ((~WX6792));
assign II14879 = ((~WX4644))|((~II14878));
assign WX2540 = ((~II7611))|((~II7612));
assign II11540 = ((~_2170_))|((~II11538));
assign II2606 = ((~II2616))|((~II2617));
assign II31725 = ((~WX9689))|((~II31724));
assign II2741 = ((~II2731))|((~II2739));
assign WX3600 = (WX3599&WX3591);
assign II30100 = ((~WX9828))|((~WX9892));
assign II2663 = ((~II2653))|((~II2661));
assign II34810 = ((~WX11103))|((~II34802));
assign II19521 = ((~WX5811))|((~II19520));
assign II10503 = ((~II10493))|((~II10501));
assign II6271 = ((~II6273))|((~II6274));
assign WX7999 = ((~WX8762));
assign WX10062 = ((~WX10061));
assign WX3583 = ((~TM0));
assign II10682 = ((~WX3275))|((~II10680));
assign WX1859 = ((~WX2230));
assign II23638 = ((~WX7090))|((~II23637));
assign WX9541 = (WX9544&RESET);
assign WX6630 = (_2259_&WX7469);
assign II14499 = ((~WX4881))|((~WX4556));
assign II11610 = ((~_2160_))|((~II11608));
assign WX11620 = (WX11602&WX11607);
assign II6056 = ((~WX2294))|((~II6055));
assign WX3738 = ((~WX3737));
assign WX3262 = (WX2858&RESET);
assign WX3140 = ((~WX3563));
assign WX9759 = (WX9696&RESET);
assign II22252 = ((~II22228))|((~II22244));
assign WX3470 = (WX3407&RESET);
assign WX2859 = (WX2870&WX3589);
assign WX2331 = (WX2329)|(WX2328);
assign WX6261 = ((~WX6260));
assign II34710 = ((~WX11346))|((~WX11033));
assign II15621 = ((~WX4503))|((~II15620));
assign WX9420 = ((~WX9411));
assign WX7327 = (WX7264&RESET);
assign WX4927 = ((~II15146))|((~II15147));
assign WX4165 = ((~WX4164));
assign WX5434 = (WX5432)|(WX5431);
assign II30262 = ((~II30238))|((~II30254));
assign II10743 = ((~WX3588))|((~II10742));
assign WX6691 = (WX7568&WX6692);
assign WX2133 = (WX2070&RESET);
assign II14335 = ((~II14311))|((~II14327));
assign WX9629 = ((~WX10012));
assign II19585 = ((~_2229_))|((~II19583));
assign II18689 = ((~II18691))|((~II18692));
assign II6591 = ((~II6581))|((~II6589));
assign WX2205 = ((~II6388))|((~II6389));
assign WX1767 = (WX3815&WX1768);
assign WX10359 = (WX10295&WX10314);
assign WX6655 = (WX6661&WX6656);
assign WX3643 = (WX3173&WX3644);
assign WX5780 = ((~WX5748));
assign WX9585 = (WX9588&RESET);
assign WX1417 = (WX3640&WX1418);
assign II22881 = ((~WX7467))|((~WX7166));
assign II6048 = ((~II6038))|((~II6046));
assign WX5216 = (WX6184&WX5217);
assign WX1090 = ((~II3209))|((~II3210));
assign II26655 = ((~WX8635))|((~II26653));
assign II10424 = ((~II10399))|((~II10423));
assign II15492 = ((~_2188_))|((~II15484));
assign II10734 = ((~II10709))|((~II10733));
assign II10082 = ((~II10058))|((~II10074));
assign WX6297 = ((~II19294))|((~II19295));
assign WX11468 = ((~WX11467));
assign WX6401 = ((~WX6400));
assign II2677 = ((~WX753))|((~II2669));
assign WX1957 = (WX1481&RESET);
assign WX4018 = ((~WX4883));
assign II6797 = ((~II6807))|((~II6808));
assign WX8921 = ((~WX8763));
assign II22952 = ((~II22942))|((~II22950));
assign WX3695 = ((~WX3694));
assign II30481 = ((~II30471))|((~II30479));
assign II10387 = ((~WX3447))|((~II10385));
assign II35582 = ((~WX10959))|((~_2360_));
assign II30223 = ((~II30225))|((~II30226));
assign II23597 = ((~_2260_))|((~II23595));
assign WX9066 = (WX9002&WX9021);
assign WX4038 = ((~WX4029));
assign II35532 = ((~_2343_))|((~II35524));
assign WX11094 = (WX11031&RESET);
assign WX5514 = ((~WX5513));
assign II7535 = ((~_2138_))|((~II7533));
assign WX7693 = ((~WX7692));
assign WX4617 = (WX4554&RESET);
assign WX2507 = ((~WX2506));
assign WX11487 = (WX11485)|(WX11484);
assign WX984 = ((~WX910));
assign II10811 = ((~WX3347))|((~II10803));
assign WX5207 = (WX5218&WX6175);
assign WX7056 = ((~WX7024));
assign WX6201 = (WX5755&WX6202);
assign WX7535 = (WX7534&WX7470);
assign II19189 = ((~WX5761))|((~WX5675));
assign WX412 = ((~WX411));
assign WX11597 = ((~II35688))|((~II35689));
assign WX247 = ((~WX1003));
assign WX10677 = (_2343_&WX11348);
assign WX10984 = ((~WX11237));
assign WX10870 = (WX10873&RESET);
assign WX5385 = ((~WX6176));
assign WX2808 = (WX4982&WX2809);
assign WX11232 = (WX11169&RESET);
assign II18675 = ((~WX5987))|((~II18674));
assign II30758 = ((~II30734))|((~II30750));
assign II6336 = ((~WX1960))|((~II6334));
assign WX356 = ((~WX355));
assign II22238 = ((~WX7188))|((~II22237));
assign II2423 = ((~WX1001))|((~II2422));
assign WX4261 = (WX4259)|(WX4258);
assign II31127 = ((~WX9634))|((~II31126));
assign II7624 = ((~WX1919))|((~_2125_));
assign II6181 = ((~WX1950))|((~II6179));
assign WX3152 = ((~WX3523));
assign WX4876 = ((~TM0));
assign WX5025 = ((~II15328))|((~II15329));
assign II26738 = ((~WX8513))|((~II26730));
assign WX11588 = ((~II35625))|((~II35626));
assign WX4222 = (WX4233&WX4882);
assign WX10866 = (WX10869&RESET);
assign II14390 = ((~WX4676))|((~WX4740));
assign II22663 = ((~II22665))|((~II22666));
assign WX2347 = ((~WX2346));
assign WX8984 = ((~WX8763));
assign II22153 = ((~WX7246))|((~II22152));
assign II11526 = ((~_2172_))|((~II11524));
assign II2081 = ((~WX1001))|((~WX651));
assign WX7454 = ((~WX7453));
assign II34588 = ((~WX11025))|((~II34586));
assign WX5054 = (WX5053&WX4884);
assign II22944 = ((~WX7467))|((~II22943));
assign WX11018 = (WX10602&RESET);
assign WX2980 = (WX3773&WX2981);
assign WX7994 = (WX10161&WX7995);
assign WX6010 = (WX5947&RESET);
assign WX3771 = (WX3769)|(WX3768);
assign II34781 = ((~II34771))|((~II34779));
assign WX9133 = (WX11377&WX9134);
assign WX7741 = (WX7723&WX7728);
assign WX2599 = (WX2538&WX2556);
assign II19591 = ((~WX5791))|((~II19590));
assign II18566 = ((~WX6174))|((~WX5853));
assign WX6858 = (WX7000&WX7469);
assign DATA_9_23 = ((~WX1067));
assign II34137 = ((~WX11123))|((~II34136));
assign WX6032 = (WX5969&RESET);
assign WX1819 = (WX1822&RESET);
assign II30876 = ((~WX9878))|((~II30875));
assign WX6890 = ((~WX6881));
assign II34864 = ((~II34866))|((~II34867));
assign WX864 = (WX801&RESET);
assign WX3587 = ((~WX3586));
assign II15606 = ((~WX4501))|((~_2193_));
assign WX8002 = ((~WX8001));
assign WX2256 = ((~WX2255));
assign II10417 = ((~WX3385))|((~II10416));
assign WX460 = (WX2515&WX461);
assign WX10783 = ((~WX10774));
assign WX7563 = (WX7562&WX7470);
assign WX1746 = ((~WX1737));
assign WX2479 = ((~WX2478));
assign WX11378 = ((~II35145))|((~II35146));
assign WX7518 = ((~WX7517));
assign II6722 = ((~WX2112))|((~II6721));
assign WX4229 = (WX4227)|(WX4226);
assign WX110 = (WX2340&WX111);
assign II2609 = ((~WX1002))|((~II2608));
assign WX1220 = (WX1218)|(WX1217);
assign WX7115 = (WX6555&RESET);
assign WX1878 = ((~WX1846));
assign II35618 = ((~WX10964))|((~II35617));
assign WX2875 = ((~WX3589));
assign II22556 = ((~WX7272))|((~II22555));
assign WX9957 = ((~II30232))|((~II30233));
assign WX7367 = ((~II22098))|((~II22099));
assign WX3025 = ((~WX3016));
assign WX2783 = (WX3093&WX3590);
assign WX2490 = (WX1900&WX2491);
assign II6317 = ((~II6319))|((~II6320));
assign WX8375 = ((~WX8605));
assign II35673 = ((~WX10973))|((~_2346_));
assign II15684 = ((~WX4514))|((~II15683));
assign WX7771 = (WX7710&WX7728);
assign II18304 = ((~WX6027))|((~II18302));
assign WX11102 = (WX11039&RESET);
assign II6274 = ((~WX1956))|((~II6272));
assign WX5277 = (WX5288&WX6175);
assign WX9809 = (WX9746&RESET);
assign II30564 = ((~II30566))|((~II30567));
assign WX11660 = (WX11584&WX11607);
assign WX8356 = ((~WX8324));
assign WX2183 = (WX2120&RESET);
assign WX5258 = (WX6205&WX5259);
assign WX4942 = (WX4941&WX4884);
assign WX5928 = (WX5865&RESET);
assign II22998 = ((~II22988))|((~II22996));
assign II6559 = ((~WX2038))|((~II6558));
assign WX222 = (WX2396&WX223);
assign II15727 = ((~_2173_))|((~II15725));
assign II6729 = ((~II6704))|((~II6728));
assign II31655 = ((~WX9677))|((~II31654));
assign II2702 = ((~WX1002))|((~II2701));
assign WX189 = (WX200&WX1003);
assign II35326 = ((~WX10942))|((~WX10865));
assign WX7759 = (WX7715&WX7728);
assign WX3708 = (WX3706)|(WX3705);
assign II34881 = ((~WX11171))|((~II34880));
assign II3184 = ((~WX505))|((~II3182));
assign II34898 = ((~WX11045))|((~II34896));
assign WX5222 = (WX5228&WX5223);
assign WX6452 = (WX6428&WX6435);
assign II26125 = ((~II26127))|((~II26128));
assign II11075 = ((~WX3167))|((~WX3073));
assign II18320 = ((~WX5837))|((~II18318));
assign II10393 = ((~II10368))|((~II10392));
assign II6115 = ((~II6125))|((~II6126));
assign WX11436 = (WX10936&WX11437);
assign WX6634 = (WX6968&WX7469);
assign WX3769 = (WX3191&WX3770);
assign WX4705 = (WX4642&RESET);
assign II14608 = ((~WX4690))|((~II14607));
assign II14081 = ((~WX4656))|((~II14080));
assign WX5535 = ((~WX6176));
assign II6945 = ((~II6921))|((~II6937));
assign II6612 = ((~II6614))|((~II6615));
assign WX8136 = (WX8134)|(WX8133);
assign II26140 = ((~II26150))|((~II26151));
assign WX8134 = (WX10231&WX8135);
assign WX7101 = ((~WX7350));
assign II15593 = ((~WX4499))|((~II15592));
assign WX1432 = ((~WX2297));
assign WX2755 = (WX3089&WX3590);
assign WX1186 = ((~WX1185));
assign II27239 = ((~WX8350))|((~II27238));
assign II7596 = ((~WX1915))|((~_2129_));
assign II18118 = ((~WX6015))|((~II18116));
assign II3551 = ((~_2103_))|((~II3549));
assign WX333 = (_2087_&WX1004);
assign WX219 = ((~WX1003));
assign II6930 = ((~WX2062))|((~II6922));
assign WX182 = (WX180)|(WX179);
assign WX9781 = (WX9718&RESET);
assign II2841 = ((~WX827))|((~II2840));
assign II3710 = ((~WX642))|((~_2077_));
assign WX9437 = (WX9443&WX9438);
assign WX8386 = ((~WX8627));
assign II27095 = ((~WX8339))|((~WX8245));
assign WX10139 = ((~WX10138));
assign WX8747 = ((~WX8746));
assign II22827 = ((~WX7226))|((~II22826));
assign WX2395 = ((~WX2394));
assign II22253 = ((~II22228))|((~II22252));
assign WX5761 = ((~WX5729));
assign II22834 = ((~WX7290))|((~WX7354));
assign WX10465 = ((~WX11347));
assign WX9677 = ((~WX9916));
assign WX10069 = ((~WX10068));
assign WX4126 = ((~WX4882));
assign WX3904 = (WX3825&WX3849);
assign II35729 = ((~WX10982))|((~_2337_));
assign II22619 = ((~WX7340))|((~II22617));
assign II6435 = ((~WX2030))|((~II6434));
assign II19562 = ((~WX5787))|((~_2232_));
assign WX10087 = (WX9635&WX10088);
assign II10828 = ((~II10818))|((~II10826));
assign WX1376 = ((~WX2297));
assign II27227 = ((~WX8265))|((~II27225));
assign WX7229 = (WX7166&RESET);
assign WX3677 = (WX3676&WX3591);
assign WX6322 = (WX6320)|(WX6319);
assign WX7614 = ((~WX7470));
assign WX6287 = (WX6285)|(WX6284);
assign WX6307 = ((~WX6177));
assign II9998 = ((~WX3587))|((~WX3231));
assign WX5447 = ((~WX6175));
assign WX9511 = (WX11566&WX9512);
assign WX1856 = ((~WX2288));
assign WX9521 = (WX9527&WX9522);
assign II2731 = ((~II2733))|((~II2734));
assign WX8167 = ((~WX8762));
assign II34130 = ((~II34120))|((~II34128));
assign WX2354 = ((~WX2353));
assign WX9211 = ((~WX9210));
assign II30231 = ((~II30207))|((~II30223));
assign II15185 = ((~WX4468))|((~II15184));
assign II7176 = ((~WX1796))|((~II7174));
assign WX5138 = ((~II15705))|((~II15706));
assign II6193 = ((~II6195))|((~II6196));
assign II2903 = ((~WX831))|((~II2902));
assign WX2470 = ((~WX2298));
assign WX2203 = ((~II6326))|((~II6327));
assign II6170 = ((~II6146))|((~II6162));
assign WX78 = (WX84&WX79);
assign WX11503 = ((~WX11502));
assign II22159 = ((~II22135))|((~II22151));
assign WX716 = (WX653&RESET);
assign WX6840 = (_2244_&WX7469);
assign II26319 = ((~II26295))|((~II26311));
assign WX10267 = ((~II31478))|((~II31479));
assign II34694 = ((~WX11159))|((~WX11223));
assign II34114 = ((~II34104))|((~II34112));
assign WX1741 = (WX1739)|(WX1738);
assign WX588 = ((~WX556));
assign WX5253 = (_2233_&WX6176);
assign WX322 = (WX320)|(WX319);
assign WX6766 = (WX6777&WX7468);
assign II26794 = ((~WX8760))|((~II26793));
assign WX1203 = (WX1202&WX1005);
assign WX7588 = ((~WX7587));
assign WX11654 = (WX11587&WX11607);
assign WX3828 = ((~II11581))|((~II11582));
assign WX3758 = ((~WX3757));
assign WX2443 = (WX2441)|(WX2440);
assign WX6871 = (WX6869)|(WX6868);
assign WX7737 = (WX7698&WX7728);
assign WX4448 = ((~WX4822));
assign II2532 = ((~WX871))|((~II2530));
assign II2237 = ((~WX1001))|((~II2236));
assign WX3952 = ((~WX4883));
assign WX1871 = ((~WX2254));
assign WX7926 = (WX7924)|(WX7923);
assign WX1151 = ((~WX1150));
assign WX2872 = ((~WX2871));
assign WX6417 = ((~II19612))|((~II19613));
assign WX5309 = (_2229_&WX6176);
assign WX5399 = ((~WX6176));
assign II3092 = ((~WX583))|((~II3091));
assign WX9549 = (WX9552&RESET);
assign II23526 = ((~WX7104))|((~II23525));
assign WX10253 = ((~II31452))|((~II31453));
assign WX7257 = (WX7194&RESET);
assign II19703 = ((~WX5809))|((~II19702));
assign II18161 = ((~II18171))|((~II18172));
assign II6131 = ((~II6133))|((~II6134));
assign WX2171 = (WX2108&RESET);
assign WX2416 = ((~WX2415));
assign WX2960 = (WX2958)|(WX2957);
assign WX10581 = ((~WX11348));
assign II11608 = ((~WX3209))|((~_2160_));
assign WX1043 = (WX585&WX1044);
assign WX1690 = ((~WX1681));
assign WX8798 = ((~WX8797));
assign WX8225 = ((~WX8216));
assign II35145 = ((~WX10928))|((~II35144));
assign II2765 = ((~WX695))|((~II2763));
assign II30913 = ((~II30889))|((~II30905));
assign II7358 = ((~WX1824))|((~II7356));
assign WX10249 = ((~WX10056));
assign WX8098 = (WX8096)|(WX8095);
assign WX2977 = ((~WX3590));
assign II31414 = ((~WX9586))|((~II31412));
assign II18394 = ((~II18396))|((~II18397));
assign II26605 = ((~II26615))|((~II26616));
assign II26150 = ((~WX8475))|((~II26149));
assign WX7952 = (WX10140&WX7953);
assign II35198 = ((~WX10845))|((~II35196));
assign II19606 = ((~_2226_))|((~II19604));
assign II14764 = ((~WX4764))|((~II14762));
assign WX1241 = ((~II3564))|((~II3565));
assign WX6803 = (WX7624&WX6804);
assign II30023 = ((~WX10052))|((~WX9696));
assign WX9204 = ((~WX10055));
assign II18053 = ((~II18055))|((~II18056));
assign WX8109 = (WX8287&WX8762);
assign WX9990 = ((~WX9989));
assign II34516 = ((~II34491))|((~II34515));
assign WX571 = ((~WX947));
assign II23130 = ((~WX7049))|((~II23129));
assign WX9141 = ((~WX9140));
assign II14988 = ((~II14978))|((~II14986));
assign II10377 = ((~WX3319))|((~II10369));
assign WX9330 = ((~WX10055));
assign II22996 = ((~II22972))|((~II22988));
assign II14809 = ((~WX4881))|((~WX4576));
assign WX8426 = (WX7974&RESET);
assign WX9245 = (WX11433&WX9246);
assign WX283 = ((~WX1004));
assign II35457 = ((~WX10952))|((~II35456));
assign II31620 = ((~WX9672))|((~II31619));
assign II35731 = ((~_2337_))|((~II35729));
assign WX448 = (WX446)|(WX445);
assign WX8770 = ((~WX8769));
assign WX4815 = ((~WX4797));
assign II7135 = ((~WX1879))|((~WX1790));
assign WX7836 = (WX7842&WX7837);
assign WX1979 = (WX1635&RESET);
assign WX4137 = ((~WX4136));
assign II35596 = ((~WX10961))|((~_2358_));
assign II31100 = ((~WX9632))|((~WX9538));
assign II18854 = ((~II18844))|((~II18852));
assign WX10939 = ((~WX10907));
assign WX7235 = (WX7172&RESET);
assign WX7119 = (WX6583&RESET);
assign WX2318 = ((~WX2317));
assign II6955 = ((~WX2295))|((~II6954));
assign II2058 = ((~WX713))|((~II2057));
assign WX8091 = (_2279_&WX8762);
assign WX1517 = (WX1515)|(WX1514);
assign II18845 = ((~WX6174))|((~WX5871));
assign WX10819 = ((~WX11348));
assign II34949 = ((~II34925))|((~II34941));
assign WX10258 = ((~WX10257));
assign II3499 = ((~II3501))|((~II3502));
assign WX298 = (WX296)|(WX295);
assign WX6713 = (WX6711)|(WX6710);
assign WX4835 = ((~WX4807));
assign II26870 = ((~WX8585))|((~WX8649));
assign WX1983 = (WX1663&RESET);
assign II23338 = ((~WX7065))|((~II23337));
assign WX1250 = ((~II3627))|((~II3628));
assign WX1726 = ((~WX2297));
assign II35639 = ((~WX10967))|((~II35638));
assign II19243 = ((~WX5683))|((~II19241));
assign WX1600 = ((~WX2297));
assign WX3448 = (WX3385&RESET);
assign WX8877 = (WX8876&WX8763);
assign WX11322 = ((~WX11251));
assign II3621 = ((~_2093_))|((~II3619));
assign WX5754 = ((~WX5722));
assign II34321 = ((~II34323))|((~II34324));
assign WX8828 = (WX8827&WX8763);
assign WX3988 = (_2199_&WX4883);
assign WX9270 = ((~WX10054));
assign WX231 = (WX242&WX1003);
assign WX2386 = ((~WX2298));
assign WX3218 = ((~WX3463));
assign WX3729 = (WX3727)|(WX3726);
assign WX4822 = ((~WX4821));
assign II27355 = ((~WX8359))|((~WX8285));
assign II23723 = ((~_2239_))|((~II23721));
assign II22594 = ((~II22569))|((~II22593));
assign II14181 = ((~II14156))|((~II14180));
assign II26171 = ((~II26181))|((~II26182));
assign II14066 = ((~WX4880))|((~II14065));
assign WX2371 = (WX1883&WX2372);
assign WX8233 = ((~WX8762));
assign WX8186 = (WX8192&WX8187);
assign II19569 = ((~WX5788))|((~_2231_));
assign WX5722 = ((~WX6141));
assign II23194 = ((~WX7054))|((~WX6968));
assign II14125 = ((~II14135))|((~II14136));
assign II7292 = ((~WX1891))|((~II7291));
assign WX5132 = ((~II15663))|((~II15664));
assign WX4475 = ((~WX4443));
assign II10434 = ((~WX3259))|((~II10432));
assign II30202 = ((~II30192))|((~II30200));
assign WX8708 = ((~WX8683));
assign II26020 = ((~WX8403))|((~II26018));
assign WX10918 = ((~WX11297));
assign WX9601 = ((~WX10020));
assign WX10156 = (WX10155&WX10056);
assign WX6752 = (WX6763&WX7468);
assign WX10647 = ((~WX11347));
assign WX1703 = (WX1701)|(WX1700);
assign WX7076 = ((~WX7044));
assign II10795 = ((~II10771))|((~II10787));
assign WX2330 = ((~WX2298));
assign WX9339 = (WX9345&WX9340);
assign WX5248 = ((~WX5247));
assign WX6864 = (WX6875&WX7468);
assign WX8758 = ((~TM1));
assign WX8659 = ((~II26072))|((~II26073));
assign WX1442 = ((~WX2296));
assign WX1115 = (WX1113)|(WX1112);
assign WX7239 = (WX7176&RESET);
assign II27665 = ((~_2282_))|((~II27663));
assign WX1037 = ((~WX1005));
assign WX955 = ((~WX954));
assign WX2652 = (WX2650)|(WX2649);
assign II2717 = ((~WX819))|((~II2716));
assign WX9528 = (WX9598&WX10055);
assign WX8911 = ((~II27356))|((~II27357));
assign WX6107 = ((~WX6106));
assign WX2816 = ((~WX2815));
assign II30845 = ((~WX9876))|((~II30844));
assign II18295 = ((~WX5899))|((~II18294));
assign WX5790 = ((~WX6021));
assign WX2498 = ((~WX2298));
assign WX4462 = ((~WX4430));
assign II30442 = ((~WX9850))|((~II30441));
assign WX4735 = (WX4672&RESET);
assign WX9188 = (_2325_&WX10055);
assign II18358 = ((~II18348))|((~II18356));
assign II30660 = ((~WX9928))|((~II30658));
assign II14274 = ((~II14249))|((~II14273));
assign WX9477 = ((~WX9476));
assign WX3674 = ((~WX3673));
assign WX7402 = ((~WX7401));
assign II34965 = ((~WX11113))|((~II34957));
assign II30409 = ((~II30411))|((~II30412));
assign WX2011 = (WX1948&RESET);
assign WX11002 = (WX10490&RESET);
assign II22200 = ((~WX7466))|((~II22199));
assign WX1913 = ((~WX2146));
assign II15692 = ((~_2179_))|((~II15690));
assign II14281 = ((~II14283))|((~II14284));
assign II6163 = ((~WX2076))|((~WX2140));
assign II10068 = ((~WX3299))|((~II10067));
assign II22361 = ((~WX7196))|((~II22353));
assign WX1423 = (WX1421)|(WX1420);
assign II22826 = ((~WX7226))|((~II22818));
assign II19138 = ((~WX5757))|((~II19137));
assign II10689 = ((~II10679))|((~II10687));
assign II22991 = ((~WX7364))|((~II22989));
assign II31704 = ((~WX9686))|((~II31703));
assign WX10834 = (WX10837&RESET);
assign II27278 = ((~WX8353))|((~II27277));
assign WX143 = ((~WX1004));
assign II6388 = ((~II6363))|((~II6387));
assign WX5478 = (WX7610&WX5479);
assign WX1656 = ((~WX2297));
assign WX9476 = ((~WX9467));
assign WX5990 = (WX5927&RESET);
assign II6258 = ((~WX2146))|((~II6256));
assign WX5804 = ((~WX6049));
assign II35632 = ((~WX10966))|((~II35631));
assign WX11418 = ((~WX11417));
assign WX9952 = ((~II30077))|((~II30078));
assign WX3938 = ((~WX4883));
assign II3626 = ((~WX628))|((~_2091_));
assign WX2741 = (WX3087&WX3590);
assign WX6216 = ((~WX6177));
assign II22268 = ((~WX7190))|((~II22260));
assign II26290 = ((~II26280))|((~II26288));
assign II14501 = ((~WX4556))|((~II14499));
assign II2910 = ((~II2885))|((~II2909));
assign WX6860 = ((~WX7469));
assign WX3609 = ((~WX3591));
assign II22780 = ((~II22755))|((~II22779));
assign WX8933 = (WX8932&WX8763);
assign WX2238 = ((~WX2237));
assign WX6673 = (WX8854&WX6674);
assign WX5469 = ((~WX6176));
assign II34145 = ((~II34135))|((~II34143));
assign WX8859 = (WX8857)|(WX8856);
assign WX10812 = ((~WX10811));
assign II23658 = ((~WX7094))|((~_2250_));
assign WX4079 = (WX4077)|(WX4076);
assign II23576 = ((~_2263_))|((~II23574));
assign WX7708 = ((~II23603))|((~II23604));
assign WX2567 = (WX2552&WX2556);
assign II22859 = ((~II22849))|((~II22857));
assign WX8856 = (WX8855&WX8763);
assign WX3211 = ((~WX3449));
assign II23616 = ((~WX7087))|((~_2257_));
assign WX2950 = (WX2948)|(WX2947);
assign WX9294 = ((~WX9285));
assign WX7498 = ((~WX7497));
assign WX9314 = (_2316_&WX10055);
assign II30078 = ((~II30068))|((~II30076));
assign II3275 = ((~WX519))|((~II3273));
assign WX1142 = ((~WX1005));
assign WX6771 = (WX8903&WX6772);
assign WX4641 = (WX4578&RESET);
assign WX1052 = (WX1050)|(WX1049);
assign II22053 = ((~II22043))|((~II22051));
assign II22678 = ((~II22680))|((~II22681));
assign WX3922 = (WX4364&WX4883);
assign WX10433 = ((~WX10424));
assign II35722 = ((~WX10981))|((~_2338_));
assign WX10098 = ((~WX10097));
assign II2003 = ((~WX773))|((~WX837));
assign WX3637 = ((~WX3591));
assign WX6834 = ((~WX6825));
assign WX1667 = (WX1665)|(WX1664);
assign II15172 = ((~WX4467))|((~II15171));
assign WX9468 = (_2305_&WX10055);
assign WX10920 = ((~WX11301));
assign II11116 = ((~WX3079))|((~II11114));
assign WX8762 = ((~WX8755));
assign WX9711 = (WX9211&RESET);
assign WX8679 = ((~II26692))|((~II26693));
assign II26405 = ((~WX8555))|((~WX8619));
assign II22913 = ((~WX7467))|((~II22912));
assign WX11048 = (WX10812&RESET);
assign II27607 = ((~WX8378))|((~_2291_));
assign II26640 = ((~WX8443))|((~II26638));
assign WX3941 = ((~WX3940));
assign WX10166 = (WX10164)|(WX10163);
assign WX4495 = ((~WX4724));
assign WX6105 = ((~WX6104));
assign WX10654 = (WX11489&WX10655);
assign WX7036 = ((~WX7412));
assign II26578 = ((~WX8439))|((~II26576));
assign II14655 = ((~WX4881))|((~II14654));
assign WX8936 = (WX8934)|(WX8933);
assign WX8719 = ((~WX8718));
assign II30827 = ((~II30837))|((~II30838));
assign II34734 = ((~II34724))|((~II34732));
assign II30796 = ((~II30806))|((~II30807));
assign WX3579 = ((~WX3578));
assign WX5226 = (WX7484&WX5227);
assign II15516 = ((~WX4518))|((~II15515));
assign WX9195 = (WX9193)|(WX9192);
assign II6405 = ((~II6395))|((~II6403));
assign II6373 = ((~WX2026))|((~II6372));
assign WX7857 = (WX8251&WX8762);
assign WX6683 = (WX6689&WX6684);
assign WX11265 = ((~II34702))|((~II34703));
assign II2856 = ((~WX1002))|((~WX701));
assign II10454 = ((~II10430))|((~II10446));
assign WX97 = ((~WX1004));
assign WX2723 = (_2165_&WX3590);
assign II26568 = ((~II26543))|((~II26567));
assign II26699 = ((~II26701))|((~II26702));
assign II22355 = ((~WX7466))|((~II22354));
assign WX1390 = ((~WX2297));
assign WX5740 = ((~WX6113));
assign WX10327 = (WX10309&WX10314);
assign WX9608 = ((~WX10034));
assign WX10878 = (WX10881&RESET);
assign WX1492 = ((~WX2297));
assign WX2381 = ((~WX2380));
assign WX9014 = ((~II27699))|((~II27700));
assign WX2865 = ((~WX3590));
assign WX54 = (WX2312&WX55);
assign II6604 = ((~II6580))|((~II6596));
assign WX4901 = (WX4461&WX4902);
assign WX2129 = (WX2066&RESET);
assign WX2893 = ((~WX3590));
assign II31006 = ((~II30982))|((~II30998));
assign WX968 = ((~WX902));
assign II10642 = ((~II10632))|((~II10640));
assign WX8711 = ((~WX8710));
assign WX4500 = ((~WX4734));
assign WX291 = (_2090_&WX1004);
assign WX11347 = ((~WX11343));
assign WX367 = ((~WX1004));
assign II19604 = ((~WX5793))|((~_2226_));
assign II26740 = ((~II26730))|((~II26738));
assign WX5421 = (_2221_&WX6176);
assign WX7221 = (WX7158&RESET);
assign II35624 = ((~WX10965))|((~_2354_));
assign II10780 = ((~WX3345))|((~II10772));
assign II2198 = ((~II2188))|((~II2196));
assign WX10927 = ((~WX10895));
assign II18938 = ((~WX6174))|((~WX5877));
assign WX424 = (WX422)|(WX421);
assign WX4177 = (WX4175)|(WX4174);
assign WX11304 = ((~WX11274));
assign II26639 = ((~WX8760))|((~II26638));
assign II11362 = ((~WX3189))|((~II11361));
assign II3065 = ((~WX581))|((~WX487));
assign WX4771 = (WX4708&RESET);
assign WX8721 = ((~WX8720));
assign II11466 = ((~WX3197))|((~II11465));
assign WX7799 = ((~WX8762));
assign II22370 = ((~WX7260))|((~II22369));
assign II2182 = ((~WX721))|((~II2181));
assign WX6472 = (WX6420&WX6435);
assign II22368 = ((~II22370))|((~II22371));
assign WX10143 = (WX9643&WX10144);
assign WX11495 = ((~WX11494));
assign II35709 = ((~WX10979))|((~II35708));
assign II31465 = ((~WX9660))|((~II31464));
assign WX60 = (WX58)|(WX57);
assign WX10604 = (WX10610&WX10605);
assign II30667 = ((~II30657))|((~II30665));
assign WX10207 = ((~WX10056));
assign WX5416 = ((~WX5415));
assign II23495 = ((~WX7092))|((~_2268_));
assign WX8674 = ((~II26537))|((~II26538));
assign II34601 = ((~WX11153))|((~WX11217));
assign WX10260 = ((~II31465))|((~II31466));
assign WX1169 = (WX603&WX1170);
assign II15536 = ((~WX4491))|((~_2203_));
assign WX1371 = (WX1377&WX1372);
assign WX8197 = ((~WX8188));
assign WX6989 = (WX6992&RESET);
assign II19506 = ((~WX5804))|((~II19505));
assign WX7581 = ((~WX7580));
assign WX5433 = ((~WX6175));
assign II2259 = ((~II2234))|((~II2258));
assign WX814 = (WX751&RESET);
assign WX2881 = (WX3107&WX3590);
assign II18433 = ((~II18409))|((~II18425));
assign WX351 = (WX529&WX1004);
assign II31598 = ((~WX9669))|((~_2325_));
assign II22306 = ((~II22308))|((~II22309));
assign WX7954 = (WX7952)|(WX7951);
assign II22363 = ((~II22353))|((~II22361));
assign II6243 = ((~WX1954))|((~II6241));
assign WX10231 = ((~WX10230));
assign WX4028 = ((~WX4882));
assign II18583 = ((~WX6045))|((~II18581));
assign II14904 = ((~WX4582))|((~II14902));
assign WX6154 = ((~WX6081));
assign WX640 = ((~WX893));
assign II6596 = ((~II6598))|((~II6599));
assign II10518 = ((~II10508))|((~II10516));
assign WX8003 = (WX8014&WX8761);
assign WX5747 = ((~WX6127));
assign WX8015 = ((~WX8006));
assign II34207 = ((~II34197))|((~II34205));
assign WX7917 = ((~WX7908));
assign II14322 = ((~II14312))|((~II14320));
assign WX3410 = (WX3347&RESET);
assign WX1102 = ((~WX1101));
assign II30207 = ((~II30217))|((~II30218));
assign WX752 = (WX689&RESET);
assign II31591 = ((~WX9668))|((~_2326_));
assign WX10743 = (WX10754&WX11347);
assign II26375 = ((~WX8553))|((~II26374));
assign II18821 = ((~WX5933))|((~II18813));
assign II10680 = ((~WX3588))|((~WX3275));
assign WX7660 = ((~II23429))|((~II23430));
assign WX7547 = ((~WX7546));
assign WX6131 = ((~WX6130));
assign WX8116 = (WX8122&WX8117);
assign WX4226 = (_2182_&WX4883);
assign WX1057 = (WX587&WX1058);
assign WX3645 = (WX3643)|(WX3642);
assign WX6093 = ((~II18682))|((~II18683));
assign WX2766 = (WX4961&WX2767);
assign WX6985 = (WX6988&RESET);
assign WX911 = ((~II2352))|((~II2353));
assign II6155 = ((~WX2012))|((~II6147));
assign WX7643 = (WX7641)|(WX7640);
assign WX4996 = ((~WX4995));
assign WX7593 = ((~WX7470));
assign II7477 = ((~_2140_))|((~II7475));
assign II2408 = ((~WX863))|((~II2406));
assign WX1975 = (WX1607&RESET);
assign WX5050 = (WX5048)|(WX5047);
assign II7521 = ((~_2140_))|((~II7519));
assign WX4749 = (WX4686&RESET);
assign WX1737 = (WX1735)|(WX1734);
assign II30278 = ((~WX9776))|((~II30270));
assign WX3795 = ((~II11440))|((~II11441));
assign WX7504 = ((~WX7503));
assign WX7048 = ((~WX7016));
assign WX9396 = ((~WX10054));
assign WX2163 = (WX2100&RESET);
assign WX11594 = ((~II35667))|((~II35668));
assign WX5984 = (WX5921&RESET);
assign WX1001 = ((~WX1000));
assign WX11072 = (WX11009&RESET);
assign WX2071 = (WX2008&RESET);
assign WX5022 = (WX5020)|(WX5019);
assign II31677 = ((~_2313_))|((~II31675));
assign II10649 = ((~WX3588))|((~WX3273));
assign WX7868 = (WX10098&WX7869);
assign WX7881 = (_2294_&WX8762);
assign WX846 = (WX783&RESET);
assign WX1238 = ((~II3543))|((~II3544));
assign WX4118 = (WX4392&WX4883);
assign II35341 = ((~WX10867))|((~II35339));
assign WX11289 = ((~WX11288));
assign WX7057 = ((~WX7025));
assign WX4521 = ((~WX4776));
assign II30635 = ((~II30610))|((~II30634));
assign WX9863 = (WX9800&RESET);
assign II14391 = ((~WX4676))|((~II14390));
assign II22105 = ((~II22107))|((~II22108));
assign WX3772 = ((~WX3771));
assign II30402 = ((~WX9784))|((~II30394));
assign WX396 = (WX394)|(WX393);
assign WX4932 = ((~WX4931));
assign II18955 = ((~WX6069))|((~II18953));
assign II11497 = ((~_2172_))|((~II11495));
assign WX10611 = (WX10861&WX11348);
assign WX5493 = ((~WX6176));
assign II15262 = ((~WX4474))|((~WX4394));
assign WX5378 = (WX5376)|(WX5375);
assign WX11120 = (WX11057&RESET);
assign WX5084 = ((~WX4884));
assign II5993 = ((~WX2294))|((~WX1938));
assign WX7747 = (WX7720&WX7728);
assign WX766 = (WX703&RESET);
assign II30225 = ((~WX9836))|((~II30224));
assign WX2441 = (WX1893&WX2442);
assign WX11545 = ((~WX11544));
assign WX8170 = ((~WX8169));
assign II2770 = ((~WX759))|((~II2762));
assign II2460 = ((~WX739))|((~II2452));
assign WX9559 = (WX9562&RESET);
assign II6343 = ((~II6333))|((~II6341));
assign WX11664 = (WX11582&WX11607);
assign WX4111 = (WX4117&WX4112);
assign WX7191 = (WX7128&RESET);
assign WX786 = (WX723&RESET);
assign II3170 = ((~WX589))|((~II3169));
assign WX3712 = (WX3711&WX3591);
assign WX7725 = ((~II23722))|((~II23723));
assign WX5320 = (WX5326&WX5321);
assign II10911 = ((~II10913))|((~II10914));
assign DATA_9_19 = ((~WX1095));
assign II18606 = ((~II18596))|((~II18604));
assign WX8584 = (WX8521&RESET);
assign WX9381 = (WX9387&WX9382);
assign WX1915 = ((~WX2150));
assign WX2346 = ((~WX2345));
assign II18699 = ((~II18689))|((~II18697));
assign WX11066 = (WX11003&RESET);
assign II3364 = ((~WX604))|((~WX533));
assign WX3000 = (WX3006&WX3001);
assign II6203 = ((~II6193))|((~II6201));
assign II10664 = ((~WX3401))|((~WX3465));
assign WX11390 = ((~WX11389));
assign WX6797 = (WX6795)|(WX6794);
assign II34820 = ((~WX11231))|((~II34818));
assign II31230 = ((~WX9642))|((~WX9558));
assign II14036 = ((~WX4526))|((~II14034));
assign WX8725 = ((~WX8724));
assign WX2843 = ((~WX2834));
assign II26677 = ((~WX8509))|((~II26676));
assign WX2515 = ((~WX2514));
assign II14972 = ((~WX4650))|((~II14971));
assign II26094 = ((~II26096))|((~II26097));
assign II34936 = ((~II34926))|((~II34934));
assign II18411 = ((~WX6173))|((~WX5843));
assign WX9274 = ((~WX10055));
assign WX1008 = (WX580&WX1009);
assign WX335 = ((~WX1004));
assign II2129 = ((~WX845))|((~II2127));
assign WX11372 = (WX11371&WX11349);
assign WX379 = (WX533&WX1004);
assign WX2617 = (WX2529&WX2556);
assign II3606 = ((~WX624))|((~II3605));
assign II2338 = ((~II2328))|((~II2336));
assign WX434 = (WX432)|(WX431);
assign WX8027 = ((~WX8762));
assign II31362 = ((~WX9578))|((~II31360));
assign II23220 = ((~WX7056))|((~WX6972));
assign WX4108 = ((~WX4099));
assign WX8050 = (WX10189&WX8051);
assign II22687 = ((~II22662))|((~II22686));
assign II6023 = ((~II6025))|((~II6026));
assign WX5114 = ((~II15537))|((~II15538));
assign WX9040 = (WX9013&WX9021);
assign WX5540 = (WX5538)|(WX5537);
assign WX702 = (WX454&RESET);
assign II18465 = ((~II18440))|((~II18464));
assign WX2041 = (WX1978&RESET);
assign WX6859 = (WX7652&WX6860);
assign WX4101 = (WX6275&WX4102);
assign WX11032 = (WX10700&RESET);
assign WX11670 = (WX11579&WX11607);
assign WX952 = ((~WX926));
assign WX2397 = ((~II7240))|((~II7241));
assign WX10606 = (WX10604)|(WX10603);
assign WX8369 = ((~WX8337));
assign II26948 = ((~WX8760))|((~WX8463));
assign WX2218 = ((~II6791))|((~II6792));
assign II26237 = ((~WX8417))|((~II26235));
assign WX6373 = ((~WX6372));
assign II2469 = ((~WX803))|((~II2468));
assign II27580 = ((~WX8374))|((~II27579));
assign II3544 = ((~_2104_))|((~II3542));
assign WX10796 = (WX10794)|(WX10793);
assign WX2531 = ((~II7548))|((~II7549));
assign II19462 = ((~WX5782))|((~WX5717));
assign II10123 = ((~WX3587))|((~II10122));
assign II6187 = ((~WX2014))|((~II6186));
assign WX3541 = ((~WX3540));
assign WX95 = (_2104_&WX1004);
assign WX4290 = ((~WX4281));
assign II34446 = ((~WX11143))|((~WX11207));
assign II35647 = ((~_2351_))|((~II35645));
assign WX9001 = ((~II27608))|((~II27609));
assign II3078 = ((~WX582))|((~WX489));
assign WX8379 = ((~WX8613));
assign WX10663 = (_2344_&WX11348);
assign WX11362 = ((~WX11361));
assign WX5799 = ((~WX6039));
assign II7318 = ((~WX1893))|((~II7317));
assign WX5806 = ((~WX6053));
assign II34656 = ((~WX11093))|((~II34655));
assign WX3846 = ((~II11707))|((~II11708));
assign WX2938 = (WX3752&WX2939);
assign WX6012 = (WX5949&RESET);
assign WX5649 = (WX5719&WX6176);
assign II31535 = ((~WX9690))|((~_2332_));
assign WX6141 = ((~WX6140));
assign WX3739 = ((~II11336))|((~II11337));
assign WX1526 = ((~WX2296));
assign WX7031 = ((~WX7402));
assign II26513 = ((~II26515))|((~II26516));
assign WX9328 = (_2315_&WX10055);
assign WX3961 = (WX6205&WX3962);
assign WX1022 = (WX582&WX1023);
assign WX8803 = (WX8801)|(WX8800);
assign WX6557 = (WX6563&WX6558);
assign WX3076 = (WX3079&RESET);
assign WX2185 = (WX2122&RESET);
assign II6072 = ((~WX2134))|((~II6070));
assign WX8069 = ((~WX8762));
assign WX7313 = (WX7250&RESET);
assign WX4213 = (WX6331&WX4214);
assign II10818 = ((~II10820))|((~II10821));
assign WX1841 = ((~WX2258));
assign WX10396 = (WX10394)|(WX10393);
assign WX1547 = (WX2410&WX1548);
assign II10044 = ((~WX3361))|((~WX3425));
assign II15676 = ((~WX4513))|((~_2181_));
assign WX1413 = (WX1419&WX1414);
assign WX1378 = (WX1784&WX2297);
assign II27740 = ((~WX8400))|((~_2269_));
assign II30659 = ((~WX9864))|((~II30658));
assign II18986 = ((~WX6071))|((~II18984));
assign WX3116 = (WX3119&RESET);
assign WX8226 = ((~WX8225));
assign II26941 = ((~II26931))|((~II26939));
assign WX9539 = (WX9542&RESET);
assign WX8498 = (WX8435&RESET);
assign II14219 = ((~II14221))|((~II14222));
assign II2291 = ((~II2281))|((~II2289));
assign II34712 = ((~WX11033))|((~II34710));
assign WX2280 = ((~WX2279));
assign II26965 = ((~WX8655))|((~II26963));
assign II22168 = ((~WX7466))|((~WX7120));
assign II2538 = ((~II2513))|((~II2537));
assign WX7574 = ((~WX7573));
assign WX4141 = (WX4139)|(WX4138);
assign WX5834 = (WX5346&RESET);
assign II6412 = ((~WX2092))|((~II6411));
assign WX7689 = (WX7688&WX7470);
assign II11482 = ((~_2172_))|((~II11480));
assign WX9655 = ((~WX9623));
assign II18363 = ((~II18365))|((~II18366));
assign WX3290 = (WX3054&RESET);
assign WX6235 = (WX6234&WX6177);
assign WX8723 = ((~WX8722));
assign II10361 = ((~II10337))|((~II10353));
assign WX9656 = ((~WX9624));
assign II35443 = ((~WX10951))|((~WX10883));
assign WX9998 = ((~WX9997));
assign WX5801 = ((~WX6043));
assign II3145 = ((~WX499))|((~II3143));
assign WX8948 = (WX8364&WX8949);
assign II34292 = ((~WX11133))|((~II34291));
assign II10711 = ((~WX3588))|((~WX3277));
assign WX8866 = (WX8864)|(WX8863);
assign II18280 = ((~II18270))|((~II18278));
assign II23555 = ((~_2266_))|((~II23553));
assign WX10473 = ((~WX11348));
assign WX10242 = ((~WX10056));
assign WX5811 = ((~WX6063));
assign WX2155 = (WX2092&RESET);
assign WX6436 = (WX6406&WX6435);
assign WX7477 = ((~WX7476));
assign WX959 = ((~WX958));
assign II34794 = ((~II34770))|((~II34786));
assign II10000 = ((~WX3231))|((~II9998));
assign II2298 = ((~WX1001))|((~WX665));
assign WX10487 = ((~WX11348));
assign WX1833 = (WX1836&RESET);
assign II11609 = ((~WX3209))|((~II11608));
assign WX1609 = (WX1615&WX1610);
assign WX48 = ((~WX47));
assign II27524 = ((~II27514))|((~II27522));
assign WX576 = ((~WX957));
assign WX2145 = (WX2082&RESET);
assign II10789 = ((~WX3409))|((~II10788));
assign II2864 = ((~WX765))|((~II2863));
assign II35604 = ((~WX10962))|((~II35603));
assign II15145 = ((~WX4465))|((~WX4376));
assign WX1404 = ((~WX2297));
assign WX5045 = ((~WX5044));
assign II30449 = ((~II30424))|((~II30448));
assign DATA_9_12 = ((~WX1144));
assign WX6819 = (WX6817)|(WX6816);
assign WX8779 = (WX8778&WX8763);
assign II10091 = ((~WX3587))|((~WX3237));
assign WX6812 = (_2246_&WX7469);
assign WX4046 = ((~WX4883));
assign WX6612 = (WX6623&WX7468);
assign WX9847 = (WX9784&RESET);
assign WX1446 = ((~WX2297));
assign WX2324 = (WX2322)|(WX2321);
assign II27602 = ((~_2292_))|((~II27600));
assign II6001 = ((~WX2002))|((~II6000));
assign WX7411 = ((~WX7388));
assign WX2099 = (WX2036&RESET);
assign WX4681 = (WX4618&RESET);
assign WX4917 = (WX4915)|(WX4914);
assign WX2527 = ((~II7520))|((~II7521));
assign WX477 = (WX547&WX1004);
assign WX6138 = ((~WX6073));
assign WX10021 = ((~WX9954));
assign II11479 = ((~II11481))|((~II11482));
assign WX119 = (WX130&WX1003);
assign WX6251 = ((~WX6177));
assign WX4812 = ((~WX4811));
assign WX1174 = ((~II3365))|((~II3366));
assign WX10083 = ((~WX10082));
assign WX6902 = ((~WX7469));
assign WX10180 = (WX10178)|(WX10177);
assign II26854 = ((~II26856))|((~II26857));
assign WX7374 = ((~II22315))|((~II22316));
assign WX3652 = (WX3650)|(WX3649);
assign WX2852 = (WX2850)|(WX2849);
assign WX9418 = ((~WX10055));
assign WX6142 = ((~WX6075));
assign WX8020 = (WX8018)|(WX8017);
assign II10640 = ((~II10616))|((~II10632));
assign WX4884 = ((~WX4875));
assign II15407 = ((~WX4416))|((~II15405));
assign WX9321 = (WX9319)|(WX9318);
assign II14157 = ((~II14159))|((~II14160));
assign II3670 = ((~_2084_))|((~II3668));
assign II10858 = ((~II10833))|((~II10857));
assign WX4091 = (WX4975&WX4092);
assign II2546 = ((~WX1002))|((~WX681));
assign II22275 = ((~II22277))|((~II22278));
assign WX1675 = (WX1673)|(WX1672);
assign WX2305 = ((~WX2304));
assign II18859 = ((~II18861))|((~II18862));
assign II6326 = ((~II6301))|((~II6325));
assign WX6929 = (WX7687&WX6930);
assign WX10601 = ((~WX10592));
assign WX9148 = ((~WX10055));
assign WX9825 = (WX9762&RESET);
assign WX8624 = (WX8561&RESET);
assign WX11200 = (WX11137&RESET);
assign WX2489 = (WX2488&WX2298);
assign WX1616 = (WX1818&WX2297);
assign WX6077 = ((~II18186))|((~II18187));
assign WX2633 = ((~WX2624));
assign WX9117 = (WX9115)|(WX9114);
assign WX2352 = (WX2350)|(WX2349);
assign II22104 = ((~II22114))|((~II22115));
assign WX1533 = (WX2403&WX1534);
assign WX4788 = ((~II14305))|((~II14306));
assign WX5474 = (WX5480&WX5475);
assign II18471 = ((~II18481))|((~II18482));
assign II10369 = ((~II10371))|((~II10372));
assign II3340 = ((~WX529))|((~II3338));
assign WX6179 = (WX6178&WX6177);
assign WX7808 = (WX7814&WX7809);
assign II26909 = ((~II26884))|((~II26908));
assign II22604 = ((~WX7148))|((~II22602));
assign WX3535 = ((~WX3534));
assign II26361 = ((~WX8425))|((~II26359));
assign II2563 = ((~WX873))|((~II2561));
assign WX9899 = (WX9836&RESET);
assign II14537 = ((~WX4622))|((~II14529));
assign II34340 = ((~WX11009))|((~II34338));
assign II14528 = ((~II14538))|((~II14539));
assign WX1588 = (WX1814&WX2297);
assign WX608 = ((~WX576));
assign WX581 = ((~WX549));
assign WX11592 = ((~II35653))|((~II35654));
assign WX10124 = (WX10122)|(WX10121);
assign WX252 = (WX250)|(WX249);
assign WX1017 = (WX1015)|(WX1014);
assign WX2830 = ((~WX2829));
assign II22873 = ((~II22848))|((~II22872));
assign WX5629 = ((~WX6175));
assign II18769 = ((~WX6057))|((~II18767));
assign II18480 = ((~WX5911))|((~II18472));
assign WX7463 = ((~TM0));
assign II23286 = ((~WX7061))|((~II23285));
assign WX8296 = (WX8299&RESET);
assign II34409 = ((~II34399))|((~II34407));
assign WX4852 = ((~WX4851));
assign WX481 = ((~WX472));
assign WX3498 = ((~II10393))|((~II10394));
assign WX6509 = (WX7477&WX6510);
assign WX8344 = ((~WX8312));
assign WX9166 = ((~WX10055));
assign WX8041 = ((~WX8762));
assign WX5708 = (WX5711&RESET);
assign WX2226 = ((~WX2225));
assign WX8442 = (WX8086&RESET);
assign II14856 = ((~WX4706))|((~II14855));
assign WX1592 = ((~WX1583));
assign II10370 = ((~WX3587))|((~WX3255));
assign WX2480 = ((~WX2479));
assign II34068 = ((~II34058))|((~II34066));
assign WX5872 = (WX5612&RESET);
assign II30548 = ((~II30558))|((~II30559));
assign II23261 = ((~WX6978))|((~II23259));
assign WX10462 = ((~WX10461));
assign WX3205 = ((~WX3437));
assign II22789 = ((~WX7467))|((~II22788));
assign II2932 = ((~II2934))|((~II2935));
assign II18263 = ((~WX5897))|((~II18255));
assign WX7940 = (WX7938)|(WX7937);
assign WX10972 = ((~WX11213));
assign WX7853 = (_2296_&WX8762);
assign WX3934 = ((~WX4883));
assign II30650 = ((~WX9800))|((~II30642));
assign II19667 = ((~WX5803))|((~_2216_));
assign WX890 = (WX827&RESET);
assign WX7383 = ((~II22594))|((~II22595));
assign WX7219 = (WX7156&RESET);
assign II34169 = ((~WX11189))|((~II34167));
assign WX8241 = ((~WX8243));
assign WX10270 = ((~WX10056));
assign WX11052 = (WX10989&RESET);
assign WX4567 = (WX4235&RESET);
assign WX4182 = ((~WX4882));
assign II7489 = ((~II7491))|((~II7492));
assign II6395 = ((~II6397))|((~II6398));
assign WX4577 = (WX4305&RESET);
assign WX156 = (DATA_9_23&WX157);
assign WX1191 = ((~WX1005));
assign WX4072 = (_2193_&WX4883);
assign WX124 = (WX2347&WX125);
assign WX7551 = ((~WX7470));
assign WX10509 = (_2355_&WX11348);
assign WX3049 = (WX3131&WX3590);
assign WX496 = (WX499&RESET);
assign WX9496 = (_2303_&WX10055);
assign WX10001 = ((~WX9976));
assign WX6087 = ((~II18496))|((~II18497));
assign WX7329 = (WX7266&RESET);
assign II14840 = ((~WX4881))|((~WX4578));
assign II15704 = ((~WX4517))|((~_2177_));
assign WX71 = (WX489&WX1004);
assign II26747 = ((~WX8577))|((~II26746));
assign II22089 = ((~II22091))|((~II22092));
assign WX2571 = (WX2550&WX2556);
assign II34347 = ((~II34337))|((~II34345));
assign II26180 = ((~WX8477))|((~II26172));
assign WX10387 = (WX10829&WX11348);
assign WX8080 = (WX8078)|(WX8077);
assign WX329 = (WX340&WX1003);
assign WX1078 = (WX590&WX1079);
assign WX1144 = ((~WX1143));
assign WX6589 = (WX8812&WX6590);
assign II30365 = ((~WX10052))|((~II30364));
assign WX595 = ((~WX563));
assign II14687 = ((~WX4568))|((~II14685));
assign WX8311 = ((~WX8733));
assign WX6080 = ((~II18279))|((~II18280));
assign WX11626 = (WX11599&WX11607);
assign II10797 = ((~II10787))|((~II10795));
assign II3493 = ((~_2087_))|((~II3492));
assign WX5107 = ((~WX5106));
assign II22169 = ((~WX7466))|((~II22168));
assign II6038 = ((~II6040))|((~II6041));
assign II35524 = ((~II35526))|((~II35527));
assign WX10198 = (WX10197&WX10056);
assign WX1661 = (WX1659)|(WX1658);
assign II23129 = ((~WX7049))|((~WX6958));
assign WX3800 = ((~WX3799));
assign WX1507 = (WX1505)|(WX1504);
assign II10448 = ((~WX3387))|((~II10447));
assign II10440 = ((~WX3323))|((~II10439));
assign WX5759 = ((~WX5727));
assign II18287 = ((~WX6173))|((~WX5835));
assign WX938 = ((~WX919));
assign WX1244 = ((~II3585))|((~II3586));
assign II26118 = ((~WX8473))|((~II26110));
assign WX7421 = ((~WX7393));
assign II35224 = ((~WX10849))|((~II35222));
assign II2446 = ((~II2436))|((~II2444));
assign WX8971 = (WX8969)|(WX8968);
assign WX7157 = (WX6849&RESET);
assign WX4491 = ((~WX4716));
assign WX5127 = ((~II15628))|((~II15629));
assign WX4939 = ((~WX4938));
assign WX6805 = (WX6803)|(WX6802);
assign WX7910 = (WX10119&WX7911);
assign WX7978 = (WX7976)|(WX7975);
assign WX6358 = ((~WX6357));
assign WX8702 = ((~WX8680));
assign WX7026 = ((~WX7456));
assign II3105 = ((~WX584))|((~II3104));
assign II34274 = ((~II34284))|((~II34285));
assign II3117 = ((~WX585))|((~WX495));
assign WX7812 = (WX10070&WX7813);
assign WX6284 = (WX6283&WX6177);
assign WX4947 = ((~WX4946));
assign II6295 = ((~II6270))|((~II6294));
assign II14446 = ((~II14436))|((~II14444));
assign WX4185 = (WX6317&WX4186);
assign WX3625 = ((~WX3624));
assign WX5612 = ((~WX5611));
assign II34431 = ((~WX11345))|((~WX11015));
assign II22417 = ((~WX7466))|((~II22416));
assign II14237 = ((~WX4730))|((~II14235));
assign WX166 = (WX2368&WX167);
assign WX6742 = (_2251_&WX7469);
assign WX7083 = ((~WX7314));
assign WX10106 = ((~II31179))|((~II31180));
assign WX1848 = ((~WX2272));
assign II2330 = ((~WX1001))|((~II2329));
assign WX1696 = (_2114_&WX2297);
assign WX2837 = ((~WX3590));
assign II31336 = ((~WX9574))|((~II31334));
assign WX10005 = ((~WX9978));
assign II26159 = ((~WX8603))|((~II26157));
assign II19717 = ((~WX5812))|((~II19716));
assign II6846 = ((~WX2120))|((~II6845));
assign WX11315 = ((~WX11314));
assign WX10459 = ((~WX11348));
assign WX3975 = (WX6212&WX3976);
assign WX373 = ((~WX1003));
assign WX5838 = (WX5374&RESET);
assign II26187 = ((~II26189))|((~II26190));
assign WX10380 = (WX10386&WX10381);
assign WX3035 = (WX3129&WX3590);
assign WX216 = ((~WX215));
assign WX2563 = (WX2553&WX2556);
assign WX9618 = ((~WX9990));
assign II30302 = ((~WX10052))|((~WX9714));
assign II19710 = ((~WX5810))|((~II19709));
assign WX1809 = (WX1812&RESET);
assign II23403 = ((~WX7070))|((~II23402));
assign WX5547 = (_2212_&WX6176);
assign WX8688 = ((~II26971))|((~II26972));
assign WX6000 = (WX5937&RESET);
assign WX7470 = ((~WX7461));
assign WX6897 = (WX8966&WX6898);
assign II22797 = ((~II22787))|((~II22795));
assign WX9662 = ((~WX9630));
assign WX4099 = (WX4097)|(WX4096);
assign WX10550 = (WX10548)|(WX10547);
assign II6690 = ((~WX2110))|((~WX2174));
assign WX2739 = ((~WX3590));
assign II10898 = ((~WX3588))|((~II10897));
assign WX1491 = (WX2382&WX1492);
assign WX10557 = ((~WX11348));
assign II2300 = ((~WX665))|((~II2298));
assign II11245 = ((~WX3180))|((~II11244));
assign II14346 = ((~WX4546))|((~II14344));
assign II2863 = ((~WX765))|((~II2855));
assign II6907 = ((~WX2124))|((~WX2188));
assign WX7982 = (WX7980)|(WX7979);
assign WX3420 = (WX3357&RESET);
assign II2732 = ((~WX1002))|((~WX693));
assign II15517 = ((~_2204_))|((~II15515));
assign II6644 = ((~WX2295))|((~WX1980));
assign WX7283 = (WX7220&RESET);
assign WX3917 = (WX3915)|(WX3914);
assign WX8918 = ((~II27369))|((~II27370));
assign II26445 = ((~II26435))|((~II26443));
assign WX6891 = ((~WX6890));
assign WX2702 = (WX2700)|(WX2699);
assign WX2967 = ((~WX3590));
assign WX3632 = ((~WX3631));
assign WX5075 = (WX5074&WX4884);
assign WX6601 = (WX6599)|(WX6598);
assign II35716 = ((~WX10980))|((~II35715));
assign WX1366 = ((~WX2297));
assign WX7819 = ((~WX7810));
assign WX9947 = (WX9884&RESET);
assign WX5151 = (WX5112&WX5142);
assign WX7933 = (WX7944&WX8761);
assign II27369 = ((~WX8360))|((~II27368));
assign WX4906 = ((~II15107))|((~II15108));
assign WX10480 = (WX10478)|(WX10477);
assign II18574 = ((~WX5917))|((~II18573));
assign WX3812 = ((~WX3591));
assign WX5574 = (WX5572)|(WX5571);
assign II26547 = ((~WX8437))|((~II26545));
assign WX10685 = ((~WX10676));
assign WX3894 = (WX3830&WX3849);
assign II18690 = ((~WX6174))|((~WX5861));
assign WX9388 = (WX9578&WX10055);
assign WX8782 = (WX8780)|(WX8779);
assign WX4006 = (WX4376&WX4883);
assign WX3216 = ((~WX3459));
assign II14670 = ((~WX4694))|((~II14669));
assign DATA_9_3 = ((~WX1207));
assign WX3069 = ((~WX3071));
assign WX3432 = (WX3369&RESET);
assign WX1683 = (WX3773&WX1684);
assign WX1652 = ((~WX2296));
assign WX1967 = (WX1551&RESET);
assign WX7720 = ((~II23687))|((~II23688));
assign WX3749 = ((~WX3591));
assign II14376 = ((~WX4880))|((~II14375));
assign WX3831 = ((~II11602))|((~II11603));
assign WX3566 = ((~WX3494));
assign WX8698 = ((~WX8678));
assign WX8336 = ((~WX8719));
assign II10214 = ((~II10216))|((~II10217));
assign WX3760 = ((~II11375))|((~II11376));
assign WX1774 = ((~WX1765));
assign II34073 = ((~II34075))|((~II34076));
assign WX1670 = ((~WX2297));
assign WX3062 = (WX3060)|(WX3059);
assign WX11454 = ((~WX11453));
assign WX4240 = (_2181_&WX4883);
assign WX8231 = (_2269_&WX8762);
assign WX3472 = (WX3409&RESET);
assign II30373 = ((~II30363))|((~II30371));
assign II27735 = ((~_2270_))|((~II27733));
assign II18180 = ((~WX6019))|((~II18178));
assign WX9605 = ((~WX10028));
assign II2167 = ((~II2157))|((~II2165));
assign II6658 = ((~II6660))|((~II6661));
assign II23233 = ((~WX7057))|((~WX6974));
assign II11671 = ((~WX3220))|((~_2149_));
assign II27136 = ((~WX8251))|((~II27134));
assign WX1777 = (WX1780&RESET);
assign WX11548 = (WX10952&WX11549);
assign WX5840 = (WX5388&RESET);
assign WX3480 = (WX3417&RESET);
assign WX6351 = ((~WX6350));
assign II14957 = ((~II14947))|((~II14955));
assign WX1558 = ((~WX2297));
assign WX2365 = ((~WX2298));
assign II31662 = ((~WX9679))|((~II31661));
assign II2079 = ((~II2089))|((~II2090));
assign WX6048 = (WX5985&RESET);
assign II27644 = ((~_2286_))|((~II27642));
assign WX7267 = (WX7204&RESET);
assign WX2111 = (WX2048&RESET);
assign II15393 = ((~WX4484))|((~II15392));
assign II11706 = ((~WX3226))|((~_2143_));
assign II34494 = ((~WX11345))|((~II34493));
assign II30335 = ((~WX9716))|((~II30333));
assign II26438 = ((~WX8621))|((~II26436));
assign WX7667 = ((~II23442))|((~II23443));
assign II22695 = ((~WX7467))|((~WX7154));
assign WX8341 = ((~WX8309));
assign WX5625 = ((~WX5616));
assign WX7416 = ((~WX7415));
assign II6859 = ((~II6869))|((~II6870));
assign WX8288 = (WX8291&RESET);
assign II11650 = ((~WX3216))|((~_2153_));
assign II27593 = ((~WX8376))|((~_2293_));
assign II26474 = ((~II26450))|((~II26466));
assign WX7948 = (WX7954&WX7949);
assign WX6182 = (WX6180)|(WX6179);
assign WX9058 = (WX9006&WX9021);
assign WX5353 = ((~WX6176));
assign II23575 = ((~WX7081))|((~II23574));
assign WX9020 = ((~II27741))|((~II27742));
assign WX7001 = (WX7004&RESET);
assign WX4433 = ((~WX4856));
assign II26499 = ((~WX8561))|((~II26498));
assign II22331 = ((~WX7194))|((~II22330));
assign II35483 = ((~WX10954))|((~II35482));
assign II30953 = ((~WX10053))|((~WX9756));
assign WX1314 = (WX1241&WX1263);
assign WX8538 = (WX8475&RESET);
assign II31087 = ((~WX9631))|((~WX9536));
assign WX5774 = ((~WX5742));
assign WX4387 = (WX4390&RESET);
assign II10170 = ((~WX3433))|((~II10168));
assign WX7542 = (WX7541&WX7470);
assign WX10191 = (WX10190&WX10056);
assign II19190 = ((~WX5761))|((~II19189));
assign WX8350 = ((~WX8318));
assign WX8518 = (WX8455&RESET);
assign WX3173 = ((~WX3141));
assign WX11356 = ((~WX11355));
assign WX540 = (WX543&RESET);
assign WX5940 = (WX5877&RESET);
assign II30440 = ((~II30442))|((~II30443));
assign II18148 = ((~WX5953))|((~II18147));
assign WX9577 = (WX9580&RESET);
assign WX8182 = (WX8180)|(WX8179);
assign WX11412 = ((~WX11411));
assign II10656 = ((~WX3337))|((~II10648));
assign WX6935 = (WX6941&WX6936);
assign WX3816 = ((~RESET));
assign WX5466 = (WX5464)|(WX5463);
assign WX7650 = (WX7648)|(WX7647);
assign WX3575 = ((~WX3574));
assign II14575 = ((~II14577))|((~II14578));
assign WX1073 = (WX1071)|(WX1070);
assign II19464 = ((~WX5717))|((~II19462));
assign II34522 = ((~II34532))|((~II34533));
assign WX1063 = (WX1062&WX1005);
assign WX5620 = (WX5618)|(WX5617);
assign WX1868 = ((~WX2248));
assign II22562 = ((~II22538))|((~II22554));
assign II22222 = ((~II22197))|((~II22221));
assign WX7393 = ((~II22904))|((~II22905));
assign II35471 = ((~WX10887))|((~II35469));
assign WX4829 = ((~WX4804));
assign II22631 = ((~II22641))|((~II22642));
assign WX607 = ((~WX575));
assign II11166 = ((~WX3174))|((~WX3087));
assign WX1659 = (WX2466&WX1660);
assign WX908 = ((~II2259))|((~II2260));
assign WX1999 = (WX1775&RESET);
assign WX2685 = (WX3079&WX3590);
assign WX4159 = (WX4157)|(WX4156);
assign WX1133 = (WX1132&WX1005);
assign II2042 = ((~II2017))|((~II2041));
assign II30486 = ((~II30496))|((~II30497));
assign WX11571 = (WX11569)|(WX11568);
assign WX7688 = ((~II23481))|((~II23482));
assign WX6567 = (WX6565)|(WX6564);
assign WX7877 = (WX7888&WX8761);
assign II14632 = ((~II14622))|((~II14630));
assign WX3552 = ((~WX3487));
assign II19655 = ((~_2218_))|((~II19653));
assign WX4234 = ((~WX4225));
assign II26593 = ((~WX8631))|((~II26591));
assign II2670 = ((~WX1002))|((~WX689));
assign II22199 = ((~WX7466))|((~WX7122));
assign II14282 = ((~WX4880))|((~WX4542));
assign WX7619 = (WX7618&WX7470);
assign WX1719 = ((~WX1718));
assign WX2707 = ((~WX3589));
assign WX10110 = (WX10108)|(WX10107);
assign WX3811 = (WX3197&WX3812);
assign II11615 = ((~WX3210))|((~_2159_));
assign WX6272 = ((~WX6177));
assign WX10011 = ((~WX9981));
assign WX11632 = (WX11597&WX11607);
assign WX5608 = (WX6380&WX5609);
assign WX10695 = (WX10873&WX11348);
assign II10565 = ((~II10555))|((~II10563));
assign II2951 = ((~WX707))|((~II2949));
assign WX5731 = ((~WX6159));
assign WX41 = ((~WX1004));
assign II27433 = ((~WX8365))|((~WX8297));
assign WX1562 = ((~WX2297));
assign WX6755 = (WX6753)|(WX6752);
assign WX8634 = (WX8571&RESET);
assign II14700 = ((~WX4696))|((~WX4760));
assign WX2819 = ((~WX3589));
assign WX3126 = (WX3129&RESET);
assign II18341 = ((~II18316))|((~II18340));
assign WX1551 = ((~WX1550));
assign WX3972 = ((~WX4882));
assign II26801 = ((~WX8517))|((~II26800));
assign WX11556 = ((~WX11349));
assign WX928 = ((~II2879))|((~II2880));
assign WX1850 = ((~WX2276));
assign II35518 = ((~_2348_))|((~II35517));
assign WX9669 = ((~WX9900));
assign DATA_9_20 = ((~WX1088));
assign WX2906 = (WX5031&WX2907);
assign WX4150 = ((~WX4141));
assign WX4795 = ((~II14522))|((~II14523));
assign WX6363 = ((~WX6177));
assign WX10862 = (WX10865&RESET);
assign WX11552 = ((~WX11551));
assign II31607 = ((~_2324_))|((~II31605));
assign II18271 = ((~WX5961))|((~WX6025));
assign II6823 = ((~II6813))|((~II6821));
assign WX9231 = (WX11426&WX9232);
assign WX7165 = (WX6905&RESET);
assign II18202 = ((~WX5893))|((~II18201));
assign WX11333 = ((~WX11332));
assign WX1439 = ((~WX1438));
assign II6367 = ((~WX1962))|((~II6365));
assign II3676 = ((~WX636))|((~II3675));
assign WX1903 = ((~WX1871));
assign II2839 = ((~II2841))|((~II2842));
assign WX3334 = (WX3271&RESET);
assign II15223 = ((~WX4471))|((~WX4388));
assign WX10279 = ((~WX10278));
assign WX3051 = ((~WX3590));
assign II2321 = ((~II2296))|((~II2320));
assign WX5068 = (WX5067&WX4884);
assign WX3995 = (WX3993)|(WX3992);
assign II3472 = ((~_2108_))|((~II3470));
assign II22012 = ((~II22014))|((~II22015));
assign WX4960 = ((~WX4959));
assign WX5336 = (WX5334)|(WX5333);
assign WX8472 = (WX8409&RESET);
assign WX5454 = (WX6303&WX5455);
assign WX9644 = ((~WX9612));
assign WX947 = ((~WX946));
assign II27572 = ((~WX8373))|((~_2296_));
assign II26962 = ((~II26964))|((~II26965));
assign WX5018 = ((~II15315))|((~II15316));
assign WX7532 = ((~WX7531));
assign WX8592 = (WX8529&RESET);
assign WX2039 = (WX1976&RESET);
assign II34501 = ((~WX11083))|((~II34500));
assign WX7681 = ((~II23468))|((~II23469));
assign WX7054 = ((~WX7022));
assign II2523 = ((~WX743))|((~II2522));
assign WX2414 = ((~WX2298));
assign II6738 = ((~WX2295))|((~II6737));
assign II30922 = ((~WX10053))|((~WX9754));
assign II18319 = ((~WX6173))|((~II18318));
assign II26671 = ((~WX8445))|((~II26669));
assign II10558 = ((~WX3267))|((~II10556));
assign WX11214 = (WX11151&RESET);
assign II10472 = ((~II10462))|((~II10470));
assign WX4272 = (WX4414&WX4883);
assign WX4819 = ((~WX4799));
assign II6582 = ((~WX2295))|((~WX1976));
assign II30217 = ((~WX9772))|((~II30216));
assign II2622 = ((~II2624))|((~II2625));
assign WX10440 = (DATA_0_27&WX10441);
assign WX11293 = ((~WX11292));
assign WX10071 = ((~II31114))|((~II31115));
assign WX10517 = ((~WX10508));
assign WX7828 = (WX7826)|(WX7825);
assign WX7876 = ((~WX7875));
assign WX10449 = (WX10460&WX11347);
assign WX8737 = ((~WX8736));
assign WX1576 = ((~WX2297));
assign II30603 = ((~II30579))|((~II30595));
assign WX730 = (WX667&RESET);
assign II14987 = ((~II14962))|((~II14986));
assign WX8189 = (_2272_&WX8762);
assign WX5526 = (WX5524)|(WX5523);
assign WX5968 = (WX5905&RESET);
assign WX1730 = ((~WX2297));
assign II10541 = ((~WX3393))|((~II10540));
assign II6863 = ((~WX1994))|((~II6861));
assign WX6618 = ((~WX7469));
assign WX3314 = (WX3251&RESET);
assign WX617 = ((~WX847));
assign WX7989 = (WX8000&WX8761);
assign WX6661 = (WX6659)|(WX6658);
assign II27539 = ((~II27529))|((~II27537));
assign WX7892 = (WX7898&WX7893);
assign WX8887 = (WX8885)|(WX8884);
assign II18898 = ((~II18874))|((~II18890));
assign II3479 = ((~II3469))|((~II3477));
assign WX10587 = ((~WX10578));
assign WX8872 = ((~WX8763));
assign WX10421 = (WX10432&WX11347);
assign WX6167 = ((~WX6166));
assign II34515 = ((~II34491))|((~II34507));
assign WX7492 = ((~II23117))|((~II23118));
assign WX6066 = (WX6003&RESET);
assign WX2882 = (WX3724&WX2883);
assign II6077 = ((~II6053))|((~II6069));
assign II34231 = ((~WX11193))|((~II34229));
assign WX4800 = ((~II14677))|((~II14678));
assign WX5440 = (WX6296&WX5441);
assign II22647 = ((~II22649))|((~II22650));
assign WX4198 = (_2184_&WX4883);
assign WX5954 = (WX5891&RESET);
assign II34122 = ((~WX11345))|((~II34121));
assign II18102 = ((~WX6173))|((~II18101));
assign WX160 = ((~WX159));
assign II10293 = ((~WX3377))|((~II10292));
assign WX974 = ((~WX905));
assign WX11563 = ((~WX11349));
assign II19519 = ((~II19521))|((~II19522));
assign II19152 = ((~WX5669))|((~II19150));
assign WX614 = ((~WX841));
assign WX10804 = (DATA_0_1&WX10805);
assign WX8906 = (WX8358&WX8907);
assign WX11176 = (WX11113&RESET);
assign WX2287 = ((~WX2208));
assign WX10510 = (DATA_0_22&WX10511);
assign WX8982 = (WX8981&WX8763);
assign II27579 = ((~WX8374))|((~_2295_));
assign WX10774 = (WX10772)|(WX10771);
assign II18536 = ((~WX6174))|((~II18535));
assign WX6639 = ((~WX6638));
assign II7582 = ((~WX1913))|((~_2131_));
assign WX11504 = ((~II35379))|((~II35380));
assign WX3821 = ((~II11532))|((~II11533));
assign WX3958 = ((~WX4882));
assign II34243 = ((~II34253))|((~II34254));
assign II26832 = ((~WX8519))|((~II26831));
assign II34128 = ((~WX11059))|((~II34120));
assign II26886 = ((~WX8760))|((~WX8459));
assign II6568 = ((~WX2166))|((~II6566));
assign II14452 = ((~WX4680))|((~WX4744));
assign II10020 = ((~II9996))|((~II10012));
assign WX2312 = ((~WX2311));
assign WX2601 = (WX2537&WX2556);
assign II14895 = ((~II14885))|((~II14893));
assign WX6722 = ((~WX6713));
assign WX11599 = ((~II35702))|((~II35703));
assign WX4976 = ((~II15237))|((~II15238));
assign WX11244 = ((~II34051))|((~II34052));
assign II26016 = ((~II26026))|((~II26027));
assign WX8928 = ((~WX8763));
assign II14863 = ((~II14838))|((~II14862));
assign II6132 = ((~WX2074))|((~WX2138));
assign WX10179 = ((~WX10056));
assign WX11234 = (WX11171&RESET);
assign WX1341 = ((~WX1340));
assign II10046 = ((~WX3425))|((~II10044));
assign WX3181 = ((~WX3149));
assign II23156 = ((~WX7051))|((~II23155));
assign WX8825 = ((~WX8824));
assign II27108 = ((~WX8340))|((~WX8247));
assign II2958 = ((~II2948))|((~II2956));
assign II14298 = ((~WX4670))|((~II14297));
assign WX4066 = ((~WX4057));
assign WX4207 = ((~WX4206));
assign WX11284 = ((~WX11264));
assign WX4200 = ((~WX4883));
assign WX6427 = ((~II19682))|((~II19683));
assign WX209 = ((~WX1004));
assign WX9415 = (WX9413)|(WX9412);
assign WX2644 = (WX3605&WX2645);
assign II34935 = ((~WX11111))|((~II34934));
assign WX3222 = ((~WX3471));
assign II3502 = ((~_2108_))|((~II3500));
assign WX1109 = ((~WX1108));
assign II10929 = ((~WX3588))|((~II10928));
assign II10589 = ((~WX3269))|((~II10587));
assign WX11218 = (WX11155&RESET);
assign II18528 = ((~II18518))|((~II18526));
assign WX10771 = (WX10782&WX11347);
assign WX455 = (WX466&WX1003);
assign WX11401 = (WX10931&WX11402);
assign WX9120 = ((~WX10055));
assign II3579 = ((~_2099_))|((~II3577));
assign WX8323 = ((~WX8693));
assign WX8248 = (WX8251&RESET);
assign WX4551 = (WX4123&RESET);
assign WX9939 = (WX9876&RESET);
assign WX11278 = ((~WX11261));
assign WX2265 = ((~WX2197));
assign II6443 = ((~WX2094))|((~II6442));
assign WX7514 = (WX7513&WX7470);
assign WX4452 = ((~WX4830));
assign II7548 = ((~WX1908))|((~II7547));
assign II22408 = ((~II22383))|((~II22407));
assign WX5382 = (WX5380)|(WX5379);
assign II10199 = ((~WX3371))|((~WX3435));
assign II2468 = ((~WX803))|((~WX867));
assign WX7173 = (WX7110&RESET);
assign II2430 = ((~WX737))|((~II2429));
assign II18504 = ((~WX6174))|((~WX5849));
assign WX9440 = (_2307_&WX10055);
assign WX3487 = ((~II10052))|((~II10053));
assign II30629 = ((~WX9926))|((~II30627));
assign WX3513 = ((~II10858))|((~II10859));
assign II30641 = ((~II30651))|((~II30652));
assign WX10119 = ((~WX10118));
assign WX11606 = ((~II35751))|((~II35752));
assign II30767 = ((~WX10053))|((~WX9744));
assign II26127 = ((~WX8537))|((~II26126));
assign WX1569 = (WX1567)|(WX1566);
assign II22285 = ((~II22275))|((~II22283));
assign WX8237 = ((~WX8762));
assign WX132 = ((~WX131));
assign II34154 = ((~WX10997))|((~II34152));
assign WX1468 = (WX1479&WX2296);
assign WX3082 = (WX3085&RESET);
assign WX4836 = ((~WX4835));
assign WX5273 = ((~WX6176));
assign II2437 = ((~WX801))|((~WX865));
assign WX8221 = (WX8303&WX8762);
assign WX11557 = (WX11555)|(WX11554);
assign WX3464 = (WX3401&RESET);
assign WX8147 = (_2275_&WX8762);
assign WX10428 = (WX10426)|(WX10425);
assign II23181 = ((~WX7053))|((~WX6966));
assign II23363 = ((~WX7067))|((~WX6994));
assign II22144 = ((~WX7182))|((~II22136));
assign II31206 = ((~WX9554))|((~II31204));
assign II18141 = ((~II18131))|((~II18139));
assign II22790 = ((~WX7160))|((~II22788));
assign WX10760 = (WX10758)|(WX10757);
assign WX2924 = (WX3745&WX2925);
assign II2245 = ((~II2235))|((~II2243));
assign WX4445 = ((~WX4816));
assign II34236 = ((~II34212))|((~II34228));
assign II11297 = ((~WX3184))|((~II11296));
assign II10182 = ((~II10192))|((~II10193));
assign II31571 = ((~WX9665))|((~II31570));
assign II11441 = ((~WX3129))|((~II11439));
assign WX4723 = (WX4660&RESET);
assign WX2734 = (WX2740&WX2735);
assign WX5389 = (WX5400&WX6175);
assign WX9643 = ((~WX9611));
assign WX6190 = ((~WX6189));
assign WX553 = ((~WX975));
assign WX11484 = (WX11483&WX11349);
assign WX10525 = ((~WX11348));
assign WX6381 = ((~II19450))|((~II19451));
assign WX2691 = (WX2702&WX3589);
assign WX7639 = ((~II23390))|((~II23391));
assign WX7539 = ((~WX7538));
assign II34966 = ((~WX11113))|((~II34965));
assign II11568 = ((~_2166_))|((~II11566));
assign WX2528 = ((~II7527))|((~II7528));
assign WX4969 = ((~II15224))|((~II15225));
assign II31167 = ((~WX9548))|((~II31165));
assign II18223 = ((~II18233))|((~II18234));
assign WX9104 = (_2331_&WX10055);
assign II26731 = ((~WX8760))|((~WX8449));
assign WX382 = (WX380)|(WX379);
assign WX5726 = ((~WX6149));
assign II34035 = ((~WX11053))|((~II34027));
assign II15133 = ((~WX4464))|((~II15132));
assign II10548 = ((~II10523))|((~II10547));
assign WX3948 = ((~WX4883));
assign WX8140 = (WX8138)|(WX8137);
assign II2414 = ((~II2389))|((~II2413));
assign II2026 = ((~WX711))|((~II2018));
assign WX4089 = (WX4087)|(WX4086);
assign II11617 = ((~_2159_))|((~II11615));
assign WX7565 = ((~WX7470));
assign WX5994 = (WX5931&RESET);
assign II2096 = ((~WX779))|((~WX843));
assign II14072 = ((~WX4592))|((~II14064));
assign II26977 = ((~II26987))|((~II26988));
assign II30914 = ((~II30889))|((~II30913));
assign II34817 = ((~II34819))|((~II34820));
assign II10523 = ((~II10533))|((~II10534));
assign WX10864 = (WX10867&RESET);
assign WX2857 = ((~WX2848));
assign II22554 = ((~II22556))|((~II22557));
assign II18526 = ((~II18502))|((~II18518));
assign II14079 = ((~II14081))|((~II14082));
assign WX10750 = (WX10748)|(WX10747);
assign WX9344 = ((~WX10055));
assign WX8665 = ((~II26258))|((~II26259));
assign WX6494 = (WX6409&WX6435);
assign II22075 = ((~WX7466))|((~WX7114));
assign II3455 = ((~WX611))|((~WX547));
assign WX7099 = ((~WX7346));
assign II18738 = ((~WX6055))|((~II18736));
assign WX8370 = ((~WX8595));
assign WX9152 = ((~WX10055));
assign WX3736 = (WX3734)|(WX3733);
assign WX10056 = ((~WX10047));
assign II19646 = ((~WX5800))|((~_2219_));
assign II18170 = ((~WX5891))|((~II18162));
assign WX6781 = (WX6787&WX6782);
assign II7710 = ((~_2110_))|((~II7708));
assign WX364 = (WX362)|(WX361);
assign II15379 = ((~WX4483))|((~WX4412));
assign II10960 = ((~WX3588))|((~II10959));
assign WX7997 = (WX8271&WX8762);
assign II34665 = ((~WX11221))|((~II34663));
assign WX10591 = ((~WX11347));
assign II7137 = ((~WX1790))|((~II7135));
assign II27720 = ((~WX8396))|((~II27719));
assign II27447 = ((~WX8366))|((~II27446));
assign WX7452 = ((~WX7451));
assign II18891 = ((~WX6001))|((~WX6065));
assign WX2492 = (WX2490)|(WX2489);
assign II18365 = ((~WX5967))|((~II18364));
assign II14267 = ((~WX4668))|((~II14266));
assign II26653 = ((~WX8571))|((~WX8635));
assign II30900 = ((~II30890))|((~II30898));
assign II22588 = ((~WX7338))|((~II22586));
assign WX3165 = ((~WX3549));
assign WX5015 = (WX5013)|(WX5012);
assign II7513 = ((~_2112_))|((~II7512));
assign WX1722 = ((~WX2296));
assign II2700 = ((~II2702))|((~II2703));
assign WX1092 = (WX592&WX1093);
assign WX3823 = ((~II11546))|((~II11547));
assign WX10520 = (WX10526&WX10521);
assign WX8424 = (WX7960&RESET);
assign WX9455 = (WX11538&WX9456);
assign WX1036 = (WX584&WX1037);
assign II2879 = ((~II2854))|((~II2878));
assign WX4039 = ((~WX4038));
assign WX2654 = (WX4905&WX2655);
assign II34112 = ((~II34088))|((~II34104));
assign WX10892 = ((~WX11309));
assign WX11206 = (WX11143&RESET);
assign WX9727 = (WX9323&RESET);
assign WX6249 = (WX6248&WX6177);
assign WX1852 = ((~WX2280));
assign II6490 = ((~WX2295))|((~II6489));
assign WX4012 = (WX4023&WX4882);
assign II30782 = ((~WX9872))|((~WX9936));
assign II7111 = ((~WX1786))|((~II7109));
assign II2870 = ((~II2872))|((~II2873));
assign II27516 = ((~WX8390))|((~II27515));
assign II3537 = ((~_2105_))|((~II3535));
assign WX3836 = ((~II11637))|((~II11638));
assign WX2299 = ((~II7058))|((~II7059));
assign WX4929 = (WX4465&WX4930);
assign II10501 = ((~WX3327))|((~II10493));
assign WX8788 = ((~WX8763));
assign II34957 = ((~II34959))|((~II34960));
assign II6218 = ((~WX2016))|((~II6217));
assign WX1419 = (WX1417)|(WX1416);
assign II18682 = ((~II18657))|((~II18681));
assign WX10767 = ((~WX11348));
assign WX10645 = (WX10656&WX11347);
assign WX7526 = ((~WX7525));
assign WX9261 = (WX9259)|(WX9258);
assign WX4019 = (WX4017)|(WX4016);
assign WX9068 = (WX9001&WX9021);
assign II26212 = ((~WX8479))|((~II26211));
assign WX4864 = ((~WX4863));
assign II30776 = ((~II30766))|((~II30774));
assign II34987 = ((~II34997))|((~II34998));
assign II10868 = ((~WX3287))|((~II10866));
assign WX10809 = ((~WX11348));
assign II10626 = ((~WX3335))|((~II10625));
assign WX8923 = ((~WX8922));
assign WX7460 = ((~WX7459));
assign II11561 = ((~_2167_))|((~II11559));
assign II15628 = ((~WX4504))|((~II15627));
assign WX2625 = (_2172_&WX3590);
assign WX7992 = (WX7990)|(WX7989);
assign WX2195 = ((~II6078))|((~II6079));
assign WX2333 = ((~WX2332));
assign WX8093 = ((~WX8762));
assign WX1634 = ((~WX1625));
assign WX10091 = ((~WX10090));
assign WX5105 = ((~WX4884));
assign WX9088 = ((~WX10054));
assign II31452 = ((~WX9659))|((~II31451));
assign II11271 = ((~WX3182))|((~II11270));
assign II15197 = ((~WX4469))|((~WX4384));
assign WX436 = (DATA_9_3&WX437);
assign WX9306 = ((~WX10055));
assign WX6761 = (WX7603&WX6762);
assign WX5436 = (WX7589&WX5437);
assign II2607 = ((~II2609))|((~II2610));
assign II26879 = ((~II26869))|((~II26877));
assign WX5509 = (WX5699&WX6176);
assign WX3052 = (WX3050)|(WX3049);
assign II34943 = ((~WX11175))|((~II34942));
assign WX6122 = ((~WX6097));
assign WX6693 = (WX6691)|(WX6690);
assign WX5375 = (WX5386&WX6175);
assign WX6263 = (WX6262&WX6177);
assign WX11634 = (WX11596&WX11607);
assign WX2986 = (WX2992&WX2987);
assign WX1480 = ((~WX1471));
assign WX2757 = ((~WX3590));
assign WX5503 = ((~WX6175));
assign II31373 = ((~WX9653))|((~WX9580));
assign II3684 = ((~_2082_))|((~II3682));
assign WX4032 = ((~WX4883));
assign II14878 = ((~WX4644))|((~II14870));
assign II26662 = ((~II26652))|((~II26660));
assign II10804 = ((~WX3588))|((~WX3283));
assign II2926 = ((~WX769))|((~II2925));
assign WX10776 = (DATA_0_3&WX10777);
assign WX6520 = ((~WX7469));
assign II23365 = ((~WX6994))|((~II23363));
assign WX10435 = (WX10446&WX11347);
assign II22532 = ((~II22507))|((~II22531));
assign II19215 = ((~WX5763))|((~WX5679));
assign WX10929 = ((~WX10897));
assign DATA_9_8 = ((~WX1172));
assign WX87 = ((~WX1004));
assign WX8014 = (WX8012)|(WX8011);
assign II34586 = ((~WX11346))|((~WX11025));
assign II7462 = ((~WX1840))|((~II7460));
assign WX5083 = (WX4487&WX5084);
assign WX5597 = ((~WX5588));
assign II10787 = ((~II10789))|((~II10790));
assign WX11438 = (WX11436)|(WX11435);
assign WX9138 = ((~WX10055));
assign II10415 = ((~II10417))|((~II10418));
assign II30992 = ((~WX9822))|((~II30991));
assign WX9986 = ((~WX9985));
assign II6799 = ((~WX2295))|((~WX1990));
assign II26337 = ((~II26327))|((~II26335));
assign WX4920 = ((~II15133))|((~II15134));
assign WX1489 = (WX1487)|(WX1486);
assign WX4497 = ((~WX4728));
assign II26345 = ((~WX8615))|((~II26343));
assign II27685 = ((~WX8391))|((~II27684));
assign WX3818 = ((~II11503))|((~II11504));
assign WX7351 = (WX7288&RESET);
assign WX7117 = (WX6569&RESET);
assign WX5738 = ((~WX6109));
assign II18218 = ((~II18208))|((~II18216));
assign WX10325 = (WX10310&WX10314);
assign WX1873 = ((~WX1841));
assign WX4263 = ((~WX4262));
assign II34247 = ((~WX11003))|((~II34245));
assign WX2019 = (WX1956&RESET);
assign II18775 = ((~II18750))|((~II18774));
assign II23390 = ((~WX7069))|((~II23389));
assign II23077 = ((~WX7045))|((~WX6950));
assign WX6034 = (WX5971&RESET);
assign II22197 = ((~II22207))|((~II22208));
assign II14756 = ((~II14746))|((~II14754));
assign II3067 = ((~WX487))|((~II3065));
assign II2028 = ((~II2018))|((~II2026));
assign WX11110 = (WX11047&RESET);
assign II10826 = ((~II10802))|((~II10818));
assign WX2806 = (WX2804)|(WX2803);
assign WX10301 = ((~II31662))|((~II31663));
assign WX6208 = (WX5756&WX6209);
assign WX10781 = ((~WX11348));
assign WX8909 = ((~WX8908));
assign WX3150 = ((~WX3519));
assign WX3666 = (WX3664)|(WX3663);
assign WX4146 = (WX4396&WX4883);
assign WX5078 = (WX5076)|(WX5075);
assign WX7014 = ((~WX7432));
assign WX4637 = (WX4574&RESET);
assign II27317 = ((~WX8356))|((~II27316));
assign II7715 = ((~WX1935))|((~_2109_));
assign II7617 = ((~WX1918))|((~_2126_));
assign II34216 = ((~WX11001))|((~II34214));
assign WX3027 = (WX3038&WX3589);
assign II30102 = ((~WX9892))|((~II30100));
assign II10192 = ((~WX3307))|((~II10191));
assign WX3966 = ((~WX4883));
assign WX1761 = ((~WX1760));
assign WX4116 = ((~WX4883));
assign WX5056 = ((~WX4884));
assign II27719 = ((~WX8396))|((~_2273_));
assign WX6786 = ((~WX7469));
assign WX4841 = ((~WX4810));
assign II22895 = ((~II22897))|((~II22898));
assign WX5516 = (WX5522&WX5517);
assign WX4205 = (WX4203)|(WX4202);
assign II22383 = ((~II22393))|((~II22394));
assign II6195 = ((~WX2078))|((~II6194));
assign WX2761 = (WX2772&WX3589);
assign WX9869 = (WX9806&RESET);
assign WX10740 = (WX10738)|(WX10737);
assign WX10426 = (DATA_0_28&WX10427);
assign WX11603 = ((~II35730))|((~II35731));
assign WX6474 = (WX6419&WX6435);
assign WX10679 = ((~WX11348));
assign WX5205 = (WX5114&WX5142);
assign WX999 = ((~TM1));
assign WX1874 = ((~WX1842));
assign WX4898 = ((~WX4897));
assign WX5293 = ((~WX6175));
assign II34438 = ((~WX11079))|((~II34430));
assign II11623 = ((~WX3211))|((~II11622));
assign WX10913 = ((~WX11287));
assign WX407 = (WX537&WX1004);
assign WX2462 = (WX1896&WX2463);
assign WX11046 = (WX10798&RESET);
assign II14198 = ((~II14188))|((~II14196));
assign WX6971 = (WX6974&RESET);
assign WX9587 = (WX9590&RESET);
assign WX6096 = ((~II18775))|((~II18776));
assign WX4874 = ((~WX4873));
assign WX10076 = ((~WX10075));
assign II35534 = ((~II35524))|((~II35532));
assign II14585 = ((~II14575))|((~II14583));
assign II34370 = ((~WX11345))|((~II34369));
assign II10306 = ((~II10316))|((~II10317));
assign WX10308 = ((~II31711))|((~II31712));
assign II26025 = ((~WX8467))|((~II26017));
assign WX3160 = ((~WX3539));
assign II35236 = ((~WX10935))|((~II35235));
assign WX9929 = (WX9866&RESET);
assign II11102 = ((~WX3169))|((~II11101));
assign WX7440 = ((~WX7439));
assign WX112 = (WX110)|(WX109);
assign WX297 = ((~WX1004));
assign WX3919 = (WX6184&WX3920);
assign II18084 = ((~II18086))|((~II18087));
assign WX380 = (DATA_9_7&WX381);
assign II22231 = ((~WX7466))|((~II22230));
assign WX1257 = ((~II3676))|((~II3677));
assign WX5639 = ((~WX5630));
assign WX1126 = (WX1125&WX1005);
assign WX6511 = (WX6509)|(WX6508);
assign WX4895 = ((~WX4884));
assign II23686 = ((~WX7099))|((~_2245_));
assign WX10727 = ((~WX10718));
assign WX10676 = (WX10674)|(WX10673);
assign II27727 = ((~WX8398))|((~II27726));
assign II22120 = ((~II22122))|((~II22123));
assign II14213 = ((~II14203))|((~II14211));
assign WX4232 = ((~WX4883));
assign WX10948 = ((~WX10916));
assign WX5197 = (WX5118&WX5142);
assign WX9281 = ((~WX9280));
assign WX3568 = ((~WX3495));
assign WX9807 = (WX9744&RESET);
assign II18967 = ((~II18977))|((~II18978));
assign II11426 = ((~WX3194))|((~WX3127));
assign WX3141 = ((~WX3565));
assign WX9731 = (WX9351&RESET);
assign II18427 = ((~WX5971))|((~II18426));
assign II18040 = ((~WX6173))|((~II18039));
assign WX3705 = (WX3704&WX3591);
assign WX3352 = (WX3289&RESET);
assign WX9169 = ((~WX9168));
assign WX10547 = (WX10558&WX11347);
assign II7666 = ((~WX1927))|((~_2117_));
assign WX5238 = (WX5236)|(WX5235);
assign WX3780 = ((~WX3779));
assign WX1823 = (WX1826&RESET);
assign WX10701 = (WX10712&WX11347);
assign II14793 = ((~WX4702))|((~WX4766));
assign II2708 = ((~WX755))|((~II2700));
assign II2833 = ((~WX763))|((~II2832));
assign WX2995 = ((~WX3590));
assign WX9955 = ((~II30170))|((~II30171));
assign WX3743 = (WX3741)|(WX3740);
assign WX6341 = (WX5775&WX6342);
assign WX6944 = ((~WX7469));
assign WX224 = (WX222)|(WX221);
assign II30062 = ((~WX9762))|((~II30061));
assign II14638 = ((~WX4692))|((~WX4756));
assign WX10817 = (_2333_&WX11348);
assign II22492 = ((~II22494))|((~II22495));
assign WX9394 = (WX9405&WX10054);
assign II19280 = ((~WX5768))|((~WX5689));
assign WX1162 = (WX602&WX1163);
assign WX2404 = ((~II7253))|((~II7254));
assign WX4989 = ((~WX4988));
assign II34469 = ((~WX11081))|((~II34461));
assign II30859 = ((~II30861))|((~II30862));
assign WX7893 = ((~WX8761));
assign II14693 = ((~WX4632))|((~II14692));
assign II26630 = ((~II26605))|((~II26629));
assign WX9160 = (_2327_&WX10055);
assign WX1512 = ((~WX2296));
assign WX1343 = (WX1349&WX1344);
assign II10402 = ((~WX3587))|((~II10401));
assign WX9491 = ((~WX9490));
assign WX462 = (WX460)|(WX459);
assign WX2292 = ((~TM1));
assign II10896 = ((~II10898))|((~II10899));
assign II2734 = ((~WX693))|((~II2732));
assign WX4251 = (WX4257&WX4252);
assign WX3294 = (WX3231&RESET);
assign II27705 = ((~WX8394))|((~_2275_));
assign II26986 = ((~WX8529))|((~II26978));
assign II3287 = ((~WX598))|((~II3286));
assign WX2085 = (WX2022&RESET);
assign II34879 = ((~II34881))|((~II34882));
assign WX4659 = (WX4596&RESET);
assign WX10959 = ((~WX11187));
assign WX8401 = ((~WX8657));
assign WX9311 = (WX9317&WX9312);
assign WX8890 = ((~II27317))|((~II27318));
assign II18704 = ((~II18706))|((~II18707));
assign II34152 = ((~WX11345))|((~WX10997));
assign II30705 = ((~WX10053))|((~WX9740));
assign WX6207 = (WX6206&WX6177);
assign WX9301 = (WX11461&WX9302);
assign WX6223 = ((~WX6177));
assign II2228 = ((~II2203))|((~II2227));
assign WX8124 = (WX8931&WX8125);
assign WX5323 = (_2228_&WX6176);
assign II19564 = ((~_2232_))|((~II19562));
assign WX7848 = ((~WX7847));
assign WX8175 = (_2273_&WX8762);
assign WX5484 = (WX5482)|(WX5481);
assign WX1298 = (WX1249&WX1263);
assign WX4631 = (WX4568&RESET);
assign II34925 = ((~II34935))|((~II34936));
assign II23376 = ((~WX7068))|((~WX6996));
assign II31564 = ((~WX9664))|((~II31563));
assign II2105 = ((~II2095))|((~II2103));
assign II7148 = ((~WX1880))|((~WX1792));
assign WX9791 = (WX9728&RESET);
assign WX1959 = (WX1495&RESET);
assign WX7337 = (WX7274&RESET);
assign II2825 = ((~WX1002))|((~WX699));
assign WX10038 = ((~WX10037));
assign II22098 = ((~II22073))|((~II22097));
assign II22175 = ((~WX7184))|((~II22167));
assign II14955 = ((~II14931))|((~II14947));
assign II6921 = ((~II6931))|((~II6932));
assign WX5317 = ((~WX5308));
assign WX8155 = ((~WX8146));
assign WX8104 = (WX8102)|(WX8101);
assign II34199 = ((~WX11127))|((~II34198));
assign II11454 = ((~WX3131))|((~II11452));
assign WX11526 = (WX11525&WX11349);
assign WX9269 = (WX9275&WX9270);
assign II2638 = ((~II2640))|((~II2641));
assign WX623 = ((~WX859));
assign WX7969 = (WX8267&WX8762);
assign WX7509 = ((~WX7470));
assign WX4665 = (WX4602&RESET);
assign WX10187 = (WX10185)|(WX10184);
assign WX9424 = ((~WX10054));
assign WX4480 = ((~WX4448));
assign WX2089 = (WX2026&RESET);
assign WX3196 = ((~WX3164));
assign WX1664 = (WX1675&WX2296);
assign WX9537 = (WX9540&RESET);
assign WX1403 = (WX3633&WX1404);
assign WX6706 = ((~WX7469));
assign WX5783 = ((~WX5751));
assign WX2201 = ((~II6264))|((~II6265));
assign II19164 = ((~WX5759))|((~II19163));
assign WX6431 = ((~II19710))|((~II19711));
assign II22439 = ((~II22414))|((~II22438));
assign WX1619 = (WX1617)|(WX1616);
assign WX3607 = (WX3606&WX3591);
assign II23247 = ((~WX7058))|((~II23246));
assign II2235 = ((~II2237))|((~II2238));
assign II35590 = ((~WX10960))|((~II35589));
assign WX9422 = (WX9433&WX10054);
assign WX11384 = ((~WX11383));
assign WX6546 = (_2265_&WX7469);
assign WX8849 = (WX8848&WX8763);
assign II26466 = ((~II26468))|((~II26469));
assign WX1768 = ((~WX2297));
assign WX6620 = (WX6966&WX7469);
assign WX2236 = ((~WX2235));
assign II26685 = ((~WX8573))|((~II26684));
assign II14919 = ((~WX4774))|((~II14917));
assign WX8039 = (WX8277&WX8762);
assign II15237 = ((~WX4472))|((~II15236));
assign II10477 = ((~II10479))|((~II10480));
assign WX7965 = (_2288_&WX8762);
assign II18785 = ((~WX5867))|((~II18783));
assign WX8840 = ((~WX8839));
assign II34486 = ((~II34476))|((~II34484));
assign II14885 = ((~II14887))|((~II14888));
assign WX3615 = (WX3169&WX3616);
assign WX7377 = ((~II22408))|((~II22409));
assign II19578 = ((~_2230_))|((~II19576));
assign WX11188 = (WX11125&RESET);
assign II18079 = ((~II18069))|((~II18077));
assign II7499 = ((~II7489))|((~II7497));
assign WX5369 = (WX5679&WX6176);
assign II15634 = ((~WX4505))|((~_2189_));
assign II10710 = ((~II10712))|((~II10713));
assign WX5233 = ((~WX5224));
assign WX8208 = (WX8973&WX8209);
assign WX4464 = ((~WX4432));
assign II6280 = ((~WX2020))|((~II6279));
assign WX2113 = (WX2050&RESET);
assign WX9639 = ((~WX9607));
assign II18038 = ((~II18040))|((~II18041));
assign II11284 = ((~WX3183))|((~II11283));
assign WX3312 = (WX3249&RESET);
assign WX5619 = ((~WX6176));
assign II22432 = ((~WX7264))|((~II22431));
assign WX5214 = (WX5212)|(WX5211);
assign WX10251 = ((~WX10250));
assign WX2948 = (WX5052&WX2949);
assign WX2835 = (_2157_&WX3590);
assign WX8035 = (_2283_&WX8762);
assign WX2943 = (WX2954&WX3589);
assign WX10491 = (WX10502&WX11347);
assign WX9983 = ((~WX9967));
assign WX7435 = ((~WX7368));
assign WX7042 = ((~WX7424));
assign WX10498 = (WX10496)|(WX10495);
assign WX2669 = ((~WX3590));
assign II22462 = ((~WX7266))|((~WX7330));
assign II2361 = ((~WX1001))|((~II2360));
assign WX11471 = (WX10941&WX11472);
assign II26249 = ((~II26251))|((~II26252));
assign WX10802 = (WX10800)|(WX10799);
assign WX6296 = ((~WX6295));
assign WX1985 = (WX1677&RESET);
assign WX4904 = ((~WX4903));
assign WX4287 = (WX5073&WX4288);
assign WX8055 = ((~WX8762));
assign II18134 = ((~WX5825))|((~II18132));
assign WX7984 = (WX8861&WX7985);
assign WX7092 = ((~WX7332));
assign WX2240 = ((~WX2239));
assign WX6534 = ((~WX7469));
assign II11400 = ((~WX3192))|((~WX3123));
assign II10131 = ((~II10121))|((~II10129));
assign II15559 = ((~_2200_))|((~II15557));
assign WX10625 = (WX10863&WX11348);
assign WX1627 = (WX3745&WX1628);
assign WX4882 = ((~WX4878));
assign WX5097 = (WX4489&WX5098);
assign WX9839 = (WX9776&RESET);
assign II31578 = ((~WX9666))|((~II31577));
assign II27499 = ((~II27501))|((~II27502));
assign II19528 = ((~_2208_))|((~II19527));
assign WX7674 = ((~II23455))|((~II23456));
assign WX6732 = (WX6982&WX7469);
assign II6622 = ((~II6612))|((~II6620));
assign WX7255 = (WX7192&RESET);
assign II30455 = ((~II30465))|((~II30466));
assign II6093 = ((~WX2008))|((~II6085));
assign WX6535 = (WX6533)|(WX6532);
assign II15431 = ((~WX4487))|((~WX4420));
assign WX654 = (WX118&RESET);
assign WX772 = (WX709&RESET);
assign II19725 = ((~_2206_))|((~II19723));
assign WX303 = ((~WX1003));
assign II26590 = ((~II26592))|((~II26593));
assign II15578 = ((~WX4497))|((~_2197_));
assign II3352 = ((~WX603))|((~II3351));
assign WX8734 = ((~WX8664));
assign WX3526 = ((~WX3506));
assign WX10113 = ((~II31192))|((~II31193));
assign WX6158 = ((~WX6083));
assign WX8685 = ((~II26878))|((~II26879));
assign II30094 = ((~II30084))|((~II30092));
assign II3132 = ((~WX497))|((~II3130));
assign WX11395 = ((~WX11349));
assign II30605 = ((~II30595))|((~II30603));
assign WX9019 = ((~II27734))|((~II27735));
assign WX6826 = (_2245_&WX7469);
assign II11693 = ((~WX3223))|((~II11692));
assign WX6768 = ((~WX7468));
assign II7561 = ((~WX1910))|((~_2134_));
assign II10005 = ((~WX3295))|((~II9997));
assign WX9703 = (WX9155&RESET);
assign WX4428 = ((~WX4846));
assign II22890 = ((~II22880))|((~II22888));
assign WX10141 = ((~II31244))|((~II31245));
assign II31504 = ((~II31506))|((~II31507));
assign WX5061 = (WX5060&WX4884);
assign WX10876 = (WX10879&RESET);
assign WX5000 = ((~WX4884));
assign II2305 = ((~WX729))|((~II2297));
assign WX5752 = ((~WX5720));
assign WX6932 = ((~WX6923));
assign WX1641 = (WX3752&WX1642);
assign WX3016 = (WX3014)|(WX3013);
assign II10409 = ((~WX3321))|((~II10408));
assign II31322 = ((~WX9649))|((~II31321));
assign II18009 = ((~WX6173))|((~II18008));
assign II2191 = ((~WX849))|((~II2189));
assign WX1355 = ((~WX1354));
assign WX5240 = (WX7491&WX5241);
assign WX6385 = (WX6383)|(WX6382);
assign WX10922 = ((~WX11305));
assign II22926 = ((~II22928))|((~II22929));
assign II2947 = ((~II2957))|((~II2958));
assign WX6502 = ((~WX7468));
assign II30676 = ((~WX9738))|((~II30674));
assign II2312 = ((~II2314))|((~II2315));
assign II11322 = ((~WX3186))|((~WX3111));
assign WX852 = (WX789&RESET);
assign II34135 = ((~II34137))|((~II34138));
assign WX7499 = ((~II23130))|((~II23131));
assign II22771 = ((~II22773))|((~II22774));
assign WX6644 = (_2258_&WX7469);
assign WX4477 = ((~WX4445));
assign II22539 = ((~II22541))|((~II22542));
assign WX7074 = ((~WX7042));
assign WX11004 = (WX10504&RESET);
assign WX4436 = ((~WX4862));
assign WX1155 = (WX601&WX1156);
assign II30543 = ((~II30533))|((~II30541));
assign II14025 = ((~II14001))|((~II14017));
assign II26522 = ((~WX8499))|((~II26521));
assign WX10565 = (_2351_&WX11348);
assign WX10225 = ((~II31400))|((~II31401));
assign II10089 = ((~II10099))|((~II10100));
assign II18875 = ((~II18877))|((~II18878));
assign II3195 = ((~WX591))|((~WX507));
assign WX4139 = (WX4145&WX4140);
assign WX4057 = (WX4055)|(WX4054);
assign II19549 = ((~WX5785))|((~II19548));
assign WX2845 = (WX2856&WX3589);
assign WX1586 = ((~WX2297));
assign II22610 = ((~WX7212))|((~II22609));
assign WX58 = (DATA_9_30&WX59);
assign WX7928 = (WX8833&WX7929);
assign WX3238 = (WX2690&RESET);
assign WX2427 = (WX1891&WX2428);
assign WX6232 = ((~WX6231));
assign WX10832 = (WX10835&RESET);
assign II26957 = ((~II26947))|((~II26955));
assign II10456 = ((~II10446))|((~II10454));
assign II19583 = ((~WX5790))|((~_2229_));
assign II34563 = ((~WX11087))|((~II34562));
assign II3196 = ((~WX591))|((~II3195));
assign II7702 = ((~WX1933))|((~II7701));
assign II2206 = ((~WX1001))|((~II2205));
assign II2345 = ((~WX795))|((~II2344));
assign II22911 = ((~II22913))|((~II22914));
assign II35431 = ((~WX10950))|((~II35430));
assign WX327 = ((~WX318));
assign II22299 = ((~WX7192))|((~II22291));
assign II18456 = ((~II18458))|((~II18459));
assign WX3720 = (WX3184&WX3721);
assign WX7034 = ((~WX7408));
assign WX11640 = (WX11575&WX11607);
assign II18714 = ((~II18704))|((~II18712));
assign WX2433 = (WX2432&WX2298);
assign WX6901 = (WX7673&WX6902);
assign WX11510 = ((~WX11509));
assign II31008 = ((~II30998))|((~II31006));
assign II30843 = ((~II30845))|((~II30846));
assign WX7706 = ((~II23589))|((~II23590));
assign II34448 = ((~WX11207))|((~II34446));
assign WX5427 = ((~WX6176));
assign WX8704 = ((~WX8681));
assign II35172 = ((~WX10841))|((~II35170));
assign WX5459 = (WX5470&WX6175);
assign II6108 = ((~II6084))|((~II6100));
assign WX11508 = (WX11506)|(WX11505);
assign WX2828 = (WX2826)|(WX2825);
assign WX4737 = (WX4674&RESET);
assign WX3688 = ((~WX3687));
assign II11090 = ((~WX3075))|((~II11088));
assign WX8792 = ((~II27135))|((~II27136));
assign II18644 = ((~WX5985))|((~II18643));
assign WX5118 = ((~II15565))|((~II15566));
assign WX5581 = ((~WX6176));
assign II34339 = ((~WX11345))|((~II34338));
assign II22066 = ((~II22042))|((~II22058));
assign WX2979 = (WX3121&WX3590);
assign WX144 = (WX142)|(WX141);
assign WX3924 = ((~WX4883));
assign II22573 = ((~WX7146))|((~II22571));
assign WX8799 = ((~II27148))|((~II27149));
assign II35738 = ((~_2335_))|((~II35736));
assign WX9296 = (WX9307&WX10054);
assign II2925 = ((~WX769))|((~II2917));
assign II31613 = ((~WX9671))|((~II31612));
assign WX6675 = (WX6673)|(WX6672);
assign WX1654 = (_2117_&WX2297);
assign WX4178 = ((~WX4169));
assign WX10247 = (WX10246&WX10056);
assign WX9517 = (WX9515)|(WX9514);
assign WX3943 = (WX3949&WX3944);
assign WX403 = (_2082_&WX1004);
assign WX1467 = ((~WX1466));
assign II34360 = ((~II34336))|((~II34352));
assign WX5615 = ((~WX6175));
assign II18061 = ((~II18037))|((~II18053));
assign II18723 = ((~WX5863))|((~II18721));
assign II15485 = ((~WX4506))|((~_2204_));
assign II2792 = ((~II2802))|((~II2803));
assign II26149 = ((~WX8475))|((~II26141));
assign WX8695 = ((~WX8694));
assign WX2390 = ((~II7227))|((~II7228));
assign II26637 = ((~II26639))|((~II26640));
assign WX10214 = ((~WX10056));
assign WX6670 = ((~WX7468));
assign II10403 = ((~WX3257))|((~II10401));
assign WX2661 = ((~WX2652));
assign II18837 = ((~II18812))|((~II18836));
assign WX11497 = ((~II35366))|((~II35367));
assign II30852 = ((~II30827))|((~II30851));
assign II27213 = ((~WX8348))|((~II27212));
assign WX62 = ((~WX61));
assign II22857 = ((~WX7228))|((~II22849));
assign II22820 = ((~WX7467))|((~II22819));
assign II18356 = ((~WX5903))|((~II18348));
assign II11114 = ((~WX3170))|((~WX3079));
assign II23618 = ((~_2257_))|((~II23616));
assign WX2952 = (WX3759&WX2953);
assign WX10430 = (WX11377&WX10431);
assign WX1973 = (WX1593&RESET);
assign WX6188 = ((~WX6177));
assign II2083 = ((~WX651))|((~II2081));
assign WX4509 = ((~WX4752));
assign WX10540 = (WX10538)|(WX10537);
assign WX6685 = (WX6683)|(WX6682);
assign WX4959 = (WX4957)|(WX4956);
assign WX358 = (WX364&WX359);
assign WX6109 = ((~WX6108));
assign WX4169 = (WX4167)|(WX4166);
assign II6126 = ((~II6116))|((~II6124));
assign WX2508 = ((~WX2507));
assign II14166 = ((~WX4598))|((~II14165));
assign WX8764 = ((~II27083))|((~II27084));
assign II23311 = ((~WX7063))|((~WX6986));
assign WX6390 = (WX5782&WX6391);
assign WX9407 = ((~WX9406));
assign II35724 = ((~_2338_))|((~II35722));
assign II34369 = ((~WX11345))|((~WX11011));
assign II3325 = ((~WX601))|((~WX527));
assign WX6773 = (WX6771)|(WX6770);
assign WX5414 = (WX5412)|(WX5411);
assign II2919 = ((~WX1002))|((~II2918));
assign WX11349 = ((~WX11340));
assign II34190 = ((~WX11063))|((~II34182));
assign WX9479 = (WX9485&WX9480);
assign WX2863 = (_2155_&WX3590);
assign WX5403 = (WX5414&WX6175);
assign II26745 = ((~II26747))|((~II26748));
assign WX3693 = ((~WX3591));
assign WX2891 = (_2153_&WX3590);
assign II14187 = ((~II14197))|((~II14198));
assign WX4356 = (WX4426&WX4883);
assign WX3672 = ((~WX3591));
assign WX126 = (WX124)|(WX123);
assign WX10916 = ((~WX11293));
assign WX5768 = ((~WX5736));
assign WX1193 = ((~WX1192));
assign WX11458 = ((~WX11349));
assign WX4502 = ((~WX4738));
assign WX1754 = ((~WX2297));
assign WX4810 = ((~II14987))|((~II14988));
assign WX2772 = (WX2770)|(WX2769);
assign II14910 = ((~WX4646))|((~II14909));
assign WX6379 = ((~WX6378));
assign WX3687 = (WX3685)|(WX3684);
assign II30665 = ((~II30641))|((~II30657));
assign II18518 = ((~II18520))|((~II18521));
assign WX6285 = (WX5767&WX6286);
assign WX9508 = ((~WX10054));
assign WX1699 = (WX1697)|(WX1696);
assign II30567 = ((~WX9922))|((~II30565));
assign WX7406 = ((~WX7405));
assign WX3044 = (WX3042)|(WX3041);
assign II6016 = ((~II5991))|((~II6015));
assign WX2779 = (_2161_&WX3590);
assign WX56 = (WX54)|(WX53);
assign II22673 = ((~II22663))|((~II22671));
assign II22182 = ((~II22184))|((~II22185));
assign II19372 = ((~WX5775))|((~II19371));
assign II6720 = ((~II6722))|((~II6723));
assign WX7365 = ((~II22036))|((~II22037));
assign WX1748 = (WX1759&WX2296);
assign WX8126 = (WX8124)|(WX8123);
assign WX9197 = ((~WX9196));
assign WX6862 = ((~WX6853));
assign II35380 = ((~WX10873))|((~II35378));
assign II30722 = ((~WX9932))|((~II30720));
assign II15538 = ((~_2203_))|((~II15536));
assign II6630 = ((~WX2170))|((~II6628));
assign WX9159 = (WX9157)|(WX9156);
assign WX8480 = (WX8417&RESET);
assign II2858 = ((~WX701))|((~II2856));
assign WX10652 = (WX10650)|(WX10649);
assign II22836 = ((~WX7354))|((~II22834));
assign II23351 = ((~WX7066))|((~II23350));
assign WX343 = (WX354&WX1003);
assign WX11306 = ((~WX11275));
assign II26624 = ((~WX8633))|((~II26622));
assign WX1494 = ((~WX1485));
assign WX10209 = ((~WX10208));
assign WX2860 = (WX2866&WX2861);
assign WX7409 = ((~WX7387));
assign II6460 = ((~WX1968))|((~II6458));
assign WX317 = ((~WX1003));
assign II23708 = ((~WX7102))|((~II23707));
assign WX9366 = (WX9377&WX10054);
assign WX8500 = (WX8437&RESET);
assign WX7601 = (WX7599)|(WX7598);
assign WX4940 = ((~WX4939));
assign WX9091 = (WX11356&WX9092);
assign WX10212 = (WX10211&WX10056);
assign II34050 = ((~II34026))|((~II34042));
assign II6637 = ((~II6627))|((~II6635));
assign II10687 = ((~WX3339))|((~II10679));
assign II34851 = ((~WX11233))|((~II34849));
assign WX7592 = (WX7062&WX7593);
assign WX5530 = (WX5536&WX5531);
assign WX3843 = ((~II11686))|((~II11687));
assign II6224 = ((~II6226))|((~II6227));
assign WX7223 = (WX7160&RESET);
assign II34185 = ((~WX10999))|((~II34183));
assign II10093 = ((~WX3237))|((~II10091));
assign WX1206 = (WX1204)|(WX1203);
assign II23350 = ((~WX7066))|((~WX6992));
assign II15342 = ((~WX4406))|((~II15340));
assign WX5445 = (WX5456&WX6175);
assign WX2477 = ((~WX2298));
assign WX2147 = (WX2084&RESET);
assign WX832 = (WX769&RESET);
assign II10648 = ((~II10650))|((~II10651));
assign II31001 = ((~WX9950))|((~II30999));
assign WX310 = (DATA_9_12&WX311);
assign WX5165 = (WX5111&WX5142);
assign II35378 = ((~WX10946))|((~WX10873));
assign WX9246 = ((~WX10055));
assign II27394 = ((~WX8362))|((~WX8291));
assign WX3767 = ((~II11388))|((~II11389));
assign WX11666 = (WX11581&WX11607);
assign WX2474 = ((~II7383))|((~II7384));
assign WX7446 = ((~WX7445));
assign II22975 = ((~WX7467))|((~II22974));
assign WX4070 = ((~WX4882));
assign WX1059 = (WX1057)|(WX1056);
assign II34307 = ((~WX11345))|((~WX11007));
assign II10594 = ((~WX3333))|((~II10586));
assign WX5491 = (_2216_&WX6176);
assign WX9350 = ((~WX9341));
assign WX3789 = (WX3788&WX3591);
assign WX2676 = ((~WX2675));
assign WX3989 = (WX6219&WX3990);
assign WX1146 = ((~II3313))|((~II3314));
assign WX9252 = ((~WX9243));
assign WX2969 = ((~WX2960));
assign WX3187 = ((~WX3155));
assign WX5255 = ((~WX6176));
assign II30889 = ((~II30899))|((~II30900));
assign II34887 = ((~II34863))|((~II34879));
assign WX8138 = (WX8938&WX8139);
assign WX3639 = ((~WX3638));
assign II10904 = ((~WX3353))|((~II10896));
assign WX10137 = ((~WX10056));
assign II15698 = ((~WX4516))|((~II15697));
assign II6333 = ((~II6335))|((~II6336));
assign WX11434 = ((~II35249))|((~II35250));
assign WX9616 = ((~WX9986));
assign WX9439 = (WX9437)|(WX9436);
assign WX992 = ((~WX914));
assign II30131 = ((~WX9830))|((~WX9894));
assign WX9174 = (_2326_&WX10055);
assign II30955 = ((~WX9756))|((~II30953));
assign II6830 = ((~WX2295))|((~WX1992));
assign WX5129 = ((~II15642))|((~II15643));
assign WX1236 = ((~II3529))|((~II3530));
assign WX8836 = (WX8348&WX8837);
assign II3508 = ((~_2080_))|((~II3507));
assign II30025 = ((~WX9696))|((~II30023));
assign WX3630 = ((~WX3591));
assign WX5537 = (WX5703&WX6176);
assign WX6412 = ((~II19577))|((~II19578));
assign WX9765 = (WX9702&RESET);
assign WX8172 = (WX8178&WX8173);
assign WX4820 = ((~WX4819));
assign WX11154 = (WX11091&RESET);
assign WX2379 = ((~WX2298));
assign II26280 = ((~II26282))|((~II26283));
assign II7188 = ((~WX1883))|((~II7187));
assign II6932 = ((~II6922))|((~II6930));
assign WX233 = ((~WX1003));
assign WX6133 = ((~WX6132));
assign WX7765 = (WX7713&WX7728);
assign WX892 = (WX829&RESET);
assign WX5329 = ((~WX6176));
assign WX10269 = (WX9661&WX10270);
assign WX8745 = ((~WX8744));
assign WX121 = ((~WX1003));
assign II30551 = ((~WX10053))|((~II30550));
assign WX3756 = ((~WX3591));
assign WX9213 = (WX9219&WX9214);
assign II2281 = ((~II2283))|((~II2284));
assign WX7427 = ((~WX7396));
assign WX4707 = (WX4644&RESET);
assign WX8713 = ((~WX8712));
assign II34076 = ((~WX11183))|((~II34074));
assign II30549 = ((~II30551))|((~II30552));
assign II26707 = ((~WX8511))|((~II26699));
assign WX8953 = ((~II27434))|((~II27435));
assign II7490 = ((~WX1925))|((~_2140_));
assign WX4338 = (_2174_&WX4883);
assign WX6238 = (WX6236)|(WX6235);
assign WX8998 = ((~II27587))|((~II27588));
assign WX6873 = (WX7659&WX6874);
assign WX5886 = (WX5823&RESET);
assign II27501 = ((~WX8385))|((~II27500));
assign WX1434 = (WX1792&WX2297);
assign II23590 = ((~_2261_))|((~II23588));
assign WX3390 = (WX3327&RESET);
assign II6334 = ((~WX2294))|((~WX1960));
assign II30977 = ((~II30967))|((~II30975));
assign WX3504 = ((~II10579))|((~II10580));
assign WX180 = (WX2375&WX181);
assign II18843 = ((~II18853))|((~II18854));
assign II10516 = ((~II10492))|((~II10508));
assign WX11096 = (WX11033&RESET);
assign WX5279 = ((~WX6175));
assign WX4677 = (WX4614&RESET);
assign II7150 = ((~WX1792))|((~II7148));
assign WX5482 = (WX6317&WX5483);
assign WX7739 = (WX7724&WX7728);
assign WX10402 = (WX11363&WX10403);
assign WX7599 = (WX7063&WX7600);
assign II35393 = ((~WX10875))|((~II35391));
assign II34896 = ((~WX11346))|((~WX11045));
assign WX3699 = (WX3181&WX3700);
assign WX2249 = ((~WX2221));
assign II6776 = ((~WX2052))|((~II6775));
assign WX1219 = ((~WX1005));
assign WX5387 = ((~WX5378));
assign WX9034 = (WX9016&WX9021);
assign WX4335 = (WX4341&WX4336);
assign II35131 = ((~WX10927))|((~WX10835));
assign II35598 = ((~_2358_))|((~II35596));
assign WX6883 = (WX8959&WX6884);
assign II34223 = ((~II34213))|((~II34221));
assign II3366 = ((~WX533))|((~II3364));
assign WX5428 = (WX5426)|(WX5425);
assign WX11431 = (WX11429)|(WX11428);
assign II30579 = ((~II30589))|((~II30590));
assign II3404 = ((~WX607))|((~II3403));
assign WX10614 = (WX10612)|(WX10611);
assign WX4621 = (WX4558&RESET);
assign II30830 = ((~WX10053))|((~II30829));
assign II30820 = ((~II30796))|((~II30812));
assign WX10456 = (WX10454)|(WX10453);
assign WX3827 = ((~II11574))|((~II11575));
assign WX11515 = (WX11513)|(WX11512);
assign II26312 = ((~WX8549))|((~WX8613));
assign II22455 = ((~WX7202))|((~II22454));
assign II6364 = ((~II6366))|((~II6367));
assign WX5286 = (WX6219&WX5287);
assign II22166 = ((~II22176))|((~II22177));
assign II18829 = ((~WX5997))|((~WX6061));
assign II3628 = ((~_2091_))|((~II3626));
assign II2679 = ((~II2669))|((~II2677));
assign WX1045 = (WX1043)|(WX1042);
assign WX10992 = (WX10420&RESET);
assign WX1624 = ((~WX2296));
assign II34960 = ((~WX11049))|((~II34958));
assign II30404 = ((~II30394))|((~II30402));
assign WX5404 = (WX5410&WX5405);
assign WX3755 = (WX3189&WX3756);
assign WX9202 = (_2324_&WX10055);
assign WX5217 = ((~WX6176));
assign II3501 = ((~WX639))|((~II3500));
assign WX6916 = ((~WX7469));
assign WX5260 = (WX5258)|(WX5257);
assign WX2555 = ((~II7716))|((~II7717));
assign WX426 = ((~WX425));
assign WX10085 = ((~II31140))|((~II31141));
assign II2693 = ((~II2668))|((~II2692));
assign WX9978 = ((~II30883))|((~II30884));
assign WX7533 = ((~WX7532));
assign WX7785 = (WX7703&WX7728);
assign II7590 = ((~WX1914))|((~II7589));
assign II34641 = ((~II34631))|((~II34639));
assign II18441 = ((~II18443))|((~II18444));
assign WX5307 = ((~WX6175));
assign WX8946 = ((~II27421))|((~II27422));
assign WX2388 = ((~WX2387));
assign WX6277 = (WX6276&WX6177);
assign WX4949 = (WX4948&WX4884);
assign WX6403 = ((~II19498))|((~II19499));
assign WX2383 = ((~II7214))|((~II7215));
assign WX7237 = (WX7174&RESET);
assign WX2496 = (WX2495&WX2298);
assign WX11656 = (WX11586&WX11607);
assign WX5745 = ((~WX6123));
assign II34719 = ((~II34709))|((~II34717));
assign II3530 = ((~_2106_))|((~II3528));
assign II19178 = ((~WX5673))|((~II19176));
assign WX9625 = ((~WX10004));
assign WX10824 = (WX10822)|(WX10821);
assign WX6842 = ((~WX7469));
assign WX3902 = (WX3826&WX3849);
assign WX5568 = (WX5566)|(WX5565);
assign WX8321 = ((~WX8753));
assign WX3538 = ((~WX3512));
assign WX8875 = ((~WX8874));
assign WX1184 = ((~WX1005));
assign WX285 = ((~WX276));
assign WX884 = (WX821&RESET);
assign WX6866 = ((~WX7468));
assign WX11392 = ((~II35171))|((~II35172));
assign WX9996 = ((~WX9995));
assign WX8388 = ((~WX8631));
assign II27742 = ((~_2269_))|((~II27740));
assign WX8881 = ((~WX8880));
assign WX7400 = ((~WX7399));
assign WX1153 = ((~II3326))|((~II3327));
assign II7604 = ((~WX1916))|((~II7603));
assign II6953 = ((~II6955))|((~II6956));
assign WX6118 = ((~WX6095));
assign II10229 = ((~II10231))|((~II10232));
assign WX3518 = ((~WX3502));
assign II34355 = ((~WX11201))|((~II34353));
assign WX11420 = ((~II35223))|((~II35224));
assign WX1729 = (WX2501&WX1730);
assign WX7243 = (WX7180&RESET);
assign II6761 = ((~II6751))|((~II6759));
assign WX8408 = (WX7848&RESET);
assign WX3180 = ((~WX3148));
assign WX6399 = (WX6397)|(WX6396);
assign WX2173 = (WX2110&RESET);
assign WX4805 = ((~II14832))|((~II14833));
assign II31412 = ((~WX9656))|((~WX9586));
assign II26173 = ((~WX8759))|((~WX8413));
assign II10113 = ((~II10089))|((~II10105));
assign II19359 = ((~WX5774))|((~II19358));
assign II27122 = ((~WX8341))|((~II27121));
assign WX950 = ((~WX925));
assign WX10638 = (WX10636)|(WX10635);
assign WX2870 = (WX2868)|(WX2867);
assign WX4767 = (WX4704&RESET);
assign WX320 = (WX2445&WX321);
assign WX1743 = (WX2508&WX1744);
assign WX4162 = ((~WX4883));
assign II14771 = ((~II14761))|((~II14769));
assign WX276 = (WX274)|(WX273);
assign WX10132 = ((~WX10131));
assign WX10943 = ((~WX10911));
assign WX9430 = (WX9584&WX10055);
assign WX8029 = ((~WX8020));
assign WX1276 = (WX1258&WX1263);
assign WX6875 = (WX6873)|(WX6872);
assign II2630 = ((~II2606))|((~II2622));
assign WX9209 = (WX9207)|(WX9206);
assign II26392 = ((~WX8427))|((~II26390));
assign WX8848 = ((~II27239))|((~II27240));
assign WX7521 = (WX7520&WX7470);
assign II10672 = ((~II10647))|((~II10671));
assign II26281 = ((~WX8547))|((~WX8611));
assign II30984 = ((~WX10053))|((~WX9758));
assign WX6428 = ((~II19689))|((~II19690));
assign WX9707 = (WX9183&RESET);
assign WX7249 = (WX7186&RESET);
assign WX8716 = ((~WX8687));
assign II23169 = ((~WX7052))|((~II23168));
assign II31308 = ((~WX9648))|((~WX9570));
assign WX1892 = ((~WX1860));
assign WX5413 = ((~WX6176));
assign WX7390 = ((~II22811))|((~II22812));
assign WX1139 = ((~II3300))|((~II3301));
assign II34894 = ((~II34904))|((~II34905));
assign WX10846 = (WX10849&RESET);
assign WX6476 = (WX6418&WX6435);
assign WX9819 = (WX9756&RESET);
assign WX5261 = ((~WX5252));
assign WX10914 = ((~WX11289));
assign WX141 = (WX499&WX1004);
assign II26894 = ((~WX8523))|((~II26893));
assign II10773 = ((~WX3588))|((~WX3281));
assign II27459 = ((~WX8367))|((~WX8301));
assign II2027 = ((~WX711))|((~II2026));
assign WX4206 = ((~WX4197));
assign WX4825 = ((~WX4802));
assign WX9434 = ((~WX9425));
assign WX10975 = ((~WX11219));
assign WX3158 = ((~WX3535));
assign WX5892 = (WX5829&RESET);
assign II18823 = ((~II18813))|((~II18821));
assign WX7225 = (WX7162&RESET);
assign WX10312 = ((~II31739))|((~II31740));
assign WX5388 = ((~WX5387));
assign WX10477 = (WX10488&WX11347);
assign WX11178 = (WX11115&RESET);
assign WX9763 = (WX9700&RESET);
assign WX2453 = ((~II7344))|((~II7345));
assign WX3697 = ((~II11258))|((~II11259));
assign II14227 = ((~WX4602))|((~II14219));
assign WX10140 = ((~WX10139));
assign WX2607 = (WX2534&WX2556);
assign WX5332 = ((~WX5331));
assign WX486 = (WX489&RESET);
assign II2344 = ((~WX795))|((~WX859));
assign WX5784 = ((~WX6009));
assign WX9337 = ((~WX9336));
assign II2756 = ((~II2746))|((~II2754));
assign WX3690 = ((~II11245))|((~II11246));
assign WX2061 = (WX1998&RESET);
assign WX2421 = ((~WX2298));
assign WX11288 = ((~WX11266));
assign WX2402 = ((~WX2401));
assign II35352 = ((~WX10944))|((~WX10869));
assign II10849 = ((~II10851))|((~II10852));
assign WX1209 = ((~II3430))|((~II3431));
assign WX1396 = ((~WX1387));
assign WX9352 = (WX9363&WX10054);
assign WX5130 = ((~II15649))|((~II15650));
assign II18396 = ((~WX5969))|((~II18395));
assign WX349 = ((~WX1004));
assign WX9215 = (WX9213)|(WX9212);
assign WX7569 = ((~II23260))|((~II23261));
assign WX1757 = (WX2515&WX1758);
assign WX11472 = ((~WX11349));
assign WX2200 = ((~II6233))|((~II6234));
assign II34600 = ((~II34602))|((~II34603));
assign II31310 = ((~WX9570))|((~II31308));
assign II30154 = ((~WX9768))|((~II30146));
assign WX3183 = ((~WX3151));
assign WX5274 = (WX5272)|(WX5271);
assign II27396 = ((~WX8291))|((~II27394));
assign WX8165 = (WX8295&WX8762);
assign II7370 = ((~WX1897))|((~II7369));
assign WX10621 = (_2347_&WX11348);
assign WX1934 = ((~WX2188));
assign WX1048 = ((~II3131))|((~II3132));
assign WX245 = (WX256&WX1003);
assign WX997 = ((~TM0));
assign WX11650 = (WX11589&WX11607);
assign WX10827 = ((~WX10829));
assign II10665 = ((~WX3401))|((~II10664));
assign WX2446 = ((~II7331))|((~II7332));
assign II11603 = ((~_2161_))|((~II11601));
assign II6179 = ((~WX2294))|((~WX1950));
assign WX1930 = ((~WX2180));
assign WX8092 = (WX10210&WX8093);
assign II14559 = ((~II14569))|((~II14570));
assign WX7604 = ((~II23325))|((~II23326));
assign WX5259 = ((~WX6176));
assign WX8127 = ((~WX8118));
assign II10224 = ((~II10214))|((~II10222));
assign II34502 = ((~II34492))|((~II34500));
assign II14941 = ((~WX4648))|((~II14940));
assign WX9335 = (WX9333)|(WX9332);
assign WX2303 = (WX2301)|(WX2300);
assign WX4814 = ((~WX4813));
assign WX2811 = (WX3097&WX3590);
assign II30208 = ((~II30210))|((~II30211));
assign II19704 = ((~_2210_))|((~II19702));
assign WX1351 = (WX2312&WX1352);
assign II27552 = ((~WX8370))|((~II27551));
assign WX10628 = (WX10626)|(WX10625);
assign II34617 = ((~WX11346))|((~WX11027));
assign II6937 = ((~II6939))|((~II6940));
assign II34222 = ((~WX11065))|((~II34221));
assign WX3786 = ((~WX3785));
assign WX4498 = ((~WX4730));
assign II19423 = ((~WX5779))|((~WX5711));
assign WX9172 = ((~WX10054));
assign WX3215 = ((~WX3457));
assign WX3765 = ((~WX3764));
assign WX11432 = ((~WX11431));
assign WX10946 = ((~WX10914));
assign II34858 = ((~II34848))|((~II34856));
assign II22879 = ((~II22889))|((~II22890));
assign II22014 = ((~WX7466))|((~II22013));
assign WX8192 = (WX8190)|(WX8189);
assign WX5686 = (WX5689&RESET);
assign WX2964 = (WX2962)|(WX2961);
assign WX10309 = ((~II31718))|((~II31719));
assign WX10908 = ((~WX11277));
assign WX1125 = ((~II3274))|((~II3275));
assign WX1207 = ((~WX1206));
assign II7344 = ((~WX1895))|((~II7343));
assign WX7703 = ((~II23568))|((~II23569));
assign WX11441 = ((~II35262))|((~II35263));
assign II10603 = ((~WX3397))|((~II10602));
assign WX11410 = (WX11408)|(WX11407);
assign II27559 = ((~WX8371))|((~II27558));
assign WX3802 = ((~II11453))|((~II11454));
assign II14377 = ((~WX4548))|((~II14375));
assign WX1863 = ((~WX2238));
assign WX5488 = (WX5494&WX5489);
assign WX6170 = ((~TM0));
assign WX1189 = (WX1188&WX1005);
assign II14786 = ((~WX4638))|((~II14785));
assign WX8145 = ((~WX8761));
assign WX10609 = ((~WX11348));
assign II2390 = ((~II2392))|((~II2393));
assign WX2472 = ((~WX2471));
assign II2524 = ((~II2514))|((~II2522));
assign WX7289 = (WX7226&RESET);
assign WX9611 = ((~WX10040));
assign II6382 = ((~WX2154))|((~II6380));
assign WX9219 = (WX9217)|(WX9216);
assign II6208 = ((~II6218))|((~II6219));
assign II22228 = ((~II22238))|((~II22239));
assign WX82 = (WX2326&WX83);
assign II18922 = ((~WX6003))|((~WX6067));
assign II2715 = ((~II2717))|((~II2718));
assign WX3356 = (WX3293&RESET);
assign WX4956 = (WX4955&WX4884);
assign II18196 = ((~WX5829))|((~II18194));
assign II19087 = ((~WX5659))|((~II19085));
assign II31711 = ((~WX9687))|((~II31710));
assign WX5266 = (WX5264)|(WX5263);
assign WX6550 = (WX6956&WX7469);
assign II26175 = ((~WX8413))|((~II26173));
assign WX1621 = ((~WX1620));
assign WX4123 = ((~WX4122));
assign WX4444 = ((~WX4814));
assign II35751 = ((~WX10986))|((~II35750));
assign II30076 = ((~II30052))|((~II30068));
assign II15106 = ((~WX4462))|((~WX4370));
assign II7512 = ((~_2112_))|((~II7504));
assign WX7583 = ((~II23286))|((~II23287));
assign WX7855 = ((~WX8762));
assign II34509 = ((~WX11147))|((~II34508));
assign II26266 = ((~WX8759))|((~WX8419));
assign WX1827 = (WX1830&RESET);
assign WX6448 = (WX6430&WX6435);
assign WX8005 = ((~WX8761));
assign II22352 = ((~II22362))|((~II22363));
assign II10740 = ((~II10750))|((~II10751));
assign WX6847 = (WX6845)|(WX6844);
assign WX6222 = (WX5758&WX6223);
assign WX5305 = (WX5316&WX6175);
assign II14862 = ((~II14838))|((~II14854));
assign WX2485 = (WX2483)|(WX2482);
assign WX10135 = (WX10134&WX10056);
assign II2885 = ((~II2895))|((~II2896));
assign II30745 = ((~II30735))|((~II30743));
assign II22929 = ((~WX7360))|((~II22927));
assign WX2679 = ((~WX3589));
assign WX10066 = (WX9632&WX10067);
assign WX8162 = (WX10245&WX8163);
assign WX10117 = (WX10115)|(WX10114);
assign II22617 = ((~WX7276))|((~WX7340));
assign WX11604 = ((~II35737))|((~II35738));
assign WX8179 = (WX8297&WX8762);
assign II14601 = ((~II14591))|((~II14599));
assign WX375 = (_2084_&WX1004);
assign WX10457 = (WX10839&WX11348);
assign WX10775 = (_2336_&WX11348);
assign WX6100 = ((~II18899))|((~II18900));
assign II2826 = ((~WX1002))|((~II2825));
assign WX4011 = ((~WX4010));
assign WX4450 = ((~WX4826));
assign WX10228 = ((~WX10056));
assign WX8430 = (WX8002&RESET);
assign WX10263 = ((~WX10056));
assign WX2344 = ((~WX2298));
assign II31179 = ((~WX9638))|((~II31178));
assign II6567 = ((~WX2102))|((~II6566));
assign II10790 = ((~WX3473))|((~II10788));
assign II22696 = ((~WX7467))|((~II22695));
assign WX5481 = (WX5695&WX6176);
assign II35653 = ((~WX10969))|((~II35652));
assign II19563 = ((~WX5787))|((~II19562));
assign II2639 = ((~WX1002))|((~WX687));
assign WX1694 = ((~WX2296));
assign WX5534 = (WX7638&WX5535);
assign WX4945 = (WX4943)|(WX4942);
assign WX6279 = ((~WX6177));
assign WX7104 = ((~WX7356));
assign WX11136 = (WX11073&RESET);
assign WX5456 = (WX5454)|(WX5453);
assign II11259 = ((~WX3101))|((~II11257));
assign II2872 = ((~WX829))|((~II2871));
assign WX6210 = (WX6208)|(WX6207);
assign II19513 = ((~_2215_))|((~II19512));
assign WX10099 = ((~II31166))|((~II31167));
assign WX2314 = (WX2313&WX2298);
assign WX2223 = ((~II6946))|((~II6947));
assign WX1969 = (WX1565&RESET);
assign WX8530 = (WX8467&RESET);
assign II27614 = ((~WX8379))|((~_2290_));
assign II22936 = ((~II22926))|((~II22934));
assign II34919 = ((~II34894))|((~II34918));
assign WX4160 = (WX4398&WX4883);
assign WX235 = (_2094_&WX1004);
assign WX10254 = (WX10253&WX10056);
assign WX5692 = (WX5695&RESET);
assign WX9785 = (WX9722&RESET);
assign II3093 = ((~WX491))|((~II3091));
assign II18342 = ((~II18332))|((~II18340));
assign WX130 = (WX128)|(WX127);
assign WX11270 = ((~II34857))|((~II34858));
assign WX360 = (WX358)|(WX357);
assign II10657 = ((~WX3337))|((~II10656));
assign WX10820 = (WX10818)|(WX10817);
assign II15418 = ((~WX4486))|((~WX4418));
assign WX10092 = ((~II31153))|((~II31154));
assign II6893 = ((~WX2295))|((~II6892));
assign WX9626 = ((~WX10006));
assign WX281 = (WX519&WX1004);
assign II22191 = ((~II22166))|((~II22190));
assign II35591 = ((~_2359_))|((~II35589));
assign II26420 = ((~II26422))|((~II26423));
assign WX2553 = ((~II7702))|((~II7703));
assign II23246 = ((~WX7058))|((~WX6976));
assign II15566 = ((~_2199_))|((~II15564));
assign II2462 = ((~II2452))|((~II2460));
assign WX3326 = (WX3263&RESET);
assign II10694 = ((~II10696))|((~II10697));
assign WX7404 = ((~WX7403));
assign II26436 = ((~WX8557))|((~WX8621));
assign II30541 = ((~II30517))|((~II30533));
assign WX11511 = ((~II35392))|((~II35393));
assign WX7017 = ((~WX7438));
assign WX4439 = ((~WX4868));
assign WX8696 = ((~WX8677));
assign II18876 = ((~WX6174))|((~WX5873));
assign WX9448 = ((~WX9439));
assign II26559 = ((~II26561))|((~II26562));
assign II22037 = ((~II22027))|((~II22035));
assign II18719 = ((~II18729))|((~II18730));
assign II10100 = ((~II10090))|((~II10098));
assign II6069 = ((~II6071))|((~II6072));
assign II7688 = ((~WX1930))|((~II7687));
assign II10974 = ((~WX3421))|((~WX3485));
assign II10967 = ((~WX3357))|((~II10966));
assign II18976 = ((~WX5943))|((~II18968));
assign WX6383 = (WX5781&WX6384);
assign WX1226 = ((~WX1005));
assign II26314 = ((~WX8613))|((~II26312));
assign II14291 = ((~II14281))|((~II14289));
assign WX8528 = (WX8465&RESET);
assign II10547 = ((~II10523))|((~II10539));
assign WX488 = (WX491&RESET);
assign WX2467 = ((~II7370))|((~II7371));
assign II19216 = ((~WX5763))|((~II19215));
assign WX421 = (WX539&WX1004);
assign II26583 = ((~WX8503))|((~II26575));
assign WX8916 = ((~WX8915));
assign WX8955 = (WX8365&WX8956);
assign II15236 = ((~WX4472))|((~WX4390));
assign II11715 = ((~_2142_))|((~II11713));
assign II31605 = ((~WX9670))|((~_2324_));
assign II30657 = ((~II30659))|((~II30660));
assign II22681 = ((~WX7344))|((~II22679));
assign II15250 = ((~WX4473))|((~II15249));
assign WX1745 = (WX1743)|(WX1742);
assign II6970 = ((~WX2128))|((~II6969));
assign WX6867 = (WX6865)|(WX6864);
assign II19676 = ((~_2214_))|((~II19674));
assign WX9857 = (WX9794&RESET);
assign II2367 = ((~WX733))|((~II2359));
assign WX946 = ((~WX923));
assign WX2399 = (WX1887&WX2400);
assign II22058 = ((~II22060))|((~II22061));
assign WX6566 = ((~WX7469));
assign II7279 = ((~WX1890))|((~II7278));
assign WX11309 = ((~WX11308));
assign WX1025 = ((~WX1024));
assign WX6888 = ((~WX7469));
assign II34205 = ((~II34181))|((~II34197));
assign WX5617 = (_2207_&WX6176);
assign WX4054 = (WX4065&WX4882);
assign II18458 = ((~WX5973))|((~II18457));
assign WX754 = (WX691&RESET);
assign WX353 = ((~WX1004));
assign II10007 = ((~II9997))|((~II10005));
assign WX11350 = ((~II35093))|((~II35094));
assign WX7311 = (WX7248&RESET);
assign WX1628 = ((~WX2297));
assign WX8854 = ((~WX8853));
assign WX306 = (WX2438&WX307);
assign WX318 = (WX316)|(WX315);
assign DATA_9_27 = ((~WX1039));
assign WX3649 = (WX3648&WX3591);
assign WX2651 = ((~WX3589));
assign II14437 = ((~WX4880))|((~WX4552));
assign WX10296 = ((~II31627))|((~II31628));
assign WX6184 = ((~WX6183));
assign II22121 = ((~WX7244))|((~WX7308));
assign II22340 = ((~WX7322))|((~II22338));
assign WX8743 = ((~WX8742));
assign II34464 = ((~WX11017))|((~II34462));
assign WX4571 = (WX4263&RESET);
assign II22973 = ((~II22975))|((~II22976));
assign II26729 = ((~II26739))|((~II26740));
assign WX2781 = ((~WX3590));
assign II30534 = ((~WX9856))|((~WX9920));
assign II6032 = ((~WX2004))|((~II6031));
assign WX8871 = (WX8353&WX8872);
assign WX3633 = ((~WX3632));
assign WX11479 = ((~WX11349));
assign II30851 = ((~II30827))|((~II30843));
assign WX10412 = (DATA_0_29&WX10413);
assign WX11425 = ((~WX11424));
assign II35667 = ((~WX10972))|((~II35666));
assign WX3138 = ((~WX3559));
assign WX9463 = ((~WX9462));
assign II6119 = ((~WX1946))|((~II6117));
assign WX4096 = (WX4107&WX4882);
assign II18007 = ((~II18009))|((~II18010));
assign WX9192 = (WX9550&WX10055);
assign WX3400 = (WX3337&RESET);
assign WX784 = (WX721&RESET);
assign WX5249 = (WX5260&WX6175);
assign II34626 = ((~II34616))|((~II34624));
assign WX5120 = ((~II15579))|((~II15580));
assign II27199 = ((~WX8347))|((~WX8261));
assign II18712 = ((~II18688))|((~II18704));
assign II31683 = ((~WX9682))|((~II31682));
assign WX5606 = (WX5604)|(WX5603);
assign WX2385 = (WX1885&WX2386);
assign WX1288 = (WX1253&WX1263);
assign WX3380 = (WX3317&RESET);
assign II14005 = ((~WX4524))|((~II14003));
assign II26621 = ((~II26623))|((~II26624));
assign II14438 = ((~WX4880))|((~II14437));
assign WX7507 = (WX7506&WX7470);
assign WX3671 = (WX3177&WX3672);
assign WX286 = ((~WX285));
assign II11673 = ((~_2149_))|((~II11671));
assign WX4346 = ((~WX4337));
assign WX2898 = (WX2896)|(WX2895);
assign II27264 = ((~WX8352))|((~WX8271));
assign WX9811 = (WX9748&RESET);
assign WX4555 = (WX4151&RESET);
assign II2513 = ((~II2523))|((~II2524));
assign WX1653 = (WX1651)|(WX1650);
assign WX9715 = (WX9239&RESET);
assign II27342 = ((~WX8358))|((~WX8283));
assign II2482 = ((~II2492))|((~II2493));
assign II11257 = ((~WX3181))|((~WX3101));
assign WX11106 = (WX11043&RESET);
assign WX1272 = (WX1233&WX1263);
assign WX7203 = (WX7140&RESET);
assign II2529 = ((~II2531))|((~II2532));
assign WX8727 = ((~WX8726));
assign II3351 = ((~WX603))|((~WX531));
assign WX2615 = (WX2530&WX2556);
assign WX8440 = (WX8072&RESET);
assign WX8640 = (WX8577&RESET);
assign II34316 = ((~II34306))|((~II34314));
assign WX4518 = ((~WX4770));
assign WX10538 = (DATA_0_20&WX10539);
assign II30675 = ((~WX10053))|((~II30674));
assign II18753 = ((~WX6174))|((~II18752));
assign WX3100 = (WX3103&RESET);
assign WX6580 = ((~WX7469));
assign II34083 = ((~II34073))|((~II34081));
assign II7584 = ((~_2131_))|((~II7582));
assign WX11269 = ((~II34826))|((~II34827));
assign WX7901 = ((~WX8762));
assign WX6525 = (WX6523)|(WX6522);
assign II26351 = ((~II26326))|((~II26350));
assign WX9471 = (WX9469)|(WX9468);
assign II14167 = ((~II14157))|((~II14165));
assign II31718 = ((~WX9688))|((~II31717));
assign II31584 = ((~WX9667))|((~_2327_));
assign WX359 = ((~WX1003));
assign WX6638 = ((~WX6629));
assign II34664 = ((~WX11157))|((~II34663));
assign WX2434 = (WX1892&WX2435);
assign II10077 = ((~WX3427))|((~II10075));
assign WX6879 = (WX6885&WX6880);
assign WX6913 = (WX6911)|(WX6910);
assign II26096 = ((~WX8535))|((~II26095));
assign WX4679 = (WX4616&RESET);
assign II7331 = ((~WX1894))|((~II7330));
assign WX11521 = ((~WX11349));
assign II2204 = ((~II2206))|((~II2207));
assign WX3284 = (WX3012&RESET);
assign II18645 = ((~WX6049))|((~II18643));
assign WX11407 = (WX11406&WX11349);
assign WX8812 = ((~WX8811));
assign WX4413 = (WX4416&RESET);
assign WX9299 = (WX9297)|(WX9296);
assign II26342 = ((~II26344))|((~II26345));
assign WX273 = (WX284&WX1003);
assign WX6377 = ((~WX6177));
assign WX5250 = (WX5256&WX5251);
assign WX9176 = ((~WX10055));
assign II23117 = ((~WX7048))|((~II23116));
assign II10735 = ((~II10725))|((~II10733));
assign WX9198 = (WX9209&WX10054);
assign WX9228 = ((~WX10054));
assign WX3454 = (WX3391&RESET);
assign II6265 = ((~II6255))|((~II6263));
assign II23377 = ((~WX7068))|((~II23376));
assign II14383 = ((~WX4612))|((~II14382));
assign WX11429 = (WX10935&WX11430);
assign WX1515 = (WX3689&WX1516);
assign WX8709 = ((~WX8708));
assign WX1182 = (WX1181&WX1005);
assign WX10218 = ((~II31387))|((~II31388));
assign WX3006 = (WX3004)|(WX3003);
assign II14873 = ((~WX4580))|((~II14871));
assign WX1041 = ((~II3118))|((~II3119));
assign II18048 = ((~II18038))|((~II18046));
assign WX9291 = (WX10161&WX9292);
assign II10322 = ((~II10324))|((~II10325));
assign WX3808 = ((~WX3807));
assign WX4485 = ((~WX4453));
assign WX50 = (WX56&WX51);
assign II34362 = ((~II34352))|((~II34360));
assign WX4459 = ((~WX4427));
assign II2382 = ((~II2358))|((~II2374));
assign WX10711 = ((~WX11348));
assign WX10659 = (WX10670&WX11347);
assign II2327 = ((~II2337))|((~II2338));
assign WX9345 = (WX9343)|(WX9342);
assign II26413 = ((~II26388))|((~II26412));
assign WX1895 = ((~WX1863));
assign II19584 = ((~WX5790))|((~II19583));
assign WX57 = (WX487&WX1004);
assign WX8671 = ((~II26444))|((~II26445));
assign II2103 = ((~II2079))|((~II2095));
assign WX4210 = ((~WX4882));
assign WX9474 = ((~WX10055));
assign II23611 = ((~_2258_))|((~II23609));
assign II35589 = ((~WX10960))|((~_2359_));
assign II34290 = ((~II34292))|((~II34293));
assign WX9993 = ((~WX9972));
assign II18520 = ((~WX5977))|((~II18519));
assign WX2533 = ((~II7562))|((~II7563));
assign WX8326 = ((~WX8699));
assign WX11499 = (WX10945&WX11500);
assign WX11644 = (WX11592&WX11607);
assign WX2983 = ((~WX2974));
assign II27500 = ((~WX8385))|((~_2300_));
assign WX9010 = ((~II27671))|((~II27672));
assign WX858 = (WX795&RESET);
assign WX10564 = (WX10562)|(WX10561);
assign WX5793 = ((~WX6027));
assign II14553 = ((~II14528))|((~II14552));
assign II7423 = ((~WX1834))|((~II7421));
assign WX8502 = (WX8439&RESET);
assign WX4471 = ((~WX4439));
assign II2113 = ((~WX1001))|((~II2112));
assign II27507 = ((~_2284_))|((~II27499));
assign WX7494 = (WX7048&WX7495);
assign II34159 = ((~WX11061))|((~II34151));
assign WX7077 = ((~WX7302));
assign WX340 = (WX338)|(WX337);
assign II18815 = ((~WX6174))|((~II18814));
assign WX2954 = (WX2952)|(WX2951);
assign WX9044 = (WX8990&WX9021);
assign WX6144 = ((~WX6076));
assign II6008 = ((~WX2066))|((~WX2130));
assign WX3462 = (WX3399&RESET);
assign II15225 = ((~WX4388))|((~II15223));
assign II10355 = ((~WX3381))|((~II10354));
assign WX8394 = ((~WX8643));
assign II35418 = ((~WX10949))|((~II35417));
assign WX5918 = (WX5855&RESET);
assign WX2157 = (WX2094&RESET);
assign II27522 = ((~_2279_))|((~II27514));
assign WX10493 = ((~WX11347));
assign II35640 = ((~_2352_))|((~II35638));
assign WX962 = ((~WX931));
assign WX8111 = ((~WX8762));
assign II2699 = ((~II2709))|((~II2710));
assign II2669 = ((~II2671))|((~II2672));
assign WX2500 = ((~WX2499));
assign II35197 = ((~WX10932))|((~II35196));
assign WX4131 = (WX4129)|(WX4128);
assign II22960 = ((~WX7362))|((~II22958));
assign II27637 = ((~_2287_))|((~II27635));
assign WX8847 = ((~WX8846));
assign II14964 = ((~WX4881))|((~WX4586));
assign WX6117 = ((~WX6116));
assign WX1056 = (WX1055&WX1005);
assign II30511 = ((~II30486))|((~II30510));
assign II6792 = ((~II6782))|((~II6790));
assign WX6537 = (WX7491&WX6538);
assign WX3043 = ((~WX3589));
assign WX7376 = ((~II22377))|((~II22378));
assign WX3224 = ((~WX3475));
assign WX3935 = (WX3933)|(WX3932);
assign WX983 = ((~WX982));
assign WX1574 = (WX1812&WX2297);
assign II6574 = ((~II6549))|((~II6573));
assign II2072 = ((~II2048))|((~II2064));
assign WX10709 = (WX10875&WX11348);
assign WX6559 = (WX6557)|(WX6556);
assign WX8077 = (_2280_&WX8762);
assign WX2429 = (WX2427)|(WX2426);
assign WX65 = ((~WX1003));
assign II34299 = ((~II34274))|((~II34298));
assign WX192 = (WX190)|(WX189);
assign II34788 = ((~WX11165))|((~II34787));
assign II26778 = ((~WX8579))|((~II26777));
assign WX9671 = ((~WX9904));
assign WX5637 = ((~WX6176));
assign WX6438 = (WX6434&WX6435);
assign II26388 = ((~II26398))|((~II26399));
assign II2267 = ((~WX1001))|((~WX663));
assign WX3611 = ((~WX3610));
assign WX10724 = (WX11524&WX10725);
assign WX7459 = ((~WX7380));
assign II22042 = ((~II22052))|((~II22053));
assign WX5746 = ((~WX6125));
assign II6584 = ((~WX1976))|((~II6582));
assign II26032 = ((~II26034))|((~II26035));
assign II18077 = ((~WX5885))|((~II18069));
assign WX5864 = (WX5556&RESET);
assign WX84 = (WX82)|(WX81);
assign WX1296 = (WX1231&WX1263);
assign II18162 = ((~II18164))|((~II18165));
assign WX7052 = ((~WX7020));
assign WX2270 = ((~WX2269));
assign II31648 = ((~WX9676))|((~II31647));
assign WX200 = (WX198)|(WX197);
assign WX3020 = (WX3018)|(WX3017);
assign WX4753 = (WX4690&RESET);
assign WX7107 = ((~WX7362));
assign WX10725 = ((~WX11348));
assign II15608 = ((~_2193_))|((~II15606));
assign WX1953 = (WX1453&RESET);
assign WX3521 = ((~WX3520));
assign WX10439 = (_2360_&WX11348);
assign II6427 = ((~WX2294))|((~WX1966));
assign WX8031 = (WX8042&WX8761);
assign WX6411 = ((~II19570))|((~II19571));
assign WX2087 = (WX2024&RESET);
assign II18940 = ((~WX5877))|((~II18938));
assign WX2282 = ((~WX2281));
assign WX8650 = (WX8587&RESET);
assign WX2970 = ((~WX2969));
assign WX1451 = (WX1449)|(WX1448);
assign II11502 = ((~_2151_))|((~II11494));
assign WX746 = (WX683&RESET);
assign II31191 = ((~WX9639))|((~WX9552));
assign WX7355 = (WX7292&RESET);
assign WX6714 = (_2253_&WX7469);
assign II22400 = ((~WX7262))|((~WX7326));
assign II3249 = ((~WX515))|((~II3247));
assign II10121 = ((~II10123))|((~II10124));
assign II34593 = ((~WX11089))|((~II34585));
assign WX2279 = ((~WX2204));
assign WX3640 = ((~WX3639));
assign WX5094 = ((~WX5093));
assign II23646 = ((~_2253_))|((~II23644));
assign II3403 = ((~WX607))|((~WX539));
assign WX6610 = ((~WX6601));
assign WX459 = (_2078_&WX1004);
assign II35638 = ((~WX10967))|((~_2352_));
assign II6868 = ((~WX2058))|((~II6860));
assign WX1614 = ((~WX2297));
assign WX6947 = ((~WX6946));
assign WX8052 = (WX8050)|(WX8049);
assign WX9310 = (WX9321&WX10054);
assign WX2083 = (WX2020&RESET);
assign II22438 = ((~II22414))|((~II22430));
assign WX5373 = ((~WX5364));
assign II30698 = ((~II30688))|((~II30696));
assign II30193 = ((~WX9834))|((~WX9898));
assign II10285 = ((~WX3313))|((~II10284));
assign WX1164 = (WX1162)|(WX1161);
assign WX10503 = ((~WX10494));
assign WX8733 = ((~WX8732));
assign II26327 = ((~II26329))|((~II26330));
assign WX3199 = ((~WX3425));
assign II14143 = ((~WX4660))|((~II14142));
assign II30232 = ((~II30207))|((~II30231));
assign II10309 = ((~WX3587))|((~II10308));
assign II10099 = ((~WX3301))|((~II10098));
assign WX7845 = ((~WX8762));
assign II7626 = ((~_2125_))|((~II7624));
assign WX3663 = (WX3662&WX3591);
assign II18426 = ((~WX5971))|((~WX6035));
assign II23624 = ((~WX7088))|((~II23623));
assign II26981 = ((~WX8465))|((~II26979));
assign WX1444 = (_2132_&WX2297);
assign WX9371 = (WX11496&WX9372);
assign II30309 = ((~WX9778))|((~II30301));
assign II7476 = ((~WX1920))|((~II7475));
assign WX9631 = ((~WX9599));
assign WX479 = ((~WX1004));
assign II26840 = ((~WX8583))|((~II26839));
assign WX1119 = (WX1118&WX1005);
assign II31243 = ((~WX9643))|((~WX9560));
assign II15433 = ((~WX4420))|((~II15431));
assign WX9236 = ((~WX10055));
assign WX1815 = (WX1818&RESET);
assign II10866 = ((~WX3588))|((~WX3287));
assign WX7478 = ((~II23091))|((~II23092));
assign WX1482 = (WX1493&WX2296);
assign II3312 = ((~WX600))|((~WX525));
assign II26972 = ((~II26962))|((~II26970));
assign WX259 = (WX270&WX1003);
assign II11657 = ((~WX3217))|((~_2152_));
assign WX10397 = (_2363_&WX11348);
assign WX10955 = ((~WX10923));
assign II35328 = ((~WX10865))|((~II35326));
assign II14305 = ((~II14280))|((~II14304));
assign WX3252 = (WX2788&RESET);
assign WX1594 = (WX1605&WX2296);
assign WX5426 = (WX6289&WX5427);
assign WX207 = (_2096_&WX1004);
assign II7483 = ((~_2124_))|((~II7482));
assign WX6687 = (WX8861&WX6688);
assign WX6678 = ((~WX7469));
assign II6062 = ((~WX2006))|((~II6054));
assign II34927 = ((~WX11346))|((~WX11047));
assign WX4531 = (WX3983&RESET);
assign WX4085 = (WX4083)|(WX4082);
assign WX8205 = ((~WX8762));
assign WX4635 = (WX4572&RESET);
assign II14539 = ((~II14529))|((~II14537));
assign WX2272 = ((~WX2271));
assign WX250 = (WX2410&WX251);
assign WX2946 = (WX2944)|(WX2943);
assign WX10158 = ((~WX10056));
assign WX5376 = (WX5382&WX5377);
assign WX10807 = (WX10889&WX11348);
assign WX3162 = ((~WX3543));
assign WX6407 = ((~II19542))|((~II19543));
assign WX10705 = (_2341_&WX11348);
assign II7215 = ((~WX1802))|((~II7213));
assign II2389 = ((~II2399))|((~II2400));
assign WX8400 = ((~WX8655));
assign II18992 = ((~II18967))|((~II18991));
assign WX2664 = (WX2670&WX2665);
assign II30510 = ((~II30486))|((~II30502));
assign II2832 = ((~WX763))|((~II2824));
assign WX2672 = (WX3619&WX2673);
assign WX6206 = ((~II19125))|((~II19126));
assign WX11301 = ((~WX11300));
assign WX4203 = (WX5031&WX4204);
assign II6753 = ((~WX2114))|((~II6752));
assign II6041 = ((~WX2132))|((~II6039));
assign II19425 = ((~WX5711))|((~II19423));
assign WX139 = ((~WX1004));
assign WX4844 = ((~WX4843));
assign WX6874 = ((~WX7469));
assign II18326 = ((~WX5901))|((~II18325));
assign WX2235 = ((~WX2214));
assign WX5231 = ((~WX6176));
assign WX2255 = ((~WX2224));
assign WX7436 = ((~WX7435));
assign II15446 = ((~WX4422))|((~II15444));
assign WX5234 = ((~WX5233));
assign II7408 = ((~WX1900))|((~WX1832));
assign WX6895 = (WX6893)|(WX6892);
assign WX7914 = (WX8826&WX7915);
assign WX9569 = (WX9572&RESET);
assign WX10600 = (WX10598)|(WX10597);
assign II22480 = ((~WX7140))|((~II22478));
assign II23443 = ((~WX7006))|((~II23441));
assign II15712 = ((~WX4519))|((~II15711));
assign II3662 = ((~WX634))|((~II3661));
assign WX5145 = (WX5141&WX5142);
assign WX1532 = (WX1806&WX2297);
assign II15158 = ((~WX4466))|((~WX4378));
assign WX1587 = (WX1585)|(WX1584);
assign II2896 = ((~II2886))|((~II2894));
assign WX2658 = (WX3612&WX2659);
assign II34895 = ((~II34897))|((~II34898));
assign WX4285 = (WX4283)|(WX4282);
assign WX7676 = (WX7074&WX7677);
assign II30300 = ((~II30310))|((~II30311));
assign II10906 = ((~II10896))|((~II10904));
assign II2786 = ((~II2761))|((~II2785));
assign WX2931 = ((~WX3589));
assign WX10541 = (WX10851&WX11348);
assign WX4721 = (WX4658&RESET);
assign II23509 = ((~II23511))|((~II23512));
assign II34571 = ((~WX11151))|((~II34570));
assign II34562 = ((~WX11087))|((~II34554));
assign WX6121 = ((~WX6120));
assign WX5326 = (WX5324)|(WX5323);
assign II22666 = ((~WX7152))|((~II22664));
assign WX2461 = (WX2460&WX2298);
assign WX264 = (WX2417&WX265);
assign WX6843 = (WX6841)|(WX6840);
assign WX1668 = (_2116_&WX2297);
assign WX7462 = ((~TM0));
assign WX660 = (WX160&RESET);
assign WX7046 = ((~WX7014));
assign WX1326 = (WX1235&WX1263);
assign WX2681 = (_2168_&WX3590);
assign WX7654 = (WX7653&WX7470);
assign II26808 = ((~WX8581))|((~WX8645));
assign WX11226 = (WX11163&RESET);
assign WX3148 = ((~WX3579));
assign WX9632 = ((~WX9600));
assign II14468 = ((~WX4880))|((~WX4554));
assign II14043 = ((~II14033))|((~II14041));
assign WX3860 = (WX3845&WX3849);
assign WX2876 = (WX2874)|(WX2873);
assign II19334 = ((~WX5697))|((~II19332));
assign II2470 = ((~WX867))|((~II2468));
assign WX10619 = ((~WX11347));
assign WX11252 = ((~II34299))|((~II34300));
assign WX7615 = (WX7613)|(WX7612);
assign WX6266 = (WX6264)|(WX6263);
assign WX1876 = ((~WX1844));
assign WX3029 = ((~WX3589));
assign WX8095 = (WX8285&WX8762);
assign WX6892 = (WX6903&WX7468);
assign WX3128 = (WX3131&RESET);
assign WX100 = (DATA_9_27&WX101);
assign II6201 = ((~II6177))|((~II6193));
assign WX637 = ((~WX887));
assign WX470 = (WX476&WX471);
assign II18598 = ((~WX6174))|((~II18597));
assign WX11464 = (WX10940&WX11465);
assign WX7699 = ((~II23540))|((~II23541));
assign II11089 = ((~WX3168))|((~II11088));
assign WX4191 = (WX4189)|(WX4188);
assign WX9164 = (WX9546&WX10055);
assign WX8945 = ((~WX8944));
assign II27134 = ((~WX8342))|((~WX8251));
assign WX10234 = (WX9656&WX10235);
assign II22308 = ((~WX7256))|((~II22307));
assign WX6282 = ((~WX6281));
assign WX7450 = ((~WX7449));
assign WX7609 = ((~WX7608));
assign WX4316 = ((~WX4883));
assign WX10302 = ((~II31669))|((~II31670));
assign II19450 = ((~WX5781))|((~II19449));
assign WX8176 = (WX10252&WX8177);
assign WX4344 = ((~WX4883));
assign II18404 = ((~II18394))|((~II18402));
assign II22587 = ((~WX7274))|((~II22586));
assign WX8215 = ((~WX8761));
assign WX4609 = (WX4546&RESET);
assign II11720 = ((~WX3228))|((~_2141_));
assign WX6772 = ((~WX7469));
assign WX10032 = ((~WX10031));
assign WX6621 = (WX7533&WX6622);
assign WX2211 = ((~II6574))|((~II6575));
assign WX7998 = (WX8868&WX7999);
assign WX10167 = ((~WX10166));
assign II2692 = ((~II2668))|((~II2684));
assign WX4846 = ((~WX4845));
assign WX5570 = ((~WX5569));
assign WX109 = (_2103_&WX1004);
assign WX2363 = (WX2362&WX2298);
assign WX2115 = (WX2052&RESET);
assign WX9972 = ((~II30697))|((~II30698));
assign WX3826 = ((~II11567))|((~II11568));
assign II18487 = ((~II18489))|((~II18490));
assign WX5592 = (WX5590)|(WX5589);
assign II27329 = ((~WX8357))|((~WX8281));
assign II7661 = ((~_2118_))|((~II7659));
assign WX9660 = ((~WX9628));
assign II27544 = ((~WX8401))|((~_2300_));
assign II18892 = ((~WX6001))|((~II18891));
assign WX10365 = (WX10292&WX10314);
assign WX9390 = ((~WX10055));
assign II15636 = ((~_2189_))|((~II15634));
assign WX1477 = (WX2375&WX1478);
assign WX2747 = (WX2758&WX3589);
assign WX6997 = (WX7000&RESET);
assign WX8864 = (WX8352&WX8865);
assign II14320 = ((~WX4608))|((~II14312));
assign WX6464 = (WX6423&WX6435);
assign II6683 = ((~WX2046))|((~II6682));
assign WX9893 = (WX9830&RESET);
assign WX988 = ((~WX912));
assign II2601 = ((~II2591))|((~II2599));
assign WX4362 = ((~WX4364));
assign WX642 = ((~WX897));
assign WX2856 = (WX2854)|(WX2853);
assign WX3701 = (WX3699)|(WX3698);
assign II34422 = ((~II34398))|((~II34414));
assign WX9182 = ((~WX9173));
assign WX9507 = (WX9513&WX9508);
assign WX8152 = (WX8945&WX8153);
assign WX9022 = (WX8992&WX9021);
assign WX10039 = ((~WX9963));
assign WX5073 = ((~WX5072));
assign WX7967 = ((~WX8762));
assign II27545 = ((~WX8401))|((~II27544));
assign WX5008 = (WX5006)|(WX5005);
assign WX7431 = ((~WX7366));
assign WX5211 = (_2236_&WX6176);
assign WX2804 = (WX2810&WX2805);
assign WX4921 = (WX4920&WX4884);
assign II22301 = ((~II22291))|((~II22299));
assign II34285 = ((~II34275))|((~II34283));
assign WX75 = ((~WX66));
assign WX4331 = (WX4329)|(WX4328);
assign WX6303 = ((~WX6302));
assign II2314 = ((~WX793))|((~II2313));
assign WX260 = (WX266&WX261);
assign WX2759 = ((~WX2750));
assign II35366 = ((~WX10945))|((~II35365));
assign II18800 = ((~WX6059))|((~II18798));
assign WX115 = ((~WX1004));
assign II7519 = ((~WX1936))|((~_2140_));
assign WX10081 = ((~WX10056));
assign WX9987 = ((~WX9969));
assign WX8067 = (WX8281&WX8762);
assign WX1414 = ((~WX2296));
assign DATA_9_1 = ((~WX1221));
assign WX10054 = ((~WX10050));
assign WX1255 = ((~II3662))|((~II3663));
assign II34709 = ((~II34711))|((~II34712));
assign WX292 = (WX2431&WX293);
assign WX6648 = (WX6970&WX7469);
assign WX2992 = (WX2990)|(WX2989);
assign II35406 = ((~WX10877))|((~II35404));
assign WX11020 = (WX10616&RESET);
assign WX6933 = ((~WX6932));
assign WX3968 = ((~WX3959));
assign II2662 = ((~II2637))|((~II2661));
assign II14513 = ((~II14515))|((~II14516));
assign WX7866 = (WX7864)|(WX7863);
assign WX1147 = (WX1146&WX1005);
assign II10524 = ((~II10526))|((~II10527));
assign WX3292 = (WX3068&RESET);
assign II35555 = ((~WX10987))|((~II35554));
assign WX3396 = (WX3333&RESET);
assign WX1500 = (_2128_&WX2297);
assign WX7562 = ((~II23247))|((~II23248));
assign WX969 = ((~WX968));
assign WX9255 = (WX9261&WX9256);
assign II30597 = ((~WX9860))|((~II30596));
assign WX2105 = (WX2042&RESET);
assign WX1130 = ((~WX1129));
assign WX6110 = ((~WX6091));
assign WX9980 = ((~II30945))|((~II30946));
assign II27686 = ((~_2278_))|((~II27684));
assign WX4871 = ((~WX4793));
assign WX2409 = ((~WX2408));
assign WX1312 = (WX1242&WX1263);
assign WX4711 = (WX4648&RESET);
assign WX7695 = ((~RESET));
assign WX6963 = (WX6966&RESET);
assign WX8831 = (WX8829)|(WX8828);
assign WX2017 = (WX1954&RESET);
assign WX3733 = (WX3732&WX3591);
assign II26047 = ((~II26057))|((~II26058));
assign WX6574 = (_2263_&WX7469);
assign WX1881 = ((~WX1849));
assign II26026 = ((~WX8467))|((~II26025));
assign WX387 = ((~WX1003));
assign II18736 = ((~WX5991))|((~WX6055));
assign WX4369 = (WX4372&RESET);
assign II14389 = ((~II14391))|((~II14392));
assign WX6014 = (WX5951&RESET);
assign WX3618 = ((~WX3617));
assign WX10090 = ((~WX10089));
assign II30712 = ((~WX9804))|((~II30704));
assign WX8159 = ((~WX8761));
assign II23700 = ((~WX7101))|((~_2243_));
assign II6705 = ((~II6707))|((~II6708));
assign WX1705 = ((~WX1704));
assign WX432 = (WX2501&WX433);
assign II18495 = ((~II18471))|((~II18487));
assign WX7397 = ((~WX7381));
assign WX5053 = ((~II15380))|((~II15381));
assign II22982 = ((~WX7236))|((~II22981));
assign II34052 = ((~II34042))|((~II34050));
assign WX9689 = ((~WX9940));
assign WX4138 = (WX4149&WX4882);
assign II30388 = ((~II30378))|((~II30386));
assign II2592 = ((~WX811))|((~WX875));
assign WX3562 = ((~WX3492));
assign WX5723 = ((~WX6143));
assign II15159 = ((~WX4466))|((~II15158));
assign II2871 = ((~WX829))|((~WX893));
assign WX6293 = ((~WX6177));
assign WX1763 = (WX1769&WX1764);
assign II23104 = ((~WX7047))|((~II23103));
assign WX10390 = (WX10388)|(WX10387);
assign II18070 = ((~WX6173))|((~WX5821));
assign WX10405 = ((~WX10396));
assign WX3963 = (WX3961)|(WX3960);
assign II18596 = ((~II18598))|((~II18599));
assign II10573 = ((~WX3459))|((~II10571));
assign WX9305 = (WX10168&WX9306);
assign WX2628 = (WX2626)|(WX2625);
assign II23679 = ((~WX7098))|((~_2246_));
assign II30356 = ((~II30331))|((~II30355));
assign WX8228 = (WX8234&WX8229);
assign WX5328 = (WX6240&WX5329);
assign II34213 = ((~II34215))|((~II34216));
assign II10981 = ((~II10957))|((~II10973));
assign WX9212 = (WX9223&WX10054);
assign II6885 = ((~II6875))|((~II6883));
assign II2358 = ((~II2368))|((~II2369));
assign WX5296 = (WX7519&WX5297);
assign II6146 = ((~II6156))|((~II6157));
assign II30620 = ((~WX9798))|((~II30619));
assign II30970 = ((~WX9948))|((~II30968));
assign II30456 = ((~II30458))|((~II30459));
assign WX8059 = (WX8070&WX8761);
assign WX7716 = ((~II23659))|((~II23660));
assign II2608 = ((~WX1002))|((~WX685));
assign II23610 = ((~WX7086))|((~II23609));
assign WX11387 = (WX10929&WX11388);
assign WX5518 = (WX5516)|(WX5515);
assign WX11084 = (WX11021&RESET);
assign II14842 = ((~WX4578))|((~II14840));
assign WX3278 = (WX2970&RESET);
assign II26995 = ((~WX8593))|((~II26994));
assign WX1011 = ((~WX1010));
assign WX7072 = ((~WX7040));
assign II26166 = ((~II26156))|((~II26164));
assign II2594 = ((~WX875))|((~II2592));
assign WX9953 = ((~II30108))|((~II30109));
assign II35509 = ((~II35511))|((~II35512));
assign II30347 = ((~II30349))|((~II30350));
assign II18550 = ((~WX5979))|((~WX6043));
assign II6196 = ((~WX2142))|((~II6194));
assign WX808 = (WX745&RESET);
assign WX9488 = ((~WX10055));
assign WX5004 = ((~II15289))|((~II15290));
assign WX9454 = (_2306_&WX10055);
assign WX443 = ((~WX1003));
assign WX6953 = (WX6956&RESET);
assign II34958 = ((~WX11346))|((~WX11049));
assign WX5088 = ((~II15445))|((~II15446));
assign II15690 = ((~WX4515))|((~_2179_));
assign WX7480 = (WX7046&WX7481);
assign WX1825 = (WX1828&RESET);
assign II14981 = ((~WX4778))|((~II14979));
assign WX10461 = ((~WX10452));
assign WX4342 = (WX4424&WX4883);
assign II10508 = ((~II10510))|((~II10511));
assign WX8284 = (WX8287&RESET);
assign WX1331 = (WX1329)|(WX1328);
assign II31514 = ((~II31504))|((~II31512));
assign WX2692 = (WX2698&WX2693);
assign II22114 = ((~WX7180))|((~II22113));
assign II18412 = ((~WX6173))|((~II18411));
assign WX11228 = (WX11165&RESET);
assign II30068 = ((~II30070))|((~II30071));
assign II2761 = ((~II2771))|((~II2772));
assign WX8240 = ((~WX8239));
assign WX5012 = (WX5011&WX4884);
assign WX944 = ((~WX922));
assign WX2362 = ((~II7175))|((~II7176));
assign WX11224 = (WX11161&RESET);
assign II18552 = ((~WX6043))|((~II18550));
assign WX3824 = ((~II11553))|((~II11554));
assign WX7487 = (WX7047&WX7488);
assign WX11255 = ((~II34392))|((~II34393));
assign II30226 = ((~WX9900))|((~II30224));
assign WX8903 = ((~WX8902));
assign II6226 = ((~WX2080))|((~II6225));
assign II27588 = ((~_2294_))|((~II27586));
assign II11664 = ((~WX3219))|((~_2150_));
assign WX1801 = (WX1804&RESET);
assign WX11544 = ((~WX11543));
assign WX2412 = (WX2411&WX2298);
assign II22076 = ((~WX7466))|((~II22075));
assign WX3176 = ((~WX3144));
assign II30378 = ((~II30380))|((~II30381));
assign WX3122 = (WX3125&RESET);
assign WX9690 = ((~WX9942));
assign WX11610 = (WX11606&WX11607);
assign WX9392 = ((~WX9383));
assign WX2686 = (WX3626&WX2687);
assign WX1947 = (WX1411&RESET);
assign WX125 = ((~WX1004));
assign II1987 = ((~II1989))|((~II1990));
assign WX5189 = (WX5122&WX5142);
assign WX639 = ((~WX891));
assign WX11550 = (WX11548)|(WX11547);
assign WX10761 = (_2337_&WX11348);
assign II23454 = ((~WX7074))|((~WX7008));
assign WX5472 = ((~WX5471));
assign II34500 = ((~WX11083))|((~II34492));
assign WX3745 = ((~WX3744));
assign WX7335 = (WX7272&RESET);
assign WX6423 = ((~II19654))|((~II19655));
assign WX5684 = (WX5687&RESET);
assign II2584 = ((~WX747))|((~II2576));
assign WX11343 = ((~TM1));
assign WX5820 = (WX5248&RESET);
assign II22851 = ((~WX7467))|((~II22850));
assign WX8823 = ((~WX8763));
assign WX6652 = ((~WX6643));
assign II6413 = ((~WX2156))|((~II6411));
assign WX9445 = (WX10238&WX9446);
assign II34819 = ((~WX11167))|((~II34818));
assign WX7425 = ((~WX7395));
assign II22135 = ((~II22145))|((~II22146));
assign WX7127 = (WX6639&RESET);
assign WX1245 = ((~II3592))|((~II3593));
assign WX2231 = ((~WX2212));
assign WX7630 = ((~WX7629));
assign WX240 = (DATA_9_17&WX241);
assign WX612 = ((~WX837));
assign II11439 = ((~WX3195))|((~WX3129));
assign WX3874 = (WX3839&WX3849);
assign WX6667 = ((~WX6666));
assign II14429 = ((~II14404))|((~II14428));
assign WX1399 = (WX1405&WX1400);
assign WX5319 = (WX5330&WX6175);
assign II26120 = ((~II26110))|((~II26118));
assign II14408 = ((~WX4550))|((~II14406));
assign II10028 = ((~II10030))|((~II10031));
assign II34097 = ((~WX11057))|((~II34089));
assign WX7879 = ((~WX8761));
assign II22802 = ((~II22804))|((~II22805));
assign II22526 = ((~WX7334))|((~II22524));
assign WX4966 = (WX4964)|(WX4963);
assign II22315 = ((~II22290))|((~II22314));
assign WX6914 = (WX7008&WX7469);
assign WX9369 = (WX9367)|(WX9366);
assign II30218 = ((~II30208))|((~II30216));
assign WX10765 = (WX10883&WX11348);
assign WX6649 = (WX7547&WX6650);
assign II26760 = ((~II26770))|((~II26771));
assign II10873 = ((~WX3351))|((~II10865));
assign WX2075 = (WX2012&RESET);
assign II10092 = ((~WX3587))|((~II10091));
assign II26669 = ((~WX8760))|((~WX8445));
assign WX830 = (WX767&RESET);
assign WX7171 = (WX6947&RESET);
assign II30030 = ((~WX9760))|((~II30022));
assign II10155 = ((~WX3241))|((~II10153));
assign WX1470 = ((~WX2296));
assign WX979 = ((~WX978));
assign WX1456 = ((~WX2296));
assign WX1369 = ((~WX1368));
assign WX3990 = ((~WX4883));
assign WX7495 = ((~WX7470));
assign WX8987 = ((~WX8986));
assign II18652 = ((~II18642))|((~II18650));
assign II10720 = ((~II10710))|((~II10718));
assign II22084 = ((~II22074))|((~II22082));
assign WX7874 = (WX7872)|(WX7871);
assign II6542 = ((~II6518))|((~II6534));
assign II10022 = ((~II10012))|((~II10020));
assign WX8392 = ((~WX8639));
assign WX8693 = ((~WX8692));
assign II18115 = ((~II18117))|((~II18118));
assign WX904 = ((~II2135))|((~II2136));
assign II34462 = ((~WX11345))|((~WX11017));
assign II2320 = ((~II2296))|((~II2312));
assign WX8976 = (WX8368&WX8977);
assign WX4284 = ((~WX4883));
assign WX4839 = ((~WX4809));
assign WX8302 = (WX8305&RESET);
assign WX3194 = ((~WX3162));
assign WX8804 = ((~WX8803));
assign WX11276 = ((~WX11260));
assign WX6060 = (WX5997&RESET);
assign WX2695 = (_2167_&WX3590);
assign II7605 = ((~_2128_))|((~II7603));
assign II34553 = ((~II34563))|((~II34564));
assign WX11334 = ((~WX11257));
assign WX2350 = (WX1880&WX2351);
assign II30806 = ((~WX9810))|((~II30805));
assign WX3658 = ((~WX3591));
assign WX6708 = ((~WX6699));
assign II31599 = ((~WX9669))|((~II31598));
assign WX3135 = ((~WX3553));
assign II2160 = ((~WX847))|((~II2158));
assign WX575 = ((~WX955));
assign II35120 = ((~WX10833))|((~II35118));
assign II26660 = ((~II26636))|((~II26652));
assign II15522 = ((~_2176_))|((~II15514));
assign WX6660 = ((~WX7469));
assign II23092 = ((~WX6952))|((~II23090));
assign WX6729 = (WX8882&WX6730);
assign II26019 = ((~WX8759))|((~II26018));
assign WX10194 = (WX10192)|(WX10191);
assign II18165 = ((~WX5827))|((~II18163));
assign WX3570 = ((~WX3496));
assign WX2905 = (_2152_&WX3590);
assign WX9121 = (WX9119)|(WX9118);
assign WX11398 = ((~WX11397));
assign II2966 = ((~WX899))|((~II2964));
assign WX4302 = ((~WX4883));
assign WX1364 = (WX1782&WX2297);
assign II30210 = ((~WX10052))|((~II30209));
assign WX2790 = (WX2796&WX2791);
assign II34121 = ((~WX11345))|((~WX10995));
assign II30589 = ((~WX9796))|((~II30588));
assign WX6397 = (WX5783&WX6398);
assign WX11313 = ((~WX11312));
assign WX4713 = (WX4650&RESET);
assign WX7686 = ((~WX7685));
assign WX3949 = (WX3947)|(WX3946);
assign WX6762 = ((~WX7469));
assign WX3512 = ((~II10827))|((~II10828));
assign II19256 = ((~WX5685))|((~II19254));
assign WX8063 = (_2281_&WX8762);
assign II2686 = ((~WX817))|((~II2685));
assign II2477 = ((~II2467))|((~II2475));
assign WX8883 = ((~II27304))|((~II27305));
assign WX8187 = ((~WX8761));
assign II35379 = ((~WX10946))|((~II35378));
assign WX6413 = ((~II19584))|((~II19585));
assign WX4792 = ((~II14429))|((~II14430));
assign II30046 = ((~II30021))|((~II30045));
assign WX5970 = (WX5907&RESET);
assign WX4806 = ((~II14863))|((~II14864));
assign WX2902 = (WX2908&WX2903);
assign II26221 = ((~WX8607))|((~II26219));
assign II34826 = ((~II34801))|((~II34825));
assign WX11564 = (WX11562)|(WX11561);
assign II10912 = ((~WX3417))|((~WX3481));
assign WX274 = (WX280&WX275);
assign WX4296 = (_2177_&WX4883);
assign II30751 = ((~WX9870))|((~WX9934));
assign WX8234 = (WX8232)|(WX8231);
assign WX6721 = (WX6719)|(WX6718);
assign WX7652 = ((~WX7651));
assign II18650 = ((~II18626))|((~II18642));
assign II15458 = ((~WX4489))|((~II15457));
assign WX3807 = ((~WX3806));
assign II34300 = ((~II34290))|((~II34298));
assign II7304 = ((~WX1892))|((~WX1816));
assign WX6615 = (WX6613)|(WX6612);
assign II30496 = ((~WX9790))|((~II30495));
assign II7317 = ((~WX1893))|((~WX1818));
assign II2710 = ((~II2700))|((~II2708));
assign II14616 = ((~II14606))|((~II14614));
assign WX1058 = ((~WX1005));
assign II34804 = ((~WX11346))|((~II34803));
assign II27530 = ((~WX8397))|((~_2300_));
assign II34742 = ((~WX11346))|((~II34741));
assign WX1700 = (WX1830&WX2297);
assign WX3438 = (WX3375&RESET);
assign II19683 = ((~_2213_))|((~II19681));
assign WX2302 = ((~WX2298));
assign WX3564 = ((~WX3493));
assign WX7062 = ((~WX7030));
assign WX2419 = (WX2418&WX2298);
assign WX4881 = ((~WX4877));
assign WX8558 = (WX8495&RESET);
assign WX6181 = ((~WX6177));
assign WX1333 = (WX3598&WX1334);
assign WX726 = (WX663&RESET);
assign WX732 = (WX669&RESET);
assign WX2581 = (WX2546&WX2556);
assign WX4992 = (WX4474&WX4993);
assign II30286 = ((~WX9840))|((~WX9904));
assign WX8363 = ((~WX8331));
assign WX7317 = (WX7254&RESET);
assign II26220 = ((~WX8543))|((~II26219));
assign WX9747 = (WX9463&RESET);
assign II31746 = ((~WX9693))|((~II31745));
assign WX650 = (WX90&RESET);
assign WX5288 = (WX5286)|(WX5285);
assign II18798 = ((~WX5995))|((~WX6059));
assign WX10822 = (WX11573&WX10823);
assign WX5406 = (WX5404)|(WX5403);
assign WX9103 = (WX9101)|(WX9100);
assign II23735 = ((~WX7107))|((~_2237_));
assign II14739 = ((~II14714))|((~II14738));
assign WX7888 = (WX7886)|(WX7885);
assign WX7731 = (WX7727&WX7728);
assign WX8767 = ((~WX8763));
assign II26251 = ((~WX8545))|((~II26250));
assign II3585 = ((~WX621))|((~II3584));
assign II26753 = ((~II26729))|((~II26745));
assign II10586 = ((~II10588))|((~II10589));
assign WX8898 = (WX8897&WX8763);
assign WX2577 = (WX2547&WX2556);
assign WX6807 = ((~WX6806));
assign WX3932 = (_2203_&WX4883);
assign II34507 = ((~II34509))|((~II34510));
assign II22742 = ((~WX7284))|((~II22741));
assign II23155 = ((~WX7051))|((~WX6962));
assign WX4975 = ((~WX4974));
assign WX10130 = ((~WX10056));
assign WX1384 = (WX1395&WX2296);
assign WX2889 = ((~WX3589));
assign WX7829 = (WX8247&WX8762);
assign WX8568 = (WX8505&RESET);
assign WX2458 = ((~WX2457));
assign II18420 = ((~II18410))|((~II18418));
assign WX9646 = ((~WX9614));
assign II3313 = ((~WX600))|((~II3312));
assign WX10419 = ((~WX10410));
assign WX2488 = ((~II7409))|((~II7410));
assign II19681 = ((~WX5806))|((~_2213_));
assign WX238 = (WX236)|(WX235);
assign WX389 = (_2083_&WX1004);
assign WX9682 = ((~WX9926));
assign WX5775 = ((~WX5743));
assign II19599 = ((~_2227_))|((~II19597));
assign II11179 = ((~WX3175))|((~WX3089));
assign WX10786 = (WX10792&WX10787);
assign WX8482 = (WX8419&RESET);
assign II30242 = ((~WX9710))|((~II30240));
assign II18838 = ((~II18828))|((~II18836));
assign II6642 = ((~II6652))|((~II6653));
assign WX8964 = (WX8962)|(WX8961);
assign II30348 = ((~WX9844))|((~WX9908));
assign II18559 = ((~II18549))|((~II18557));
assign WX3220 = ((~WX3467));
assign WX5461 = ((~WX6175));
assign II34440 = ((~II34430))|((~II34438));
assign WX5272 = (WX6212&WX5273);
assign WX2193 = ((~II6016))|((~II6017));
assign WX8105 = (_2278_&WX8762);
assign WX9052 = (WX9008&WX9021);
assign WX7668 = (WX7667&WX7470);
assign WX5067 = ((~II15406))|((~II15407));
assign WX2704 = ((~WX2703));
assign WX11507 = ((~WX11349));
assign WX6334 = (WX5774&WX6335);
assign WX2315 = (WX1875&WX2316);
assign II34974 = ((~WX11177))|((~II34973));
assign II30418 = ((~II30393))|((~II30417));
assign WX6056 = (WX5993&RESET);
assign WX3424 = (WX3361&RESET);
assign WX1308 = (WX1244&WX1263);
assign WX9941 = (WX9878&RESET);
assign WX912 = ((~II2383))|((~II2384));
assign WX7469 = ((~WX7462));
assign II2393 = ((~WX671))|((~II2391));
assign WX1791 = (WX1794&RESET);
assign WX10714 = ((~WX10713));
assign WX2357 = (WX1881&WX2358);
assign WX2826 = (WX3696&WX2827);
assign II2098 = ((~WX843))|((~II2096));
assign WX7626 = (WX7625&WX7470);
assign II11504 = ((~II11494))|((~II11502));
assign II6673 = ((~II6683))|((~II6684));
assign II2655 = ((~WX815))|((~II2654));
assign WX7347 = (WX7284&RESET);
assign II10074 = ((~II10076))|((~II10077));
assign WX7457 = ((~WX7379));
assign II11701 = ((~_2145_))|((~II11699));
assign WX1524 = (WX1535&WX2296);
assign WX11524 = ((~WX11523));
assign II26536 = ((~II26512))|((~II26528));
assign II15420 = ((~WX4418))|((~II15418));
assign II10146 = ((~II10136))|((~II10144));
assign II35011 = ((~II34987))|((~II35003));
assign II22795 = ((~WX7224))|((~II22787));
assign II7563 = ((~_2134_))|((~II7561));
assign WX3426 = (WX3363&RESET);
assign WX6247 = ((~WX6246));
assign II2780 = ((~WX887))|((~II2778));
assign WX405 = ((~WX1004));
assign WX568 = ((~WX941));
assign II23415 = ((~WX7071))|((~WX7002));
assign II6900 = ((~WX2060))|((~II6899));
assign WX684 = (WX328&RESET);
assign II10555 = ((~II10557))|((~II10558));
assign WX10589 = (WX10600&WX11347);
assign WX630 = ((~WX873));
assign II15173 = ((~WX4380))|((~II15171));
assign WX2556 = ((~WX2523));
assign II1997 = ((~II1987))|((~II1995));
assign WX4022 = ((~WX4883));
assign II10895 = ((~II10905))|((~II10906));
assign WX6312 = (WX6311&WX6177);
assign WX9042 = (WX9012&WX9021);
assign WX951 = ((~WX950));
assign WX964 = ((~WX900));
assign II15289 = ((~WX4476))|((~II15288));
assign WX10980 = ((~WX11229));
assign WX11403 = (WX11401)|(WX11400);
assign WX10201 = (WX10199)|(WX10198);
assign II10348 = ((~II10338))|((~II10346));
assign II34314 = ((~WX11071))|((~II34306));
assign WX7871 = (WX8253&WX8762);
assign WX9833 = (WX9770&RESET);
assign WX10643 = ((~WX10634));
assign WX7906 = (WX7912&WX7907);
assign WX4529 = (WX3969&RESET);
assign WX626 = ((~WX865));
assign WX37 = ((~WX1003));
assign WX7659 = ((~WX7658));
assign II2290 = ((~II2265))|((~II2289));
assign WX10514 = (WX11419&WX10515);
assign WX8939 = ((~II27408))|((~II27409));
assign WX5650 = (WX6401&WX5651);
assign II35703 = ((~_2341_))|((~II35701));
assign II18916 = ((~II18906))|((~II18914));
assign WX1731 = (WX1729)|(WX1728);
assign II31204 = ((~WX9640))|((~WX9554));
assign II6908 = ((~WX2124))|((~II6907));
assign WX917 = ((~II2538))|((~II2539));
assign WX2880 = (WX2878)|(WX2877);
assign WX6738 = (WX6749&WX7468);
assign II35517 = ((~_2348_))|((~II35509));
assign WX10010 = ((~WX10009));
assign II14459 = ((~II14435))|((~II14451));
assign WX9723 = (WX9295&RESET);
assign WX2728 = (WX3647&WX2729);
assign WX1839 = (WX1776&RESET);
assign WX1405 = (WX1403)|(WX1402);
assign II22323 = ((~WX7466))|((~WX7130));
assign II3689 = ((~WX638))|((~_2081_));
assign II6296 = ((~II6286))|((~II6294));
assign WX3008 = (WX3787&WX3009);
assign WX909 = ((~II2290))|((~II2291));
assign WX3832 = ((~II11609))|((~II11610));
assign WX4375 = (WX4378&RESET);
assign II2019 = ((~WX1001))|((~WX647));
assign WX2613 = (WX2531&WX2556);
assign II6870 = ((~II6860))|((~II6868));
assign II2143 = ((~WX1001))|((~WX655));
assign WX3226 = ((~WX3479));
assign WX179 = (_2098_&WX1004);
assign WX6119 = ((~WX6118));
assign II26917 = ((~WX8760))|((~WX8461));
assign II10191 = ((~WX3307))|((~II10183));
assign WX6740 = ((~WX7468));
assign WX8929 = (WX8927)|(WX8926);
assign WX1630 = (WX1820&WX2297);
assign WX2646 = (WX2644)|(WX2643);
assign WX1294 = (WX1250&WX1263);
assign WX8668 = ((~II26351))|((~II26352));
assign II23248 = ((~WX6976))|((~II23246));
assign II14702 = ((~WX4760))|((~II14700));
assign II3478 = ((~_2092_))|((~II3477));
assign II2135 = ((~II2110))|((~II2134));
assign WX6569 = ((~WX6568));
assign WX11391 = ((~WX11390));
assign WX6046 = (WX5983&RESET);
assign WX4853 = ((~WX4784));
assign WX5800 = ((~WX6041));
assign II30238 = ((~II30248))|((~II30249));
assign WX5349 = ((~WX6175));
assign WX1543 = (WX3703&WX1544);
assign II6472 = ((~II6474))|((~II6475));
assign II3118 = ((~WX585))|((~II3117));
assign WX7305 = (WX7242&RESET);
assign WX176 = (WX182&WX177);
assign II10511 = ((~WX3455))|((~II10509));
assign II10850 = ((~WX3413))|((~WX3477));
assign WX1479 = (WX1477)|(WX1476);
assign WX6112 = ((~WX6092));
assign II30341 = ((~WX9780))|((~II30340));
assign WX8930 = ((~WX8929));
assign II30861 = ((~WX10053))|((~II30860));
assign II30162 = ((~WX9832))|((~WX9896));
assign WX3304 = (WX3241&RESET);
assign WX2209 = ((~II6512))|((~II6513));
assign WX2015 = (WX1952&RESET);
assign II27529 = ((~II27531))|((~II27532));
assign WX7597 = ((~II23312))|((~II23313));
assign WX295 = (WX521&WX1004);
assign II18032 = ((~II18022))|((~II18030));
assign WX5143 = (WX5113&WX5142);
assign WX3689 = ((~WX3688));
assign II18534 = ((~II18536))|((~II18537));
assign II30466 = ((~II30456))|((~II30464));
assign II22270 = ((~II22260))|((~II22268));
assign WX6606 = (WX6964&WX7469);
assign WX8180 = (WX8959&WX8181);
assign WX6225 = ((~WX6224));
assign WX5621 = (WX5715&WX6176);
assign II35526 = ((~WX10976))|((~II35525));
assign II26368 = ((~II26358))|((~II26366));
assign WX11376 = ((~WX11375));
assign WX2025 = (WX1962&RESET);
assign II2306 = ((~WX729))|((~II2305));
assign WX401 = ((~WX1003));
assign WX3650 = (WX3174&WX3651);
assign II22385 = ((~WX7466))|((~WX7134));
assign WX4751 = (WX4688&RESET);
assign WX1682 = (_2115_&WX2297);
assign WX2754 = (WX2752)|(WX2751);
assign II30037 = ((~II30039))|((~II30040));
assign WX7417 = ((~WX7391));
assign WX8312 = ((~WX8735));
assign II14825 = ((~WX4704))|((~II14824));
assign II18185 = ((~II18161))|((~II18177));
assign WX11192 = (WX11129&RESET);
assign WX6598 = (WX6609&WX7468);
assign WX11040 = (WX10756&RESET);
assign WX9925 = (WX9862&RESET);
assign II15487 = ((~_2204_))|((~II15485));
assign WX4065 = (WX4063)|(WX4062);
assign WX7540 = ((~WX7539));
assign II34105 = ((~WX11121))|((~WX11185));
assign WX2915 = (WX2926&WX3589);
assign II30146 = ((~II30148))|((~II30149));
assign WX10898 = ((~WX11321));
assign II2817 = ((~II2792))|((~II2816));
assign WX5736 = ((~WX6105));
assign WX8914 = ((~WX8763));
assign II27303 = ((~WX8355))|((~WX8277));
assign WX4747 = (WX4684&RESET);
assign WX6642 = ((~WX7468));
assign WX170 = (DATA_9_22&WX171);
assign II35696 = ((~_2342_))|((~II35694));
assign II3572 = ((~_2100_))|((~II3570));
assign WX7622 = (WX7620)|(WX7619);
assign II34687 = ((~WX11095))|((~II34686));
assign II10556 = ((~WX3588))|((~WX3267));
assign II23568 = ((~WX7080))|((~II23567));
assign WX590 = ((~WX558));
assign WX603 = ((~WX571));
assign DATA_9_6 = ((~WX1186));
assign WX3054 = ((~WX3053));
assign WX8349 = ((~WX8317));
assign II6860 = ((~II6862))|((~II6863));
assign WX10610 = (WX10608)|(WX10607);
assign II34795 = ((~II34770))|((~II34794));
assign II3690 = ((~WX638))|((~II3689));
assign WX1538 = (WX1549&WX2296);
assign WX3553 = ((~WX3552));
assign II3405 = ((~WX539))|((~II3403));
assign II34237 = ((~II34212))|((~II34236));
assign WX6405 = ((~II19528))|((~II19529));
assign WX6098 = ((~II18837))|((~II18838));
assign WX7069 = ((~WX7037));
assign WX6591 = (WX6589)|(WX6588);
assign WX4797 = ((~II14584))|((~II14585));
assign WX10553 = ((~WX11348));
assign WX558 = ((~WX985));
assign II14730 = ((~II14732))|((~II14733));
assign WX7444 = ((~WX7443));
assign WX11601 = ((~II35716))|((~II35717));
assign WX5085 = (WX5083)|(WX5082);
assign WX1353 = (WX1351)|(WX1350);
assign WX3547 = ((~WX3546));
assign II10959 = ((~WX3588))|((~WX3293));
assign WX7590 = ((~II23299))|((~II23300));
assign II22424 = ((~WX7200))|((~II22423));
assign WX8794 = (WX8342&WX8795);
assign WX3001 = ((~WX3589));
assign WX2716 = (WX2714)|(WX2713);
assign WX8755 = ((~TM0));
assign II14748 = ((~WX4881))|((~II14747));
assign II26908 = ((~II26884))|((~II26900));
assign WX6560 = (_2264_&WX7469);
assign II30642 = ((~II30644))|((~II30645));
assign WX6274 = ((~WX6273));
assign II6379 = ((~II6381))|((~II6382));
assign II11588 = ((~WX3206))|((~II11587));
assign II3158 = ((~WX501))|((~II3156));
assign WX1360 = (_2138_&WX2297);
assign II2672 = ((~WX689))|((~II2670));
assign WX5603 = (_2208_&WX6176);
assign II27407 = ((~WX8363))|((~WX8293));
assign WX1104 = ((~II3235))|((~II3236));
assign II15315 = ((~WX4478))|((~II15314));
assign WX10552 = (DATA_0_19&WX10553);
assign WX10210 = ((~WX10209));
assign II6358 = ((~II6348))|((~II6356));
assign WX190 = (WX196&WX191);
assign II18419 = ((~WX5907))|((~II18418));
assign II15586 = ((~WX4498))|((~II15585));
assign WX2774 = ((~WX2773));
assign WX9694 = ((~WX9950));
assign WX2656 = (WX2654)|(WX2653);
assign WX10688 = (WX10694&WX10689);
assign II26955 = ((~WX8527))|((~II26947));
assign WX698 = (WX426&RESET);
assign II18791 = ((~WX5931))|((~II18790));
assign II2794 = ((~WX1002))|((~WX697));
assign II30410 = ((~WX9848))|((~WX9912));
assign WX6756 = (_2250_&WX7469);
assign WX5523 = (WX5701&WX6176);
assign II22347 = ((~II22337))|((~II22345));
assign WX7818 = (WX7816)|(WX7815);
assign WX920 = ((~II2631))|((~II2632));
assign WX93 = ((~WX1003));
assign WX2795 = ((~WX3590));
assign WX11296 = ((~WX11270));
assign II19386 = ((~WX5705))|((~II19384));
assign WX10559 = ((~WX10550));
assign II2623 = ((~WX813))|((~WX877));
assign WX4987 = (WX4985)|(WX4984);
assign II10136 = ((~II10138))|((~II10139));
assign WX826 = (WX763&RESET);
assign WX9602 = ((~WX10022));
assign WX10223 = ((~WX10222));
assign II34572 = ((~WX11215))|((~II34570));
assign II10882 = ((~WX3415))|((~II10881));
assign WX9903 = (WX9840&RESET);
assign WX4154 = ((~WX4882));
assign II3443 = ((~WX610))|((~II3442));
assign II26714 = ((~II26716))|((~II26717));
assign II23582 = ((~WX7082))|((~II23581));
assign II2544 = ((~II2554))|((~II2555));
assign WX10176 = ((~II31309))|((~II31310));
assign WX6165 = ((~WX6164));
assign II14289 = ((~WX4606))|((~II14281));
assign WX8524 = (WX8461&RESET);
assign WX6083 = ((~II18372))|((~II18373));
assign II18767 = ((~WX5993))|((~WX6057));
assign II3469 = ((~II3471))|((~II3472));
assign II2653 = ((~II2655))|((~II2656));
assign II27693 = ((~_2277_))|((~II27691));
assign II11324 = ((~WX3111))|((~II11322));
assign II34183 = ((~WX11345))|((~WX10999));
assign II26853 = ((~II26863))|((~II26864));
assign II22865 = ((~WX7292))|((~WX7356));
assign WX596 = ((~WX564));
assign WX4114 = (_2190_&WX4883);
assign WX9114 = (WX9125&WX10054);
assign WX7472 = (WX7471&WX7470);
assign WX46 = (WX44)|(WX43);
assign II14173 = ((~WX4662))|((~WX4726));
assign II26492 = ((~II26482))|((~II26490));
assign II18954 = ((~WX6005))|((~II18953));
assign WX73 = ((~WX1004));
assign WX7949 = ((~WX8761));
assign II10461 = ((~II10471))|((~II10472));
assign WX6924 = (_2238_&WX7469);
assign WX5846 = (WX5430&RESET);
assign WX10241 = (WX9657&WX10242);
assign WX7199 = (WX7136&RESET);
assign II23222 = ((~WX6972))|((~II23220));
assign II14352 = ((~WX4610))|((~II14351));
assign II18340 = ((~II18316))|((~II18332));
assign WX10880 = (WX10883&RESET);
assign II6513 = ((~II6503))|((~II6511));
assign WX10094 = (WX9636&WX10095);
assign WX9500 = (WX9594&WX10055);
assign WX9497 = (WX11559&WX9498);
assign II14492 = ((~II14482))|((~II14490));
assign WX2153 = (WX2090&RESET);
assign WX4591 = (WX4528&RESET);
assign WX500 = (WX503&RESET);
assign WX2934 = (WX5045&WX2935);
assign II6652 = ((~WX2044))|((~II6651));
assign WX3376 = (WX3313&RESET);
assign WX10181 = ((~WX10180));
assign II23469 = ((~WX7010))|((~II23467));
assign WX4421 = (WX4424&RESET);
assign WX7261 = (WX7198&RESET);
assign WX1005 = ((~WX996));
assign II22464 = ((~WX7330))|((~II22462));
assign II15550 = ((~WX4493))|((~_2201_));
assign WX876 = (WX813&RESET);
assign WX7838 = (WX7836)|(WX7835);
assign II18410 = ((~II18412))|((~II18413));
assign WX7724 = ((~II23715))|((~II23716));
assign WX3969 = ((~WX3968));
assign WX3296 = (WX3233&RESET);
assign WX1530 = ((~WX2297));
assign WX10952 = ((~WX10920));
assign II23533 = ((~_2240_))|((~II23532));
assign WX4789 = ((~II14336))|((~II14337));
assign WX1505 = (WX2389&WX1506);
assign II10167 = ((~II10169))|((~II10170));
assign WX3978 = (WX4372&WX4883);
assign WX3499 = ((~II10424))|((~II10425));
assign II26746 = ((~WX8577))|((~WX8641));
assign WX1733 = ((~WX1732));
assign WX7979 = (_2287_&WX8762);
assign WX3065 = ((~WX3590));
assign II30116 = ((~WX10052))|((~WX9702));
assign WX9284 = ((~WX10054));
assign II2012 = ((~II2002))|((~II2010));
assign WX3336 = (WX3273&RESET);
assign WX1171 = (WX1169)|(WX1168);
assign II19613 = ((~_2225_))|((~II19611));
assign WX2392 = (WX1886&WX2393);
assign II35119 = ((~WX10926))|((~II35118));
assign WX9147 = (WX11384&WX9148);
assign WX2949 = ((~WX3590));
assign WX4893 = (WX4892&WX4884);
assign II26823 = ((~II26825))|((~II26826));
assign WX8149 = ((~WX8762));
assign II18907 = ((~WX6174))|((~WX5875));
assign WX9323 = ((~WX9322));
assign WX6699 = (WX6697)|(WX6696);
assign WX9855 = (WX9792&RESET);
assign II10726 = ((~WX3405))|((~WX3469));
assign II14475 = ((~WX4618))|((~II14467));
assign II10611 = ((~II10601))|((~II10609));
assign WX8974 = ((~II27473))|((~II27474));
assign WX10432 = (WX10430)|(WX10429);
assign WX6885 = (WX6883)|(WX6882);
assign WX11126 = (WX11063&RESET);
assign WX1123 = ((~WX1122));
assign II10718 = ((~WX3341))|((~II10710));
assign WX10696 = (WX11510&WX10697);
assign II30317 = ((~WX9842))|((~WX9906));
assign WX1310 = (WX1243&WX1263);
assign WX5110 = ((~II15493))|((~II15494));
assign WX2911 = ((~WX3590));
assign II30707 = ((~WX9740))|((~II30705));
assign WX6528 = (WX6539&WX7468);
assign WX5810 = ((~WX6061));
assign WX1449 = (WX2361&WX1450);
assign WX1711 = (WX3787&WX1712);
assign II19411 = ((~WX5778))|((~II19410));
assign WX6364 = (WX6362)|(WX6361);
assign WX11140 = (WX11077&RESET);
assign WX704 = (WX468&RESET);
assign WX5037 = ((~WX5036));
assign WX6079 = ((~II18248))|((~II18249));
assign II18140 = ((~WX5889))|((~II18139));
assign WX5122 = ((~II15593))|((~II15594));
assign WX3206 = ((~WX3439));
assign II10775 = ((~WX3281))|((~II10773));
assign WX8057 = ((~WX8048));
assign WX9406 = ((~WX9397));
assign II30837 = ((~WX9812))|((~II30836));
assign WX3492 = ((~II10207))|((~II10208));
assign II23609 = ((~WX7086))|((~_2258_));
assign WX6825 = (WX6823)|(WX6822);
assign WX546 = (WX483&RESET);
assign WX9095 = (WX10063&WX9096);
assign WX10122 = (WX9640&WX10123);
assign WX6242 = (WX6241&WX6177);
assign WX5758 = ((~WX5726));
assign WX1389 = (WX3626&WX1390);
assign II23539 = ((~WX7108))|((~_2268_));
assign WX6850 = (WX6861&WX7468);
assign II31663 = ((~_2315_))|((~II31661));
assign WX391 = ((~WX1004));
assign WX10129 = (WX9641&WX10130);
assign II34398 = ((~II34408))|((~II34409));
assign WX2247 = ((~WX2220));
assign II22656 = ((~II22631))|((~II22655));
assign WX6927 = (WX6925)|(WX6924);
assign II23511 = ((~WX7097))|((~II23510));
assign II18389 = ((~II18379))|((~II18387));
assign II11296 = ((~WX3184))|((~WX3107));
assign WX1176 = (WX604&WX1177);
assign WX165 = (_2099_&WX1004);
assign II18482 = ((~II18472))|((~II18480));
assign WX927 = ((~II2848))|((~II2849));
assign II35469 = ((~WX10953))|((~WX10887));
assign WX935 = ((~WX934));
assign WX7939 = ((~WX8762));
assign WX7524 = (WX7522)|(WX7521);
assign II2141 = ((~II2151))|((~II2152));
assign WX4918 = ((~WX4917));
assign WX4325 = (WX6387&WX4326);
assign WX2341 = ((~II7136))|((~II7137));
assign WX6433 = ((~II19724))|((~II19725));
assign WX5562 = (WX7652&WX5563);
assign WX10454 = (DATA_0_26&WX10455);
assign WX2529 = ((~II7534))|((~II7535));
assign WX756 = (WX693&RESET);
assign WX4865 = ((~WX4790));
assign WX3661 = ((~WX3660));
assign WX10998 = (WX10462&RESET);
assign II26855 = ((~WX8760))|((~WX8457));
assign II30734 = ((~II30744))|((~II30745));
assign II35211 = ((~WX10847))|((~II35209));
assign WX9535 = (WX9538&RESET);
assign WX9505 = ((~WX9504));
assign WX4215 = (WX4213)|(WX4212);
assign WX6813 = (WX8924&WX6814);
assign II34981 = ((~II34956))|((~II34980));
assign II30425 = ((~II30427))|((~II30428));
assign II15529 = ((~WX4522))|((~_2204_));
assign WX9737 = (WX9393&RESET);
assign II26716 = ((~WX8575))|((~II26715));
assign II6264 = ((~II6239))|((~II6263));
assign WX4323 = (WX4321)|(WX4320);
assign WX4003 = (WX6226&WX4004);
assign II15499 = ((~II15501))|((~II15502));
assign II3130 = ((~WX586))|((~WX497));
assign WX2908 = (WX2906)|(WX2905);
assign WX5337 = (_2227_&WX6176);
assign WX10472 = (WX11398&WX10473);
assign WX4457 = ((~WX4840));
assign WX2836 = (WX4996&WX2837);
assign II26691 = ((~II26667))|((~II26683));
assign WX9651 = ((~WX9619));
assign WX7086 = ((~WX7320));
assign WX8891 = (WX8890&WX8763);
assign WX3918 = (_2204_&WX4883);
assign II27600 = ((~WX8377))|((~_2292_));
assign II14715 = ((~II14717))|((~II14718));
assign WX7570 = (WX7569&WX7470);
assign II27251 = ((~WX8351))|((~WX8269));
assign WX490 = (WX493&RESET);
assign WX8738 = ((~WX8666));
assign WX9416 = (WX9582&WX10055);
assign WX6370 = ((~WX6177));
assign II30610 = ((~II30620))|((~II30621));
assign II11594 = ((~WX3207))|((~_2162_));
assign II11525 = ((~WX3229))|((~II11524));
assign WX7729 = (WX7699&WX7728);
assign WX5229 = (WX5659&WX6176);
assign II26156 = ((~II26158))|((~II26159));
assign WX1662 = ((~WX1653));
assign WX3716 = ((~WX3715));
assign WX6050 = (WX5987&RESET);
assign II35562 = ((~WX10956))|((~II35561));
assign II7709 = ((~WX1934))|((~II7708));
assign WX150 = (WX148)|(WX147);
assign WX4557 = (WX4165&RESET);
assign WX4060 = ((~WX4883));
assign WX3820 = ((~II11525))|((~II11526));
assign II34951 = ((~II34941))|((~II34949));
assign WX2520 = (WX2518)|(WX2517);
assign WX4782 = ((~II14119))|((~II14120));
assign WX1465 = (WX1463)|(WX1462);
assign II34770 = ((~II34780))|((~II34781));
assign II31712 = ((~_2307_))|((~II31710));
assign WX3627 = ((~II11128))|((~II11129));
assign II22290 = ((~II22300))|((~II22301));
assign II18155 = ((~II18130))|((~II18154));
assign WX5890 = (WX5827&RESET);
assign II27253 = ((~WX8269))|((~II27251));
assign WX370 = ((~WX369));
assign WX1916 = ((~WX2152));
assign DATA_9_17 = ((~WX1109));
assign WX10049 = ((~TM0));
assign WX11517 = ((~WX11516));
assign II35367 = ((~WX10871))|((~II35365));
assign II2282 = ((~WX791))|((~WX855));
assign WX7895 = (_2293_&WX8762);
assign II3565 = ((~_2101_))|((~II3563));
assign WX11591 = ((~II35646))|((~II35647));
assign WX8206 = (WX8204)|(WX8203);
assign WX4075 = (WX4073)|(WX4072);
assign WX10027 = ((~WX9957));
assign II26233 = ((~II26243))|((~II26244));
assign II22748 = ((~II22724))|((~II22740));
assign II15557 = ((~WX4494))|((~_2200_));
assign II10486 = ((~II10461))|((~II10485));
assign WX10293 = ((~II31606))|((~II31607));
assign WX10926 = ((~WX10894));
assign II7696 = ((~_2113_))|((~II7694));
assign WX10108 = (WX9638&WX10109);
assign II18443 = ((~WX6173))|((~II18442));
assign WX10531 = ((~WX10522));
assign II31192 = ((~WX9639))|((~II31191));
assign WX9523 = (WX9521)|(WX9520);
assign II19668 = ((~WX5803))|((~II19667));
assign WX5551 = (WX5705&WX6176);
assign WX11409 = ((~WX11349));
assign II22261 = ((~WX7466))|((~WX7126));
assign II6327 = ((~II6317))|((~II6325));
assign II18720 = ((~II18722))|((~II18723));
assign WX7941 = (WX8263&WX8762);
assign WX6835 = ((~WX6834));
assign II3054 = ((~WX485))|((~II3052));
assign WX9674 = ((~WX9910));
assign II2516 = ((~WX1002))|((~II2515));
assign WX7970 = (WX8854&WX7971);
assign WX5706 = (WX5709&RESET);
assign II7576 = ((~WX1912))|((~II7575));
assign II7526 = ((~WX1905))|((~_2139_));
assign II22021 = ((~WX7174))|((~II22020));
assign II19555 = ((~WX5786))|((~_2233_));
assign WX10102 = ((~WX10056));
assign II19550 = ((~_2234_))|((~II19548));
assign II26079 = ((~II26081))|((~II26082));
assign WX6137 = ((~WX6136));
assign WX10385 = ((~WX11348));
assign II14314 = ((~WX4880))|((~II14313));
assign WX3246 = (WX2746&RESET);
assign WX620 = ((~WX853));
assign WX8771 = ((~II27096))|((~II27097));
assign WX9139 = (WX9137)|(WX9136);
assign WX6799 = (WX8917&WX6800);
assign WX3167 = ((~WX3135));
assign II11652 = ((~_2153_))|((~II11650));
assign WX10573 = ((~WX10564));
assign II18094 = ((~II18084))|((~II18092));
assign WX10331 = (WX10307&WX10314);
assign II6442 = ((~WX2094))|((~WX2158));
assign WX7576 = ((~II23273))|((~II23274));
assign WX415 = ((~WX1003));
assign WX11283 = ((~WX11282));
assign WX2984 = ((~WX2983));
assign WX6196 = (WX6194)|(WX6193);
assign II31593 = ((~_2326_))|((~II31591));
assign II6487 = ((~II6497))|((~II6498));
assign WX6212 = ((~WX6211));
assign WX9654 = ((~WX9622));
assign WX9775 = (WX9712&RESET);
assign WX6237 = ((~WX6177));
assign WX3665 = ((~WX3591));
assign WX7414 = ((~WX7413));
assign II14694 = ((~II14684))|((~II14692));
assign II30744 = ((~WX9806))|((~II30743));
assign WX398 = ((~WX397));
assign WX6500 = (WX6511&WX7468);
assign WX10836 = (WX10839&RESET);
assign II23285 = ((~WX7061))|((~WX6982));
assign WX10798 = ((~WX10797));
assign II14568 = ((~WX4624))|((~II14560));
assign WX4233 = (WX4231)|(WX4230);
assign II15249 = ((~WX4473))|((~WX4392));
assign II2253 = ((~WX853))|((~II2251));
assign WX10732 = (WX10730)|(WX10729);
assign II11141 = ((~WX3172))|((~II11140));
assign WX11366 = (WX10926&WX11367);
assign WX9589 = (WX9592&RESET);
assign II26561 = ((~WX8565))|((~II26560));
assign II31257 = ((~WX9644))|((~II31256));
assign II18071 = ((~WX6173))|((~II18070));
assign II10802 = ((~II10812))|((~II10813));
assign II3635 = ((~_2090_))|((~II3633));
assign WX7646 = ((~II23403))|((~II23404));
assign WX6325 = ((~II19346))|((~II19347));
assign II23687 = ((~WX7099))|((~II23686));
assign II15656 = ((~WX4509))|((~II15655));
assign WX4043 = (WX4041)|(WX4040);
assign WX7831 = ((~WX8762));
assign WX8012 = (WX8875&WX8013);
assign WX9411 = (WX9409)|(WX9408);
assign WX1781 = (WX1784&RESET);
assign WX1924 = ((~WX2168));
assign II7619 = ((~_2126_))|((~II7617));
assign WX7956 = (WX8847&WX7957);
assign II6086 = ((~WX2294))|((~WX1944));
assign WX4034 = (WX4380&WX4883);
assign WX1681 = (WX1679)|(WX1678);
assign II2049 = ((~II2051))|((~II2052));
assign WX10977 = ((~WX11223));
assign II23680 = ((~WX7098))|((~II23679));
assign WX1842 = ((~WX2260));
assign WX11624 = (WX11600&WX11607);
assign WX7386 = ((~II22687))|((~II22688));
assign WX1410 = ((~WX1401));
assign II26732 = ((~WX8760))|((~II26731));
assign WX3596 = (WX3594)|(WX3593);
assign II18730 = ((~II18720))|((~II18728));
assign WX10739 = ((~WX11348));
assign II31551 = ((~_2332_))|((~II31549));
assign II30729 = ((~II30719))|((~II30727));
assign II30117 = ((~WX10052))|((~II30116));
assign WX8630 = (WX8567&RESET);
assign WX4595 = (WX4532&RESET);
assign WX8068 = (WX8903&WX8069);
assign WX5643 = ((~WX6175));
assign WX8510 = (WX8447&RESET);
assign WX4266 = ((~WX4882));
assign WX2169 = (WX2106&RESET);
assign WX7016 = ((~WX7436));
assign II22569 = ((~II22579))|((~II22580));
assign II26516 = ((~WX8435))|((~II26514));
assign WX6659 = (WX8847&WX6660);
assign WX3647 = ((~WX3646));
assign WX8118 = (WX8116)|(WX8115);
assign WX3778 = (WX3776)|(WX3775);
assign WX11361 = (WX11359)|(WX11358);
assign II18729 = ((~WX5927))|((~II18728));
assign II7555 = ((~WX1909))|((~II7554));
assign WX1548 = ((~WX2297));
assign WX3597 = ((~WX3596));
assign II18589 = ((~II18564))|((~II18588));
assign WX8371 = ((~WX8597));
assign II30784 = ((~WX9936))|((~II30782));
assign WX1499 = (WX1497)|(WX1496);
assign WX1014 = (WX1013&WX1005);
assign II2331 = ((~WX667))|((~II2329));
assign WX5587 = ((~WX6175));
assign II27421 = ((~WX8364))|((~II27420));
assign II10704 = ((~II10694))|((~II10702));
assign II6963 = ((~II6953))|((~II6961));
assign WX6387 = ((~WX6386));
assign WX1591 = (WX1589)|(WX1588);
assign II23602 = ((~WX7085))|((~_2259_));
assign II35547 = ((~_2336_))|((~II35539));
assign II6645 = ((~WX2295))|((~II6644));
assign WX3680 = (WX3678)|(WX3677);
assign II26359 = ((~WX8759))|((~WX8425));
assign WX2510 = (WX2509&WX2298);
assign WX768 = (WX705&RESET);
assign WX7023 = ((~WX7450));
assign WX1510 = (WX1521&WX2296);
assign WX10912 = ((~WX11285));
assign II22549 = ((~II22539))|((~II22547));
assign WX1605 = (WX1603)|(WX1602);
assign WX9861 = (WX9798&RESET);
assign II26236 = ((~WX8759))|((~II26235));
assign WX4171 = (WX6310&WX4172);
assign WX10145 = (WX10143)|(WX10142);
assign WX1377 = (WX1375)|(WX1374);
assign II35093 = ((~WX10924))|((~II35092));
assign II27514 = ((~II27516))|((~II27517));
assign WX2879 = ((~WX3590));
assign II19125 = ((~WX5756))|((~II19124));
assign II3299 = ((~WX599))|((~WX523));
assign WX7822 = (WX7828&WX7823);
assign WX694 = (WX398&RESET);
assign II22593 = ((~II22569))|((~II22585));
assign II14244 = ((~II14234))|((~II14242));
assign WX8980 = ((~WX8979));
assign II14196 = ((~WX4600))|((~II14188));
assign II14058 = ((~II14048))|((~II14056));
assign WX6800 = ((~WX7469));
assign WX8087 = (WX8098&WX8761);
assign II26203 = ((~II26205))|((~II26206));
assign WX1566 = (WX1577&WX2296);
assign WX11481 = ((~WX11480));
assign WX8532 = (WX8469&RESET);
assign II2585 = ((~WX747))|((~II2584));
assign WX990 = ((~WX913));
assign WX1490 = (WX1800&WX2297);
assign II30396 = ((~WX10052))|((~II30395));
assign II18635 = ((~WX5921))|((~II18627));
assign WX6349 = ((~WX6177));
assign WX1554 = ((~WX2296));
assign WX6354 = (WX6353&WX6177);
assign WX6553 = (WX6551)|(WX6550);
assign WX2721 = ((~WX3589));
assign II26963 = ((~WX8591))|((~WX8655));
assign II31309 = ((~WX9648))|((~II31308));
assign WX7009 = (WX7012&RESET);
assign II18372 = ((~II18347))|((~II18371));
assign WX3456 = (WX3393&RESET);
assign II6599 = ((~WX2168))|((~II6597));
assign WX5021 = ((~WX4884));
assign WX7988 = ((~WX7987));
assign WX10216 = ((~WX10215));
assign WX9128 = (WX9139&WX10054);
assign WX5854 = (WX5486&RESET);
assign WX4911 = ((~WX4910));
assign II30890 = ((~II30892))|((~II30893));
assign WX5798 = ((~WX6037));
assign WX11593 = ((~II35660))|((~II35661));
assign WX7745 = (WX7721&WX7728);
assign WX8008 = (WX10168&WX8009);
assign WX1023 = ((~WX1005));
assign WX3997 = ((~WX3996));
assign II22547 = ((~WX7208))|((~II22539));
assign II6078 = ((~II6053))|((~II6077));
assign WX10905 = ((~WX11335));
assign WX9961 = ((~II30356))|((~II30357));
assign II18580 = ((~II18582))|((~II18583));
assign II18931 = ((~II18921))|((~II18929));
assign WX7502 = ((~WX7470));
assign WX3170 = ((~WX3138));
assign WX6152 = ((~WX6080));
assign WX4254 = (_2180_&WX4883);
assign WX7981 = ((~WX8762));
assign II18697 = ((~WX5925))|((~II18689));
assign WX3796 = (WX3795&WX3591);
assign WX3026 = ((~WX3025));
assign WX5858 = (WX5514&RESET);
assign WX4318 = ((~WX4309));
assign WX4358 = ((~WX4883));
assign II26419 = ((~II26429))|((~II26430));
assign WX7577 = (WX7576&WX7470);
assign II18668 = ((~II18658))|((~II18666));
assign II34385 = ((~WX11139))|((~II34384));
assign II31284 = ((~WX9566))|((~II31282));
assign II18349 = ((~WX6173))|((~WX5839));
assign WX10337 = (WX10283&WX10314);
assign WX7959 = ((~WX7950));
assign II31732 = ((~WX9691))|((~II31731));
assign II22402 = ((~WX7326))|((~II22400));
assign WX10273 = ((~WX10272));
assign II31592 = ((~WX9668))|((~II31591));
assign II18659 = ((~WX6174))|((~WX5859));
assign II14095 = ((~II14097))|((~II14098));
assign II6699 = ((~II6689))|((~II6697));
assign II10765 = ((~II10740))|((~II10764));
assign II10316 = ((~WX3315))|((~II10315));
assign WX9008 = ((~II27657))|((~II27658));
assign II19073 = ((~WX5752))|((~II19072));
assign WX6016 = (WX5953&RESET);
assign II35682 = ((~_2345_))|((~II35680));
assign II34345 = ((~WX11073))|((~II34337));
assign WX2213 = ((~II6636))|((~II6637));
assign II23730 = ((~_2238_))|((~II23728));
assign WX2545 = ((~II7646))|((~II7647));
assign WX10793 = (WX10887&WX11348);
assign WX5874 = (WX5626&RESET);
assign WX2788 = ((~WX2787));
assign WX4522 = ((~WX4778));
assign WX3474 = (WX3411&RESET);
assign WX4147 = (WX5003&WX4148);
assign WX2635 = (WX2646&WX3589);
assign WX7361 = (WX7298&RESET);
assign II30969 = ((~WX9884))|((~II30968));
assign II14640 = ((~WX4756))|((~II14638));
assign WX6626 = (WX6637&WX7468);
assign WX10445 = ((~WX11348));
assign WX1072 = ((~WX1005));
assign WX5569 = ((~WX5560));
assign II14932 = ((~II14934))|((~II14935));
assign WX11327 = ((~WX11326));
assign WX5074 = ((~II15419))|((~II15420));
assign WX868 = (WX805&RESET);
assign II34758 = ((~WX11227))|((~II34756));
assign WX6518 = (_2267_&WX7469);
assign WX3354 = (WX3291&RESET);
assign II31295 = ((~WX9647))|((~WX9568));
assign II31439 = ((~WX9658))|((~II31438));
assign II7239 = ((~WX1887))|((~WX1806));
assign WX2264 = ((~WX2263));
assign WX5809 = ((~WX6059));
assign WX9093 = (WX9091)|(WX9090);
assign WX6788 = (WX6990&WX7469);
assign WX211 = (WX509&WX1004);
assign II14725 = ((~II14715))|((~II14723));
assign WX10042 = ((~WX10041));
assign WX5647 = ((~WX6176));
assign II27628 = ((~WX8381))|((~_2288_));
assign WX1596 = ((~WX2296));
assign WX2309 = ((~WX2298));
assign II30324 = ((~II30300))|((~II30316));
assign II14035 = ((~WX4880))|((~II14034));
assign WX5103 = (WX5102&WX4884);
assign II10291 = ((~II10293))|((~II10294));
assign II26040 = ((~II26016))|((~II26032));
assign II22694 = ((~II22696))|((~II22697));
assign II19504 = ((~II19506))|((~II19507));
assign WX10745 = ((~WX11347));
assign WX7661 = (WX7660&WX7470);
assign WX9288 = ((~WX10055));
assign II6707 = ((~WX2295))|((~II6706));
assign WX10770 = ((~WX10769));
assign WX3384 = (WX3321&RESET);
assign WX8412 = (WX7876&RESET);
assign WX6680 = ((~WX6671));
assign WX3192 = ((~WX3160));
assign II27671 = ((~WX8388))|((~II27670));
assign II27616 = ((~_2290_))|((~II27614));
assign WX6360 = ((~II19411))|((~II19412));
assign WX7209 = (WX7146&RESET);
assign WX5654 = ((~WX5653));
assign II26268 = ((~WX8419))|((~II26266));
assign II35625 = ((~WX10965))|((~II35624));
assign WX7066 = ((~WX7034));
assign WX7412 = ((~WX7411));
assign II34584 = ((~II34594))|((~II34595));
assign II7293 = ((~WX1814))|((~II7291));
assign DATA_9_25 = ((~WX1053));
assign WX8065 = ((~WX8762));
assign WX11000 = (WX10476&RESET);
assign WX2465 = ((~WX2464));
assign WX1076 = ((~II3183))|((~II3184));
assign II22966 = ((~II22941))|((~II22965));
assign WX4383 = (WX4386&RESET);
assign II15514 = ((~II15516))|((~II15517));
assign II6063 = ((~WX2006))|((~II6062));
assign II30310 = ((~WX9778))|((~II30309));
assign II6481 = ((~II6456))|((~II6480));
assign II2484 = ((~WX1002))|((~WX677));
assign WX7912 = (WX7910)|(WX7909);
assign II26273 = ((~WX8483))|((~II26265));
assign WX1963 = (WX1523&RESET);
assign II2066 = ((~WX777))|((~II2065));
assign II26305 = ((~WX8485))|((~II26304));
assign II14398 = ((~II14373))|((~II14397));
assign WX6759 = (WX6757)|(WX6756);
assign WX10966 = ((~WX11201));
assign II18614 = ((~WX6047))|((~II18612));
assign WX6671 = (WX6669)|(WX6668);
assign II19674 = ((~WX5805))|((~_2214_));
assign WX7038 = ((~WX7416));
assign WX2666 = (WX2664)|(WX2663);
assign II30200 = ((~II30176))|((~II30192));
assign II23581 = ((~WX7082))|((~_2262_));
assign II2369 = ((~II2359))|((~II2367));
assign II22872 = ((~II22848))|((~II22864));
assign II22154 = ((~WX7310))|((~II22152));
assign WX7815 = (WX8245&WX8762);
assign WX1649 = ((~WX1648));
assign II22184 = ((~WX7248))|((~II22183));
assign WX423 = ((~WX1004));
assign WX11460 = ((~WX11459));
assign WX4868 = ((~WX4867));
assign WX4629 = (WX4566&RESET);
assign WX6682 = (WX6693&WX7468);
assign WX2874 = (WX2880&WX2875);
assign II27266 = ((~WX8271))|((~II27264));
assign WX6845 = (WX7645&WX6846);
assign WX2069 = (WX2006&RESET);
assign II18978 = ((~II18968))|((~II18976));
assign WX10470 = (WX10468)|(WX10467);
assign WX4653 = (WX4590&RESET);
assign WX1907 = ((~WX2134));
assign II34090 = ((~WX11345))|((~WX10993));
assign II27344 = ((~WX8283))|((~II27342));
assign II6256 = ((~WX2082))|((~WX2146));
assign II30464 = ((~WX9788))|((~II30456));
assign II30293 = ((~II30269))|((~II30285));
assign WX11352 = (WX10924&WX11353);
assign WX227 = ((~WX1004));
assign WX1328 = (WX1339&WX2296);
assign II30799 = ((~WX10053))|((~II30798));
assign II30071 = ((~WX9890))|((~II30069));
assign II14584 = ((~II14559))|((~II14583));
assign WX6869 = (WX8952&WX6870);
assign WX10050 = ((~TM1));
assign II15380 = ((~WX4483))|((~II15379));
assign WX2274 = ((~WX2273));
assign WX316 = (WX322&WX317);
assign WX8238 = (WX8236)|(WX8235);
assign II31684 = ((~_2312_))|((~II31682));
assign WX3880 = (WX3836&WX3849);
assign WX1688 = ((~WX2297));
assign WX2792 = (WX2790)|(WX2789);
assign WX5042 = ((~WX4884));
assign II26910 = ((~II26900))|((~II26908));
assign WX11272 = ((~II34919))|((~II34920));
assign WX77 = (WX88&WX1003);
assign WX1486 = (_2129_&WX2297);
assign II30853 = ((~II30843))|((~II30851));
assign WX1217 = (WX1216&WX1005);
assign II34663 = ((~WX11157))|((~WX11221));
assign II31347 = ((~WX9651))|((~WX9576));
assign WX9974 = ((~II30759))|((~II30760));
assign II34639 = ((~II34615))|((~II34631));
assign WX5585 = (WX5596&WX6175);
assign WX1702 = ((~WX2297));
assign II23524 = ((~II23526))|((~II23527));
assign II26296 = ((~II26298))|((~II26299));
assign II10162 = ((~II10152))|((~II10160));
assign II22704 = ((~II22694))|((~II22702));
assign WX69 = ((~WX1004));
assign II26609 = ((~WX8441))|((~II26607));
assign II18867 = ((~II18843))|((~II18859));
assign WX11423 = ((~WX11349));
assign WX6316 = ((~WX6315));
assign WX7019 = ((~WX7442));
assign II15355 = ((~WX4408))|((~II15353));
assign WX4902 = ((~WX4884));
assign WX7712 = ((~II23631))|((~II23632));
assign WX2081 = (WX2018&RESET);
assign WX1274 = (WX1259&WX1263);
assign II10496 = ((~WX3263))|((~II10494));
assign WX9835 = (WX9772&RESET);
assign WX8720 = ((~WX8689));
assign II22354 = ((~WX7466))|((~WX7132));
assign II19254 = ((~WX5766))|((~WX5685));
assign WX9465 = (WX9471&WX9466);
assign WX8754 = ((~TM0));
assign WX9248 = (WX9558&WX10055);
assign II34283 = ((~WX11069))|((~II34275));
assign WX2107 = (WX2044&RESET);
assign WX3635 = (WX3634&WX3591);
assign WX822 = (WX759&RESET);
assign WX1195 = ((~II3404))|((~II3405));
assign WX9951 = ((~II30046))|((~II30047));
assign WX7201 = (WX7138&RESET);
assign II35391 = ((~WX10947))|((~WX10875));
assign WX11536 = (WX11534)|(WX11533);
assign II22688 = ((~II22678))|((~II22686));
assign WX4504 = ((~WX4742));
assign WX5241 = ((~WX6176));
assign WX1585 = (WX3724&WX1586);
assign WX2377 = (WX2376&WX2298);
assign II18813 = ((~II18815))|((~II18816));
assign II26397 = ((~WX8491))|((~II26389));
assign WX9713 = (WX9225&RESET);
assign WX2813 = ((~WX3590));
assign WX1651 = (WX1657&WX1652);
assign WX8810 = (WX8808)|(WX8807);
assign WX3360 = (WX3297&RESET);
assign WX10848 = (WX10851&RESET);
assign WX9293 = (WX9291)|(WX9290);
assign II34526 = ((~WX11021))|((~II34524));
assign II23659 = ((~WX7094))|((~II23658));
assign WX9222 = ((~WX10055));
assign II10844 = ((~II10834))|((~II10842));
assign WX8814 = (WX8813&WX8763);
assign WX4153 = (WX4159&WX4154);
assign II14871 = ((~WX4881))|((~WX4580));
assign II10880 = ((~II10882))|((~II10883));
assign II2112 = ((~WX1001))|((~WX653));
assign WX1374 = (_2137_&WX2297);
assign II10278 = ((~WX3587))|((~II10277));
assign II27609 = ((~_2291_))|((~II27607));
assign II2887 = ((~WX1002))|((~WX703));
assign WX362 = (WX2466&WX363);
assign WX4573 = (WX4277&RESET);
assign II2360 = ((~WX1001))|((~WX669));
assign II10749 = ((~WX3343))|((~II10741));
assign WX3197 = ((~WX3165));
assign WX6496 = (WX6408&WX6435);
assign II35263 = ((~WX10855))|((~II35261));
assign WX6949 = (WX6952&RESET);
assign WX10500 = (WX11412&WX10501);
assign WX8853 = ((~WX8852));
assign WX9341 = (WX9339)|(WX9338);
assign II22477 = ((~II22479))|((~II22480));
assign II11076 = ((~WX3167))|((~II11075));
assign II10075 = ((~WX3363))|((~WX3427));
assign WX10202 = ((~WX10201));
assign WX1622 = (WX1633&WX2296);
assign II31440 = ((~WX9590))|((~II31438));
assign WX4391 = (WX4394&RESET);
assign WX8710 = ((~WX8684));
assign WX8957 = (WX8955)|(WX8954);
assign WX11142 = (WX11079&RESET);
assign II6853 = ((~II6828))|((~II6852));
assign WX52 = (WX50)|(WX49);
assign WX1642 = ((~WX2297));
assign WX10586 = (WX10584)|(WX10583);
assign WX6931 = (WX6929)|(WX6928);
assign WX4765 = (WX4702&RESET);
assign WX2674 = (WX2672)|(WX2671);
assign WX11513 = (WX10947&WX11514);
assign II18351 = ((~WX5839))|((~II18349));
assign II2383 = ((~II2358))|((~II2382));
assign WX3912 = (WX3821&WX3849);
assign WX7617 = ((~WX7616));
assign WX10452 = (WX10450)|(WX10449);
assign II19522 = ((~_2236_))|((~II19520));
assign II2855 = ((~II2857))|((~II2858));
assign WX4194 = (WX4205&WX4882);
assign WX9404 = ((~WX10055));
assign II23630 = ((~WX7089))|((~_2255_));
assign WX9499 = (WX9497)|(WX9496);
assign WX3785 = (WX3783)|(WX3782);
assign WX10410 = (WX10408)|(WX10407);
assign II6891 = ((~II6893))|((~II6894));
assign WX2974 = (WX2972)|(WX2971);
assign WX4517 = ((~WX4768));
assign WX7922 = (WX7920)|(WX7919);
assign WX8673 = ((~II26506))|((~II26507));
assign WX886 = (WX823&RESET);
assign WX326 = (WX324)|(WX323);
assign WX5276 = ((~WX5275));
assign WX9999 = ((~WX9975));
assign WX10919 = ((~WX11299));
assign II14777 = ((~II14779))|((~II14780));
assign II2119 = ((~WX717))|((~II2111));
assign WX1759 = (WX1757)|(WX1756);
assign II35159 = ((~WX10839))|((~II35157));
assign WX9312 = ((~WX10054));
assign WX11646 = (WX11591&WX11607);
assign WX9851 = (WX9788&RESET);
assign WX2956 = ((~WX2955));
assign WX11298 = ((~WX11271));
assign WX3310 = (WX3247&RESET);
assign WX624 = ((~WX861));
assign WX1231 = ((~II3478))|((~II3479));
assign II14817 = ((~WX4640))|((~II14816));
assign WX6402 = ((~RESET));
assign WX9783 = (WX9720&RESET);
assign II26481 = ((~II26491))|((~II26492));
assign II10805 = ((~WX3588))|((~II10804));
assign WX8878 = (WX8354&WX8879);
assign II14273 = ((~II14249))|((~II14265));
assign WX7842 = (WX7840)|(WX7839);
assign WX3282 = (WX2998&RESET);
assign II14832 = ((~II14807))|((~II14831));
assign WX7719 = ((~II23680))|((~II23681));
assign WX9200 = ((~WX10054));
assign II27713 = ((~WX8395))|((~II27712));
assign WX4473 = ((~WX4441));
assign WX6215 = (WX5757&WX6216);
assign WX5411 = (WX5685&WX6176);
assign II30750 = ((~II30752))|((~II30753));
assign II2212 = ((~WX723))|((~II2204));
assign II26329 = ((~WX8759))|((~II26328));
assign II3327 = ((~WX527))|((~II3325));
assign WX10443 = (WX10837&WX11348);
assign WX3753 = ((~II11362))|((~II11363));
assign II34192 = ((~II34182))|((~II34190));
assign WX10310 = ((~II31725))|((~II31726));
assign WX237 = ((~WX1004));
assign WX5263 = (WX5274&WX6175);
assign WX7990 = (WX7996&WX7991);
assign II34268 = ((~II34243))|((~II34267));
assign II26390 = ((~WX8759))|((~WX8427));
assign II22284 = ((~II22259))|((~II22283));
assign WX11652 = (WX11588&WX11607);
assign II18952 = ((~II18954))|((~II18955));
assign II6465 = ((~WX2032))|((~II6457));
assign WX9354 = ((~WX10054));
assign WX10162 = ((~II31283))|((~II31284));
assign WX8113 = ((~WX8104));
assign WX3750 = (WX3748)|(WX3747);
assign WX6218 = ((~WX6217));
assign WX6881 = (WX6879)|(WX6878);
assign WX10314 = ((~WX10281));
assign II3273 = ((~WX597))|((~WX519));
assign II26143 = ((~WX8759))|((~II26142));
assign II7638 = ((~WX1922))|((~_2122_));
assign WX8884 = (WX8883&WX8763);
assign II14656 = ((~WX4566))|((~II14654));
assign WX8676 = ((~II26599))|((~II26600));
assign WX2423 = ((~WX2422));
assign II34619 = ((~WX11027))|((~II34617));
assign WX1855 = ((~WX2286));
assign II31102 = ((~WX9538))|((~II31100));
assign II22510 = ((~WX7467))|((~II22509));
assign II7227 = ((~WX1886))|((~II7226));
assign WX7733 = (WX7726&WX7728);
assign WX1243 = ((~II3578))|((~II3579));
assign DATA_9_24 = ((~WX1060));
assign WX1385 = (WX1391&WX1386);
assign WX2444 = ((~WX2443));
assign WX9362 = ((~WX10055));
assign II10431 = ((~II10433))|((~II10434));
assign II34254 = ((~II34244))|((~II34252));
assign II10821 = ((~WX3475))|((~II10819));
assign WX67 = (_2106_&WX1004);
assign WX3728 = ((~WX3591));
assign II18333 = ((~WX5965))|((~WX6029));
assign II6177 = ((~II6187))|((~II6188));
assign WX7849 = (WX7860&WX8761);
assign II10107 = ((~WX3365))|((~II10106));
assign II15544 = ((~WX4492))|((~II15543));
assign II23518 = ((~_2247_))|((~II23517));
assign II10926 = ((~II10936))|((~II10937));
assign WX5423 = ((~WX6176));
assign WX9436 = (WX9447&WX10054);
assign II26862 = ((~WX8521))|((~II26854));
assign II22741 = ((~WX7284))|((~WX7348));
assign II22207 = ((~WX7186))|((~II22206));
assign II35736 = ((~WX10984))|((~_2335_));
assign WX5395 = ((~WX6176));
assign II19230 = ((~WX5681))|((~II19228));
assign WX4411 = (WX4414&RESET);
assign II31427 = ((~WX9588))|((~II31425));
assign WX8606 = (WX8543&RESET);
assign WX2417 = ((~WX2416));
assign WX5688 = (WX5691&RESET);
assign WX2609 = (WX2533&WX2556);
assign II14063 = ((~II14073))|((~II14074));
assign WX10114 = (WX10113&WX10056);
assign WX7050 = ((~WX7018));
assign II18497 = ((~II18487))|((~II18495));
assign II3431 = ((~WX543))|((~II3429));
assign WX5228 = (WX5226)|(WX5225);
assign II34856 = ((~II34832))|((~II34848));
assign WX3856 = (WX3846&WX3849);
assign WX10930 = ((~WX10898));
assign WX271 = ((~WX262));
assign WX1728 = (WX1834&WX2297);
assign WX2981 = ((~WX3590));
assign II18123 = ((~II18099))|((~II18115));
assign WX7043 = ((~WX7426));
assign WX9155 = ((~WX9154));
assign II31634 = ((~WX9674))|((~II31633));
assign II2917 = ((~II2919))|((~II2920));
assign WX9217 = (WX11419&WX9218);
assign WX8396 = ((~WX8647));
assign WX347 = (_2086_&WX1004);
assign WX7919 = (WX7930&WX8761);
assign WX6849 = ((~WX6848));
assign II35133 = ((~WX10835))|((~II35131));
assign WX9991 = ((~WX9971));
assign WX11443 = (WX10937&WX11444);
assign WX7767 = (WX7712&WX7728);
assign II14823 = ((~II14825))|((~II14826));
assign WX7098 = ((~WX7344));
assign II30022 = ((~II30024))|((~II30025));
assign II7631 = ((~WX1921))|((~_2123_));
assign II1986 = ((~II1996))|((~II1997));
assign WX5291 = (WX5302&WX6175);
assign WX10623 = ((~WX11348));
assign II26250 = ((~WX8545))|((~WX8609));
assign WX278 = (WX2424&WX279);
assign II34595 = ((~II34585))|((~II34593));
assign II2779 = ((~WX823))|((~II2778));
assign II2522 = ((~WX743))|((~II2514));
assign WX11430 = ((~WX11349));
assign WX11190 = (WX11127&RESET);
assign WX1149 = ((~WX1005));
assign WX5252 = (WX5250)|(WX5249);
assign WX2387 = (WX2385)|(WX2384);
assign II2431 = ((~II2421))|((~II2429));
assign WX4673 = (WX4610&RESET);
assign WX7671 = (WX7669)|(WX7668);
assign II14869 = ((~II14879))|((~II14880));
assign WX7339 = (WX7276&RESET);
assign WX2478 = (WX2476)|(WX2475);
assign WX2744 = (WX2742)|(WX2741);
assign WX80 = (WX78)|(WX77);
assign WX7263 = (WX7200&RESET);
assign WX1932 = ((~WX2184));
assign II6558 = ((~WX2038))|((~II6550));
assign WX9241 = (WX9247&WX9242);
assign II18233 = ((~WX5895))|((~II18232));
assign WX9813 = (WX9750&RESET);
assign WX4348 = (WX4359&WX4882);
assign WX3358 = (WX3295&RESET);
assign WX4427 = ((~WX4844));
assign WX7663 = ((~WX7470));
assign WX10593 = (_2349_&WX11348);
assign WX10424 = (WX10422)|(WX10421);
assign II10153 = ((~WX3587))|((~WX3241));
assign WX8353 = ((~WX8321));
assign II10634 = ((~WX3399))|((~II10633));
assign WX4823 = ((~WX4801));
assign WX2245 = ((~WX2219));
assign WX243 = ((~WX234));
assign WX10265 = ((~WX10264));
assign II10836 = ((~WX3588))|((~II10835));
assign II31478 = ((~WX9661))|((~II31477));
assign WX1205 = ((~WX1005));
assign WX2897 = ((~WX3590));
assign II27460 = ((~WX8367))|((~II27459));
assign WX11416 = ((~WX11349));
assign II35302 = ((~WX10861))|((~II35300));
assign II2920 = ((~WX705))|((~II2918));
assign WX11528 = ((~WX11349));
assign II22580 = ((~II22570))|((~II22578));
assign WX6194 = (WX5754&WX6195);
assign II11415 = ((~WX3125))|((~II11413));
assign WX9187 = (WX9185)|(WX9184);
assign II26257 = ((~II26233))|((~II26249));
assign WX7701 = ((~II23554))|((~II23555));
assign II31491 = ((~WX9662))|((~II31490));
assign WX2534 = ((~II7569))|((~II7570));
assign WX1158 = ((~WX1157));
assign II3106 = ((~WX493))|((~II3104));
assign WX10057 = ((~II31088))|((~II31089));
assign II15564 = ((~WX4495))|((~_2199_));
assign II34081 = ((~II34057))|((~II34073));
assign WX578 = ((~WX961));
assign WX7795 = ((~WX8761));
assign II19228 = ((~WX5764))|((~WX5681));
assign WX185 = ((~WX1004));
assign WX1817 = (WX1820&RESET);
assign WX5744 = ((~WX6121));
assign WX10546 = ((~WX10545));
assign II3557 = ((~WX617))|((~II3556));
assign WX4193 = ((~WX4192));
assign II3378 = ((~WX605))|((~II3377));
assign II26482 = ((~II26484))|((~II26485));
assign WX6006 = (WX5943&RESET);
assign WX4121 = (WX4119)|(WX4118);
assign II34261 = ((~WX11131))|((~II34260));
assign II18056 = ((~WX6011))|((~II18054));
assign WX1258 = ((~II3683))|((~II3684));
assign II6273 = ((~WX2294))|((~II6272));
assign WX10633 = ((~WX11347));
assign II10982 = ((~II10957))|((~II10981));
assign WX4333 = ((~WX4332));
assign WX8143 = (WX8154&WX8761);
assign WX377 = ((~WX1004));
assign II30536 = ((~WX9920))|((~II30534));
assign II30086 = ((~WX10052))|((~II30085));
assign II15523 = ((~_2176_))|((~II15522));
assign WX1394 = ((~WX2297));
assign II2050 = ((~WX1001))|((~WX649));
assign WX5135 = ((~II15684))|((~II15685));
assign WX7585 = (WX7061&WX7586);
assign WX1890 = ((~WX1858));
assign WX6150 = ((~WX6079));
assign WX5424 = (WX5422)|(WX5421);
assign WX8160 = (WX8158)|(WX8157);
assign II15329 = ((~WX4404))|((~II15327));
assign WX9793 = (WX9730&RESET);
assign WX11501 = (WX11499)|(WX11498);
assign WX10379 = (WX10390&WX11347);
assign WX7149 = (WX6793&RESET);
assign II30176 = ((~II30186))|((~II30187));
assign WX9179 = (WX10105&WX9180);
assign WX4080 = ((~WX4071));
assign II10014 = ((~WX3359))|((~II10013));
assign WX10816 = (WX10814)|(WX10813);
assign II31128 = ((~WX9542))|((~II31126));
assign WX89 = ((~WX80));
assign II15108 = ((~WX4370))|((~II15106));
assign II35275 = ((~WX10938))|((~II35274));
assign WX4954 = ((~WX4953));
assign II26297 = ((~WX8759))|((~WX8421));
assign WX10825 = ((~WX10816));
assign II10742 = ((~WX3588))|((~WX3279));
assign WX385 = (WX396&WX1003);
assign II34655 = ((~WX11093))|((~II34647));
assign II10651 = ((~WX3273))|((~II10649));
assign II7681 = ((~WX1929))|((~II7680));
assign WX1770 = (WX1840&WX2297);
assign WX9519 = ((~WX9518));
assign II18983 = ((~II18985))|((~II18986));
assign II3260 = ((~WX596))|((~WX517));
assign II2823 = ((~II2833))|((~II2834));
assign II6939 = ((~WX2126))|((~II6938));
assign WX7610 = ((~WX7609));
assign II34834 = ((~WX11346))|((~WX11041));
assign WX6466 = (WX6422&WX6435);
assign WX2487 = ((~WX2486));
assign WX5734 = ((~WX6165));
assign II2641 = ((~WX687))|((~II2639));
assign WX2221 = ((~II6884))|((~II6885));
assign II6728 = ((~II6704))|((~II6720));
assign WX2767 = ((~WX3590));
assign WX5224 = (WX5222)|(WX5221);
assign WX8943 = (WX8941)|(WX8940);
assign WX10133 = ((~WX10132));
assign II2755 = ((~II2730))|((~II2754));
assign WX11259 = ((~II34516))|((~II34517));
assign WX4833 = ((~WX4806));
assign WX6102 = ((~II18961))|((~II18962));
assign WX7538 = (WX7536)|(WX7535);
assign WX11138 = (WX11075&RESET);
assign WX2261 = ((~WX2195));
assign WX3642 = (WX3641&WX3591);
assign II2646 = ((~WX751))|((~II2638));
assign WX345 = ((~WX1003));
assign WX5556 = ((~WX5555));
assign WX5766 = ((~WX5734));
assign II18924 = ((~WX6067))|((~II18922));
assign WX5448 = (WX5446)|(WX5445);
assign WX3704 = ((~II11271))|((~II11272));
assign II2972 = ((~II2947))|((~II2971));
assign WX4166 = (WX4177&WX4882);
assign WX8131 = ((~WX8761));
assign II14948 = ((~WX4712))|((~WX4776));
assign WX9461 = (WX9459)|(WX9458);
assign II10372 = ((~WX3255))|((~II10370));
assign II3705 = ((~_2078_))|((~II3703));
assign WX1253 = ((~II3648))|((~II3649));
assign II26506 = ((~II26481))|((~II26505));
assign II14808 = ((~II14810))|((~II14811));
assign II18194 = ((~WX6173))|((~WX5829));
assign WX4405 = (WX4408&RESET);
assign WX1572 = ((~WX2297));
assign WX9709 = (WX9197&RESET);
assign WX2228 = ((~WX2227));
assign WX10408 = (WX10414&WX10409);
assign II34772 = ((~WX11346))|((~WX11037));
assign WX1829 = (WX1832&RESET);
assign WX6394 = ((~WX6393));
assign WX6690 = (WX6976&WX7469);
assign WX1747 = ((~WX1746));
assign WX7783 = (WX7704&WX7728);
assign II30882 = ((~II30858))|((~II30874));
assign WX6245 = (WX6243)|(WX6242);
assign II10464 = ((~WX3587))|((~II10463));
assign WX6268 = ((~WX6267));
assign WX262 = (WX260)|(WX259);
assign WX1639 = (WX1637)|(WX1636);
assign WX4277 = ((~WX4276));
assign WX6999 = (WX7002&RESET);
assign WX3849 = ((~WX3816));
assign WX10052 = ((~WX10051));
assign WX3953 = (WX3951)|(WX3950);
assign WX4016 = (_2197_&WX4883);
assign II10610 = ((~II10585))|((~II10609));
assign WX2400 = ((~WX2298));
assign II10332 = ((~II10322))|((~II10330));
assign WX5347 = (WX5358&WX6175);
assign WX3862 = (WX3844&WX3849);
assign WX7929 = ((~WX8762));
assign WX7697 = ((~II23518))|((~II23519));
assign II35185 = ((~WX10843))|((~II35183));
assign II30264 = ((~II30254))|((~II30262));
assign WX1693 = (WX1699&WX1694);
assign WX1522 = ((~WX1513));
assign WX5632 = (WX7687&WX5633);
assign WX3146 = ((~WX3575));
assign WX3155 = ((~WX3529));
assign II30595 = ((~II30597))|((~II30598));
assign II14795 = ((~WX4766))|((~II14793));
assign II14012 = ((~II14002))|((~II14010));
assign II19438 = ((~WX5713))|((~II19436));
assign WX6940 = ((~WX7469));
assign II26970 = ((~II26946))|((~II26962));
assign II15601 = ((~_2194_))|((~II15599));
assign II2888 = ((~WX1002))|((~II2887));
assign WX7307 = (WX7244&RESET);
assign II2802 = ((~WX761))|((~II2801));
assign WX3022 = (WX3794&WX3023);
assign WX2551 = ((~II7688))|((~II7689));
assign WX6764 = ((~WX6755));
assign WX9343 = (WX11482&WX9344);
assign WX10753 = ((~WX11348));
assign WX6530 = ((~WX7468));
assign II11722 = ((~_2141_))|((~II11720));
assign II23548 = ((~_2267_))|((~II23546));
assign II6125 = ((~WX2010))|((~II6124));
assign WX199 = ((~WX1004));
assign WX5511 = ((~WX6176));
assign WX9000 = ((~II27601))|((~II27602));
assign WX10059 = (WX9631&WX10060);
assign WX4925 = ((~WX4924));
assign WX4013 = (WX4019&WX4014);
assign WX8967 = ((~II27460))|((~II27461));
assign II34391 = ((~II34367))|((~II34383));
assign WX3605 = ((~WX3604));
assign II30790 = ((~II30765))|((~II30789));
assign II18379 = ((~II18381))|((~II18382));
assign II11194 = ((~WX3091))|((~II11192));
assign II6140 = ((~II6115))|((~II6139));
assign WX6782 = ((~WX7468));
assign WX8661 = ((~II26134))|((~II26135));
assign II11180 = ((~WX3175))|((~II11179));
assign WX8428 = (WX7988&RESET);
assign WX5281 = (_2231_&WX6176);
assign WX7357 = (WX7294&RESET);
assign WX6108 = ((~WX6090));
assign II31586 = ((~_2327_))|((~II31584));
assign WX3731 = ((~WX3730));
assign WX1190 = (WX606&WX1191);
assign II34548 = ((~II34538))|((~II34546));
assign WX355 = ((~WX346));
assign WX10987 = ((~WX11243));
assign WX1847 = ((~WX2270));
assign WX10742 = ((~WX10741));
assign WX4314 = (WX4420&WX4883);
assign II7506 = ((~WX1932))|((~II7505));
assign WX3840 = ((~II11665))|((~II11666));
assign II30714 = ((~II30704))|((~II30712));
assign WX1234 = ((~II3515))|((~II3516));
assign WX8588 = (WX8525&RESET);
assign II34424 = ((~II34414))|((~II34422));
assign WX6646 = ((~WX7469));
assign WX4611 = (WX4548&RESET);
assign WX2045 = (WX1982&RESET);
assign WX6299 = (WX5769&WX6300);
assign II35288 = ((~WX10939))|((~II35287));
assign WX7600 = ((~WX7470));
assign WX5101 = ((~WX5100));
assign II7252 = ((~WX1888))|((~WX1808));
assign WX6961 = (WX6964&RESET);
assign WX4816 = ((~WX4815));
assign II11601 = ((~WX3208))|((~_2161_));
assign II18489 = ((~WX5975))|((~II18488));
assign WX1870 = ((~WX2252));
assign WX4923 = ((~WX4884));
assign WX10986 = ((~WX11241));
assign WX4255 = (WX6352&WX4256);
assign II34646 = ((~II34656))|((~II34657));
assign WX8991 = ((~II27538))|((~II27539));
assign II19332 = ((~WX5772))|((~WX5697));
assign II34764 = ((~II34739))|((~II34763));
assign II14088 = ((~II14063))|((~II14087));
assign WX10367 = (WX10291&WX10314);
assign WX7835 = (WX7846&WX8761);
assign WX2802 = ((~WX2801));
assign WX8097 = ((~WX8762));
assign II35661 = ((~_2349_))|((~II35659));
assign WX4943 = (WX4467&WX4944);
assign WX5027 = (WX4479&WX5028);
assign II15622 = ((~_2191_))|((~II15620));
assign WX1452 = ((~WX1443));
assign WX10329 = (WX10308&WX10314);
assign II23467 = ((~WX7075))|((~WX7010));
assign WX6523 = (WX7484&WX6524);
assign WX2410 = ((~WX2409));
assign WX2854 = (WX3710&WX2855);
assign WX9891 = (WX9828&RESET);
assign II23337 = ((~WX7065))|((~WX6990));
assign II10875 = ((~II10865))|((~II10873));
assign WX464 = (DATA_9_1&WX465);
assign II15719 = ((~WX4520))|((~II15718));
assign WX728 = (WX665&RESET);
assign II14707 = ((~II14683))|((~II14699));
assign WX3586 = ((~TM1));
assign II26785 = ((~II26760))|((~II26784));
assign II14211 = ((~II14187))|((~II14203));
assign WX11254 = ((~II34361))|((~II34362));
assign II34602 = ((~WX11153))|((~II34601));
assign WX2121 = (WX2058&RESET);
assign WX9257 = (WX9255)|(WX9254);
assign WX9086 = (WX9097&WX10054);
assign WX4176 = ((~WX4883));
assign WX6338 = ((~WX6337));
assign II27096 = ((~WX8339))|((~II27095));
assign WX7323 = (WX7260&RESET);
assign WX1095 = ((~WX1094));
assign II34873 = ((~WX11107))|((~II34872));
assign II30517 = ((~II30527))|((~II30528));
assign II30092 = ((~WX9764))|((~II30084));
assign WX7544 = ((~WX7470));
assign WX8960 = ((~II27447))|((~II27448));
assign WX7996 = (WX7994)|(WX7993);
assign WX2407 = ((~WX2298));
assign II2575 = ((~II2585))|((~II2586));
assign II26063 = ((~II26065))|((~II26066));
assign II30719 = ((~II30721))|((~II30722));
assign WX5721 = ((~WX6139));
assign II18069 = ((~II18071))|((~II18072));
assign WX9885 = (WX9822&RESET);
assign WX1928 = ((~WX2176));
assign WX9333 = (WX10182&WX9334);
assign II27664 = ((~WX8387))|((~II27663));
assign WX1900 = ((~WX1868));
assign WX10777 = ((~WX11348));
assign WX4478 = ((~WX4446));
assign II35539 = ((~II35541))|((~II35542));
assign WX8213 = (WX8224&WX8761);
assign WX7714 = ((~II23645))|((~II23646));
assign II22951 = ((~WX7234))|((~II22950));
assign WX6231 = (WX6229)|(WX6228);
assign WX1981 = (WX1649&RESET);
assign II2176 = ((~WX657))|((~II2174));
assign WX3616 = ((~WX3591));
assign WX10151 = ((~WX10056));
assign II26461 = ((~II26451))|((~II26459));
assign WX1106 = (WX594&WX1107);
assign II2021 = ((~WX647))|((~II2019));
assign II3591 = ((~WX622))|((~_2097_));
assign II22942 = ((~II22944))|((~II22945));
assign II19597 = ((~WX5792))|((~_2227_));
assign II10771 = ((~II10781))|((~II10782));
assign WX8018 = (WX8024&WX8019);
assign WX8833 = ((~WX8832));
assign WX5844 = (WX5416&RESET);
assign WX9263 = (WX10147&WX9264);
assign WX6582 = ((~WX6573));
assign II19397 = ((~WX5777))|((~WX5707));
assign II22051 = ((~WX7176))|((~II22043));
assign II14699 = ((~II14701))|((~II14702));
assign WX6227 = ((~II19164))|((~II19165));
assign WX5974 = (WX5911&RESET);
assign WX806 = (WX743&RESET);
assign WX782 = (WX719&RESET);
assign WX1764 = ((~WX2296));
assign WX11492 = (WX10944&WX11493);
assign II14048 = ((~II14050))|((~II14051));
assign WX9981 = ((~II30976))|((~II30977));
assign WX5006 = (WX4476&WX5007);
assign II14041 = ((~WX4590))|((~II14033));
assign WX7395 = ((~II22966))|((~II22967));
assign II14662 = ((~WX4630))|((~II14661));
assign WX10650 = (DATA_0_12&WX10651);
assign WX2336 = (WX1878&WX2337);
assign II23631 = ((~WX7089))|((~II23630));
assign WX3582 = ((~TM0));
assign WX2846 = (WX2852&WX2847);
assign II27621 = ((~WX8380))|((~_2289_));
assign WX7690 = (WX7076&WX7691);
assign WX6828 = ((~WX7469));
assign WX10937 = ((~WX10905));
assign WX7903 = ((~WX7894));
assign WX7035 = ((~WX7410));
assign WX2502 = ((~II7435))|((~II7436));
assign WX5964 = (WX5901&RESET);
assign II2637 = ((~II2647))|((~II2648));
assign WX7070 = ((~WX7038));
assign II2901 = ((~II2903))|((~II2904));
assign II18257 = ((~WX6173))|((~II18256));
assign WX4891 = ((~WX4890));
assign II10679 = ((~II10681))|((~II10682));
assign II30892 = ((~WX10053))|((~II30891));
assign WX8863 = (WX8862&WX8763);
assign WX1430 = (_2133_&WX2297);
assign II26164 = ((~II26140))|((~II26156));
assign WX2737 = (_2164_&WX3590);
assign WX7227 = (WX7164&RESET);
assign WX862 = (WX799&RESET);
assign WX1921 = ((~WX2162));
assign WX10789 = (_2335_&WX11348);
assign WX4878 = ((~TM1));
assign WX6623 = (WX6621)|(WX6620);
assign II34491 = ((~II34501))|((~II34502));
assign II14033 = ((~II14035))|((~II14036));
assign WX6541 = ((~WX6540));
assign WX8839 = ((~WX8838));
assign II14545 = ((~WX4686))|((~WX4750));
assign II2048 = ((~II2058))|((~II2059));
assign II14646 = ((~II14621))|((~II14645));
assign WX4058 = (_2194_&WX4883);
assign WX428 = (WX434&WX429);
assign II2051 = ((~WX1001))|((~II2050));
assign WX10784 = ((~WX10783));
assign II34670 = ((~II34646))|((~II34662));
assign II14420 = ((~II14422))|((~II14423));
assign II2352 = ((~II2327))|((~II2351));
assign WX4270 = ((~WX4883));
assign II22726 = ((~WX7467))|((~WX7156));
assign II19360 = ((~WX5701))|((~II19358));
assign WX3169 = ((~WX3137));
assign WX117 = ((~WX108));
assign WX9968 = ((~II30573))|((~II30574));
assign II26554 = ((~II26544))|((~II26552));
assign II23702 = ((~_2243_))|((~II23700));
assign II26049 = ((~WX8759))|((~WX8405));
assign II6436 = ((~II6426))|((~II6434));
assign WX4607 = (WX4544&RESET);
assign WX8258 = (WX8261&RESET);
assign WX3545 = ((~WX3544));
assign WX3004 = (WX5080&WX3005);
assign II2359 = ((~II2361))|((~II2362));
assign WX8432 = (WX8016&RESET);
assign WX7271 = (WX7208&RESET);
assign WX484 = (WX487&RESET);
assign WX4513 = ((~WX4760));
assign WX1408 = ((~WX2297));
assign WX5092 = (WX5090)|(WX5089);
assign II22471 = ((~II22461))|((~II22469));
assign WX4743 = (WX4680&RESET);
assign WX6905 = ((~WX6904));
assign WX8845 = (WX8843)|(WX8842);
assign WX11303 = ((~WX11302));
assign WX3763 = ((~WX3591));
assign II10230 = ((~WX3373))|((~WX3437));
assign WX2233 = ((~WX2213));
assign WX9533 = ((~WX9532));
assign WX7962 = (WX7968&WX7963);
assign WX10434 = ((~WX10433));
assign II34812 = ((~II34802))|((~II34810));
assign II14848 = ((~WX4642))|((~II14847));
assign II6053 = ((~II6063))|((~II6064));
assign WX6289 = ((~WX6288));
assign II6829 = ((~II6831))|((~II6832));
assign II34695 = ((~WX11159))|((~II34694));
assign II34417 = ((~WX11205))|((~II34415));
assign II14552 = ((~II14528))|((~II14544));
assign WX10571 = ((~WX11348));
assign II2616 = ((~WX749))|((~II2615));
assign II34609 = ((~II34584))|((~II34608));
assign II2579 = ((~WX683))|((~II2577));
assign WX9431 = (WX10231&WX9432);
assign WX1137 = ((~WX1136));
assign II27635 = ((~WX8382))|((~_2287_));
assign II2074 = ((~II2064))|((~II2072));
assign WX2290 = ((~TM0));
assign II30156 = ((~II30146))|((~II30154));
assign WX585 = ((~WX553));
assign WX4601 = (WX4538&RESET);
assign WX10657 = ((~WX10648));
assign II22091 = ((~WX7242))|((~II22090));
assign II11645 = ((~_2154_))|((~II11643));
assign WX5908 = (WX5845&RESET);
assign II26468 = ((~WX8559))|((~II26467));
assign II6553 = ((~WX1974))|((~II6551));
assign WX11329 = ((~WX11328));
assign WX1897 = ((~WX1865));
assign WX4777 = (WX4714&RESET);
assign WX6815 = (WX6813)|(WX6812);
assign WX1345 = (WX1343)|(WX1342);
assign WX6737 = ((~WX6736));
assign WX8075 = ((~WX8761));
assign II35612 = ((~_2356_))|((~II35610));
assign WX5334 = (WX5340&WX5335);
assign WX5501 = (WX5512&WX6175);
assign II7383 = ((~WX1898))|((~II7382));
assign II2269 = ((~WX663))|((~II2267));
assign II34119 = ((~II34129))|((~II34130));
assign II22454 = ((~WX7202))|((~II22446));
assign II10943 = ((~WX3419))|((~WX3483));
assign WX1887 = ((~WX1855));
assign II15614 = ((~WX4502))|((~II15613));
assign WX8199 = (WX8210&WX8761);
assign WX7863 = (WX7874&WX8761);
assign II30691 = ((~WX9930))|((~II30689));
assign WX10805 = ((~WX11348));
assign II14966 = ((~WX4586))|((~II14964));
assign WX5470 = (WX5468)|(WX5467);
assign II26776 = ((~II26778))|((~II26779));
assign WX1340 = ((~WX1331));
assign II6529 = ((~II6519))|((~II6527));
assign WX2117 = (WX2054&RESET);
assign WX6128 = ((~WX6100));
assign WX2622 = (WX2628&WX2623);
assign II2260 = ((~II2250))|((~II2258));
assign WX4461 = ((~WX4429));
assign WX4112 = ((~WX4882));
assign WX10437 = ((~WX11347));
assign II22595 = ((~II22585))|((~II22593));
assign II22214 = ((~WX7250))|((~WX7314));
assign II30673 = ((~II30675))|((~II30676));
assign II19492 = ((~_2236_))|((~II19490));
assign WX2688 = (WX2686)|(WX2685);
assign II19086 = ((~WX5753))|((~II19085));
assign WX7159 = (WX6863&RESET);
assign WX1955 = (WX1467&RESET);
assign WX3041 = (WX3052&WX3589);
assign II26869 = ((~II26871))|((~II26872));
assign WX1707 = (WX1713&WX1708);
assign II26406 = ((~WX8555))|((~II26405));
assign II23389 = ((~WX7069))|((~WX6998));
assign WX7930 = (WX7928)|(WX7927);
assign WX11474 = ((~WX11473));
assign II10208 = ((~II10198))|((~II10206));
assign II6311 = ((~WX2022))|((~II6310));
assign WX7111 = (WX6527&RESET);
assign WX1425 = ((~WX1424));
assign WX7301 = (WX7238&RESET);
assign II35458 = ((~WX10885))|((~II35456));
assign WX10882 = (WX10885&RESET);
assign II14329 = ((~WX4672))|((~II14328));
assign II30458 = ((~WX10052))|((~II30457));
assign WX474 = (WX2522&WX475);
assign II34929 = ((~WX11047))|((~II34927));
assign II30986 = ((~WX9758))|((~II30984));
assign WX4731 = (WX4668&RESET);
assign WX3569 = ((~WX3568));
assign WX6175 = ((~WX6171));
assign WX5577 = ((~WX6176));
assign II34867 = ((~WX11043))|((~II34865));
assign II30836 = ((~WX9812))|((~II30828));
assign WX6531 = (WX6529)|(WX6528);
assign WX4133 = (WX4996&WX4134);
assign II35404 = ((~WX10948))|((~WX10877));
assign WX6346 = ((~II19385))|((~II19386));
assign WX502 = (WX505&RESET);
assign WX1032 = ((~WX1031));
assign II22988 = ((~II22990))|((~II22991));
assign II30735 = ((~II30737))|((~II30738));
assign II14925 = ((~II14900))|((~II14924));
assign WX10274 = ((~II31491))|((~II31492));
assign WX10172 = ((~WX10056));
assign WX2972 = (WX2978&WX2973);
assign II10813 = ((~II10803))|((~II10811));
assign WX1161 = (WX1160&WX1005);
assign WX5912 = (WX5849&RESET);
assign WX5866 = (WX5570&RESET);
assign II22883 = ((~WX7166))|((~II22881));
assign WX710 = (WX647&RESET);
assign II26816 = ((~II26791))|((~II26815));
assign WX1484 = ((~WX2296));
assign II3457 = ((~WX547))|((~II3455));
assign WX9427 = (WX11524&WX9428);
assign WX9015 = ((~II27706))|((~II27707));
assign WX10641 = ((~WX11348));
assign WX3038 = (WX3036)|(WX3035);
assign II22502 = ((~II22492))|((~II22500));
assign II14515 = ((~WX4684))|((~II14514));
assign II27726 = ((~WX8398))|((~_2271_));
assign WX6716 = ((~WX7469));
assign WX1443 = (WX1441)|(WX1440);
assign WX4858 = ((~WX4857));
assign II30273 = ((~WX9712))|((~II30271));
assign II23502 = ((~_2252_))|((~II23494));
assign II6496 = ((~WX2034))|((~II6488));
assign WX9356 = (_2313_&WX10055);
assign WX599 = ((~WX567));
assign II15444 = ((~WX4488))|((~WX4422));
assign WX8203 = (_2271_&WX8762);
assign WX748 = (WX685&RESET);
assign WX8030 = ((~WX8029));
assign II26196 = ((~II26171))|((~II26195));
assign II22818 = ((~II22820))|((~II22821));
assign II10394 = ((~II10384))|((~II10392));
assign II35745 = ((~_2334_))|((~II35743));
assign WX8120 = (WX10224&WX8121);
assign WX3015 = ((~WX3589));
assign WX7851 = ((~WX8761));
assign WX4148 = ((~WX4883));
assign WX11245 = ((~II34082))|((~II34083));
assign II30471 = ((~II30473))|((~II30474));
assign WX10505 = (WX10516&WX11347);
assign WX10700 = ((~WX10699));
assign WX4053 = ((~WX4052));
assign WX7483 = ((~WX7482));
assign II18132 = ((~WX6173))|((~WX5825));
assign II6653 = ((~II6643))|((~II6651));
assign II23496 = ((~WX7092))|((~II23495));
assign WX4483 = ((~WX4451));
assign WX6036 = (WX5973&RESET);
assign WX6938 = (_2237_&WX7469);
assign II23694 = ((~WX7100))|((~II23693));
assign WX2944 = (WX2950&WX2945);
assign WX6292 = (WX5768&WX6293);
assign WX7102 = ((~WX7352));
assign WX2139 = (WX2076&RESET);
assign WX2933 = (_2150_&WX3590);
assign WX6172 = ((~TM1));
assign WX9234 = (WX9556&WX10055);
assign WX9136 = (WX9542&WX10055);
assign II14916 = ((~II14918))|((~II14919));
assign II6149 = ((~WX2294))|((~II6148));
assign II34181 = ((~II34191))|((~II34192));
assign WX10602 = ((~WX10601));
assign II14435 = ((~II14445))|((~II14446));
assign II11452 = ((~WX3196))|((~WX3131));
assign WX2253 = ((~WX2223));
assign WX11585 = ((~II35604))|((~II35605));
assign WX11014 = (WX10574&RESET);
assign WX11388 = ((~WX11349));
assign WX7960 = ((~WX7959));
assign WX4309 = (WX4307)|(WX4306);
assign II35314 = ((~WX10941))|((~II35313));
assign II34058 = ((~II34060))|((~II34061));
assign II26283 = ((~WX8611))|((~II26281));
assign WX10707 = ((~WX11348));
assign II18626 = ((~II18636))|((~II18637));
assign WX3031 = (_2143_&WX3590);
assign WX6409 = ((~II19556))|((~II19557));
assign II18147 = ((~WX5953))|((~WX6017));
assign II14019 = ((~WX4652))|((~II14018));
assign II18131 = ((~II18133))|((~II18134));
assign II34306 = ((~II34308))|((~II34309));
assign II18674 = ((~WX5987))|((~WX6051));
assign WX1066 = (WX1064)|(WX1063);
assign WX5303 = ((~WX5294));
assign WX5636 = (WX6394&WX5637);
assign WX549 = ((~WX967));
assign II2894 = ((~WX767))|((~II2886));
assign WX9238 = ((~WX9229));
assign II34401 = ((~WX11345))|((~II34400));
assign II22934 = ((~II22910))|((~II22926));
assign II7213 = ((~WX1885))|((~WX1802));
assign WX4701 = (WX4638&RESET);
assign II34578 = ((~II34553))|((~II34577));
assign II30169 = ((~II30145))|((~II30161));
assign WX6851 = (WX6857&WX6852);
assign WX8072 = ((~WX8071));
assign WX8309 = ((~WX8729));
assign II6429 = ((~WX1966))|((~II6427));
assign WX8638 = (WX8575&RESET);
assign WX1224 = (WX1223&WX1005);
assign II26771 = ((~II26761))|((~II26769));
assign WX10495 = (_2356_&WX11348);
assign II31113 = ((~WX9633))|((~WX9540));
assign WX2595 = (WX2540&WX2556);
assign II35106 = ((~WX10925))|((~II35105));
assign WX2494 = ((~WX2493));
assign II6070 = ((~WX2070))|((~WX2134));
assign II30450 = ((~II30440))|((~II30448));
assign II10719 = ((~WX3341))|((~II10718));
assign WX256 = (WX254)|(WX253);
assign II30907 = ((~WX9880))|((~II30906));
assign WX444 = (WX442)|(WX441);
assign WX1270 = (WX1260&WX1263);
assign II35701 = ((~WX10978))|((~_2341_));
assign II35631 = ((~WX10966))|((~_2353_));
assign WX2328 = (WX2327&WX2298);
assign WX7678 = (WX7676)|(WX7675);
assign WX10569 = (WX10855&WX11348);
assign II18878 = ((~WX5873))|((~II18876));
assign II14111 = ((~WX4658))|((~WX4722));
assign WX4201 = (WX4199)|(WX4198);
assign WX7467 = ((~WX7463));
assign WX10543 = ((~WX11348));
assign II10245 = ((~II10247))|((~II10248));
assign WX9426 = (_2308_&WX10055);
assign WX6204 = ((~WX6203));
assign II14141 = ((~II14143))|((~II14144));
assign WX8107 = ((~WX8762));
assign WX10196 = ((~WX10195));
assign II23090 = ((~WX7046))|((~WX6952));
assign II26979 = ((~WX8760))|((~WX8465));
assign II7492 = ((~_2140_))|((~II7490));
assign II34027 = ((~II34029))|((~II34030));
assign II2391 = ((~WX1001))|((~WX671));
assign WX8150 = (WX8148)|(WX8147);
assign II30130 = ((~II30132))|((~II30133));
assign WX6114 = ((~WX6093));
assign WX2373 = (WX2371)|(WX2370);
assign WX3306 = (WX3243&RESET);
assign WX7628 = ((~WX7470));
assign WX4135 = (WX4133)|(WX4132);
assign II30061 = ((~WX9762))|((~II30053));
assign II18884 = ((~WX5937))|((~II18883));
assign WX921 = ((~II2662))|((~II2663));
assign WX3724 = ((~WX3723));
assign WX7908 = (WX7906)|(WX7905);
assign II22842 = ((~II22817))|((~II22841));
assign II7058 = ((~WX1873))|((~II7057));
assign WX9142 = (WX9153&WX10054);
assign II2452 = ((~II2454))|((~II2455));
assign II14849 = ((~II14839))|((~II14847));
assign WX8932 = ((~II27395))|((~II27396));
assign WX9680 = ((~WX9922));
assign II34252 = ((~WX11067))|((~II34244));
assign WX5771 = ((~WX5739));
assign WX2951 = (WX3117&WX3590);
assign WX11230 = (WX11167&RESET);
assign II7266 = ((~WX1889))|((~II7265));
assign WX11541 = (WX10951&WX11542);
assign WX1121 = ((~WX1005));
assign WX9012 = ((~II27685))|((~II27686));
assign WX8962 = (WX8366&WX8963);
assign WX8937 = ((~WX8936));
assign WX2175 = (WX2112&RESET);
assign II11636 = ((~WX3214))|((~_2155_));
assign WX8548 = (WX8485&RESET);
assign WX2824 = (WX2822)|(WX2821);
assign II6666 = ((~II6642))|((~II6658));
assign II14104 = ((~WX4594))|((~II14103));
assign II2956 = ((~WX771))|((~II2948));
assign WX2917 = ((~WX3589));
assign WX7490 = ((~WX7489));
assign WX4373 = (WX4376&RESET);
assign WX9054 = (WX8989&WX9021);
assign II15706 = ((~_2177_))|((~II15704));
assign II1995 = ((~WX709))|((~II1987));
assign II26903 = ((~WX8651))|((~II26901));
assign II10727 = ((~WX3405))|((~II10726));
assign WX7605 = (WX7604&WX7470);
assign WX3476 = (WX3413&RESET);
assign II34557 = ((~WX11023))|((~II34555));
assign II2127 = ((~WX781))|((~WX845));
assign WX6817 = (WX7631&WX6818);
assign WX2181 = (WX2118&RESET);
assign WX2814 = (WX2812)|(WX2811);
assign WX9666 = ((~WX9894));
assign II15171 = ((~WX4467))|((~WX4380));
assign WX468 = ((~WX467));
assign WX4063 = (WX4961&WX4064);
assign II2625 = ((~WX877))|((~II2623));
assign II6675 = ((~WX2295))|((~WX1982));
assign WX563 = ((~WX995));
assign II7447 = ((~WX1903))|((~WX1838));
assign WX2648 = ((~WX2647));
assign II22292 = ((~WX7466))|((~WX7128));
assign II10539 = ((~II10541))|((~II10542));
assign WX6894 = ((~WX7468));
assign II26097 = ((~WX8599))|((~II26095));
assign II22849 = ((~II22851))|((~II22852));
assign WX4351 = (WX4349)|(WX4348);
assign WX10814 = (WX10820&WX10815);
assign II3222 = ((~WX593))|((~II3221));
assign WX10064 = ((~II31101))|((~II31102));
assign WX6327 = (WX5773&WX6328);
assign II18557 = ((~II18533))|((~II18549));
assign WX4174 = (WX4400&WX4883);
assign II22015 = ((~WX7110))|((~II22013));
assign WX7824 = (WX7822)|(WX7821);
assign WX9024 = (WX9020&WX9021);
assign WX2289 = ((~TM0));
assign II26946 = ((~II26956))|((~II26957));
assign WX8352 = ((~WX8320));
assign WX3328 = (WX3265&RESET);
assign II30582 = ((~WX10053))|((~II30581));
assign WX10931 = ((~WX10899));
assign II2005 = ((~WX837))|((~II2003));
assign WX3228 = ((~WX3483));
assign WX986 = ((~WX911));
assign WX8730 = ((~WX8662));
assign WX3656 = (WX3655&WX3591);
assign II31537 = ((~_2332_))|((~II31535));
assign II10945 = ((~WX3483))|((~II10943));
assign WX1545 = (WX1543)|(WX1542);
assign WX2962 = (WX5059&WX2963);
assign WX7021 = ((~WX7446));
assign WX8722 = ((~WX8658));
assign WX4212 = (_2183_&WX4883);
assign II30240 = ((~WX10052))|((~WX9710));
assign WX6608 = ((~WX7469));
assign WX10276 = (WX9662&WX10277);
assign WX10170 = (WX10169&WX10056);
assign WX3177 = ((~WX3145));
assign WX6562 = ((~WX7469));
assign WX2207 = ((~II6450))|((~II6451));
assign WX3884 = (WX3835&WX3849);
assign II34044 = ((~WX11117))|((~II34043));
assign II27291 = ((~WX8354))|((~II27290));
assign II26538 = ((~II26528))|((~II26536));
assign WX11569 = (WX10955&WX11570);
assign II27649 = ((~WX8384))|((~_2285_));
assign WX6906 = (WX6917&WX7468);
assign WX6653 = ((~WX6652));
assign II6380 = ((~WX2090))|((~WX2154));
assign WX9943 = (WX9880&RESET);
assign WX3422 = (WX3359&RESET);
assign WX601 = ((~WX569));
assign WX9907 = (WX9844&RESET);
assign WX11374 = ((~WX11349));
assign II10138 = ((~WX3367))|((~II10137));
assign II2599 = ((~II2575))|((~II2591));
assign WX7325 = (WX7262&RESET);
assign II3563 = ((~WX618))|((~_2101_));
assign WX102 = (WX100)|(WX99);
assign WX5652 = (WX5650)|(WX5649);
assign II6534 = ((~II6536))|((~II6537));
assign II10084 = ((~II10074))|((~II10082));
assign WX3980 = ((~WX4883));
assign II2777 = ((~II2779))|((~II2780));
assign WX7345 = (WX7282&RESET);
assign WX4585 = (WX4361&RESET);
assign II27566 = ((~WX8372))|((~II27565));
assign WX6703 = (WX6701)|(WX6700);
assign WX6106 = ((~WX6089));
assign WX8969 = (WX8367&WX8970);
assign II27677 = ((~WX8389))|((~_2280_));
assign WX8359 = ((~WX8327));
assign II18852 = ((~WX5935))|((~II18844));
assign WX10555 = (WX10853&WX11348);
assign WX7273 = (WX7210&RESET);
assign WX2797 = (WX3095&WX3590);
assign WX7986 = (WX7984)|(WX7983);
assign WX8210 = (WX8208)|(WX8207);
assign WX7389 = ((~II22780))|((~II22781));
assign WX6701 = (WX8868&WX6702);
assign WX2990 = (WX5073&WX2991);
assign WX8270 = (WX8273&RESET);
assign WX11405 = ((~WX11404));
assign II34843 = ((~II34833))|((~II34841));
assign II11488 = ((~_2156_))|((~II11487));
assign II26366 = ((~WX8489))|((~II26358));
assign WX3036 = (WX3801&WX3037);
assign II14732 = ((~WX4698))|((~II14731));
assign WX6718 = (WX6980&WX7469);
assign II30644 = ((~WX10053))|((~II30643));
assign II22325 = ((~WX7130))|((~II22323));
assign II18691 = ((~WX6174))|((~II18690));
assign WX966 = ((~WX901));
assign WX7064 = ((~WX7032));
assign WX8219 = ((~WX8762));
assign WX4799 = ((~II14646))|((~II14647));
assign II27409 = ((~WX8293))|((~II27407));
assign II14802 = ((~II14792))|((~II14800));
assign WX4001 = (WX3999)|(WX3998);
assign WX5815 = ((~WX6071));
assign II30574 = ((~II30564))|((~II30572));
assign WX5141 = ((~II15726))|((~II15727));
assign II10526 = ((~WX3588))|((~II10525));
assign II18255 = ((~II18257))|((~II18258));
assign WX7546 = ((~WX7545));
assign WX2712 = (WX2710)|(WX2709);
assign WX2929 = (WX2940&WX3589);
assign WX3555 = ((~WX3554));
assign II15508 = ((~_2183_))|((~II15507));
assign WX981 = ((~WX980));
assign WX5463 = (_2218_&WX6176);
assign II30884 = ((~II30874))|((~II30882));
assign WX2718 = ((~WX2717));
assign WX11595 = ((~II35674))|((~II35675));
assign WX10722 = (WX10720)|(WX10719);
assign WX414 = (WX420&WX415);
assign II35688 = ((~WX10975))|((~II35687));
assign II11538 = ((~WX3199))|((~_2170_));
assign WX7505 = ((~WX7504));
assign WX8691 = ((~WX8690));
assign WX6695 = ((~WX6694));
assign WX11267 = ((~II34764))|((~II34765));
assign II34030 = ((~WX10989))|((~II34028));
assign II26708 = ((~WX8511))|((~II26707));
assign WX3834 = ((~II11623))|((~II11624));
assign WX11583 = ((~II35590))|((~II35591));
assign II2810 = ((~WX825))|((~II2809));
assign WX7596 = ((~WX7595));
assign WX6332 = ((~II19359))|((~II19360));
assign WX8526 = (WX8463&RESET);
assign II2243 = ((~WX725))|((~II2235));
assign WX6711 = (WX6717&WX6712);
assign WX8347 = ((~WX8315));
assign WX2266 = ((~WX2265));
assign WX11194 = (WX11131&RESET);
assign WX2752 = (WX4954&WX2753);
assign II10324 = ((~WX3379))|((~II10323));
assign WX5601 = ((~WX6175));
assign WX9145 = (WX9143)|(WX9142);
assign WX3067 = ((~WX3058));
assign II19384 = ((~WX5776))|((~WX5705));
assign WX7624 = ((~WX7623));
assign WX6203 = (WX6201)|(WX6200);
assign II26423 = ((~WX8429))|((~II26421));
assign II35006 = ((~WX11243))|((~II35004));
assign WX174 = ((~WX173));
assign WX5187 = (WX5123&WX5142);
assign II6801 = ((~WX1990))|((~II6799));
assign WX2258 = ((~WX2257));
assign II30936 = ((~II30938))|((~II30939));
assign WX1140 = (WX1139&WX1005);
assign II6046 = ((~II6022))|((~II6038));
assign WX254 = (DATA_9_16&WX255);
assign WX5623 = ((~WX6176));
assign WX1335 = (WX1333)|(WX1332);
assign II27698 = ((~WX8393))|((~_2276_));
assign II11532 = ((~WX3198))|((~II11531));
assign WX2542 = ((~II7625))|((~II7626));
assign II19626 = ((~WX5796))|((~II19625));
assign II14594 = ((~WX4562))|((~II14592));
assign WX2197 = ((~II6140))|((~II6141));
assign II18512 = ((~WX5913))|((~II18511));
assign WX9927 = (WX9864&RESET);
assign II30559 = ((~II30549))|((~II30557));
assign II10392 = ((~II10368))|((~II10384));
assign WX5704 = (WX5707&RESET);
assign II18914 = ((~WX5939))|((~II18906));
assign WX9600 = ((~WX10018));
assign WX566 = ((~WX937));
assign WX6596 = ((~WX6587));
assign II34677 = ((~II34687))|((~II34688));
assign II22138 = ((~WX7466))|((~II22137));
assign WX915 = ((~II2476))|((~II2477));
assign WX4275 = (WX4273)|(WX4272);
assign WX972 = ((~WX904));
assign II15580 = ((~_2197_))|((~II15578));
assign WX4985 = (WX4473&WX4986);
assign II30899 = ((~WX9816))|((~II30898));
assign II7123 = ((~WX1878))|((~II7122));
assign WX4488 = ((~WX4456));
assign WX10896 = ((~WX11317));
assign II14490 = ((~II14466))|((~II14482));
assign WX6163 = ((~WX6162));
assign WX2251 = ((~WX2222));
assign II30528 = ((~II30518))|((~II30526));
assign II34383 = ((~II34385))|((~II34386));
assign WX592 = ((~WX560));
assign WX9360 = (WX9574&WX10055);
assign WX4936 = (WX4466&WX4937);
assign II34972 = ((~II34974))|((~II34975));
assign WX10523 = (_2354_&WX11348);
assign WX4733 = (WX4670&RESET);
assign WX6604 = ((~WX7469));
assign II18657 = ((~II18667))|((~II18668));
assign II2796 = ((~WX697))|((~II2794));
assign WX6366 = ((~WX6365));
assign WX7511 = ((~WX7510));
assign II26459 = ((~WX8495))|((~II26451));
assign II2809 = ((~WX825))|((~WX889));
assign WX9692 = ((~WX9946));
assign WX828 = (WX765&RESET);
assign WX1178 = (WX1176)|(WX1175);
assign WX7579 = ((~WX7470));
assign WX5785 = ((~WX6011));
assign WX5529 = (WX5540&WX6175);
assign II11559 = ((~WX3202))|((~_2167_));
assign WX6425 = ((~II19668))|((~II19669));
assign WX4441 = ((~WX4872));
assign WX7636 = (WX7634)|(WX7633);
assign WX8338 = ((~WX8306));
assign II27586 = ((~WX8375))|((~_2294_));
assign WX1382 = ((~WX1373));
assign WX2637 = ((~WX3589));
assign WX10903 = ((~WX11331));
assign WX9451 = (WX9457&WX9452);
assign WX2436 = (WX2434)|(WX2433);
assign WX7489 = (WX7487)|(WX7486);
assign WX3798 = ((~WX3591));
assign WX7105 = ((~WX7358));
assign II26227 = ((~II26202))|((~II26226));
assign WX8026 = (WX8882&WX8027);
assign II26034 = ((~WX8531))|((~II26033));
assign II19661 = ((~WX5802))|((~II19660));
assign II2531 = ((~WX807))|((~II2530));
assign WX3057 = ((~WX3589));
assign II6544 = ((~II6534))|((~II6542));
assign WX2360 = ((~WX2359));
assign II10889 = ((~II10864))|((~II10888));
assign II23143 = ((~WX7050))|((~II23142));
assign WX3088 = (WX3091&RESET);
assign II18860 = ((~WX5999))|((~WX6063));
assign WX874 = (WX811&RESET);
assign II30921 = ((~II30923))|((~II30924));
assign II26932 = ((~WX8589))|((~WX8653));
assign II26181 = ((~WX8477))|((~II26180));
assign II22517 = ((~WX7206))|((~II22516));
assign WX10463 = (WX10474&WX11347);
assign WX7554 = ((~WX7553));
assign WX696 = (WX412&RESET);
assign WX5308 = (WX5306)|(WX5305);
assign II34168 = ((~WX11125))|((~II34167));
assign WX11104 = (WX11041&RESET);
assign WX6193 = (WX6192&WX6177);
assign WX331 = ((~WX1003));
assign II2275 = ((~WX727))|((~II2274));
assign WX8365 = ((~WX8333));
assign WX393 = (WX535&WX1004);
assign II31283 = ((~WX9646))|((~II31282));
assign WX8129 = (WX8140&WX8761);
assign WX9030 = (WX8991&WX9021);
assign WX4990 = ((~II15263))|((~II15264));
assign WX10046 = ((~WX10045));
assign WX11336 = ((~WX11258));
assign WX6062 = (WX5999&RESET);
assign WX9258 = (_2320_&WX10055);
assign WX7886 = (WX8812&WX7887);
assign WX7500 = (WX7499&WX7470);
assign II14763 = ((~WX4700))|((~II14762));
assign II35261 = ((~WX10937))|((~WX10855));
assign WX450 = (DATA_9_2&WX451);
assign WX4282 = (_2178_&WX4883);
assign WX8978 = (WX8976)|(WX8975);
assign II15725 = ((~WX4521))|((~_2173_));
assign II34541 = ((~WX11213))|((~II34539));
assign WX8795 = ((~WX8763));
assign WX1044 = ((~WX1005));
assign II26616 = ((~II26606))|((~II26614));
assign II30566 = ((~WX9858))|((~II30565));
assign II34740 = ((~II34742))|((~II34743));
assign WX7482 = (WX7480)|(WX7479);
assign II11205 = ((~WX3177))|((~WX3093));
assign WX3955 = ((~WX3954));
assign WX6018 = (WX5955&RESET);
assign WX3132 = (WX3069&RESET);
assign II2221 = ((~WX787))|((~II2220));
assign II30055 = ((~WX10052))|((~II30054));
assign WX840 = (WX777&RESET);
assign WX3124 = (WX3127&RESET);
assign II2453 = ((~WX1001))|((~WX675));
assign WX9414 = ((~WX10055));
assign WX3510 = ((~II10765))|((~II10766));
assign II30178 = ((~WX10052))|((~WX9706));
assign II26701 = ((~WX8760))|((~II26700));
assign II6363 = ((~II6373))|((~II6374));
assign II7504 = ((~II7506))|((~II7507));
assign II35496 = ((~WX10955))|((~II35495));
assign WX6665 = (WX6663)|(WX6662);
assign WX7465 = ((~TM1));
assign II26670 = ((~WX8760))|((~II26669));
assign WX6697 = (WX6703&WX6698);
assign WX544 = (WX547&RESET);
assign WX8314 = ((~WX8739));
assign WX5521 = ((~WX6176));
assign WX11216 = (WX11153&RESET);
assign WX8300 = (WX8303&RESET);
assign WX1564 = ((~WX1555));
assign II3648 = ((~WX631))|((~II3647));
assign WX10698 = (WX10696)|(WX10695);
assign II18831 = ((~WX6061))|((~II18829));
assign WX1362 = ((~WX2297));
assign II19543 = ((~_2235_))|((~II19541));
assign II10169 = ((~WX3369))|((~II10168));
assign WX7422 = ((~WX7421));
assign WX4268 = (_2179_&WX4883);
assign II30619 = ((~WX9798))|((~II30611));
assign WX3500 = ((~II10455))|((~II10456));
assign II3522 = ((~WX612))|((~II3521));
assign WX8993 = ((~II27552))|((~II27553));
assign II18124 = ((~II18099))|((~II18123));
assign WX9805 = (WX9742&RESET);
assign WX10763 = ((~WX11348));
assign II22524 = ((~WX7270))|((~WX7334));
assign II11387 = ((~WX3191))|((~WX3121));
assign WX3213 = ((~WX3453));
assign WX5010 = ((~WX5009));
assign WX1779 = (WX1782&RESET);
assign WX11559 = ((~WX11558));
assign II2950 = ((~WX1002))|((~II2949));
assign WX11257 = ((~II34454))|((~II34455));
assign WX1713 = (WX1711)|(WX1710);
assign WX6305 = (WX6304&WX6177);
assign II19571 = ((~_2231_))|((~II19569));
assign WX8328 = ((~WX8703));
assign WX7632 = ((~II23377))|((~II23378));
assign WX4964 = (WX4470&WX4965);
assign WX11358 = (WX11357&WX11349);
assign WX2697 = ((~WX3590));
assign WX7125 = (WX6625&RESET);
assign WX372 = (WX378&WX373);
assign WX2900 = ((~WX2899));
assign WX8901 = (WX8899)|(WX8898);
assign II30488 = ((~WX10052))|((~WX9726));
assign II26667 = ((~II26677))|((~II26678));
assign II11518 = ((~_2144_))|((~II11517));
assign WX9097 = (WX9095)|(WX9094);
assign WX1084 = (WX1083&WX1005);
assign WX1458 = (_2131_&WX2297);
assign WX1397 = ((~WX1396));
assign WX2913 = ((~WX2904));
assign II19731 = ((~WX5814))|((~II19730));
assign II11494 = ((~II11496))|((~II11497));
assign WX9640 = ((~WX9608));
assign II2684 = ((~II2686))|((~II2687));
assign WX10996 = (WX10448&RESET);
assign WX8861 = ((~WX8860));
assign WX7611 = ((~II23338))|((~II23339));
assign II7306 = ((~WX1816))|((~II7304));
assign WX11662 = (WX11583&WX11607);
assign II6449 = ((~II6425))|((~II6441));
assign WX5564 = (WX5562)|(WX5561);
assign WX2451 = ((~WX2450));
assign II22082 = ((~WX7178))|((~II22074));
assign II11375 = ((~WX3190))|((~II11374));
assign WX5071 = (WX5069)|(WX5068);
assign WX4785 = ((~II14212))|((~II14213));
assign WX11320 = ((~WX11250));
assign II30148 = ((~WX10052))|((~II30147));
assign WX8185 = (WX8196&WX8761);
assign WX11573 = ((~WX11572));
assign WX2369 = ((~II7188))|((~II7189));
assign II34393 = ((~II34383))|((~II34391));
assign II22774 = ((~WX7350))|((~II22772));
assign II2964 = ((~WX835))|((~WX899));
assign II34555 = ((~WX11346))|((~WX11023));
assign II34454 = ((~II34429))|((~II34453));
assign II2716 = ((~WX819))|((~WX883));
assign WX2013 = (WX1950&RESET);
assign II10782 = ((~II10772))|((~II10780));
assign WX6415 = ((~II19598))|((~II19599));
assign WX4173 = (WX4171)|(WX4170);
assign II6351 = ((~WX2152))|((~II6349));
assign WX9612 = ((~WX10042));
assign WX11562 = (WX10954&WX11563);
assign WX618 = ((~WX849));
assign WX7315 = (WX7252&RESET);
assign WX2887 = (WX2898&WX3589);
assign WX5495 = (WX5697&WX6176);
assign II23666 = ((~WX7095))|((~II23665));
assign WX3270 = (WX2914&RESET);
assign WX8061 = ((~WX8761));
assign II19688 = ((~WX5807))|((~_2212_));
assign WX11509 = ((~WX11508));
assign WX11060 = (WX10997&RESET);
assign WX8985 = (WX8983)|(WX8982);
assign II34756 = ((~WX11163))|((~WX11227));
assign II14110 = ((~II14112))|((~II14113));
assign WX2123 = (WX2060&RESET);
assign II10930 = ((~WX3291))|((~II10928));
assign WX3572 = ((~WX3497));
assign WX6177 = ((~WX6168));
assign WX3992 = (WX4374&WX4883);
assign WX1028 = (WX1027&WX1005);
assign II26072 = ((~II26047))|((~II26071));
assign II19490 = ((~WX5799))|((~_2236_));
assign II14220 = ((~WX4880))|((~WX4538));
assign WX6810 = ((~WX7468));
assign WX8736 = ((~WX8665));
assign WX3872 = (WX3818&WX3849);
assign WX3986 = ((~WX4882));
assign WX9101 = (WX9107&WX9102);
assign WX6507 = (WX6505)|(WX6504);
assign WX2698 = (WX2696)|(WX2695);
assign II30249 = ((~II30239))|((~II30247));
assign II27357 = ((~WX8285))|((~II27355));
assign WX8821 = (WX8820&WX8763);
assign II30520 = ((~WX10053))|((~II30519));
assign WX5339 = ((~WX6176));
assign WX9480 = ((~WX10054));
assign II10750 = ((~WX3343))|((~II10749));
assign WX5396 = (WX5394)|(WX5393);
assign WX4804 = ((~II14801))|((~II14802));
assign WX2522 = ((~WX2521));
assign WX734 = (WX671&RESET);
assign WX2735 = ((~WX3589));
assign WX6727 = (WX6725)|(WX6724);
assign WX6837 = (WX6843&WX6838);
assign II34176 = ((~II34166))|((~II34174));
assign WX9282 = (WX9293&WX10054);
assign WX10584 = (WX11454&WX10585);
assign WX5351 = (_2226_&WX6176);
assign II30521 = ((~WX9728))|((~II30519));
assign II2165 = ((~II2141))|((~II2157));
assign II19203 = ((~WX5762))|((~II19202));
assign II6769 = ((~WX2295))|((~II6768));
assign WX4446 = ((~WX4818));
assign WX3540 = ((~WX3513));
assign WX1860 = ((~WX2232));
assign WX2583 = (WX2545&WX2556);
assign II31544 = ((~II31534))|((~II31542));
assign II1989 = ((~WX1001))|((~II1988));
assign II31492 = ((~WX9598))|((~II31490));
assign WX4715 = (WX4652&RESET);
assign WX4466 = ((~WX4434));
assign II19639 = ((~WX5798))|((~_2221_));
assign WX8590 = (WX8527&RESET);
assign WX5450 = (WX7596&WX5451);
assign II22445 = ((~II22455))|((~II22456));
assign II2284 = ((~WX855))|((~II2282));
assign WX2456 = ((~WX2298));
assign II3209 = ((~WX592))|((~II3208));
assign WX4999 = (WX4475&WX5000);
assign II15543 = ((~WX4492))|((~_2202_));
assign WX5342 = (WX6247&WX5343);
assign WX5958 = (WX5895&RESET);
assign II9999 = ((~WX3587))|((~II9998));
assign WX3186 = ((~WX3154));
assign WX6613 = (WX6619&WX6614);
assign II3182 = ((~WX590))|((~WX505));
assign WX3534 = ((~WX3510));
assign WX11311 = ((~WX11310));
assign II26857 = ((~WX8457))|((~II26855));
assign WX4661 = (WX4598&RESET);
assign WX2998 = ((~WX2997));
assign WX4972 = ((~WX4884));
assign II26792 = ((~II26794))|((~II26795));
assign II3641 = ((~WX630))|((~II3640));
assign WX7684 = ((~WX7470));
assign II30363 = ((~II30365))|((~II30366));
assign WX288 = (WX294&WX289);
assign WX11172 = (WX11109&RESET);
assign WX11281 = ((~WX11280));
assign II35540 = ((~WX10983))|((~_2364_));
assign II14577 = ((~WX4688))|((~II14576));
assign II35542 = ((~_2364_))|((~II35540));
assign WX9841 = (WX9778&RESET);
assign WX4403 = (WX4406&RESET);
assign WX6004 = (WX5941&RESET);
assign WX4962 = ((~II15211))|((~II15212));
assign II19241 = ((~WX5765))|((~WX5683));
assign WX3776 = (WX3192&WX3777);
assign WX4049 = (WX4954&WX4050);
assign II30627 = ((~WX9862))|((~WX9926));
assign II10914 = ((~WX3481))|((~II10912));
assign II2553 = ((~WX745))|((~II2545));
assign II22642 = ((~II22632))|((~II22640));
assign WX4094 = ((~WX4085));
assign WX8446 = (WX8114&RESET);
assign WX1392 = (WX1786&WX2297);
assign II35170 = ((~WX10930))|((~WX10841));
assign II10151 = ((~II10161))|((~II10162));
assign WX3981 = (WX3979)|(WX3978);
assign II26357 = ((~II26367))|((~II26368));
assign WX688 = (WX356&RESET);
assign WX6092 = ((~II18651))|((~II18652));
assign II35549 = ((~II35539))|((~II35547));
assign WX6498 = (WX6407&WX6435);
assign WX7572 = ((~WX7470));
assign WX10304 = ((~II31683))|((~II31684));
assign WX9221 = (WX10126&WX9222);
assign II15392 = ((~WX4484))|((~WX4414));
assign II10494 = ((~WX3588))|((~WX3263));
assign II2476 = ((~II2451))|((~II2475));
assign WX5270 = (WX5268)|(WX5267);
assign II14268 = ((~WX4732))|((~II14266));
assign WX4041 = (WX4047&WX4042);
assign II14894 = ((~II14869))|((~II14893));
assign II6180 = ((~WX2294))|((~II6179));
assign WX6576 = ((~WX7469));
assign II30427 = ((~WX10052))|((~II30426));
assign WX2191 = (WX2128&RESET);
assign WX6400 = ((~WX6399));
assign WX10013 = ((~WX9982));
assign II14978 = ((~II14980))|((~II14981));
assign II10696 = ((~WX3403))|((~II10695));
assign WX11475 = ((~WX11474));
assign WX3805 = ((~WX3591));
assign WX2575 = (WX2548&WX2556);
assign WX953 = ((~WX952));
assign WX8019 = ((~WX8761));
assign WX9006 = ((~II27643))|((~II27644));
assign WX2536 = ((~II7583))|((~II7584));
assign WX6790 = ((~WX7469));
assign II11510 = ((~WX3225))|((~_2172_));
assign WX9373 = (WX9371)|(WX9370);
assign WX7648 = (WX7070&WX7649);
assign WX9348 = ((~WX10055));
assign II14206 = ((~WX4728))|((~II14204));
assign WX888 = (WX825&RESET);
assign II6659 = ((~WX2108))|((~WX2172));
assign II31297 = ((~WX9568))|((~II31295));
assign II34377 = ((~WX11075))|((~II34376));
assign II14971 = ((~WX4650))|((~II14963));
assign WX1529 = (WX3696&WX1530);
assign II30960 = ((~WX9820))|((~II30952));
assign WX5898 = (WX5835&RESET);
assign WX99 = (WX493&WX1004);
assign WX7388 = ((~II22749))|((~II22750));
assign WX1844 = ((~WX2264));
assign WX4312 = ((~WX4883));
assign WX5802 = ((~WX6045));
assign WX8741 = ((~WX8740));
assign WX5439 = (WX5689&WX6176);
assign II30393 = ((~II30403))|((~II30404));
assign II10864 = ((~II10874))|((~II10875));
assign WX2746 = ((~WX2745));
assign II26676 = ((~WX8509))|((~II26668));
assign WX6628 = ((~WX7468));
assign II10852 = ((~WX3477))|((~II10850));
assign WX1911 = ((~WX2142));
assign WX11381 = ((~WX11349));
assign WX10671 = ((~WX10662));
assign WX1318 = (WX1239&WX1263);
assign II2120 = ((~WX717))|((~II2119));
assign WX2355 = ((~II7162))|((~II7163));
assign II22921 = ((~II22911))|((~II22919));
assign WX10333 = (WX10306&WX10314);
assign WX10391 = ((~WX10382));
assign WX8626 = (WX8563&RESET);
assign II27174 = ((~WX8345))|((~II27173));
assign II2219 = ((~II2221))|((~II2222));
assign WX4241 = (WX6345&WX4242);
assign WX300 = ((~WX299));
assign II2405 = ((~II2407))|((~II2408));
assign II10310 = ((~WX3251))|((~II10308));
assign II22540 = ((~WX7467))|((~WX7144));
assign WX5641 = (WX5652&WX6175);
assign II2033 = ((~II2035))|((~II2036));
assign WX6253 = ((~WX6252));
assign WX10949 = ((~WX10917));
assign II11142 = ((~WX3083))|((~II11140));
assign II6923 = ((~WX2295))|((~WX1998));
assign WX644 = (WX48&RESET);
assign II26888 = ((~WX8459))|((~II26886));
assign II3390 = ((~WX606))|((~WX537));
assign II34990 = ((~WX11346))|((~II34989));
assign II30434 = ((~WX9786))|((~II30433));
assign WX3599 = ((~II11076))|((~II11077));
assign WX3594 = (WX3166&WX3595);
assign WX9652 = ((~WX9620));
assign II35511 = ((~WX10971))|((~II35510));
assign II30387 = ((~II30362))|((~II30386));
assign II18900 = ((~II18890))|((~II18898));
assign WX1922 = ((~WX2164));
assign WX3929 = (WX3935&WX3930);
assign WX9109 = (WX10070&WX9110);
assign II26500 = ((~WX8625))|((~II26498));
assign WX10758 = (WX10764&WX10759);
assign II31641 = ((~WX9675))|((~II31640));
assign II7610 = ((~WX1917))|((~_2127_));
assign WX812 = (WX749&RESET);
assign II22338 = ((~WX7258))|((~WX7322));
assign WX8765 = (WX8764&WX8763);
assign II14134 = ((~WX4596))|((~II14126));
assign II6925 = ((~WX1998))|((~II6923));
assign WX5796 = ((~WX6033));
assign WX5972 = (WX5909&RESET);
assign WX10661 = ((~WX11347));
assign II2421 = ((~II2423))|((~II2424));
assign WX11263 = ((~II34640))|((~II34641));
assign II6489 = ((~WX2295))|((~WX1970));
assign WX10733 = (_2339_&WX11348);
assign II19346 = ((~WX5773))|((~II19345));
assign WX6802 = (WX6992&WX7469);
assign WX995 = ((~WX994));
assign WX6276 = ((~II19255))|((~II19256));
assign II18604 = ((~WX5919))|((~II18596));
assign WX3791 = ((~WX3591));
assign WX977 = ((~WX976));
assign WX5645 = (_2205_&WX6176);
assign WX3682 = ((~WX3681));
assign WX3460 = (WX3397&RESET);
assign WX910 = ((~II2321))|((~II2322));
assign WX6632 = ((~WX7469));
assign WX1248 = ((~II3613))|((~II3614));
assign WX8373 = ((~WX8601));
assign WX1603 = (WX2438&WX1604);
assign II14470 = ((~WX4554))|((~II14468));
assign II6474 = ((~WX2096))|((~II6473));
assign WX10751 = (WX10881&WX11348);
assign II26545 = ((~WX8760))|((~WX8437));
assign DATA_9_4 = ((~WX1200));
assign WX5992 = (WX5929&RESET);
assign WX3577 = ((~WX3576));
assign WX1678 = (WX1689&WX2296);
assign WX2923 = (WX3113&WX3590);
assign WX8806 = ((~II27161))|((~II27162));
assign WX9157 = (WX9163&WX9158);
assign WX1379 = (WX2326&WX1380);
assign WX6856 = ((~WX7469));
assign II26576 = ((~WX8760))|((~WX8439));
assign II10950 = ((~II10926))|((~II10942));
assign WX10044 = ((~WX10043));
assign II34066 = ((~WX11055))|((~II34058));
assign WX8190 = (WX10259&WX8191);
assign WX634 = ((~WX881));
assign II34415 = ((~WX11141))|((~WX11205));
assign II23300 = ((~WX6984))|((~II23298));
assign II2376 = ((~WX797))|((~II2375));
assign WX2760 = ((~WX2759));
assign II31505 = ((~WX9678))|((~_2332_));
assign II3619 = ((~WX626))|((~_2093_));
assign II10200 = ((~WX3371))|((~II10199));
assign II6977 = ((~II6952))|((~II6976));
assign WX6774 = (WX6988&WX7469);
assign WX2801 = ((~WX2792));
assign WX10096 = (WX10094)|(WX10093);
assign II31696 = ((~WX9685))|((~_2309_));
assign II11413 = ((~WX3193))|((~WX3125));
assign II6249 = ((~WX2018))|((~II6248));
assign II30829 = ((~WX10053))|((~WX9748));
assign II26915 = ((~II26925))|((~II26926));
assign WX1367 = (WX1365)|(WX1364);
assign II11581 = ((~WX3205))|((~II11580));
assign II26762 = ((~WX8760))|((~WX8451));
assign WX7363 = (WX7300&RESET);
assign WX1070 = (WX1069&WX1005);
assign II19557 = ((~_2233_))|((~II19555));
assign II18380 = ((~WX6173))|((~WX5841));
assign WX4597 = (WX4534&RESET);
assign II6511 = ((~II6487))|((~II6503));
assign WX1536 = ((~WX1527));
assign WX10681 = (WX10871&WX11348);
assign WX5571 = (WX5582&WX6175);
assign II6697 = ((~II6673))|((~II6689));
assign WX6731 = (WX6729)|(WX6728);
assign WX10635 = (_2346_&WX11348);
assign II30503 = ((~WX9854))|((~WX9918));
assign WX9185 = (WX9191&WX9186);
assign WX10406 = ((~WX10405));
assign II26523 = ((~II26513))|((~II26521));
assign WX10079 = (WX10078&WX10056);
assign WX213 = ((~WX1004));
assign II6620 = ((~WX2042))|((~II6612));
assign WX249 = (_2093_&WX1004);
assign WX4145 = (WX4143)|(WX4142);
assign WX6514 = (WX6525&WX7468);
assign WX6830 = (WX6996&WX7469);
assign II22733 = ((~WX7220))|((~II22725));
assign WX2215 = ((~II6698))|((~II6699));
assign II26042 = ((~II26032))|((~II26040));
assign WX10747 = (_2338_&WX11348);
assign WX3446 = (WX3383&RESET);
assign II34278 = ((~WX11005))|((~II34276));
assign WX6748 = ((~WX7469));
assign WX5541 = ((~WX5532));
assign II22044 = ((~WX7466))|((~WX7112));
assign II34836 = ((~WX11041))|((~II34834));
assign WX7177 = (WX7114&RESET);
assign II14467 = ((~II14469))|((~II14470));
assign II10268 = ((~II10244))|((~II10260));
assign WX6636 = ((~WX7469));
assign II31647 = ((~WX9676))|((~_2318_));
assign II14723 = ((~WX4634))|((~II14715));
assign WX8749 = ((~WX8748));
assign WX430 = (WX428)|(WX427);
assign WX10535 = ((~WX11347));
assign WX2067 = (WX2004&RESET);
assign WX5876 = (WX5640&RESET);
assign WX6352 = ((~WX6351));
assign II6242 = ((~WX2294))|((~II6241));
assign II7569 = ((~WX1911))|((~II7568));
assign WX7898 = (WX7896)|(WX7895);
assign II23208 = ((~WX7055))|((~II23207));
assign WX6478 = (WX6417&WX6435);
assign II26925 = ((~WX8525))|((~II26924));
assign II14097 = ((~WX4880))|((~II14096));
assign II18092 = ((~II18068))|((~II18084));
assign WX214 = (WX212)|(WX211);
assign WX11290 = ((~WX11267));
assign WX6594 = ((~WX7469));
assign WX3999 = (WX4005&WX4000);
assign WX8729 = ((~WX8728));
assign II6458 = ((~WX2294))|((~WX1968));
assign WX11612 = (WX11605&WX11607);
assign WX1261 = ((~II3704))|((~II3705));
assign WX5087 = ((~WX5086));
assign WX11427 = ((~II35236))|((~II35237));
assign WX5856 = (WX5500&RESET);
assign WX6516 = ((~WX7468));
assign WX6877 = ((~WX6876));
assign WX3200 = ((~WX3427));
assign WX1598 = (_2121_&WX2297);
assign WX2307 = (WX2306&WX2298);
assign II23325 = ((~WX7064))|((~II23324));
assign WX942 = ((~WX921));
assign WX2936 = (WX2934)|(WX2933);
assign WX3248 = (WX2760&RESET);
assign WX4549 = (WX4109&RESET);
assign II18450 = ((~WX5909))|((~II18449));
assign II18108 = ((~WX5887))|((~II18100));
assign WX11038 = (WX10742&RESET);
assign WX7722 = ((~II23701))|((~II23702));
assign II10833 = ((~II10843))|((~II10844));
assign WX4189 = (WX5024&WX4190);
assign WX6922 = ((~WX7468));
assign WX2866 = (WX2864)|(WX2863);
assign WX5322 = (WX5320)|(WX5319);
assign WX3378 = (WX3315&RESET);
assign WX8222 = (WX8980&WX8223);
assign II34774 = ((~WX11037))|((~II34772));
assign II30185 = ((~WX9770))|((~II30177));
assign II26507 = ((~II26497))|((~II26505));
assign II14050 = ((~WX4654))|((~II14049));
assign II3418 = ((~WX541))|((~II3416));
assign WX9795 = (WX9732&RESET);
assign WX4593 = (WX4530&RESET);
assign WX9441 = (WX11531&WX9442);
assign WX5371 = ((~WX6176));
assign WX1735 = (WX1741&WX1736);
assign II7319 = ((~WX1818))|((~II7317));
assign WX5791 = ((~WX6023));
assign WX6072 = ((~II18031))|((~II18032));
assign WX3338 = (WX3275&RESET);
assign WX6410 = ((~II19563))|((~II19564));
assign WX8895 = ((~WX8894));
assign WX9112 = ((~WX9103));
assign WX8718 = ((~WX8688));
assign II14683 = ((~II14693))|((~II14694));
assign WX9443 = (WX9441)|(WX9440);
assign WX10280 = ((~WX10279));
assign II11350 = ((~WX3115))|((~II11348));
assign WX3718 = ((~II11297))|((~II11298));
assign WX4187 = (WX4185)|(WX4184);
assign II2150 = ((~WX719))|((~II2142));
assign WX7474 = ((~WX7470));
assign II30814 = ((~WX9874))|((~II30813));
assign II30319 = ((~WX9906))|((~II30317));
assign II18905 = ((~II18915))|((~II18916));
assign WX5310 = (WX7526&WX5311);
assign WX3172 = ((~WX3140));
assign WX6135 = ((~WX6134));
assign II27691 = ((~WX8392))|((~_2277_));
assign II23512 = ((~_2268_))|((~II23510));
assign WX10120 = ((~II31205))|((~II31206));
assign WX3915 = (WX3921&WX3916);
assign II11531 = ((~WX3198))|((~_2171_));
assign WX307 = ((~WX1004));
assign WX1387 = (WX1385)|(WX1384);
assign WX1421 = (WX2347&WX1422);
assign II15081 = ((~WX4460))|((~II15080));
assign WX4830 = ((~WX4829));
assign II14342 = ((~II14352))|((~II14353));
assign II3486 = ((~WX632))|((~II3485));
assign II34174 = ((~II34150))|((~II34166));
assign WX4934 = ((~II15159))|((~II15160));
assign WX4784 = ((~II14181))|((~II14182));
assign II11659 = ((~_2152_))|((~II11657));
assign WX5553 = ((~WX6176));
assign WX10025 = ((~WX9956));
assign WX220 = (WX218)|(WX217);
assign II15531 = ((~_2204_))|((~II15529));
assign II11127 = ((~WX3171))|((~WX3081));
assign WX1003 = ((~WX999));
assign II30753 = ((~WX9934))|((~II30751));
assign II30114 = ((~II30124))|((~II30125));
assign II22487 = ((~II22477))|((~II22485));
assign WX9513 = (WX9511)|(WX9510);
assign WX1918 = ((~WX2156));
assign WX4224 = ((~WX4882));
assign II7528 = ((~_2139_))|((~II7526));
assign WX9325 = (WX9331&WX9326);
assign WX8652 = (WX8589&RESET);
assign WX9317 = (WX9315)|(WX9314);
assign WX7972 = (WX7970)|(WX7969);
assign II30295 = ((~II30285))|((~II30293));
assign II26825 = ((~WX8760))|((~II26824));
assign WX10868 = (WX10871&RESET);
assign WX6240 = ((~WX6239));
assign WX4855 = ((~WX4785));
assign WX7813 = ((~WX8762));
assign II22889 = ((~WX7230))|((~II22888));
assign II5994 = ((~WX2294))|((~II5993));
assign WX3208 = ((~WX3443));
assign WX3620 = ((~II11115))|((~II11116));
assign II34749 = ((~WX11099))|((~II34748));
assign II6117 = ((~WX2294))|((~WX1946));
assign WX10485 = (WX10843&WX11348);
assign II30612 = ((~WX10053))|((~WX9734));
assign WX4156 = (_2187_&WX4883);
assign WX11345 = ((~WX11344));
assign WX10691 = (_2342_&WX11348);
assign WX6584 = (WX6595&WX7468);
assign WX5031 = ((~WX5030));
assign WX8282 = (WX8285&RESET);
assign II22702 = ((~WX7218))|((~II22694));
assign WX9829 = (WX9766&RESET);
assign II26320 = ((~II26295))|((~II26319));
assign WX8141 = ((~WX8132));
assign II19321 = ((~WX5695))|((~II19319));
assign WX4236 = (WX4247&WX4882);
assign II34460 = ((~II34470))|((~II34471));
assign WX91 = (WX102&WX1003);
assign WX4655 = (WX4592&RESET);
assign II10757 = ((~WX3407))|((~WX3471));
assign WX2505 = ((~WX2298));
assign II10098 = ((~WX3301))|((~II10090));
assign WX8777 = ((~WX8776));
assign WX10183 = ((~II31322))|((~II31323));
assign WX7089 = ((~WX7326));
assign WX1865 = ((~WX2242));
assign II31521 = ((~WX9683))|((~II31520));
assign II10160 = ((~WX3305))|((~II10152));
assign WX11286 = ((~WX11265));
assign WX5112 = ((~II15523))|((~II15524));
assign II2157 = ((~II2159))|((~II2160));
assign WX7802 = (WX8770&WX7803);
assign WX3011 = ((~WX3002));
assign II23588 = ((~WX7083))|((~_2261_));
assign WX10668 = (WX11496&WX10669);
assign WX4217 = (WX5038&WX4218);
assign II30040 = ((~WX9888))|((~II30038));
assign WX629 = ((~WX871));
assign II6103 = ((~WX2136))|((~II6101));
assign WX11319 = ((~WX11318));
assign WX1407 = (WX2340&WX1408);
assign II34786 = ((~II34788))|((~II34789));
assign WX7443 = ((~WX7372));
assign II14312 = ((~II14314))|((~II14315));
assign WX5364 = (WX5362)|(WX5361);
assign WX1264 = (WX1234&WX1263);
assign II3593 = ((~_2097_))|((~II3591));
assign II10052 = ((~II10027))|((~II10051));
assign WX137 = (_2101_&WX1004);
assign WX313 = ((~WX304));
assign WX8290 = (WX8293&RESET);
assign II30945 = ((~II30920))|((~II30944));
assign WX6044 = (WX5981&RESET);
assign II10635 = ((~WX3463))|((~II10633));
assign II26134 = ((~II26109))|((~II26133));
assign WX5727 = ((~WX6151));
assign WX2641 = ((~WX3590));
assign II14599 = ((~WX4626))|((~II14591));
assign II7570 = ((~_2133_))|((~II7568));
assign II22277 = ((~WX7254))|((~II22276));
assign WX11581 = ((~II35576))|((~II35577));
assign II27187 = ((~WX8346))|((~II27186));
assign WX3531 = ((~WX3530));
assign II19399 = ((~WX5707))|((~II19397));
assign WX7088 = ((~WX7324));
assign WX9383 = (WX9381)|(WX9380);
assign II26693 = ((~II26683))|((~II26691));
assign WX2834 = (WX2832)|(WX2831);
assign II27002 = ((~II26977))|((~II27001));
assign WX8368 = ((~WX8336));
assign II14017 = ((~II14019))|((~II14020));
assign WX152 = (WX2361&WX153);
assign WX3507 = ((~II10672))|((~II10673));
assign II6785 = ((~WX2180))|((~II6783));
assign WX4952 = (WX4950)|(WX4949);
assign WX2719 = (WX2730&WX3589);
assign II30822 = ((~II30812))|((~II30820));
assign II22712 = ((~WX7346))|((~II22710));
assign II15120 = ((~WX4463))|((~II15119));
assign II7674 = ((~WX1928))|((~II7673));
assign WX4077 = (WX4968&WX4078);
assign II30867 = ((~WX9814))|((~II30859));
assign II19697 = ((~_2211_))|((~II19695));
assign II10601 = ((~II10603))|((~II10604));
assign WX8045 = (WX8056&WX8761);
assign II19295 = ((~WX5691))|((~II19293));
assign WX4107 = (WX4105)|(WX4104);
assign WX4455 = ((~WX4836));
assign II6573 = ((~II6549))|((~II6565));
assign II10713 = ((~WX3277))|((~II10711));
assign WX11534 = (WX10950&WX11535);
assign WX7958 = (WX7956)|(WX7955);
assign WX42 = (WX40)|(WX39);
assign WX10383 = (_2364_&WX11348);
assign II30473 = ((~WX9852))|((~II30472));
assign WX4745 = (WX4682&RESET);
assign WX6619 = (WX6617)|(WX6616);
assign WX8381 = ((~WX8617));
assign WX9127 = ((~WX9126));
assign WX9163 = (WX9161)|(WX9160);
assign WX4024 = ((~WX4015));
assign WX44 = (DATA_9_31&WX45);
assign II10340 = ((~WX3587))|((~II10339));
assign II18247 = ((~II18223))|((~II18239));
assign II19611 = ((~WX5794))|((~_2225_));
assign II7267 = ((~WX1810))|((~II7265));
assign WX5549 = ((~WX6176));
assign WX6099 = ((~II18868))|((~II18869));
assign II23737 = ((~_2237_))|((~II23735));
assign II19165 = ((~WX5671))|((~II19163));
assign II14810 = ((~WX4881))|((~II14809));
assign WX8940 = (WX8939&WX8763);
assign II18085 = ((~WX5949))|((~WX6013));
assign WX3629 = (WX3171&WX3630);
assign WX9272 = (_2319_&WX10055);
assign WX6314 = ((~WX6177));
assign II19268 = ((~WX5767))|((~II19267));
assign WX8458 = (WX8198&RESET);
assign WX1977 = (WX1621&RESET);
assign WX5756 = ((~WX5724));
assign II10353 = ((~II10355))|((~II10356));
assign II7083 = ((~WX1875))|((~WX1782));
assign WX758 = (WX695&RESET);
assign II14175 = ((~WX4726))|((~II14173));
assign II3052 = ((~WX580))|((~WX485));
assign II31141 = ((~WX9544))|((~II31139));
assign WX10448 = ((~WX10447));
assign II10842 = ((~WX3349))|((~II10834));
assign WX7095 = ((~WX7338));
assign WX2300 = (WX2299&WX2298);
assign II22709 = ((~II22711))|((~II22712));
assign II2763 = ((~WX1002))|((~WX695));
assign WX5770 = ((~WX5738));
assign II2297 = ((~II2299))|((~II2300));
assign II30703 = ((~II30713))|((~II30714));
assign WX6809 = (WX6815&WX6810);
assign II6212 = ((~WX1952))|((~II6210));
assign II19640 = ((~WX5798))|((~II19639));
assign II6791 = ((~II6766))|((~II6790));
assign WX1882 = ((~WX1850));
assign WX5065 = ((~WX5064));
assign II22060 = ((~WX7240))|((~II22059));
assign WX1503 = (WX1501)|(WX1500);
assign WX7943 = ((~WX8762));
assign II27650 = ((~WX8384))|((~II27649));
assign WX2097 = (WX2034&RESET);
assign II14259 = ((~WX4604))|((~II14258));
assign WX10716 = (WX10722&WX10717);
assign WX7259 = (WX7196&RESET);
assign WX4321 = (WX4327&WX4322);
assign WX2630 = (WX3598&WX2631);
assign II7654 = ((~_2120_))|((~II7652));
assign WX9672 = ((~WX9906));
assign II31739 = ((~WX9692))|((~II31738));
assign WX10961 = ((~WX11191));
assign WX7844 = (WX8791&WX7845);
assign WX11668 = (WX11580&WX11607);
assign WX8377 = ((~WX8609));
assign WX8893 = ((~WX8763));
assign WX10287 = ((~II31564))|((~II31565));
assign WX5777 = ((~WX5745));
assign WX10954 = ((~WX10922));
assign WX933 = ((~WX932));
assign DATA_9_15 = ((~WX1123));
assign WX1769 = (WX1767)|(WX1766);
assign WX6769 = (WX6767)|(WX6766);
assign WX7640 = (WX7639&WX7470);
assign WX742 = (WX679&RESET);
assign WX5922 = (WX5859&RESET);
assign WX5960 = (WX5897&RESET);
assign WX9958 = ((~II30263))|((~II30264));
assign II23604 = ((~_2259_))|((~II23602));
assign II14770 = ((~II14745))|((~II14769));
assign WX5596 = (WX5594)|(WX5593);
assign II27240 = ((~WX8267))|((~II27238));
assign WX9232 = ((~WX10055));
assign WX3939 = (WX3937)|(WX3936);
assign WX10639 = (WX10865&WX11348);
assign WX2742 = (WX3654&WX2743);
assign II6838 = ((~WX2056))|((~II6837));
assign II30696 = ((~II30672))|((~II30688));
assign II26429 = ((~WX8493))|((~II26428));
assign WX8038 = (WX8036)|(WX8035);
assign II30991 = ((~WX9822))|((~II30983));
assign WX7528 = (WX7527&WX7470);
assign WX129 = ((~WX1004));
assign WX1813 = (WX1816&RESET);
assign WX374 = (WX372)|(WX371);
assign II6279 = ((~WX2020))|((~II6271));
assign WX8110 = (WX8924&WX8111);
assign II34352 = ((~II34354))|((~II34355));
assign WX3037 = ((~WX3590));
assign WX204 = (WX210&WX205);
assign WX9278 = ((~WX10055));
assign WX9300 = (_2317_&WX10055);
assign WX7749 = (WX7719&WX7728);
assign II34942 = ((~WX11175))|((~WX11239));
assign WX2243 = ((~WX2218));
assign WX6054 = (WX5991&RESET);
assign WX10429 = (WX10835&WX11348);
assign WX9733 = (WX9365&RESET);
assign WX10970 = ((~WX11209));
assign WX11406 = ((~II35197))|((~II35198));
assign II31007 = ((~II30982))|((~II31006));
assign WX6907 = (WX6913&WX6908);
assign WX3346 = (WX3283&RESET);
assign II7461 = ((~WX1904))|((~II7460));
assign II35610 = ((~WX10963))|((~_2356_));
assign II15502 = ((~_2204_))|((~II15500));
assign WX11355 = ((~WX11354));
assign II19475 = ((~WX5783))|((~WX5719));
assign II30737 = ((~WX10053))|((~II30736));
assign WX3667 = ((~WX3666));
assign WX2338 = (WX2336)|(WX2335);
assign II34547 = ((~II34522))|((~II34546));
assign II2353 = ((~II2343))|((~II2351));
assign II10139 = ((~WX3431))|((~II10137));
assign WX8700 = ((~WX8679));
assign WX7936 = (WX7934)|(WX7933);
assign WX10675 = ((~WX11347));
assign WX8682 = ((~II26785))|((~II26786));
assign II34913 = ((~WX11237))|((~II34911));
assign WX10803 = (_2334_&WX11348);
assign II30163 = ((~WX9832))|((~II30162));
assign WX6617 = (WX8826&WX6618);
assign WX4463 = ((~WX4431));
assign WX6943 = (WX7694&WX6944);
assign WX8196 = (WX8194)|(WX8193);
assign WX9984 = ((~WX9983));
assign II14692 = ((~WX4632))|((~II14684));
assign WX6555 = ((~WX6554));
assign II6770 = ((~WX1988))|((~II6768));
assign WX4840 = ((~WX4839));
assign WX10632 = (WX10638&WX10633);
assign WX1885 = ((~WX1853));
assign WX6533 = (WX8784&WX6534);
assign WX7964 = (WX7962)|(WX7961);
assign WX2119 = (WX2056&RESET);
assign WX7041 = ((~WX7422));
assign WX2029 = (WX1966&RESET);
assign II30085 = ((~WX10052))|((~WX9700));
assign WX6543 = (WX6549&WX6544);
assign WX6430 = ((~II19703))|((~II19704));
assign WX2179 = (WX2116&RESET);
assign II22230 = ((~WX7466))|((~WX7124));
assign II22046 = ((~WX7112))|((~II22044));
assign WX324 = (DATA_9_11&WX325);
assign II30326 = ((~II30316))|((~II30324));
assign WX196 = (WX194)|(WX193);
assign II26404 = ((~II26406))|((~II26407));
assign II3066 = ((~WX581))|((~II3065));
assign WX10575 = (WX10586&WX11347);
assign WX9351 = ((~WX9350));
assign II2362 = ((~WX669))|((~II2360));
assign II6961 = ((~WX2064))|((~II6953));
assign WX7434 = ((~WX7433));
assign II26182 = ((~II26172))|((~II26180));
assign WX5725 = ((~WX6147));
assign II10418 = ((~WX3449))|((~II10416));
assign II22260 = ((~II22262))|((~II22263));
assign WX4757 = (WX4694&RESET);
assign II14888 = ((~WX4772))|((~II14886));
assign II7254 = ((~WX1808))|((~II7252));
assign WX5098 = ((~WX4884));
assign II34091 = ((~WX11345))|((~II34090));
assign WX9845 = (WX9782&RESET);
assign WX10852 = (WX10855&RESET);
assign II6915 = ((~II6890))|((~II6914));
assign WX5786 = ((~WX6013));
assign II27734 = ((~WX8399))|((~II27733));
assign II2089 = ((~WX715))|((~II2088));
assign WX9593 = (WX9596&RESET);
assign WX8156 = ((~WX8155));
assign WX10728 = ((~WX10727));
assign WX5230 = (WX6191&WX5231);
assign II14212 = ((~II14187))|((~II14211));
assign WX9490 = ((~WX9481));
assign WX232 = (WX238&WX233);
assign WX1644 = (WX1822&WX2297);
assign II35570 = ((~_2362_))|((~II35568));
assign II2196 = ((~II2172))|((~II2188));
assign WX5487 = (WX5498&WX6175);
assign II27630 = ((~_2288_))|((~II27628));
assign WX9189 = (WX11405&WX9190);
assign WX10075 = (WX10073)|(WX10072);
assign II31527 = ((~_2311_))|((~II31519));
assign II18861 = ((~WX5999))|((~II18860));
assign II14708 = ((~II14683))|((~II14707));
assign WX3274 = (WX2942&RESET);
assign WX8664 = ((~II26227))|((~II26228));
assign II23729 = ((~WX7106))|((~II23728));
assign WX1803 = (WX1806&RESET);
assign WX9280 = ((~WX9271));
assign II30672 = ((~II30682))|((~II30683));
assign WX5914 = (WX5851&RESET);
assign II27643 = ((~WX8383))|((~II27642));
assign II22345 = ((~II22321))|((~II22337));
assign WX3496 = ((~II10331))|((~II10332));
assign WX1570 = (_2123_&WX2297);
assign WX4219 = (WX4217)|(WX4216);
assign WX3024 = (WX3022)|(WX3021);
assign II27448 = ((~WX8299))|((~II27446));
assign II10616 = ((~II10626))|((~II10627));
assign WX9153 = (WX9151)|(WX9150);
assign WX9755 = (WX9519&RESET);
assign WX9520 = (WX9531&WX10054);
assign WX3706 = (WX3182&WX3707);
assign WX5634 = (WX5632)|(WX5631);
assign WX3166 = ((~WX3134));
assign WX5283 = ((~WX6176));
assign WX10800 = (WX10806&WX10801);
assign WX9358 = ((~WX10055));
assign II30107 = ((~II30083))|((~II30099));
assign II26244 = ((~II26234))|((~II26242));
assign WX10319 = (WX10312&WX10314);
assign WX8843 = (WX8349&WX8844);
assign II3523 = ((~_2107_))|((~II3521));
assign WX229 = ((~WX220));
assign WX5418 = (WX5424&WX5419);
assign II34603 = ((~WX11217))|((~II34601));
assign II22578 = ((~WX7210))|((~II22570));
assign II22294 = ((~WX7128))|((~II22292));
assign II2577 = ((~WX1002))|((~WX683));
assign II6677 = ((~WX1982))|((~II6675));
assign WX5880 = (WX5817&RESET);
assign WX2942 = ((~WX2941));
assign WX10729 = (WX10740&WX11347);
assign WX10590 = (WX10596&WX10591);
assign WX3914 = (WX3925&WX4882);
assign II26189 = ((~WX8541))|((~II26188));
assign WX8970 = ((~WX8763));
assign WX6570 = (WX6581&WX7468);
assign WX3589 = ((~WX3585));
assign II22493 = ((~WX7268))|((~WX7332));
assign II10401 = ((~WX3587))|((~WX3257));
assign WX9565 = (WX9568&RESET);
assign II30192 = ((~II30194))|((~II30195));
assign WX5764 = ((~WX5732));
assign WX10033 = ((~WX9960));
assign II26476 = ((~II26466))|((~II26474));
assign WX10702 = (WX10708&WX10703);
assign WX2611 = (WX2532&WX2556);
assign WX2807 = (_2159_&WX3590);
assign WX2901 = (WX2912&WX3589);
assign WX2135 = (WX2072&RESET);
assign WX10483 = ((~WX11348));
assign WX1064 = (WX588&WX1065);
assign II18629 = ((~WX6174))|((~II18628));
assign WX1673 = (WX2473&WX1674);
assign WX10035 = ((~WX9961));
assign II3288 = ((~WX521))|((~II3286));
assign WX2239 = ((~WX2216));
assign WX1872 = ((~WX2256));
assign WX2758 = (WX2756)|(WX2755);
assign II18807 = ((~II18797))|((~II18805));
assign WX7475 = (WX7473)|(WX7472);
assign WX9161 = (WX11391&WX9162);
assign WX2660 = (WX2658)|(WX2657);
assign II34693 = ((~II34695))|((~II34696));
assign WX9623 = ((~WX10000));
assign II6288 = ((~WX2084))|((~II6287));
assign II2648 = ((~II2638))|((~II2646));
assign WX1342 = (WX1353&WX2296);
assign II19536 = ((~_2236_))|((~II19534));
assign II22662 = ((~II22672))|((~II22673));
assign II18475 = ((~WX5847))|((~II18473));
assign WX4481 = ((~WX4449));
assign WX6692 = ((~WX7469));
assign WX8121 = ((~WX8762));
assign WX10615 = ((~WX10606));
assign II35660 = ((~WX10970))|((~II35659));
assign II6110 = ((~II6100))|((~II6108));
assign WX9636 = ((~WX9604));
assign WX8444 = (WX8100&RESET);
assign WX120 = (WX126&WX121);
assign II6878 = ((~WX2186))|((~II6876));
assign WX9402 = (WX9580&WX10055);
assign WX905 = ((~II2166))|((~II2167));
assign WX941 = ((~WX940));
assign WX3839 = ((~II11658))|((~II11659));
assign II18628 = ((~WX6174))|((~WX5857));
assign WX4569 = (WX4249&RESET);
assign WX9266 = ((~WX9257));
assign WX1613 = (WX3738&WX1614);
assign WX5614 = (WX5620&WX5615);
assign WX7285 = (WX7222&RESET);
assign WX3092 = (WX3095&RESET);
assign II26211 = ((~WX8479))|((~II26203));
assign WX1422 = ((~WX2297));
assign WX4164 = ((~WX4155));
assign WX4007 = (WX4933&WX4008);
assign WX3047 = ((~WX3590));
assign II11643 = ((~WX3215))|((~_2154_));
assign II2842 = ((~WX891))|((~II2840));
assign WX8101 = (WX8112&WX8761);
assign WX5504 = (WX5502)|(WX5501);
assign II7345 = ((~WX1822))|((~II7343));
assign II6751 = ((~II6753))|((~II6754));
assign WX6936 = ((~WX7468));
assign II22130 = ((~II22120))|((~II22128));
assign WX9385 = (WX11503&WX9386);
assign WX10097 = ((~WX10096));
assign II7497 = ((~_2119_))|((~II7489));
assign WX870 = (WX807&RESET);
assign WX5208 = (WX5214&WX5209);
assign WX6460 = (WX6425&WX6435);
assign WX9429 = (WX9427)|(WX9426);
assign II11231 = ((~WX3179))|((~WX3097));
assign II10812 = ((~WX3347))|((~II10811));
assign II2678 = ((~WX753))|((~II2677));
assign WX1213 = (WX1211)|(WX1210);
assign WX7779 = (WX7706&WX7728);
assign II18217 = ((~II18192))|((~II18216));
assign II35533 = ((~_2343_))|((~II35532));
assign II34051 = ((~II34026))|((~II34050));
assign WX8099 = ((~WX8090));
assign II26739 = ((~WX8513))|((~II26738));
assign WX965 = ((~WX964));
assign WX7761 = (WX7696&WX7728);
assign WX778 = (WX715&RESET);
assign WX11488 = ((~WX11487));
assign WX3614 = (WX3613&WX3591);
assign II22384 = ((~II22386))|((~II22387));
assign II18030 = ((~II18006))|((~II18022));
assign WX8776 = ((~WX8775));
assign WX10215 = (WX10213)|(WX10212);
assign WX296 = (DATA_9_13&WX297);
assign WX10782 = (WX10780)|(WX10779);
assign II3235 = ((~WX594))|((~II3234));
assign WX9773 = (WX9710&RESET);
assign II18776 = ((~II18766))|((~II18774));
assign II18676 = ((~WX6051))|((~II18674));
assign II34423 = ((~II34398))|((~II34422));
assign WX9484 = ((~WX10055));
assign WX4998 = (WX4997&WX4884);
assign WX4262 = ((~WX4253));
assign II15683 = ((~WX4514))|((~_2180_));
assign WX4527 = (WX3955&RESET);
assign WX11467 = ((~WX11466));
assign II34191 = ((~WX11063))|((~II34190));
assign II22557 = ((~WX7336))|((~II22555));
assign WX5117 = ((~II15558))|((~II15559));
assign WX4395 = (WX4398&RESET);
assign II10527 = ((~WX3265))|((~II10525));
assign WX1902 = ((~WX1870));
assign WX1322 = (WX1237&WX1263);
assign II10764 = ((~II10740))|((~II10756));
assign WX10394 = (WX10400&WX10395);
assign II26638 = ((~WX8760))|((~WX8443));
assign WX6993 = (WX6996&RESET);
assign II22882 = ((~WX7467))|((~II22881));
assign WX10985 = ((~WX11239));
assign WX9395 = (WX9401&WX9396);
assign WX810 = (WX747&RESET);
assign II27201 = ((~WX8261))|((~II27199));
assign WX2339 = ((~WX2338));
assign WX2736 = (WX2734)|(WX2733);
assign WX7143 = (WX6751&RESET);
assign WX9132 = (_2329_&WX10055);
assign WX8070 = (WX8068)|(WX8067);
assign WX2276 = ((~WX2275));
assign II26607 = ((~WX8760))|((~WX8441));
assign WX1481 = ((~WX1480));
assign WX338 = (DATA_9_10&WX339);
assign WX5079 = ((~WX5078));
assign WX10678 = (DATA_0_10&WX10679);
assign WX5024 = ((~WX5023));
assign II7534 = ((~WX1906))|((~II7533));
assign WX3151 = ((~WX3521));
assign WX5618 = (WX7680&WX5619);
assign II18395 = ((~WX5969))|((~WX6033));
assign II10276 = ((~II10278))|((~II10279));
assign WX8218 = (WX10273&WX8219);
assign WX7183 = (WX7120&RESET);
assign II6456 = ((~II6466))|((~II6467));
assign II2236 = ((~WX1001))|((~WX661));
assign II10627 = ((~II10617))|((~II10625));
assign II30789 = ((~II30765))|((~II30781));
assign WX1698 = ((~WX2297));
assign II34718 = ((~WX11097))|((~II34717));
assign II6357 = ((~II6332))|((~II6356));
assign II3550 = ((~WX616))|((~II3549));
assign II34672 = ((~II34662))|((~II34670));
assign WX8001 = ((~WX7992));
assign WX6168 = ((~TM0));
assign WX3525 = ((~WX3524));
assign II15635 = ((~WX4505))|((~II15634));
assign WX3436 = (WX3373&RESET);
assign WX3288 = (WX3040&RESET);
assign WX4237 = (WX4243&WX4238);
assign WX10508 = (WX10506)|(WX10505);
assign II11283 = ((~WX3183))|((~WX3105));
assign II6581 = ((~II6583))|((~II6584));
assign WX3617 = (WX3615)|(WX3614);
assign II10379 = ((~II10369))|((~II10377));
assign WX664 = (WX188&RESET);
assign II35674 = ((~WX10973))|((~II35673));
assign II7625 = ((~WX1919))|((~II7624));
assign WX4339 = (WX6394&WX4340);
assign II22904 = ((~II22879))|((~II22903));
assign II10061 = ((~WX3587))|((~II10060));
assign WX6719 = (WX7582&WX6720);
assign II22092 = ((~WX7306))|((~II22090));
assign WX10361 = (WX10294&WX10314);
assign II14082 = ((~WX4720))|((~II14080));
assign II14918 = ((~WX4710))|((~II14917));
assign WX7055 = ((~WX7023));
assign WX9599 = ((~WX10016));
assign II14306 = ((~II14296))|((~II14304));
assign WX1879 = ((~WX1847));
assign WX1223 = ((~II3456))|((~II3457));
assign WX6857 = (WX6855)|(WX6854);
assign WX3588 = ((~WX3584));
assign II22943 = ((~WX7467))|((~WX7170));
assign II7124 = ((~WX1788))|((~II7122));
assign WX1637 = (WX1643&WX1638);
assign WX5751 = ((~WX6135));
assign WX3254 = (WX2802&RESET);
assign WX8851 = ((~WX8763));
assign II19625 = ((~WX5796))|((~_2223_));
assign II35183 = ((~WX10931))|((~WX10843));
assign II14136 = ((~II14126))|((~II14134));
assign II6754 = ((~WX2178))|((~II6752));
assign WX4310 = (_2176_&WX4883);
assign II18062 = ((~II18037))|((~II18061));
assign WX7455 = ((~WX7378));
assign WX5001 = (WX4999)|(WX4998);
assign WX3868 = (WX3841&WX3849);
assign WX4377 = (WX4380&RESET);
assign WX1495 = ((~WX1494));
assign WX7441 = ((~WX7371));
assign WX6957 = (WX6960&RESET);
assign II19267 = ((~WX5767))|((~WX5687));
assign WX2250 = ((~WX2249));
assign WX2668 = (WX4912&WX2669);
assign WX4863 = ((~WX4789));
assign WX5215 = (WX5657&WX6176);
assign II6590 = ((~WX2040))|((~II6589));
assign II11220 = ((~WX3095))|((~II11218));
assign WX6792 = ((~WX6783));
assign WX2848 = (WX2846)|(WX2845);
assign WX1723 = (WX1721)|(WX1720);
assign WX111 = ((~WX1004));
assign II3392 = ((~WX537))|((~II3390));
assign II10083 = ((~II10058))|((~II10082));
assign WX9628 = ((~WX10010));
assign WX10850 = (WX10853&RESET);
assign II19592 = ((~_2228_))|((~II19590));
assign WX9084 = (WX8993&WX9021);
assign WX11262 = ((~II34609))|((~II34610));
assign II7589 = ((~WX1914))|((~_2130_));
assign WX622 = ((~WX857));
assign WX408 = (DATA_9_5&WX409);
assign WX5630 = (WX5628)|(WX5627);
assign II3649 = ((~_2088_))|((~II3647));
assign WX10153 = ((~WX10152));
assign WX2548 = ((~II7667))|((~II7668));
assign II22485 = ((~WX7204))|((~II22477));
assign WX1091 = (WX1090&WX1005);
assign II14623 = ((~WX4881))|((~WX4564));
assign WX8785 = ((~II27122))|((~II27123));
assign WX9875 = (WX9812&RESET);
assign II10027 = ((~II10037))|((~II10038));
assign WX3486 = ((~II10021))|((~II10022));
assign II18366 = ((~WX6031))|((~II18364));
assign II26521 = ((~WX8499))|((~II26513));
assign WX5057 = (WX5055)|(WX5054);
assign WX1163 = ((~WX1005));
assign WX8434 = (WX8030&RESET);
assign WX4941 = ((~II15172))|((~II15173));
assign II27487 = ((~WX8305))|((~II27485));
assign WX2491 = ((~WX2298));
assign WX3741 = (WX3187&WX3742);
assign WX6248 = ((~II19203))|((~II19204));
assign WX2762 = (WX2768&WX2763);
assign WX1851 = ((~WX2278));
assign II31726 = ((~_2305_))|((~II31724));
assign II2948 = ((~II2950))|((~II2951));
assign II26103 = ((~II26078))|((~II26102));
assign II10897 = ((~WX3588))|((~WX3289));
assign WX2841 = ((~WX3590));
assign II6272 = ((~WX2294))|((~WX1956));
assign WX4030 = (_2196_&WX4883);
assign WX2624 = (WX2622)|(WX2621);
assign WX6125 = ((~WX6124));
assign WX4134 = ((~WX4883));
assign WX3394 = (WX3331&RESET);
assign II34632 = ((~WX11155))|((~WX11219));
assign WX2405 = (WX2404&WX2298);
assign WX7700 = ((~II23547))|((~II23548));
assign WX9309 = ((~WX9308));
assign WX10960 = ((~WX11189));
assign II30775 = ((~WX9808))|((~II30774));
assign II7541 = ((~WX1907))|((~II7540));
assign II2740 = ((~WX757))|((~II2739));
assign WX6643 = (WX6641)|(WX6640);
assign WX10277 = ((~WX10056));
assign WX2506 = (WX2504)|(WX2503);
assign WX3212 = ((~WX3451));
assign II2207 = ((~WX659))|((~II2205));
assign WX11448 = ((~II35275))|((~II35276));
assign WX3584 = ((~TM0));
assign II22765 = ((~WX7222))|((~II22764));
assign II15493 = ((~_2188_))|((~II15492));
assign WX1691 = ((~WX1690));
assign WX3956 = (WX3967&WX4882);
assign WX4511 = ((~WX4756));
assign II18847 = ((~WX5871))|((~II18845));
assign WX4769 = (WX4706&RESET);
assign WX2976 = (WX5066&WX2977);
assign II23637 = ((~WX7090))|((~_2254_));
assign WX1391 = (WX1389)|(WX1388);
assign WX1766 = (_2109_&WX2297);
assign II34230 = ((~WX11129))|((~II34229));
assign WX5243 = (WX5661&WX6176);
assign II34647 = ((~II34649))|((~II34650));
assign II10733 = ((~II10709))|((~II10725));
assign II6441 = ((~II6443))|((~II6444));
assign II30263 = ((~II30238))|((~II30262));
assign II14498 = ((~II14500))|((~II14501));
assign WX1134 = (WX598&WX1135);
assign II31451 = ((~WX9659))|((~WX9592));
assign II18289 = ((~WX5835))|((~II18287));
assign WX3144 = ((~WX3571));
assign WX8514 = (WX8451&RESET);
assign WX7692 = (WX7690)|(WX7689);
assign II18611 = ((~II18613))|((~II18614));
assign WX7789 = (WX7701&WX7728);
assign WX9518 = ((~WX9509));
assign II30713 = ((~WX9804))|((~II30712));
assign II18505 = ((~WX6174))|((~II18504));
assign II10532 = ((~WX3329))|((~II10524));
assign WX7394 = ((~II22935))|((~II22936));
assign II30428 = ((~WX9722))|((~II30426));
assign WX3759 = ((~WX3758));
assign WX1418 = ((~WX2297));
assign II6055 = ((~WX2294))|((~WX1942));
assign WX10511 = ((~WX11348));
assign WX3195 = ((~WX3163));
assign WX8820 = ((~II27187))|((~II27188));
assign II6816 = ((~WX2182))|((~II6814));
assign II26947 = ((~II26949))|((~II26950));
assign II14234 = ((~II14236))|((~II14237));
assign WX6233 = ((~WX6232));
assign WX4365 = (WX4368&RESET);
assign II18239 = ((~II18241))|((~II18242));
assign WX6113 = ((~WX6112));
assign WX9889 = (WX9826&RESET);
assign WX5435 = (_2220_&WX6176);
assign WX2206 = ((~II6419))|((~II6420));
assign WX1544 = ((~WX2297));
assign WX11542 = ((~WX11349));
assign WX8169 = ((~WX8160));
assign WX714 = (WX651&RESET);
assign II22254 = ((~II22244))|((~II22252));
assign II34725 = ((~WX11161))|((~WX11225));
assign WX4098 = ((~WX4882));
assign II15620 = ((~WX4503))|((~_2191_));
assign WX8636 = (WX8573&RESET);
assign WX930 = ((~II2941))|((~II2942));
assign II26950 = ((~WX8463))|((~II26948));
assign II2126 = ((~II2128))|((~II2129));
assign WX6104 = ((~WX6088));
assign II23260 = ((~WX7059))|((~II23259));
assign WX3951 = (WX4905&WX3952);
assign II19437 = ((~WX5780))|((~II19436));
assign II6171 = ((~II6146))|((~II6170));
assign WX5384 = (WX6268&WX5385);
assign WX321 = ((~WX1004));
assign WX4779 = ((~II14026))|((~II14027));
assign WX589 = ((~WX557));
assign WX7673 = ((~WX7672));
assign WX2389 = ((~WX2388));
assign WX11323 = ((~WX11322));
assign II18836 = ((~II18812))|((~II18828));
assign WX5159 = (WX5135&WX5142);
assign WX7814 = (WX7812)|(WX7811);
assign WX7536 = (WX7054&WX7537);
assign WX1725 = (WX3794&WX1726);
assign WX10455 = ((~WX11348));
assign WX1857 = ((~WX2226));
assign WX3519 = ((~WX3518));
assign II18442 = ((~WX6173))|((~WX5845));
assign WX8224 = (WX8222)|(WX8221);
assign WX11502 = ((~WX11501));
assign II18519 = ((~WX5977))|((~WX6041));
assign WX580 = ((~WX548));
assign II26795 = ((~WX8453))|((~II26793));
assign II6365 = ((~WX2294))|((~WX1962));
assign WX2442 = ((~WX2298));
assign WX10655 = ((~WX11348));
assign II10423 = ((~II10399))|((~II10415));
assign WX7245 = (WX7182&RESET);
assign WX3694 = (WX3692)|(WX3691);
assign II7357 = ((~WX1896))|((~II7356));
assign WX9478 = (WX9489&WX10054);
assign WX8829 = (WX8347&WX8830);
assign II26311 = ((~II26313))|((~II26314));
assign II19100 = ((~WX5661))|((~II19098));
assign WX2873 = (WX2884&WX3589);
assign WX5254 = (WX7498&WX5255);
assign II22912 = ((~WX7467))|((~WX7168));
assign WX2415 = (WX2413)|(WX2412);
assign II6102 = ((~WX2072))|((~II6101));
assign WX8797 = ((~WX8796));
assign WX5714 = (WX5717&RESET);
assign WX4127 = (WX4125)|(WX4124);
assign WX6917 = (WX6915)|(WX6914);
assign II18781 = ((~II18791))|((~II18792));
assign II6047 = ((~II6022))|((~II6046));
assign WX4449 = ((~WX4824));
assign WX1740 = ((~WX2297));
assign WX7033 = ((~WX7406));
assign II22758 = ((~WX7467))|((~II22757));
assign II19202 = ((~WX5762))|((~WX5677));
assign II26993 = ((~II26995))|((~II26996));
assign II6434 = ((~WX2030))|((~II6426));
assign WX3737 = ((~WX3736));
assign WX2293 = ((~TM1));
assign WX10250 = (WX10248)|(WX10247);
assign WX9821 = (WX9758&RESET);
assign WX6470 = (WX6421&WX6435);
assign WX1753 = (WX3808&WX1754);
assign WX2603 = (WX2536&WX2556);
assign WX8322 = ((~WX8691));
assign II30125 = ((~II30115))|((~II30123));
assign II2057 = ((~WX713))|((~II2049));
assign WX11394 = (WX10930&WX11395);
assign II35730 = ((~WX10982))|((~II35729));
assign II35597 = ((~WX10961))|((~II35596));
assign WX7096 = ((~WX7340));
assign WX7420 = ((~WX7419));
assign WX449 = (WX543&WX1004);
assign II14065 = ((~WX4880))|((~WX4528));
assign WX1192 = (WX1190)|(WX1189);
assign WX5769 = ((~WX5737));
assign WX10583 = (WX10857&WX11348);
assign WX1232 = ((~II3493))|((~II3494));
assign II14686 = ((~WX4881))|((~II14685));
assign WX9013 = ((~II27692))|((~II27693));
assign II31425 = ((~WX9657))|((~WX9588));
assign WX3362 = (WX3299&RESET);
assign WX10026 = ((~WX10025));
assign WX11132 = (WX11069&RESET);
assign WX3987 = (WX3985)|(WX3984);
assign II27356 = ((~WX8359))|((~II27355));
assign II19520 = ((~WX5811))|((~_2236_));
assign II6723 = ((~WX2176))|((~II6721));
assign WX4643 = (WX4580&RESET);
assign WX5430 = ((~WX5429));
assign WX5538 = (WX6345&WX5539);
assign II30024 = ((~WX10052))|((~II30023));
assign WX9205 = (WX9203)|(WX9202);
assign WX7925 = ((~WX8762));
assign WX3768 = (WX3767&WX3591);
assign II23326 = ((~WX6988))|((~II23324));
assign WX2380 = (WX2378)|(WX2377);
assign II26151 = ((~II26141))|((~II26149));
assign II10060 = ((~WX3587))|((~WX3235));
assign WX11440 = ((~WX11439));
assign WX8876 = ((~II27291))|((~II27292));
assign WX2257 = ((~WX2193));
assign WX9743 = (WX9435&RESET);
assign II27381 = ((~WX8361))|((~WX8289));
assign II3104 = ((~WX584))|((~WX493));
assign WX344 = (WX350&WX345);
assign WX3730 = ((~WX3729));
assign WX3219 = ((~WX3465));
assign WX6418 = ((~II19619))|((~II19620));
assign WX4834 = ((~WX4833));
assign WX2317 = (WX2315)|(WX2314);
assign WX7368 = ((~II22129))|((~II22130));
assign II14716 = ((~WX4881))|((~WX4570));
assign WX10595 = ((~WX11348));
assign II27173 = ((~WX8345))|((~WX8257));
assign WX2476 = (WX1898&WX2477);
assign WX4773 = (WX4710&RESET);
assign WX6712 = ((~WX7468));
assign WX2892 = (WX5024&WX2893);
assign WX3770 = ((~WX3591));
assign WX11516 = ((~WX11515));
assign WX1347 = (WX3605&WX1348);
assign II31654 = ((~WX9677))|((~_2317_));
assign WX2471 = (WX2469)|(WX2468);
assign WX7510 = (WX7508)|(WX7507);
assign WX8894 = (WX8892)|(WX8891);
assign II31000 = ((~WX9886))|((~II30999));
assign II10408 = ((~WX3321))|((~II10400));
assign II7598 = ((~_2129_))|((~II7596));
assign WX5223 = ((~WX6175));
assign WX1120 = (WX596&WX1121);
assign II19709 = ((~WX5810))|((~_2209_));
assign WX9251 = (WX9249)|(WX9248);
assign WX8135 = ((~WX8762));
assign WX9789 = (WX9726&RESET);
assign WX8355 = ((~WX8323));
assign WX2675 = ((~WX2666));
assign WX6038 = (WX5975&RESET);
assign WX5133 = ((~II15670))|((~II15671));
assign WX1625 = (WX1623)|(WX1622);
assign II30688 = ((~II30690))|((~II30691));
assign II7136 = ((~WX1879))|((~II7135));
assign WX9438 = ((~WX10054));
assign WX10605 = ((~WX11347));
assign WX5446 = (WX5452&WX5447);
assign WX11162 = (WX11099&RESET);
assign WX11445 = (WX11443)|(WX11442);
assign II23625 = ((~_2256_))|((~II23623));
assign WX10377 = (WX10286&WX10314);
assign WX5139 = ((~II15712))|((~II15713));
assign WX3188 = ((~WX3156));
assign WX10351 = (WX10299&WX10314);
assign WX8490 = (WX8427&RESET);
assign II23142 = ((~WX7050))|((~WX6960));
assign WX10149 = (WX10148&WX10056);
assign WX11279 = ((~WX11278));
assign II6777 = ((~II6767))|((~II6775));
assign WX11457 = (WX10939&WX11458);
assign II2911 = ((~II2901))|((~II2909));
assign WX425 = ((~WX416));
assign II15353 = ((~WX4481))|((~WX4408));
assign WX7858 = (WX8798&WX7859);
assign WX7429 = ((~WX7365));
assign II26141 = ((~II26143))|((~II26144));
assign WX5181 = (WX5126&WX5142);
assign WX4349 = (WX4355&WX4350);
assign WX1129 = (WX1127)|(WX1126);
assign II22650 = ((~WX7342))|((~II22648));
assign II7597 = ((~WX1915))|((~II7596));
assign WX10624 = (WX10622)|(WX10621);
assign WX10414 = (WX10412)|(WX10411);
assign II22139 = ((~WX7118))|((~II22137));
assign WX4440 = ((~WX4870));
assign WX5124 = ((~II15607))|((~II15608));
assign II27123 = ((~WX8249))|((~II27121));
assign II27472 = ((~WX8368))|((~WX8303));
assign WX11421 = (WX11420&WX11349);
assign WX8450 = (WX8142&RESET);
assign WX2968 = (WX2966)|(WX2965);
assign WX11476 = ((~II35327))|((~II35328));
assign WX1256 = ((~II3669))|((~II3670));
assign WX7113 = (WX6541&RESET);
assign WX3710 = ((~WX3709));
assign WX3003 = (_2145_&WX3590);
assign WX10369 = (WX10290&WX10314);
assign WX3678 = (WX3178&WX3679);
assign II6505 = ((~WX2098))|((~II6504));
assign WX10266 = ((~WX10265));
assign II31522 = ((~_2332_))|((~II31520));
assign II15186 = ((~WX4382))|((~II15184));
assign WX11236 = (WX11173&RESET);
assign II15592 = ((~WX4499))|((~_2195_));
assign WX8133 = (_2276_&WX8762);
assign WX59 = ((~WX1004));
assign WX6217 = (WX6215)|(WX6214);
assign II10827 = ((~II10802))|((~II10826));
assign WX10548 = (WX10554&WX10549);
assign WX4468 = ((~WX4436));
assign WX5682 = (WX5685&RESET);
assign WX6306 = (WX5770&WX6307);
assign WX10088 = ((~WX10056));
assign II6931 = ((~WX2062))|((~II6930));
assign WX2049 = (WX1986&RESET);
assign WX1433 = (WX1431)|(WX1430);
assign WX9242 = ((~WX10054));
assign WX334 = (WX2452&WX335);
assign WX11016 = (WX10588&RESET);
assign WX6633 = (WX6631)|(WX6630);
assign WX2597 = (WX2539&WX2556);
assign WX183 = (WX505&WX1004);
assign WX1156 = ((~WX1005));
assign II7369 = ((~WX1897))|((~WX1826));
assign WX9482 = (_2304_&WX10055);
assign WX7359 = (WX7296&RESET);
assign WX7587 = (WX7585)|(WX7584);
assign II15472 = ((~WX4426))|((~II15470));
assign II6808 = ((~II6798))|((~II6806));
assign WX2227 = ((~WX2210));
assign WX145 = ((~WX136));
assign WX11439 = ((~WX11438));
assign II10433 = ((~WX3587))|((~II10432));
assign II34850 = ((~WX11169))|((~II34849));
assign WX4651 = (WX4588&RESET);
assign WX3829 = ((~II11588))|((~II11589));
assign II22766 = ((~II22756))|((~II22764));
assign II10744 = ((~WX3279))|((~II10742));
assign WX5301 = ((~WX6176));
assign WX8678 = ((~II26661))|((~II26662));
assign WX9975 = ((~II30790))|((~II30791));
assign II26724 = ((~II26714))|((~II26722));
assign II23183 = ((~WX6966))|((~II23181));
assign WX8166 = (WX8952&WX8167);
assign WX2822 = (WX4989&WX2823);
assign II22772 = ((~WX7286))|((~WX7350));
assign WX10759 = ((~WX11347));
assign WX6503 = (WX6501)|(WX6500);
assign II26435 = ((~II26437))|((~II26438));
assign II26374 = ((~WX8553))|((~WX8617));
assign WX6323 = ((~WX6322));
assign II22052 = ((~WX7176))|((~II22051));
assign WX5147 = (WX5140&WX5142);
assign II22833 = ((~II22835))|((~II22836));
assign WX9450 = (WX9461&WX10054);
assign WX686 = (WX342&RESET);
assign WX1375 = (WX3619&WX1376);
assign WX446 = (WX2508&WX447);
assign II30294 = ((~II30269))|((~II30293));
assign II2902 = ((~WX831))|((~WX895));
assign WX11587 = ((~II35618))|((~II35619));
assign WX4494 = ((~WX4722));
assign WX985 = ((~WX984));
assign II2703 = ((~WX691))|((~II2701));
assign WX3272 = (WX2928&RESET);
assign WX5452 = (WX5450)|(WX5449);
assign WX2394 = (WX2392)|(WX2391);
assign II14327 = ((~II14329))|((~II14330));
assign WX5513 = ((~WX5504));
assign WX11628 = (WX11598&WX11607);
assign II2002 = ((~II2004))|((~II2005));
assign WX8021 = (_2284_&WX8762);
assign WX6391 = ((~WX6177));
assign WX314 = ((~WX313));
assign WX7408 = ((~WX7407));
assign WX5499 = ((~WX5490));
assign II6498 = ((~II6488))|((~II6496));
assign II6342 = ((~WX2024))|((~II6341));
assign WX6126 = ((~WX6099));
assign II26631 = ((~II26621))|((~II26629));
assign II34865 = ((~WX11346))|((~WX11043));
assign II22679 = ((~WX7280))|((~WX7344));
assign II6372 = ((~WX2026))|((~II6364));
assign II11115 = ((~WX3170))|((~II11114));
assign WX357 = (WX368&WX1003);
assign WX11266 = ((~II34733))|((~II34734));
assign WX7207 = (WX7144&RESET);
assign WX7717 = ((~II23666))|((~II23667));
assign II18930 = ((~II18905))|((~II18929));
assign II14654 = ((~WX4881))|((~WX4566));
assign WX2786 = (WX2784)|(WX2783);
assign WX158 = (WX156)|(WX155);
assign II22160 = ((~II22135))|((~II22159));
assign WX4515 = ((~WX4764));
assign WX11318 = ((~WX11249));
assign II5992 = ((~II5994))|((~II5995));
assign WX3508 = ((~II10703))|((~II10704));
assign WX3190 = ((~WX3158));
assign WX3819 = ((~II11518))|((~II11519));
assign WX10206 = (WX9652&WX10207);
assign WX3638 = (WX3636)|(WX3635);
assign II35708 = ((~WX10979))|((~_2340_));
assign II14562 = ((~WX4881))|((~II14561));
assign WX6147 = ((~WX6146));
assign WX8790 = ((~WX8789));
assign II31217 = ((~WX9641))|((~WX9556));
assign WX1051 = ((~WX1005));
assign II22185 = ((~WX7312))|((~II22183));
assign II22356 = ((~WX7132))|((~II22354));
assign WX5058 = ((~WX5057));
assign WX3578 = ((~WX3500));
assign II3326 = ((~WX601))|((~II3325));
assign II35222 = ((~WX10934))|((~WX10849));
assign II27214 = ((~WX8263))|((~II27212));
assign II18862 = ((~WX6063))|((~II18860));
assign WX6187 = (WX5753&WX6188);
assign II30858 = ((~II30868))|((~II30869));
assign WX5670 = (WX5673&RESET);
assign WX7497 = ((~WX7496));
assign WX9467 = (WX9465)|(WX9464);
assign WX4157 = (WX6303&WX4158);
assign WX3942 = (WX3953&WX4882);
assign WX8990 = ((~II27523))|((~II27524));
assign II27573 = ((~WX8373))|((~II27572));
assign II2857 = ((~WX1002))|((~II2856));
assign WX2724 = (WX4940&WX2725);
assign WX383 = ((~WX374));
assign WX8410 = (WX7862&RESET);
assign WX1141 = (WX599&WX1142);
assign WX10055 = ((~WX10048));
assign II18039 = ((~WX6173))|((~WX5819));
assign II26035 = ((~WX8595))|((~II26033));
assign WX9997 = ((~WX9974));
assign II35157 = ((~WX10929))|((~WX10839));
assign II7603 = ((~WX1916))|((~_2128_));
assign WX8675 = ((~II26568))|((~II26569));
assign II19605 = ((~WX5793))|((~II19604));
assign WX9367 = (WX9373&WX9368);
assign WX958 = ((~WX929));
assign WX9349 = (WX9347)|(WX9346);
assign WX8997 = ((~II27580))|((~II27581));
assign WX6684 = ((~WX7468));
assign WX7710 = ((~II23617))|((~II23618));
assign WX9609 = ((~WX10036));
assign II23494 = ((~II23496))|((~II23497));
assign WX282 = (DATA_9_14&WX283);
assign WX526 = (WX529&RESET);
assign II14003 = ((~WX4880))|((~WX4524));
assign II2095 = ((~II2097))|((~II2098));
assign WX2862 = (WX2860)|(WX2859);
assign WX4900 = (WX4899&WX4884);
assign WX7403 = ((~WX7384));
assign WX3842 = ((~II11679))|((~II11680));
assign WX9196 = ((~WX9187));
assign II2375 = ((~WX797))|((~WX861));
assign WX3886 = (WX3834&WX3849);
assign WX11496 = ((~WX11495));
assign WX8748 = ((~WX8671));
assign WX9315 = (WX11468&WX9316);
assign II30681 = ((~WX9802))|((~II30673));
assign II11467 = ((~WX3133))|((~II11465));
assign II27485 = ((~WX8369))|((~WX8305));
assign II2486 = ((~WX677))|((~II2484));
assign DATA_9_13 = ((~WX1137));
assign WX10004 = ((~WX10003));
assign WX368 = (WX366)|(WX365);
assign II31464 = ((~WX9660))|((~WX9594));
assign II19505 = ((~WX5804))|((~_2236_));
assign WX1168 = (WX1167&WX1005);
assign II27651 = ((~_2285_))|((~II27649));
assign II2181 = ((~WX721))|((~II2173));
assign WX10144 = ((~WX10056));
assign II2197 = ((~II2172))|((~II2196));
assign WX4501 = ((~WX4736));
assign WX8935 = ((~WX8763));
assign WX1749 = (WX1755&WX1750);
assign WX2895 = (WX3109&WX3590);
assign WX5417 = (WX5428&WX6175);
assign WX11305 = ((~WX11304));
assign II3274 = ((~WX597))|((~II3273));
assign WX7798 = (WX10063&WX7799);
assign WX8390 = ((~WX8635));
assign WX7797 = (_2300_&WX8762);
assign WX3896 = (WX3829&WX3849);
assign WX10305 = ((~II31690))|((~II31691));
assign WX7580 = (WX7578)|(WX7577);
assign WX10895 = ((~WX11315));
assign II18537 = ((~WX5851))|((~II18535));
assign II19534 = ((~WX5815))|((~_2236_));
assign II14336 = ((~II14311))|((~II14335));
assign II14491 = ((~II14466))|((~II14490));
assign II6480 = ((~II6456))|((~II6472));
assign WX10259 = ((~WX10258));
assign II14182 = ((~II14172))|((~II14180));
assign WX2653 = (_2170_&WX3590);
assign WX6753 = (WX6759&WX6754);
assign WX2374 = ((~WX2373));
assign WX8644 = (WX8581&RESET);
assign II14870 = ((~II14872))|((~II14873));
assign WX2063 = (WX2000&RESET);
assign WX10224 = ((~WX10223));
assign WX4230 = (WX4408&WX4883);
assign WX10648 = (WX10646)|(WX10645);
assign II6017 = ((~II6007))|((~II6015));
assign WX3930 = ((~WX4882));
assign II10681 = ((~WX3588))|((~II10680));
assign II30583 = ((~WX9732))|((~II30581));
assign II35444 = ((~WX10951))|((~II35443));
assign II14103 = ((~WX4594))|((~II14095));
assign II2508 = ((~II2498))|((~II2506));
assign WX4821 = ((~WX4800));
assign II35512 = ((~_2364_))|((~II35510));
assign WX11419 = ((~WX11418));
assign WX11618 = (WX11603&WX11607);
assign WX4506 = ((~WX4746));
assign II15302 = ((~WX4477))|((~II15301));
assign WX9527 = (WX9525)|(WX9524);
assign WX2262 = ((~WX2261));
assign WX469 = (WX480&WX1003);
assign WX10910 = ((~WX11281));
assign WX2322 = (WX1876&WX2323);
assign WX2817 = (WX2828&WX3589);
assign II15697 = ((~WX4516))|((~_2178_));
assign WX8912 = (WX8911&WX8763);
assign II15677 = ((~WX4513))|((~II15676));
assign WX9331 = (WX9329)|(WX9328);
assign II35619 = ((~_2355_))|((~II35617));
assign II34088 = ((~II34098))|((~II34099));
assign WX7594 = (WX7592)|(WX7591);
assign II30443 = ((~WX9914))|((~II30441));
assign WX1185 = (WX1183)|(WX1182);
assign WX5546 = (WX5544)|(WX5543);
assign WX5225 = (_2235_&WX6176);
assign II23131 = ((~WX6958))|((~II23129));
assign WX4429 = ((~WX4848));
assign WX8397 = ((~WX8649));
assign II31507 = ((~_2332_))|((~II31505));
assign II22920 = ((~WX7232))|((~II22919));
assign II22672 = ((~WX7216))|((~II22671));
assign II2517 = ((~WX679))|((~II2515));
assign II6250 = ((~II6240))|((~II6248));
assign WX248 = (WX246)|(WX245);
assign II14935 = ((~WX4584))|((~II14933));
assign II7291 = ((~WX1891))|((~WX1814));
assign WX5278 = (WX5284&WX5279);
assign WX11144 = (WX11081&RESET);
assign WX1704 = ((~WX1695));
assign II31556 = ((~WX9663))|((~_2331_));
assign II11587 = ((~WX3206))|((~_2163_));
assign WX11380 = (WX10928&WX11381);
assign WX10917 = ((~WX11295));
assign WX277 = (_2091_&WX1004);
assign II31323 = ((~WX9572))|((~II31321));
assign WX11648 = (WX11590&WX11607);
assign II18296 = ((~II18286))|((~II18294));
assign II34416 = ((~WX11141))|((~II34415));
assign WX6404 = ((~II19513))|((~II19514));
assign II18449 = ((~WX5909))|((~II18441));
assign II22958 = ((~WX7298))|((~WX7362));
assign II18054 = ((~WX5947))|((~WX6011));
assign WX9265 = (WX9263)|(WX9262);
assign WX9459 = (WX10245&WX9460);
assign WX8934 = (WX8362&WX8935);
assign WX4435 = ((~WX4860));
assign WX9397 = (WX9395)|(WX9394);
assign II26606 = ((~II26608))|((~II26609));
assign II14343 = ((~II14345))|((~II14346));
assign WX3725 = ((~II11310))|((~II11311));
assign WX2961 = (_2148_&WX3590);
assign II6162 = ((~II6164))|((~II6165));
assign II6491 = ((~WX1970))|((~II6489));
assign II2918 = ((~WX1002))|((~WX705));
assign WX4675 = (WX4612&RESET);
assign WX8232 = (WX10280&WX8233);
assign II7716 = ((~WX1935))|((~II7715));
assign WX363 = ((~WX1004));
assign II34166 = ((~II34168))|((~II34169));
assign WX11078 = (WX11015&RESET);
assign WX6779 = ((~WX6778));
assign WX7073 = ((~WX7041));
assign II14275 = ((~II14265))|((~II14273));
assign II34733 = ((~II34708))|((~II34732));
assign WX142 = (DATA_9_24&WX143);
assign WX780 = (WX717&RESET);
assign WX1657 = (WX1655)|(WX1654);
assign II2730 = ((~II2740))|((~II2741));
assign WX11525 = ((~II35418))|((~II35419));
assign WX10450 = (WX10456&WX10451);
assign WX2987 = ((~WX3589));
assign II27277 = ((~WX8353))|((~WX8273));
assign II22572 = ((~WX7467))|((~II22571));
assign II23481 = ((~WX7076))|((~II23480));
assign II11219 = ((~WX3178))|((~II11218));
assign WX10248 = (WX9658&WX10249);
assign WX7707 = ((~II23596))|((~II23597));
assign WX10842 = (WX10845&RESET);
assign WX5140 = ((~II15719))|((~II15720));
assign II22967 = ((~II22957))|((~II22965));
assign II14547 = ((~WX4750))|((~II14545));
assign II23681 = ((~_2246_))|((~II23679));
assign WX6863 = ((~WX6862));
assign WX3104 = (WX3107&RESET);
assign WX2958 = (WX2964&WX2959);
assign WX6288 = ((~WX6287));
assign II34253 = ((~WX11067))|((~II34252));
assign II22201 = ((~WX7122))|((~II22199));
assign II11708 = ((~_2143_))|((~II11706));
assign WX3382 = (WX3319&RESET);
assign WX3921 = (WX3919)|(WX3918);
assign WX4181 = (WX4187&WX4182);
assign II18844 = ((~II18846))|((~II18847));
assign WX336 = (WX334)|(WX333);
assign WX5468 = (WX6310&WX5469);
assign II6255 = ((~II6257))|((~II6258));
assign WX8705 = ((~WX8704));
assign II26065 = ((~WX8533))|((~II26064));
assign WX3603 = (WX3601)|(WX3600);
assign WX8858 = ((~WX8763));
assign II14779 = ((~WX4881))|((~II14778));
assign II7240 = ((~WX1887))|((~II7239));
assign WX5245 = ((~WX6176));
assign WX11346 = ((~WX11342));
assign II18971 = ((~WX5879))|((~II18969));
assign WX6833 = (WX6831)|(WX6830);
assign WX9719 = (WX9267&RESET);
assign II6335 = ((~WX2294))|((~II6334));
assign WX3608 = (WX3168&WX3609);
assign II30255 = ((~WX9838))|((~WX9902));
assign WX3773 = ((~WX3772));
assign WX10436 = (WX10442&WX10437);
assign WX6229 = (WX5759&WX6230);
assign WX10811 = ((~WX10802));
assign WX6388 = ((~II19463))|((~II19464));
assign WX9090 = (_2332_&WX10055);
assign WX3974 = (_2200_&WX4883);
assign II34430 = ((~II34432))|((~II34433));
assign II6713 = ((~WX2048))|((~II6705));
assign WX5409 = ((~WX6176));
assign WX528 = (WX531&RESET);
assign WX6191 = ((~WX6190));
assign II3599 = ((~WX623))|((~II3598));
assign WX6074 = ((~II18093))|((~II18094));
assign WX4347 = ((~WX4346));
assign WX395 = ((~WX1004));
assign WX61 = ((~WX52));
assign WX9678 = ((~WX9918));
assign WX9493 = (WX9499&WX9494);
assign WX10008 = ((~WX10007));
assign II26112 = ((~WX8759))|((~II26111));
assign WX1867 = ((~WX2246));
assign WX482 = ((~WX481));
assign WX10909 = ((~WX11279));
assign WX6829 = (WX6827)|(WX6826);
assign WX7975 = (WX7986&WX8761);
assign WX3711 = ((~II11284))|((~II11285));
assign II35569 = ((~WX10957))|((~II35568));
assign II31691 = ((~_2310_))|((~II31689));
assign II14461 = ((~II14451))|((~II14459));
assign WX4071 = (WX4069)|(WX4068);
assign WX504 = (WX507&RESET);
assign II10144 = ((~II10120))|((~II10136));
assign WX6488 = (WX6412&WX6435);
assign WX10125 = ((~WX10124));
assign II6389 = ((~II6379))|((~II6387));
assign II10399 = ((~II10409))|((~II10410));
assign II10058 = ((~II10068))|((~II10069));
assign WX5594 = (WX6373&WX5595);
assign DATA_9_10 = ((~WX1158));
assign WX5062 = (WX4484&WX5063);
assign WX4025 = ((~WX4024));
assign WX2829 = ((~WX2820));
assign WX606 = ((~WX574));
assign WX7382 = ((~II22563))|((~II22564));
assign II19139 = ((~WX5667))|((~II19137));
assign WX8256 = (WX8259&RESET);
assign II34150 = ((~II34160))|((~II34161));
assign WX2217 = ((~II6760))|((~II6761));
assign WX10086 = (WX10085&WX10056);
assign II15565 = ((~WX4495))|((~II15564));
assign WX1666 = ((~WX2296));
assign II22788 = ((~WX7467))|((~WX7160));
assign WX7550 = (WX7056&WX7551);
assign WX1676 = ((~WX1667));
assign WX5668 = (WX5671&RESET);
assign WX155 = (WX501&WX1004);
assign II22735 = ((~II22725))|((~II22733));
assign II18288 = ((~WX6173))|((~II18287));
assign WX301 = (WX312&WX1003);
assign II10124 = ((~WX3239))|((~II10122));
assign WX11316 = ((~WX11248));
assign II30828 = ((~II30830))|((~II30831));
assign WX96 = (WX2333&WX97);
assign II30846 = ((~WX9940))|((~II30844));
assign II14824 = ((~WX4704))|((~WX4768));
assign II14677 = ((~II14652))|((~II14676));
assign WX7861 = ((~WX7852));
assign II3656 = ((~_2086_))|((~II3654));
assign WX2945 = ((~WX3589));
assign II23672 = ((~WX7096))|((~_2248_));
assign WX2921 = ((~WX3590));
assign II27741 = ((~WX8400))|((~II27740));
assign WX8280 = (WX8283&RESET);
assign WX10245 = ((~WX10244));
assign II18459 = ((~WX6037))|((~II18457));
assign WX2220 = ((~II6853))|((~II6854));
assign WX6317 = ((~WX6316));
assign II30634 = ((~II30610))|((~II30626));
assign II18706 = ((~WX5989))|((~II18705));
assign WX4140 = ((~WX4882));
assign WX8687 = ((~II26940))|((~II26941));
assign II30279 = ((~WX9776))|((~II30278));
assign II26306 = ((~II26296))|((~II26304));
assign WX10957 = ((~WX11183));
assign WX10983 = ((~WX11235));
assign II10441 = ((~II10431))|((~II10439));
assign WX2031 = (WX1968&RESET);
assign II22246 = ((~WX7252))|((~II22245));
assign II15642 = ((~WX4507))|((~II15641));
assign WX10105 = ((~WX10104));
assign WX4492 = ((~WX4718));
assign WX8761 = ((~WX8757));
assign II34833 = ((~II34835))|((~II34836));
assign II22479 = ((~WX7466))|((~II22478));
assign WX2345 = (WX2343)|(WX2342);
assign WX6380 = ((~WX6379));
assign II7639 = ((~WX1922))|((~II7638));
assign II2816 = ((~II2792))|((~II2808));
assign WX10963 = ((~WX11195));
assign II14252 = ((~WX4880))|((~II14251));
assign II14156 = ((~II14166))|((~II14167));
assign II10820 = ((~WX3411))|((~II10819));
assign II6418 = ((~II6394))|((~II6410));
assign II34376 = ((~WX11075))|((~II34368));
assign WX5038 = ((~WX5037));
assign II2400 = ((~II2390))|((~II2398));
assign II19716 = ((~WX5812))|((~_2207_));
assign WX4912 = ((~WX4911));
assign WX5033 = (WX5032&WX4884);
assign WX10388 = (WX11356&WX10389);
assign WX10282 = ((~II31513))|((~II31514));
assign WX9099 = ((~WX9098));
assign WX1081 = ((~WX1080));
assign WX3684 = (WX3683&WX3591);
assign II15082 = ((~WX4366))|((~II15080));
assign WX6854 = (_2243_&WX7469);
assign II14112 = ((~WX4658))|((~II14111));
assign WX290 = (WX288)|(WX287);
assign WX10409 = ((~WX11347));
assign II18264 = ((~WX5897))|((~II18263));
assign II30812 = ((~II30814))|((~II30815));
assign WX1593 = ((~WX1592));
assign WX4633 = (WX4570&RESET);
assign WX88 = (WX86)|(WX85);
assign II15670 = ((~WX4512))|((~II15669));
assign II18761 = ((~II18751))|((~II18759));
assign WX6321 = ((~WX6177));
assign WX3242 = (WX2718&RESET);
assign WX9347 = (WX10189&WX9348);
assign II2537 = ((~II2513))|((~II2529));
assign WX6921 = (WX6927&WX6922);
assign II14243 = ((~II14218))|((~II14242));
assign WX4322 = ((~WX4882));
assign WX472 = (WX470)|(WX469);
assign II22371 = ((~WX7324))|((~II22369));
assign II2159 = ((~WX783))|((~II2158));
assign II34905 = ((~II34895))|((~II34903));
assign WX5034 = (WX4480&WX5035);
assign WX312 = (WX310)|(WX309);
assign II18984 = ((~WX6007))|((~WX6071));
assign WX2449 = ((~WX2298));
assign WX2260 = ((~WX2259));
assign II18474 = ((~WX6173))|((~II18473));
assign II10449 = ((~WX3451))|((~II10447));
assign II2145 = ((~WX655))|((~II2143));
assign WX3372 = (WX3309&RESET);
assign WX6140 = ((~WX6074));
assign WX4409 = (WX4412&RESET);
assign WX10441 = ((~WX11348));
assign II10788 = ((~WX3409))|((~WX3473));
assign II31668 = ((~WX9680))|((~_2314_));
assign WX4533 = (WX3997&RESET);
assign WX9531 = (WX9529)|(WX9528);
assign WX3655 = ((~II11180))|((~II11181));
assign WX476 = (WX474)|(WX473);
assign WX5366 = (WX7554&WX5367);
assign II14128 = ((~WX4880))|((~II14127));
assign WX3957 = (WX3963&WX3958);
assign II14838 = ((~II14848))|((~II14849));
assign WX9859 = (WX9796&RESET);
assign II10284 = ((~WX3313))|((~II10276));
assign WX1101 = (WX1099)|(WX1098);
assign WX4914 = (WX4913&WX4884);
assign II26893 = ((~WX8523))|((~II26885));
assign II2754 = ((~II2730))|((~II2746));
assign WX6981 = (WX6984&RESET);
assign II10183 = ((~II10185))|((~II10186));
assign WX7476 = ((~WX7475));
assign WX7728 = ((~WX7695));
assign WX1441 = (WX1447&WX1442);
assign WX8648 = (WX8585&RESET);
assign II14497 = ((~II14507))|((~II14508));
assign WX4329 = (WX5094&WX4330);
assign WX9399 = (WX11510&WX9400);
assign WX7082 = ((~WX7312));
assign II6396 = ((~WX2294))|((~WX1964));
assign WX7811 = (_2299_&WX8762);
assign II23404 = ((~WX7000))|((~II23402));
assign II30479 = ((~II30455))|((~II30471));
assign WX10973 = ((~WX11215));
assign WX4623 = (WX4560&RESET);
assign WX10381 = ((~WX11347));
assign WX3013 = (WX3024&WX3589);
assign II6875 = ((~II6877))|((~II6878));
assign WX9113 = ((~WX9112));
assign II23714 = ((~WX7103))|((~_2241_));
assign II6952 = ((~II6962))|((~II6963));
assign WX9699 = (WX9127&RESET);
assign WX8048 = (WX8046)|(WX8045);
assign II27161 = ((~WX8344))|((~II27160));
assign WX2095 = (WX2032&RESET);
assign II7214 = ((~WX1885))|((~II7213));
assign WX11577 = ((~II35548))|((~II35549));
assign II14423 = ((~WX4742))|((~II14421));
assign WX6255 = ((~II19216))|((~II19217));
assign WX4832 = ((~WX4831));
assign WX1426 = (WX1437&WX2296);
assign II7097 = ((~WX1876))|((~II7096));
assign WX1114 = ((~WX1005));
assign WX10577 = ((~WX11347));
assign WX3782 = (WX3781&WX3591);
assign WX8383 = ((~WX8621));
assign WX10684 = (WX10682)|(WX10681);
assign WX9617 = ((~WX9988));
assign WX1518 = (WX1804&WX2297);
assign WX3815 = ((~WX3814));
assign WX409 = ((~WX1004));
assign II30614 = ((~WX9734))|((~II30612));
assign WX10699 = ((~WX10690));
assign II10368 = ((~II10378))|((~II10379));
assign WX5113 = ((~II15530))|((~II15531));
assign WX9327 = (WX9325)|(WX9324);
assign WX10476 = ((~WX10475));
assign II22029 = ((~WX7238))|((~II22028));
assign WX2486 = ((~WX2485));
assign II23651 = ((~WX7093))|((~_2251_));
assign WX1888 = ((~WX1856));
assign WX4997 = ((~II15276))|((~II15277));
assign WX8868 = ((~WX8867));
assign II3627 = ((~WX628))|((~II3626));
assign WX4289 = (WX4287)|(WX4286);
assign WX8395 = ((~WX8645));
assign WX1015 = (WX581&WX1016);
assign WX5479 = ((~WX6176));
assign WX4885 = ((~II15068))|((~II15069));
assign II34368 = ((~II34370))|((~II34371));
assign II18249 = ((~II18239))|((~II18247));
assign II22501 = ((~II22476))|((~II22500));
assign WX1864 = ((~WX2240));
assign II34805 = ((~WX11039))|((~II34803));
assign WX3775 = (WX3774&WX3591);
assign WX7973 = ((~WX7964));
assign II34650 = ((~WX11029))|((~II34648));
assign II18103 = ((~WX5823))|((~II18101));
assign II7187 = ((~WX1883))|((~WX1798));
assign WX9803 = (WX9740&RESET);
assign WX5400 = (WX5398)|(WX5397);
assign WX6257 = (WX5763&WX6258);
assign WX10884 = (WX10887&RESET);
assign WX9510 = (_2302_&WX10055);
assign II11128 = ((~WX3171))|((~II11127));
assign WX8572 = (WX8509&RESET);
assign II7435 = ((~WX1902))|((~II7434));
assign WX5292 = (WX5298&WX5293);
assign II34414 = ((~II34416))|((~II34417));
assign II30797 = ((~II30799))|((~II30800));
assign II3484 = ((~II3486))|((~II3487));
assign WX11247 = ((~II34144))|((~II34145));
assign WX49 = (WX60&WX1003);
assign WX3240 = (WX2704&RESET);
assign WX6745 = (WX6743)|(WX6742);
assign WX3675 = ((~WX3674));
assign WX8083 = ((~WX8762));
assign II30270 = ((~II30272))|((~II30273));
assign II26389 = ((~II26391))|((~II26392));
assign WX7642 = ((~WX7470));
assign II14669 = ((~WX4694))|((~WX4758));
assign WX11575 = ((~II35518))|((~II35519));
assign WX8043 = ((~WX8034));
assign WX10230 = ((~WX10229));
assign II35633 = ((~_2353_))|((~II35631));
assign II31705 = ((~_2308_))|((~II31703));
assign WX6512 = ((~WX6503));
assign WX2939 = ((~WX3590));
assign II30465 = ((~WX9788))|((~II30464));
assign II14026 = ((~II14001))|((~II14025));
assign WX1912 = ((~WX2144));
assign WX6629 = (WX6627)|(WX6626);
assign WX9154 = ((~WX9145));
assign WX6831 = (WX7638&WX6832);
assign WX6734 = ((~WX7469));
assign WX7805 = ((~WX7796));
assign WX586 = ((~WX554));
assign WX5256 = (WX5254)|(WX5253);
assign WX11417 = (WX11415)|(WX11414);
assign II7652 = ((~WX1924))|((~_2120_));
assign WX3202 = ((~WX3431));
assign WX11064 = (WX11001&RESET);
assign WX10533 = (WX10544&WX11347);
assign WX5850 = (WX5458&RESET);
assign II3516 = ((~_2108_))|((~II3514));
assign WX9419 = (WX9417)|(WX9416);
assign WX6149 = ((~WX6148));
assign WX1018 = ((~WX1017));
assign WX1435 = (WX2354&WX1436);
assign II6210 = ((~WX2294))|((~WX1952));
assign WX2367 = ((~WX2366));
assign WX3112 = (WX3115&RESET);
assign II31549 = ((~WX9694))|((~_2332_));
assign WX7951 = (_2289_&WX8762);
assign WX10278 = (WX10276)|(WX10275);
assign WX5934 = (WX5871&RESET);
assign WX6374 = ((~II19437))|((~II19438));
assign WX6345 = ((~WX6344));
assign WX8726 = ((~WX8660));
assign WX11260 = ((~II34547))|((~II34548));
assign II26258 = ((~II26233))|((~II26257));
assign WX10797 = ((~WX10788));
assign II35659 = ((~WX10970))|((~_2349_));
assign WX5773 = ((~WX5741));
assign WX1373 = (WX1371)|(WX1370);
assign II18542 = ((~WX5915))|((~II18534));
assign WX9973 = ((~II30728))|((~II30729));
assign WX11150 = (WX11087&RESET);
assign WX1601 = (WX1599)|(WX1598);
assign II34447 = ((~WX11143))|((~II34446));
assign WX4102 = ((~WX4883));
assign WX5268 = (WX7505&WX5269);
assign II9997 = ((~II9999))|((~II10000));
assign II18279 = ((~II18254))|((~II18278));
assign II11699 = ((~WX3224))|((~_2145_));
assign WX10521 = ((~WX11347));
assign WX10902 = ((~WX11329));
assign II14973 = ((~II14963))|((~II14971));
assign WX6899 = (WX6897)|(WX6896);
assign II31438 = ((~WX9658))|((~WX9590));
assign II2222 = ((~WX851))|((~II2220));
assign WX5049 = ((~WX4884));
assign WX4717 = (WX4654&RESET);
assign II34478 = ((~WX11145))|((~II34477));
assign II2036 = ((~WX839))|((~II2034));
assign WX8264 = (WX8267&RESET);
assign II22897 = ((~WX7294))|((~II22896));
assign II18017 = ((~II18007))|((~II18015));
assign II31387 = ((~WX9654))|((~II31386));
assign WX6784 = (_2248_&WX7469);
assign WX5108 = ((~WX5107));
assign WX9457 = (WX9455)|(WX9454);
assign WX4818 = ((~WX4817));
assign WX8456 = (WX8184&RESET);
assign II14857 = ((~WX4770))|((~II14855));
assign WX104 = ((~WX103));
assign WX9140 = ((~WX9131));
assign II26512 = ((~II26522))|((~II26523));
assign II15663 = ((~WX4510))|((~II15662));
assign WX9659 = ((~WX9627));
assign II31733 = ((~_2303_))|((~II31731));
assign WX4755 = (WX4692&RESET);
assign WX1849 = ((~WX2274));
assign WX632 = ((~WX877));
assign WX9664 = ((~WX9890));
assign II6320 = ((~WX2150))|((~II6318));
assign WX10756 = ((~WX10755));
assign II23547 = ((~WX7077))|((~II23546));
assign II6482 = ((~II6472))|((~II6480));
assign WX10738 = (WX11531&WX10739);
assign WX1251 = ((~II3634))|((~II3635));
assign II18735 = ((~II18737))|((~II18738));
assign WX10749 = ((~WX11348));
assign WX939 = ((~WX938));
assign WX9779 = (WX9716&RESET);
assign WX5862 = (WX5542&RESET);
assign II10231 = ((~WX3373))|((~II10230));
assign II3682 = ((~WX637))|((~_2082_));
assign WX10666 = (WX10664)|(WX10663);
assign WX7573 = (WX7571)|(WX7570);
assign II18265 = ((~II18255))|((~II18263));
assign II18549 = ((~II18551))|((~II18552));
assign WX9567 = (WX9570&RESET);
assign II11064 = ((~WX3071))|((~II11062));
assign WX2101 = (WX2038&RESET);
assign WX9701 = (WX9141&RESET);
assign II18241 = ((~WX5959))|((~II18240));
assign WX10290 = ((~II31585))|((~II31586));
assign WX3669 = ((~II11206))|((~II11207));
assign II6815 = ((~WX2118))|((~II6814));
assign WX8907 = ((~WX8763));
assign II3600 = ((~_2096_))|((~II3598));
assign WX1266 = (WX1262&WX1263);
assign WX10735 = ((~WX11348));
assign WX10373 = (WX10288&WX10314);
assign II27083 = ((~WX8338))|((~II27082));
assign II6022 = ((~II6032))|((~II6033));
assign WX7911 = ((~WX8762));
assign WX10938 = ((~WX10906));
assign WX8724 = ((~WX8659));
assign II22161 = ((~II22151))|((~II22159));
assign WX11500 = ((~WX11349));
assign II22416 = ((~WX7466))|((~WX7136));
assign WX1221 = ((~WX1220));
assign WX6804 = ((~WX7469));
assign II2377 = ((~WX861))|((~II2375));
assign WX215 = ((~WX206));
assign II7687 = ((~WX1930))|((~_2114_));
assign II18661 = ((~WX5859))|((~II18659));
assign II14684 = ((~II14686))|((~II14687));
assign II6186 = ((~WX2014))|((~II6178));
assign WX3983 = ((~WX3982));
assign WX3005 = ((~WX3590));
assign WX8331 = ((~WX8709));
assign II10262 = ((~WX3375))|((~II10261));
assign II22495 = ((~WX7332))|((~II22493));
assign II19507 = ((~_2236_))|((~II19505));
assign WX3622 = (WX3170&WX3623);
assign II15132 = ((~WX4464))|((~WX4374));
assign II14903 = ((~WX4881))|((~II14902));
assign WX10400 = (WX10398)|(WX10397);
assign WX218 = (WX224&WX219);
assign WX4227 = (WX6338&WX4228);
assign WX8966 = ((~WX8965));
assign II23534 = ((~II23524))|((~II23532));
assign WX3592 = ((~II11063))|((~II11064));
assign WX8536 = (WX8473&RESET);
assign II18063 = ((~II18053))|((~II18061));
assign WX7841 = ((~WX8762));
assign WX9277 = (WX10154&WX9278);
assign WX1228 = ((~WX1227));
assign WX11493 = ((~WX11349));
assign WX4243 = (WX4241)|(WX4240);
assign II34841 = ((~WX11105))|((~II34833));
assign II14203 = ((~II14205))|((~II14206));
assign II6304 = ((~WX2294))|((~II6303));
assign II15545 = ((~_2202_))|((~II15543));
assign WX8064 = (WX10196&WX8065);
assign WX1263 = ((~WX1230));
assign II18874 = ((~II18884))|((~II18885));
assign WX2329 = (WX1877&WX2330);
assign WX4047 = (WX4045)|(WX4044);
assign II15263 = ((~WX4474))|((~II15262));
assign II2407 = ((~WX799))|((~II2406));
assign WX9118 = (_2330_&WX10055);
assign II18464 = ((~II18440))|((~II18456));
assign WX11371 = ((~II35132))|((~II35133));
assign II22719 = ((~II22709))|((~II22717));
assign II18605 = ((~WX5919))|((~II18604));
assign II14569 = ((~WX4624))|((~II14568));
assign II22369 = ((~WX7260))|((~WX7324));
assign WX1175 = (WX1174&WX1005);
assign WX5576 = (WX7659&WX5577);
assign II7071 = ((~WX1874))|((~II7070));
assign II34679 = ((~WX11346))|((~WX11031));
assign II6968 = ((~II6970))|((~II6971));
assign WX11122 = (WX11059&RESET);
assign II10968 = ((~II10958))|((~II10966));
assign WX3154 = ((~WX3527));
assign WX11478 = (WX10942&WX11479);
assign II18025 = ((~WX6009))|((~II18023));
assign WX6928 = (WX7010&WX7469);
assign II2764 = ((~WX1002))|((~II2763));
assign II34493 = ((~WX11345))|((~WX11019));
assign WX3164 = ((~WX3547));
assign WX9107 = (WX9105)|(WX9104);
assign WX1002 = ((~WX998));
assign WX3404 = (WX3341&RESET);
assign II7280 = ((~WX1812))|((~II7278));
assign WX10416 = (WX11370&WX10417);
assign WX970 = ((~WX903));
assign II18768 = ((~WX5993))|((~II18767));
assign II2718 = ((~WX883))|((~II2716));
assign WX7934 = (WX7940&WX7935);
assign WX9124 = ((~WX10055));
assign WX1009 = ((~WX1005));
assign WX7373 = ((~II22284))|((~II22285));
assign WX6592 = (WX6962&WX7469);
assign WX9135 = (WX9133)|(WX9132);
assign WX796 = (WX733&RESET);
assign II26336 = ((~WX8487))|((~II26335));
assign WX5565 = (WX5707&WX6176);
assign WX4110 = (WX4121&WX4882);
assign WX5718 = (WX5655&RESET);
assign II26133 = ((~II26109))|((~II26125));
assign II34882 = ((~WX11235))|((~II34880));
assign II30526 = ((~WX9792))|((~II30518));
assign WX9378 = ((~WX9369));
assign II14755 = ((~WX4636))|((~II14754));
assign II2933 = ((~WX833))|((~WX897));
assign II11512 = ((~_2172_))|((~II11510));
assign WX2353 = ((~WX2352));
assign II10857 = ((~II10833))|((~II10849));
assign II6946 = ((~II6921))|((~II6945));
assign WX5616 = (WX5614)|(WX5613);
assign WX1785 = (WX1788&RESET);
assign II18744 = ((~II18719))|((~II18743));
assign II34408 = ((~WX11077))|((~II34407));
assign WX11280 = ((~WX11262));
assign II22542 = ((~WX7144))|((~II22540));
assign WX8922 = (WX8920)|(WX8919);
assign II19345 = ((~WX5773))|((~WX5699));
assign WX676 = (WX272&RESET);
assign II22151 = ((~II22153))|((~II22154));
assign II2562 = ((~WX809))|((~II2561));
assign II22362 = ((~WX7196))|((~II22361));
assign WX11022 = (WX10630&RESET);
assign WX9879 = (WX9816&RESET);
assign WX7791 = (WX7700&WX7728);
assign WX708 = (WX645&RESET);
assign WX4040 = (WX4051&WX4882);
assign II11207 = ((~WX3093))|((~II11205));
assign WX3344 = (WX3281&RESET);
assign WX1108 = (WX1106)|(WX1105);
assign WX2348 = ((~II7149))|((~II7150));
assign II22108 = ((~WX7116))|((~II22106));
assign II10487 = ((~II10477))|((~II10485));
assign WX4828 = ((~WX4827));
assign WX2643 = (WX3073&WX3590);
assign II22407 = ((~II22383))|((~II22399));
assign II3300 = ((~WX599))|((~II3299));
assign WX2199 = ((~II6202))|((~II6203));
assign WX439 = ((~WX430));
assign WX3059 = (_2141_&WX3590);
assign II2329 = ((~WX1001))|((~WX667));
assign WX3574 = ((~WX3498));
assign II18868 = ((~II18843))|((~II18867));
assign WX7556 = (WX7555&WX7470);
assign WX11044 = (WX10784&RESET);
assign WX8183 = ((~WX8174));
assign II26934 = ((~WX8653))|((~II26932));
assign II18970 = ((~WX6174))|((~II18969));
assign WX530 = (WX533&RESET);
assign II18146 = ((~II18148))|((~II18149));
assign II14592 = ((~WX4881))|((~WX4562));
assign WX10349 = (WX10300&WX10314);
assign WX720 = (WX657&RESET);
assign II6310 = ((~WX2022))|((~II6302));
assign II34029 = ((~WX11345))|((~II34028));
assign II11567 = ((~WX3203))|((~II11566));
assign II10337 = ((~II10347))|((~II10348));
assign WX9915 = (WX9852&RESET);
assign II18303 = ((~WX5963))|((~II18302));
assign II31088 = ((~WX9631))|((~II31087));
assign II22237 = ((~WX7188))|((~II22229));
assign WX11174 = (WX11111&RESET);
assign II31245 = ((~WX9560))|((~II31243));
assign WX5680 = (WX5683&RESET);
assign II14280 = ((~II14290))|((~II14291));
assign WX4389 = (WX4392&RESET);
assign WX1474 = ((~WX2297));
assign WX3130 = (WX3133&RESET);
assign II35470 = ((~WX10953))|((~II35469));
assign II23430 = ((~WX7004))|((~II23428));
assign WX8983 = (WX8369&WX8984);
assign II30364 = ((~WX10052))|((~WX9718));
assign II22123 = ((~WX7308))|((~II22121));
assign II11685 = ((~WX3222))|((~_2147_));
assign WX11414 = (WX11413&WX11349);
assign II6767 = ((~II6769))|((~II6770));
assign WX7634 = (WX7068&WX7635);
assign II22693 = ((~II22703))|((~II22704));
assign WX9004 = ((~II27629))|((~II27630));
assign WX3945 = (WX3943)|(WX3942);
assign WX9649 = ((~WX9617));
assign II34997 = ((~WX11115))|((~II34996));
assign WX9074 = (WX8998&WX9021);
assign WX8886 = ((~WX8763));
assign II19662 = ((~_2217_))|((~II19660));
assign WX8580 = (WX8517&RESET);
assign II6783 = ((~WX2116))|((~WX2180));
assign WX1718 = ((~WX1709));
assign II34200 = ((~WX11191))|((~II34198));
assign WX554 = ((~WX977));
assign II10255 = ((~II10245))|((~II10253));
assign II3494 = ((~II3484))|((~II3492));
assign WX4158 = ((~WX4883));
assign WX6359 = ((~WX6358));
assign WX6271 = (WX5765&WX6272);
assign WX9642 = ((~WX9610));
assign II10935 = ((~WX3355))|((~II10927));
assign WX4442 = ((~WX4874));
assign WX6020 = (WX5957&RESET);
assign II10571 = ((~WX3395))|((~WX3459));
assign WX11338 = ((~WX11259));
assign WX7275 = (WX7212&RESET);
assign WX7884 = (WX7882)|(WX7881);
assign WX10506 = (WX10512&WX10507);
assign WX512 = (WX515&RESET);
assign WX11485 = (WX10943&WX11486);
assign WX3086 = (WX3089&RESET);
assign WX5335 = ((~WX6175));
assign II14415 = ((~II14405))|((~II14413));
assign II11665 = ((~WX3219))|((~II11664));
assign WX11553 = ((~II35470))|((~II35471));
assign II30053 = ((~II30055))|((~II30056));
assign II6040 = ((~WX2068))|((~II6039));
assign II3698 = ((~_2079_))|((~II3696));
assign WX135 = ((~WX1003));
assign II34624 = ((~WX11091))|((~II34616));
assign WX5016 = ((~WX5015));
assign DATA_9_22 = ((~WX1074));
assign WX7175 = (WX7112&RESET);
assign WX7638 = ((~WX7637));
assign WX3928 = (WX3939&WX4882);
assign II31542 = ((~_2304_))|((~II31534));
assign WX1563 = (WX1561)|(WX1560);
assign WX10566 = (DATA_0_18&WX10567);
assign II18203 = ((~II18193))|((~II18201));
assign II14901 = ((~II14903))|((~II14904));
assign II30133 = ((~WX9894))|((~II30131));
assign II15607 = ((~WX4501))|((~II15606));
assign WX9486 = (WX9592&WX10055);
assign WX6991 = (WX6994&RESET);
assign WX5393 = (_2223_&WX6176);
assign II30139 = ((~II30114))|((~II30138));
assign WX10072 = (WX10071&WX10056);
assign WX9965 = ((~II30480))|((~II30481));
assign II30766 = ((~II30768))|((~II30769));
assign WX4086 = (_2192_&WX4883);
assign II14032 = ((~II14042))|((~II14043));
assign WX3286 = (WX3026&RESET);
assign II22376 = ((~II22352))|((~II22368));
assign WX10112 = ((~WX10111));
assign II10549 = ((~II10539))|((~II10547));
assign WX11036 = (WX10728&RESET);
assign WX452 = (WX450)|(WX449);
assign II14345 = ((~WX4880))|((~II14344));
assign WX6664 = ((~WX7469));
assign II31153 = ((~WX9636))|((~II31152));
assign WX6564 = (WX6958&WX7469);
assign WX7564 = (WX7058&WX7565);
assign WX9614 = ((~WX10046));
assign WX2918 = (WX2916)|(WX2915);
assign II6744 = ((~WX2050))|((~II6736));
assign WX1965 = (WX1537&RESET);
assign WX2639 = (_2171_&WX3590);
assign WX10163 = (WX10162&WX10056);
assign WX3870 = (WX3840&WX3849);
assign II10890 = ((~II10880))|((~II10888));
assign II30155 = ((~WX9768))|((~II30154));
assign WX616 = ((~WX845));
assign WX10941 = ((~WX10909));
assign II11155 = ((~WX3085))|((~II11153));
assign WX11365 = (WX11364&WX11349);
assign WX1358 = ((~WX2296));
assign WX5299 = (WX5669&WX6176);
assign II6007 = ((~II6009))|((~II6010));
assign WX2204 = ((~II6357))|((~II6358));
assign WX4306 = (WX4317&WX4882);
assign WX4709 = (WX4646&RESET);
assign II14451 = ((~II14453))|((~II14454));
assign II6821 = ((~II6797))|((~II6813));
assign WX611 = ((~WX579));
assign WX461 = ((~WX1004));
assign WX7309 = (WX7246&RESET);
assign II11694 = ((~_2146_))|((~II11692));
assign WX1520 = ((~WX2297));
assign WX7020 = ((~WX7444));
assign WX6611 = ((~WX6610));
assign II31747 = ((~_2301_))|((~II31745));
assign II6739 = ((~WX1986))|((~II6737));
assign II6536 = ((~WX2100))|((~II6535));
assign WX3034 = (WX3032)|(WX3031);
assign II14160 = ((~WX4534))|((~II14158));
assign WX948 = ((~WX924));
assign II14530 = ((~WX4881))|((~WX4558));
assign II14297 = ((~WX4670))|((~WX4734));
assign II34042 = ((~II34044))|((~II34045));
assign II10471 = ((~WX3325))|((~II10470));
assign WX4787 = ((~II14274))|((~II14275));
assign II2941 = ((~II2916))|((~II2940));
assign WX6262 = ((~II19229))|((~II19230));
assign II31577 = ((~WX9666))|((~_2328_));
assign II19632 = ((~WX5797))|((~_2222_));
assign WX8554 = (WX8491&RESET);
assign WX5557 = (WX5568&WX6175);
assign II7384 = ((~WX1828))|((~II7382));
assign II7708 = ((~WX1934))|((~_2110_));
assign WX2696 = (WX4926&WX2697);
assign WX1409 = (WX1407)|(WX1406);
assign WX6725 = (WX6731&WX6726);
assign WX2769 = (WX3091&WX3590);
assign II34354 = ((~WX11137))|((~II34353));
assign WX8925 = ((~II27382))|((~II27383));
assign WX1330 = ((~WX2296));
assign WX1086 = ((~WX1005));
assign II34789 = ((~WX11229))|((~II34787));
assign WX8979 = ((~WX8978));
assign WX4105 = (WX4982&WX4106);
assign WX10084 = ((~WX10083));
assign WX8808 = (WX8344&WX8809);
assign WX9207 = (WX10119&WX9208);
assign WX5732 = ((~WX6161));
assign WX2311 = ((~WX2310));
assign WX3762 = (WX3190&WX3763);
assign II6691 = ((~WX2110))|((~II6690));
assign WX6945 = (WX6943)|(WX6942);
assign II10186 = ((~WX3243))|((~II10184));
assign II2545 = ((~II2547))|((~II2548));
assign II34123 = ((~WX10995))|((~II34121));
assign II11481 = ((~WX3213))|((~II11480));
assign WX3276 = (WX2956&RESET);
assign WX7491 = ((~WX7490));
assign II19598 = ((~WX5792))|((~II19597));
assign WX5443 = ((~WX5434));
assign WX1453 = ((~WX1452));
assign II34338 = ((~WX11345))|((~WX11009));
assign II18316 = ((~II18326))|((~II18327));
assign II3471 = ((~WX627))|((~II3470));
assign II34153 = ((~WX11345))|((~II34152));
assign WX10171 = (WX9647&WX10172);
assign WX3516 = ((~II10951))|((~II10952));
assign WX3746 = ((~II11349))|((~II11350));
assign II11546 = ((~WX3200))|((~II11545));
assign II3612 = ((~WX625))|((~_2094_));
assign WX8992 = ((~II27545))|((~II27546));
assign II2175 = ((~WX1001))|((~II2174));
assign WX8826 = ((~WX8825));
assign WX2632 = (WX2630)|(WX2629);
assign II35750 = ((~WX10986))|((~_2333_));
assign II30727 = ((~II30703))|((~II30719));
assign II19293 = ((~WX5769))|((~WX5691));
assign WX5527 = ((~WX5518));
assign II18125 = ((~II18115))|((~II18123));
assign WX5696 = (WX5699&RESET);
assign WX2885 = ((~WX2876));
assign WX11598 = ((~II35695))|((~II35696));
assign WX1380 = ((~WX2297));
assign II22843 = ((~II22833))|((~II22841));
assign WX11168 = (WX11105&RESET);
assign II30588 = ((~WX9796))|((~II30580));
assign WX163 = ((~WX1003));
assign WX2051 = (WX1988&RESET);
assign WX3536 = ((~WX3511));
assign WX4667 = (WX4604&RESET);
assign WX8999 = ((~II27594))|((~II27595));
assign WX7515 = (WX7051&WX7516);
assign II6450 = ((~II6425))|((~II6449));
assign WX4780 = ((~II14057))|((~II14058));
assign WX5550 = (WX5548)|(WX5547);
assign WX7484 = ((~WX7483));
assign II34681 = ((~WX11031))|((~II34679));
assign II14366 = ((~II14342))|((~II14358));
assign WX4246 = ((~WX4883));
assign II34036 = ((~WX11053))|((~II34035));
assign WX6505 = (WX8770&WX6506);
assign WX1462 = (WX1796&WX2297);
assign WX6656 = ((~WX7468));
assign WX6911 = (WX8973&WX6912);
assign WX7656 = ((~WX7470));
assign WX10518 = ((~WX10517));
assign WX11196 = (WX11133&RESET);
assign WX4525 = (WX3941&RESET);
assign II34246 = ((~WX11345))|((~II34245));
assign II14404 = ((~II14414))|((~II14415));
assign WX5080 = ((~WX5079));
assign II15615 = ((~_2192_))|((~II15613));
assign WX5497 = ((~WX6176));
assign II14529 = ((~II14531))|((~II14532));
assign II6518 = ((~II6528))|((~II6529));
assign WX9365 = ((~WX9364));
assign WX7682 = (WX7681&WX7470);
assign WX4982 = ((~WX4981));
assign WX2585 = (WX2544&WX2556);
assign II26484 = ((~WX8759))|((~II26483));
assign WX559 = ((~WX987));
assign II27538 = ((~_2272_))|((~II27537));
assign II22447 = ((~WX7466))|((~WX7138));
assign WX11114 = (WX11051&RESET);
assign II31557 = ((~WX9663))|((~II31556));
assign II34324 = ((~WX11199))|((~II34322));
assign II22649 = ((~WX7278))|((~II22648));
assign II18334 = ((~WX5965))|((~II18333));
assign II15146 = ((~WX4465))|((~II15145));
assign WX2539 = ((~II7604))|((~II7605));
assign II23079 = ((~WX6950))|((~II23077));
assign II15290 = ((~WX4398))|((~II15288));
assign WX5381 = ((~WX6176));
assign WX8867 = ((~WX8866));
assign WX8042 = (WX8040)|(WX8039);
assign WX8315 = ((~WX8741));
assign II26382 = ((~II26357))|((~II26381));
assign WX4587 = (WX4524&RESET);
assign WX10221 = ((~WX10056));
assign WX10528 = (WX11426&WX10529);
assign WX8362 = ((~WX8330));
assign WX9089 = (WX9087)|(WX9086);
assign II22634 = ((~WX7467))|((~II22633));
assign II11101 = ((~WX3169))|((~WX3077));
assign II34523 = ((~II34525))|((~II34526));
assign II6521 = ((~WX2295))|((~II6520));
assign WX1400 = ((~WX2296));
assign WX9843 = (WX9780&RESET);
assign WX10673 = (WX10684&WX11347);
assign WX6967 = (WX6970&RESET);
assign II23234 = ((~WX7057))|((~II23233));
assign WX3050 = (WX3808&WX3051);
assign WX932 = ((~WX916));
assign WX4069 = (WX4075&WX4070);
assign WX11535 = ((~WX11349));
assign II22393 = ((~WX7198))|((~II22392));
assign WX1550 = ((~WX1541));
assign WX11570 = ((~WX11349));
assign WX1436 = ((~WX2297));
assign WX4092 = ((~WX4883));
assign WX2296 = ((~WX2292));
assign WX5465 = ((~WX6176));
assign WX2439 = ((~II7318))|((~II7319));
assign II22097 = ((~II22073))|((~II22089));
assign WX8260 = (WX8263&RESET);
assign WX9921 = (WX9858&RESET);
assign WX9018 = ((~II27727))|((~II27728));
assign WX6198 = ((~WX6197));
assign WX2530 = ((~II7541))|((~II7542));
assign WX4971 = (WX4471&WX4972);
assign II26592 = ((~WX8567))|((~II26591));
assign II30441 = ((~WX9850))|((~WX9914));
assign WX3217 = ((~WX3461));
assign WX8816 = ((~WX8763));
assign WX1527 = (WX1525)|(WX1524);
assign WX5040 = (WX5039&WX4884);
assign WX11330 = ((~WX11255));
assign II22564 = ((~II22554))|((~II22562));
assign WX8751 = ((~WX8750));
assign WX5600 = (WX5606&WX5601);
assign WX5357 = ((~WX6176));
assign WX202 = ((~WX201));
assign WX11451 = ((~WX11349));
assign II35301 = ((~WX10940))|((~II35300));
assign II30371 = ((~WX9782))|((~II30363));
assign II26073 = ((~II26063))|((~II26071));
assign WX9686 = ((~WX9934));
assign WX1469 = (WX1475&WX1470);
assign II34533 = ((~II34523))|((~II34531));
assign WX6689 = (WX6687)|(WX6686);
assign II10578 = ((~II10554))|((~II10570));
assign WX4292 = (WX4303&WX4882);
assign II22914 = ((~WX7168))|((~II22912));
assign WX11551 = ((~WX11550));
assign WX1290 = (WX1252&WX1263);
assign II11638 = ((~_2155_))|((~II11636));
assign WX1365 = (WX2319&WX1366);
assign WX8230 = (WX8228)|(WX8227);
assign WX10343 = (WX10302&WX10314);
assign WX5361 = (WX5372&WX6175);
assign II30495 = ((~WX9790))|((~II30487));
assign II31258 = ((~WX9562))|((~II31256));
assign WX8628 = (WX8565&RESET);
assign WX10015 = ((~WX9951));
assign II6852 = ((~II6828))|((~II6844));
assign WX10226 = (WX10225&WX10056);
assign WX4214 = ((~WX4883));
assign WX2714 = (WX3640&WX2715);
assign WX6330 = ((~WX6329));
assign II23716 = ((~_2241_))|((~II23714));
assign II10921 = ((~II10911))|((~II10919));
assign WX4035 = (WX4947&WX4036);
assign II31536 = ((~WX9690))|((~II31535));
assign WX646 = (WX62&RESET);
assign WX5312 = (WX5310)|(WX5309);
assign WX106 = (WX112&WX107);
assign II30557 = ((~WX9794))|((~II30549));
assign WX168 = (WX166)|(WX165);
assign II3339 = ((~WX602))|((~II3338));
assign WX8306 = ((~WX8723));
assign II30860 = ((~WX10053))|((~WX9750));
assign II15303 = ((~WX4400))|((~II15301));
assign WX10190 = ((~II31335))|((~II31336));
assign WX7153 = (WX6821&RESET);
assign II18226 = ((~WX6173))|((~II18225));
assign WX8236 = (WX8987&WX8237);
assign WX9225 = ((~WX9224));
assign WX2733 = (WX2744&WX3589);
assign II3675 = ((~WX636))|((~_2083_));
assign WX7629 = (WX7627)|(WX7626);
assign WX4796 = ((~II14553))|((~II14554));
assign WX2775 = (WX2786&WX3589);
assign II6319 = ((~WX2086))|((~II6318));
assign II11552 = ((~WX3201))|((~_2168_));
assign II2152 = ((~II2142))|((~II2150));
assign II6660 = ((~WX2108))|((~II6659));
assign WX6705 = (WX7575&WX6706);
assign WX900 = ((~II2011))|((~II2012));
assign WX4847 = ((~WX4781));
assign WX2996 = (WX2994)|(WX2993);
assign WX736 = (WX673&RESET);
assign II2772 = ((~II2762))|((~II2770));
assign WX3434 = (WX3371&RESET);
assign WX7945 = ((~WX7936));
assign WX6161 = ((~WX6160));
assign II30930 = ((~WX9818))|((~II30929));
assign WX7123 = (WX6611&RESET);
assign II27672 = ((~_2281_))|((~II27670));
assign WX8897 = ((~II27330))|((~II27331));
assign WX1908 = ((~WX2136));
assign WX1337 = (WX2305&WX1338);
assign WX9046 = (WX9011&WX9021);
assign WX7503 = (WX7501)|(WX7500);
assign II18962 = ((~II18952))|((~II18960));
assign WX7065 = ((~WX7033));
assign WX10186 = ((~WX10056));
assign WX1805 = (WX1808&RESET);
assign WX5026 = (WX5025&WX4884);
assign WX1534 = ((~WX2297));
assign DATA_9_2 = ((~WX1214));
assign WX11274 = ((~II34981))|((~II34982));
assign WX4689 = (WX4626&RESET);
assign II10215 = ((~WX3587))|((~WX3245));
assign WX7343 = (WX7280&RESET);
assign WX11292 = ((~WX11268));
assign II23170 = ((~WX6964))|((~II23168));
assign WX1578 = ((~WX1569));
assign WX561 = ((~WX991));
assign WX2682 = (WX4919&WX2683);
assign WX10890 = (WX10827&RESET);
assign II14621 = ((~II14631))|((~II14632));
assign II22440 = ((~II22430))|((~II22438));
assign WX3466 = (WX3403&RESET);
assign WX4430 = ((~WX4850));
assign WX8333 = ((~WX8713));
assign WX3558 = ((~WX3490));
assign II10961 = ((~WX3293))|((~II10959));
assign II15094 = ((~WX4461))|((~II15093));
assign WX1773 = (WX1771)|(WX1770);
assign WX3308 = (WX3245&RESET);
assign II6636 = ((~II6611))|((~II6635));
assign WX6155 = ((~WX6154));
assign WX3223 = ((~WX3473));
assign II26940 = ((~II26915))|((~II26939));
assign WX6602 = (_2261_&WX7469);
assign WX2793 = (_2160_&WX3590);
assign WX8520 = (WX8457&RESET);
assign WX10205 = (WX10204&WX10056);
assign WX4196 = ((~WX4882));
assign WX6094 = ((~II18713))|((~II18714));
assign WX8468 = (WX8405&RESET);
assign WX1557 = (WX3710&WX1558);
assign WX680 = (WX300&RESET);
assign II7397 = ((~WX1830))|((~II7395));
assign II26646 = ((~WX8507))|((~II26645));
assign WX1943 = (WX1383&RESET);
assign II30893 = ((~WX9752))|((~II30891));
assign II26543 = ((~II26553))|((~II26554));
assign II26831 = ((~WX8519))|((~II26823));
assign WX400 = (WX406&WX401);
assign WX7878 = (WX7884&WX7879);
assign WX854 = (WX791&RESET);
assign II7449 = ((~WX1838))|((~II7447));
assign II19463 = ((~WX5782))|((~II19462));
assign II34061 = ((~WX10991))|((~II34059));
assign II31676 = ((~WX9681))|((~II31675));
assign II15394 = ((~WX4414))|((~II15392));
assign II2455 = ((~WX675))|((~II2453));
assign II22805 = ((~WX7352))|((~II22803));
assign WX1738 = (_2111_&WX2297);
assign WX7448 = ((~WX7447));
assign WX975 = ((~WX974));
assign WX10893 = ((~WX11311));
assign II30334 = ((~WX10052))|((~II30333));
assign II26529 = ((~WX8563))|((~WX8627));
assign WX6369 = (WX5779&WX6370);
assign WX1901 = ((~WX1869));
assign II34471 = ((~II34461))|((~II34469));
assign WX8024 = (WX8022)|(WX8021);
assign II14189 = ((~WX4880))|((~WX4536));
assign II6088 = ((~WX1944))|((~II6086));
assign WX2519 = ((~WX2298));
assign II6202 = ((~II6177))|((~II6201));
assign WX4273 = (WX5066&WX4274);
assign WX7909 = (_2292_&WX8762);
assign WX1280 = (WX1256&WX1263);
assign WX6462 = (WX6424&WX6435);
assign II26764 = ((~WX8451))|((~II26762));
assign II10495 = ((~WX3588))|((~II10494));
assign WX1302 = (WX1247&WX1263);
assign WX10048 = ((~TM0));
assign WX5352 = (WX7547&WX5353);
assign II22648 = ((~WX7278))|((~WX7342));
assign II30938 = ((~WX9882))|((~II30937));
assign II14484 = ((~WX4682))|((~II14483));
assign II26454 = ((~WX8431))|((~II26452));
assign WX5543 = (WX5554&WX6175);
assign II35004 = ((~WX11179))|((~WX11243));
assign II2315 = ((~WX857))|((~II2313));
assign II23561 = ((~WX7079))|((~II23560));
assign WX7875 = ((~WX7866));
assign WX8317 = ((~WX8745));
assign II2724 = ((~II2699))|((~II2723));
assign WX4869 = ((~WX4792));
assign WX8910 = ((~WX8909));
assign II10036 = ((~WX3297))|((~II10028));
assign WX7804 = (WX7802)|(WX7801);
assign WX8345 = ((~WX8313));
assign WX11547 = (WX11546&WX11349);
assign WX4860 = ((~WX4859));
assign II11678 = ((~WX3221))|((~_2148_));
assign WX6746 = (WX6984&WX7469);
assign WX9606 = ((~WX10030));
assign WX8783 = ((~WX8782));
assign WX1497 = (WX1503&WX1498);
assign II14197 = ((~WX4600))|((~II14196));
assign WX4909 = ((~WX4884));
assign II27370 = ((~WX8287))|((~II27368));
assign WX3061 = ((~WX3590));
assign WX7013 = ((~WX7430));
assign WX10924 = ((~WX10892));
assign II27684 = ((~WX8391))|((~_2278_));
assign WX4360 = ((~WX4351));
assign WX2424 = ((~WX2423));
assign WX7777 = (WX7707&WX7728);
assign II30875 = ((~WX9878))|((~WX9942));
assign II15685 = ((~_2180_))|((~II15683));
assign II2082 = ((~WX1001))|((~II2081));
assign WX10300 = ((~II31655))|((~II31656));
assign WX1488 = ((~WX2297));
assign II22880 = ((~II22882))|((~II22883));
assign WX3256 = (WX2816&RESET);
assign WX6209 = ((~WX6177));
assign WX6590 = ((~WX7469));
assign WX10403 = ((~WX11348));
assign II2017 = ((~II2027))|((~II2028));
assign II23209 = ((~WX6970))|((~II23207));
assign WX4259 = (WX5059&WX4260);
assign II35689 = ((~_2344_))|((~II35687));
assign II26599 = ((~II26574))|((~II26598));
assign WX4017 = (WX6233&WX4018);
assign WX5119 = ((~II15572))|((~II15573));
assign WX10746 = (WX10744)|(WX10743);
assign WX8841 = ((~II27226))|((~II27227));
assign WX11385 = ((~II35158))|((~II35159));
assign WX9180 = ((~WX10055));
assign WX1618 = ((~WX2297));
assign WX8566 = (WX8503&RESET);
assign WX9985 = ((~WX9968));
assign WX7513 = ((~II23156))|((~II23157));
assign WX1344 = ((~WX2296));
assign WX5515 = (WX5526&WX6175);
assign WX5236 = (WX5242&WX5237);
assign II10330 = ((~II10306))|((~II10322));
assign WX7091 = ((~WX7330));
assign II10416 = ((~WX3385))|((~WX3449));
assign WX7840 = (WX10084&WX7841);
assign WX5628 = (WX5634&WX5629);
assign II7583 = ((~WX1913))|((~II7582));
assign WX6200 = (WX6199&WX6177);
assign II2671 = ((~WX1002))|((~II2670));
assign WX8200 = (WX8206&WX8201);
assign II11401 = ((~WX3192))|((~II11400));
assign II6444 = ((~WX2158))|((~II6442));
assign II23441 = ((~WX7073))|((~WX7006));
assign II22470 = ((~II22445))|((~II22469));
assign II26636 = ((~II26646))|((~II26647));
assign II7226 = ((~WX1886))|((~WX1804));
assign II2244 = ((~WX725))|((~II2243));
assign II2694 = ((~II2684))|((~II2692));
assign II18072 = ((~WX5821))|((~II18070));
assign WX7401 = ((~WX7383));
assign WX10420 = ((~WX10419));
assign II10193 = ((~II10183))|((~II10191));
assign II10766 = ((~II10756))|((~II10764));
assign WX10147 = ((~WX10146));
assign WX6295 = ((~WX6294));
assign WX11250 = ((~II34237))|((~II34238));
assign WX10838 = (WX10841&RESET);
assign WX4379 = (WX4382&RESET);
assign II7122 = ((~WX1878))|((~WX1788));
assign WX11589 = ((~II35632))|((~II35633));
assign WX3019 = ((~WX3590));
assign WX1760 = ((~WX1751));
assign WX5294 = (WX5292)|(WX5291);
assign II26082 = ((~WX8407))|((~II26080));
assign II31565 = ((~_2330_))|((~II31563));
assign II10130 = ((~WX3303))|((~II10129));
assign II18774 = ((~II18750))|((~II18766));
assign WX5003 = ((~WX5002));
assign II34104 = ((~II34106))|((~II34107));
assign WX3142 = ((~WX3567));
assign WX1904 = ((~WX1872));
assign WX440 = ((~WX439));
assign WX2512 = ((~WX2298));
assign II27318 = ((~WX8279))|((~II27316));
assign WX10363 = (WX10293&WX10314);
assign II34476 = ((~II34478))|((~II34479));
assign II34215 = ((~WX11345))|((~II34214));
assign II26686 = ((~WX8637))|((~II26684));
assign WX10780 = (WX11552&WX10781);
assign WX9082 = (WX8994&WX9021);
assign II6194 = ((~WX2078))|((~WX2142));
assign WX3965 = (WX4912&WX3966);
assign WX2463 = ((~WX2298));
assign II34429 = ((~II34439))|((~II34440));
assign WX7453 = ((~WX7377));
assign II15579 = ((~WX4497))|((~II15578));
assign WX1038 = (WX1036)|(WX1035);
assign WX9919 = (WX9856&RESET);
assign II15551 = ((~WX4493))|((~II15550));
assign II26213 = ((~II26203))|((~II26211));
assign WX304 = (WX302)|(WX301);
assign II34587 = ((~WX11346))|((~II34586));
assign II6094 = ((~WX2008))|((~II6093));
assign WX10886 = (WX10889&RESET);
assign WX284 = (WX282)|(WX281);
assign II22945 = ((~WX7170))|((~II22943));
assign WX10526 = (WX10524)|(WX10523);
assign WX6770 = (_2249_&WX7469);
assign WX113 = (WX495&WX1004);
assign WX10947 = ((~WX10915));
assign II22533 = ((~II22523))|((~II22531));
assign II31520 = ((~WX9683))|((~_2332_));
assign WX6421 = ((~II19640))|((~II19641));
assign II10650 = ((~WX3588))|((~II10649));
assign II27383 = ((~WX8289))|((~II27381));
assign II22099 = ((~II22089))|((~II22097));
assign II22570 = ((~II22572))|((~II22573));
assign WX9683 = ((~WX9928));
assign II26078 = ((~II26088))|((~II26089));
assign II11616 = ((~WX3210))|((~II11615));
assign WX506 = (WX509&RESET);
assign WX7053 = ((~WX7021));
assign II19647 = ((~WX5800))|((~II19646));
assign WX4031 = (WX6240&WX4032);
assign WX7566 = (WX7564)|(WX7563);
assign II26833 = ((~II26823))|((~II26831));
assign II15558 = ((~WX4494))|((~II15557));
assign WX3850 = (WX3820&WX3849);
assign WX9393 = ((~WX9392));
assign WX5437 = ((~WX6176));
assign WX8436 = (WX8044&RESET);
assign WX5374 = ((~WX5373));
assign WX8889 = ((~WX8888));
assign WX3601 = (WX3167&WX3602);
assign II22601 = ((~II22603))|((~II22604));
assign II14516 = ((~WX4748))|((~II14514));
assign WX11540 = (WX11539&WX11349);
assign WX2547 = ((~II7660))|((~II7661));
assign II11575 = ((~_2165_))|((~II11573));
assign WX3418 = (WX3355&RESET);
assign WX11532 = ((~II35431))|((~II35432));
assign WX5237 = ((~WX6175));
assign WX10568 = (WX10566)|(WX10565);
assign WX9456 = ((~WX10055));
assign II7632 = ((~WX1921))|((~II7631));
assign II10905 = ((~WX3353))|((~II10904));
assign WX8512 = (WX8449&RESET);
assign II15432 = ((~WX4487))|((~II15431));
assign WX6586 = ((~WX7468));
assign II2656 = ((~WX879))|((~II2654));
assign WX10155 = ((~II31270))|((~II31271));
assign II2097 = ((~WX779))|((~II2096));
assign II35583 = ((~WX10959))|((~II35582));
assign II11589 = ((~_2163_))|((~II11587));
assign II30982 = ((~II30992))|((~II30993));
assign II14625 = ((~WX4564))|((~II14623));
assign WX2493 = ((~WX2492));
assign II19113 = ((~WX5663))|((~II19111));
assign WX4088 = ((~WX4883));
assign II18599 = ((~WX5855))|((~II18597));
assign WX1939 = (WX1355&RESET);
assign WX5247 = ((~WX5238));
assign II14073 = ((~WX4592))|((~II14072));
assign WX7560 = ((~WX7559));
assign WX10539 = ((~WX11348));
assign II18890 = ((~II18892))|((~II18893));
assign WX6123 = ((~WX6122));
assign II22074 = ((~II22076))|((~II22077));
assign WX7991 = ((~WX8761));
assign WX3612 = ((~WX3611));
assign WX1853 = ((~WX2282));
assign WX2403 = ((~WX2402));
assign WX267 = (WX517&WX1004);
assign WX3735 = ((~WX3591));
assign WX2127 = (WX2064&RESET);
assign WX1183 = (WX605&WX1184);
assign II18270 = ((~II18272))|((~II18273));
assign WX6115 = ((~WX6114));
assign WX5213 = ((~WX6176));
assign WX10646 = (WX10652&WX10647);
assign WX6159 = ((~WX6158));
assign WX8546 = (WX8483&RESET);
assign WX2591 = (WX2542&WX2556);
assign II22781 = ((~II22771))|((~II22779));
assign WX10490 = ((~WX10489));
assign II30923 = ((~WX10053))|((~II30922));
assign II27728 = ((~_2271_))|((~II27726));
assign WX6641 = (WX6647&WX6642);
assign WX7399 = ((~WX7382));
assign WX2626 = (WX4891&WX2627);
assign WX4367 = (WX4370&RESET);
assign WX4319 = ((~WX4318));
assign WX1577 = (WX1575)|(WX1574);
assign WX7757 = (WX7716&WX7728);
assign II7474 = ((~II7476))|((~II7477));
assign II3247 = ((~WX595))|((~WX515));
assign WX8787 = (WX8341&WX8788);
assign II10625 = ((~WX3335))|((~II10617));
assign WX7139 = (WX6723&RESET);
assign II2709 = ((~WX755))|((~II2708));
assign II34634 = ((~WX11219))|((~II34632));
assign WX2334 = ((~II7123))|((~II7124));
assign II11285 = ((~WX3105))|((~II11283));
assign WX11400 = (WX11399&WX11349);
assign II6270 = ((~II6280))|((~II6281));
assign WX967 = ((~WX966));
assign II30783 = ((~WX9872))|((~II30782));
assign II26654 = ((~WX8571))|((~II26653));
assign WX8905 = (WX8904&WX8763);
assign WX638 = ((~WX889));
assign II2957 = ((~WX771))|((~II2956));
assign WX1925 = ((~WX2170));
assign WX1635 = ((~WX1634));
assign WX342 = ((~WX341));
assign WX2295 = ((~WX2291));
assign WX437 = ((~WX1004));
assign II10067 = ((~WX3299))|((~II10059));
assign II14963 = ((~II14965))|((~II14966));
assign WX4249 = ((~WX4248));
assign II31374 = ((~WX9653))|((~II31373));
assign WX6915 = (WX7680&WX6916);
assign WX2310 = (WX2308)|(WX2307);
assign WX8924 = ((~WX8923));
assign II6404 = ((~WX2028))|((~II6403));
assign WX8216 = (WX8214)|(WX8213);
assign WX6951 = (WX6954&RESET);
assign WX1471 = (WX1469)|(WX1468);
assign II10045 = ((~WX3361))|((~II10044));
assign WX9307 = (WX9305)|(WX9304);
assign WX8600 = (WX8537&RESET);
assign WX7024 = ((~WX7452));
assign II34113 = ((~II34088))|((~II34112));
assign WX3392 = (WX3329&RESET);
assign WX6995 = (WX6998&RESET);
assign II10803 = ((~II10805))|((~II10806));
assign II35695 = ((~WX10977))|((~II35694));
assign WX9130 = ((~WX10054));
assign II30123 = ((~WX9766))|((~II30115));
assign WX6884 = ((~WX7469));
assign WX1951 = (WX1439&RESET);
assign WX7582 = ((~WX7581));
assign II2234 = ((~II2244))|((~II2245));
assign II18784 = ((~WX6174))|((~II18783));
assign II2927 = ((~II2917))|((~II2925));
assign WX1132 = ((~II3287))|((~II3288));
assign II10867 = ((~WX3588))|((~II10866));
assign WX11108 = (WX11045&RESET);
assign II30257 = ((~WX9902))|((~II30255));
assign WX2455 = (WX1895&WX2456);
assign II34956 = ((~II34966))|((~II34967));
assign II30967 = ((~II30969))|((~II30970));
assign II14266 = ((~WX4668))|((~WX4732));
assign II30976 = ((~II30951))|((~II30975));
assign WX1513 = (WX1511)|(WX1510);
assign II22755 = ((~II22765))|((~II22766));
assign WX7832 = (WX7830)|(WX7829);
assign WX11325 = ((~WX11324));
assign WX7525 = ((~WX7524));
assign II6057 = ((~WX1942))|((~II6055));
assign II18666 = ((~WX5923))|((~II18658));
assign II3703 = ((~WX641))|((~_2078_));
assign II3515 = ((~WX643))|((~II3514));
assign II18364 = ((~WX5967))|((~WX6031));
assign WX7694 = ((~WX7693));
assign II22208 = ((~II22198))|((~II22206));
assign II30038 = ((~WX9824))|((~WX9888));
assign WX11180 = (WX11117&RESET);
assign WX5330 = (WX5328)|(WX5327);
assign WX2237 = ((~WX2215));
assign WX8079 = ((~WX8762));
assign WX1349 = (WX1347)|(WX1346);
assign WX4299 = (WX4297)|(WX4296);
assign WX6823 = (WX6829&WX6824);
assign WX2278 = ((~WX2277));
assign WX475 = ((~WX1004));
assign II26871 = ((~WX8585))|((~II26870));
assign WX147 = (WX158&WX1003);
assign II19163 = ((~WX5759))|((~WX5671));
assign WX3094 = (WX3097&RESET);
assign WX9801 = (WX9738&RESET);
assign WX10854 = (WX10857&RESET);
assign II34229 = ((~WX11129))|((~WX11193));
assign WX7894 = (WX7892)|(WX7891);
assign II14886 = ((~WX4708))|((~WX4772));
assign WX2241 = ((~WX2217));
assign WX2753 = ((~WX3590));
assign II15500 = ((~WX4511))|((~_2204_));
assign WX7392 = ((~II22873))|((~II22874));
assign WX5598 = ((~WX5597));
assign II26878 = ((~II26853))|((~II26877));
assign II35617 = ((~WX10964))|((~_2355_));
assign WX2202 = ((~II6295))|((~II6296));
assign II19654 = ((~WX5801))|((~II19653));
assign WX6934 = (WX6945&WX7468);
assign II22027 = ((~II22029))|((~II22030));
assign WX10844 = (WX10847&RESET);
assign II10300 = ((~II10275))|((~II10299));
assign WX6545 = (WX6543)|(WX6542);
assign WX9956 = ((~II30201))|((~II30202));
assign WX9963 = ((~II30418))|((~II30419));
assign II14570 = ((~II14560))|((~II14568));
assign WX1062 = ((~II3157))|((~II3158));
assign II15484 = ((~II15486))|((~II15487));
assign II2265 = ((~II2275))|((~II2276));
assign II2346 = ((~WX859))|((~II2344));
assign WX6068 = (WX6005&RESET);
assign WX7847 = ((~WX7838));
assign WX10921 = ((~WX11303));
assign II15368 = ((~WX4410))|((~II15366));
assign WX7378 = ((~II22439))|((~II22440));
assign II31570 = ((~WX9665))|((~_2329_));
assign WX6872 = (WX7002&WX7469);
assign WX4988 = ((~WX4987));
assign WX11572 = ((~WX11571));
assign WX1665 = (WX1671&WX1666);
assign II34920 = ((~II34910))|((~II34918));
assign II19477 = ((~WX5719))|((~II19475));
assign WX5848 = (WX5444&RESET);
assign II10455 = ((~II10430))|((~II10454));
assign II31349 = ((~WX9576))|((~II31347));
assign WX7379 = ((~II22470))|((~II22471));
assign WX10427 = ((~WX11348));
assign WX8054 = (WX8896&WX8055);
assign WX4691 = (WX4628&RESET);
assign WX6406 = ((~II19535))|((~II19536));
assign II11595 = ((~WX3207))|((~II11594));
assign WX7651 = ((~WX7650));
assign WX7966 = (WX10147&WX7967);
assign II30752 = ((~WX9870))|((~II30751));
assign WX10915 = ((~WX11291));
assign WX5916 = (WX5853&RESET);
assign WX9230 = (_2322_&WX10055);
assign WX6733 = (WX7589&WX6734);
assign WX3348 = (WX3285&RESET);
assign II30998 = ((~II31000))|((~II31001));
assign II6862 = ((~WX2295))|((~II6861));
assign WX4897 = ((~WX4896));
assign WX10704 = (WX10702)|(WX10701);
assign WX2655 = ((~WX3590));
assign II10492 = ((~II10502))|((~II10503));
assign WX5096 = (WX5095&WX4884);
assign WX8194 = (WX8966&WX8195);
assign WX8835 = (WX8834&WX8763);
assign II22239 = ((~II22229))|((~II22237));
assign WX4288 = ((~WX4883));
assign II15585 = ((~WX4498))|((~_2196_));
assign WX10497 = ((~WX11348));
assign II26206 = ((~WX8415))|((~II26204));
assign WX3971 = (WX3977&WX3972);
assign II30083 = ((~II30093))|((~II30094));
assign WX4465 = ((~WX4433));
assign II26956 = ((~WX8527))|((~II26955));
assign II3620 = ((~WX626))|((~II3619));
assign WX6536 = (WX6954&WX7469);
assign WX6340 = (WX6339&WX6177);
assign II27700 = ((~_2276_))|((~II27698));
assign II18551 = ((~WX5979))|((~II18550));
assign WX744 = (WX681&RESET);
assign II6621 = ((~WX2042))|((~II6620));
assign WX1783 = (WX1786&RESET);
assign WX5962 = (WX5899&RESET);
assign WX10222 = (WX10220)|(WX10219);
assign WX8731 = ((~WX8730));
assign WX10592 = (WX10590)|(WX10589);
assign WX5091 = ((~WX4884));
assign WX1632 = ((~WX2297));
assign II14590 = ((~II14600))|((~II14601));
assign WX410 = (WX408)|(WX407);
assign WX3045 = (_2142_&WX3590);
assign WX6432 = ((~II19717))|((~II19718));
assign WX7825 = (_2298_&WX8762);
assign WX8036 = (WX10182&WX8037);
assign WX8076 = (WX8074)|(WX8073);
assign WX8090 = (WX8088)|(WX8087);
assign WX10967 = ((~WX11203));
assign WX3149 = ((~WX3581));
assign WX8033 = ((~WX8761));
assign WX6909 = (WX6907)|(WX6906);
assign WX8950 = (WX8948)|(WX8947);
assign II34138 = ((~WX11187))|((~II34136));
assign WX8598 = (WX8535&RESET);
assign II3353 = ((~WX531))|((~II3351));
assign II35576 = ((~WX10958))|((~II35575));
assign II2515 = ((~WX1002))|((~WX679));
assign WX3606 = ((~II11089))|((~II11090));
assign II22626 = ((~II22616))|((~II22624));
assign WX7602 = ((~WX7601));
assign WX10801 = ((~WX11347));
assign II2570 = ((~II2560))|((~II2568));
assign WX11034 = (WX10714&RESET);
assign II26600 = ((~II26590))|((~II26598));
assign II18681 = ((~II18657))|((~II18673));
assign WX2927 = ((~WX2918));
assign II34298 = ((~II34274))|((~II34290));
assign WX4842 = ((~WX4841));
assign WX11539 = ((~II35444))|((~II35445));
assign II22888 = ((~WX7230))|((~II22880));
assign II19306 = ((~WX5770))|((~WX5693));
assign II11560 = ((~WX3202))|((~II11559));
assign WX9400 = ((~WX10055));
assign WX2858 = ((~WX2857));
assign II14792 = ((~II14794))|((~II14795));
assign II26128 = ((~WX8601))|((~II26126));
assign II14637 = ((~II14639))|((~II14640));
assign WX9753 = (WX9505&RESET);
assign II18428 = ((~WX6035))|((~II18426));
assign WX149 = ((~WX1003));
assign II6611 = ((~II6621))|((~II6622));
assign II3377 = ((~WX605))|((~WX535));
assign WX2820 = (WX2818)|(WX2817);
assign WX4010 = ((~WX4001));
assign II30179 = ((~WX10052))|((~II30178));
assign II19098 = ((~WX5754))|((~WX5661));
assign WX2677 = (WX2688&WX3589);
assign II34439 = ((~WX11079))|((~II34438));
assign WX5788 = ((~WX6017));
assign WX2966 = (WX3766&WX2967);
assign II34649 = ((~WX11346))|((~II34648));
assign II6876 = ((~WX2122))|((~WX2186));
assign WX5269 = ((~WX6176));
assign II10509 = ((~WX3391))|((~WX3455));
assign WX2670 = (WX2668)|(WX2667);
assign II30101 = ((~WX9828))|((~II30100));
assign WX4231 = (WX5045&WX4232);
assign WX3748 = (WX3188&WX3749);
assign II22896 = ((~WX7294))|((~WX7358));
assign II11335 = ((~WX3187))|((~WX3113));
assign WX10142 = (WX10141&WX10056);
assign WX8995 = ((~II27566))|((~II27567));
assign WX9168 = ((~WX9159));
assign II26560 = ((~WX8565))|((~WX8629));
assign WX6787 = (WX6785)|(WX6784);
assign WX2940 = (WX2938)|(WX2937);
assign II2834 = ((~II2824))|((~II2832));
assign WX9739 = (WX9407&RESET);
assign WX3837 = ((~II11644))|((~II11645));
assign II2733 = ((~WX1002))|((~II2732));
assign WX2284 = ((~WX2283));
assign II19281 = ((~WX5768))|((~II19280));
assign II3677 = ((~_2083_))|((~II3675));
assign II18968 = ((~II18970))|((~II18971));
assign II18805 = ((~II18781))|((~II18797));
assign WX4896 = (WX4894)|(WX4893);
assign II27446 = ((~WX8366))|((~WX8299));
assign WX5485 = ((~WX5476));
assign II35144 = ((~WX10928))|((~WX10837));
assign WX5106 = (WX5104)|(WX5103);
assign WX6298 = (WX6297&WX6177);
assign WX6979 = (WX6982&RESET);
assign WX8209 = ((~WX8762));
assign II34198 = ((~WX11127))|((~WX11191));
assign WX463 = (WX545&WX1004);
assign II6426 = ((~II6428))|((~II6429));
assign WX9268 = (WX9279&WX10054);
assign WX1083 = ((~II3196))|((~II3197));
assign II14375 = ((~WX4880))|((~WX4548));
assign WX5203 = (WX5115&WX5142);
assign II34897 = ((~WX11346))|((~II34896));
assign WX11010 = (WX10546&RESET);
assign WX5573 = ((~WX6175));
assign WX11453 = ((~WX11452));
assign II3091 = ((~WX583))|((~WX491));
assign WX5368 = (WX5366)|(WX5365);
assign WX6760 = (WX6986&WX7469);
assign WX1098 = (WX1097&WX1005);
assign WX6965 = (WX6968&RESET);
assign II26242 = ((~WX8481))|((~II26234));
assign WX4888 = ((~WX4884));
assign II7667 = ((~WX1927))|((~II7666));
assign II26089 = ((~II26079))|((~II26087));
assign WX8154 = (WX8152)|(WX8151);
assign WX3676 = ((~II11219))|((~II11220));
assign II19497 = ((~_2220_))|((~II19489));
assign WX5690 = (WX5693&RESET);
assign WX2281 = ((~WX2205));
assign WX8773 = (WX8339&WX8774);
assign WX6264 = (WX5764&WX6265);
assign WX8103 = ((~WX8761));
assign II26987 = ((~WX8529))|((~II26986));
assign WX5257 = (WX5663&WX6176);
assign II18590 = ((~II18580))|((~II18588));
assign II35327 = ((~WX10942))|((~II35326));
assign II23596 = ((~WX7084))|((~II23595));
assign WX9492 = (WX9503&WX10054);
assign II2020 = ((~WX1001))|((~II2019));
assign WX8402 = (WX7806&RESET);
assign II27706 = ((~WX8394))|((~II27705));
assign WX3193 = ((~WX3161));
assign WX8174 = (WX8172)|(WX8171);
assign WX1611 = (WX1609)|(WX1608);
assign II22756 = ((~II22758))|((~II22759));
assign WX3506 = ((~II10641))|((~II10642));
assign WX417 = (_2081_&WX1004);
assign II18031 = ((~II18006))|((~II18030));
assign II30573 = ((~II30548))|((~II30572));
assign II18705 = ((~WX5989))|((~WX6053));
assign II6883 = ((~II6859))|((~II6875));
assign II11246 = ((~WX3099))|((~II11244));
assign WX4535 = (WX4011&RESET);
assign WX1329 = (WX1335&WX1330);
assign II3286 = ((~WX598))|((~WX521));
assign II22725 = ((~II22727))|((~II22728));
assign WX9591 = (WX9594&RESET);
assign II27636 = ((~WX8382))|((~II27635));
assign WX4928 = (WX4927&WX4884);
assign II3262 = ((~WX517))|((~II3260));
assign II26467 = ((~WX8559))|((~WX8623));
assign WX10726 = (WX10724)|(WX10723);
assign WX3660 = ((~WX3659));
assign WX1671 = (WX1669)|(WX1668);
assign WX8123 = (WX8289&WX8762);
assign II18728 = ((~WX5927))|((~II18720));
assign II14001 = ((~II14011))|((~II14012));
assign WX10208 = (WX10206)|(WX10205);
assign WX2868 = (WX3717&WX2869);
assign WX9408 = (WX9419&WX10054);
assign WX5429 = ((~WX5420));
assign II10542 = ((~WX3457))|((~II10540));
assign II27238 = ((~WX8350))|((~WX8267));
assign WX294 = (WX292)|(WX291);
assign WX2306 = ((~II7071))|((~II7072));
assign II14560 = ((~II14562))|((~II14563));
assign II6565 = ((~II6567))|((~II6568));
assign WX9158 = ((~WX10054));
assign WX2784 = (WX3675&WX2785);
assign II11465 = ((~WX3197))|((~WX3133));
assign WX5930 = (WX5867&RESET);
assign II14600 = ((~WX4626))|((~II14599));
assign II2183 = ((~II2173))|((~II2181));
assign WX9624 = ((~WX10002));
assign WX10217 = ((~WX10216));
assign WX2861 = ((~WX3589));
assign WX11580 = ((~II35569))|((~II35570));
assign II10238 = ((~II10213))|((~II10237));
assign WX760 = (WX697&RESET);
assign WX2516 = ((~II7461))|((~II7462));
assign WX4170 = (_2186_&WX4883);
assign WX1211 = (WX609&WX1212);
assign II35723 = ((~WX10981))|((~II35722));
assign WX5580 = (WX6366&WX5581);
assign WX5483 = ((~WX6176));
assign WX9970 = ((~II30635))|((~II30636));
assign WX11498 = (WX11497&WX11349);
assign WX11348 = ((~WX11341));
assign WX5672 = (WX5675&RESET);
assign II34863 = ((~II34873))|((~II34874));
assign WX8714 = ((~WX8686));
assign WX4875 = ((~TM0));
assign DATA_9_29 = ((~WX1025));
assign II18643 = ((~WX5985))|((~WX6049));
assign WX10268 = (WX10267&WX10056);
assign WX9638 = ((~WX9606));
assign II10307 = ((~II10309))|((~II10310));
assign II22664 = ((~WX7467))|((~WX7152));
assign WX524 = (WX527&RESET);
assign WX5324 = (WX7533&WX5325);
assign WX3631 = (WX3629)|(WX3628);
assign WX8800 = (WX8799&WX8763);
assign WX1143 = (WX1141)|(WX1140);
assign II6257 = ((~WX2082))|((~II6256));
assign II15406 = ((~WX4485))|((~II15405));
assign WX10037 = ((~WX9962));
assign II27175 = ((~WX8257))|((~II27173));
assign II2687 = ((~WX881))|((~II2685));
assign WX8694 = ((~WX8676));
assign WX9210 = ((~WX9201));
assign II19358 = ((~WX5774))|((~WX5701));
assign WX5306 = (WX5312&WX5307);
assign WX4220 = ((~WX4211));
assign WX6189 = (WX6187)|(WX6186);
assign WX319 = (_2088_&WX1004);
assign II26577 = ((~WX8760))|((~II26576));
assign II14004 = ((~WX4880))|((~II14003));
assign WX10030 = ((~WX10029));
assign II3711 = ((~WX642))|((~II3710));
assign II22972 = ((~II22982))|((~II22983));
assign II6294 = ((~II6270))|((~II6286));
assign WX6324 = ((~WX6323));
assign WX5506 = (WX7624&WX5507);
assign II23312 = ((~WX7063))|((~II23311));
assign WX5658 = (WX5661&RESET);
assign II22585 = ((~II22587))|((~II22588));
assign WX246 = (WX252&WX247);
assign WX10165 = ((~WX10056));
assign WX427 = (WX438&WX1003);
assign WX9831 = (WX9768&RESET);
assign II14911 = ((~II14901))|((~II14909));
assign WX3673 = (WX3671)|(WX3670);
assign WX10070 = ((~WX10069));
assign II6015 = ((~II5991))|((~II6007));
assign II23468 = ((~WX7075))|((~II23467));
assign II23567 = ((~WX7080))|((~_2264_));
assign WX10077 = ((~WX10076));
assign II14180 = ((~II14156))|((~II14172));
assign WX4486 = ((~WX4454));
assign WX2103 = (WX2040&RESET);
assign WX6286 = ((~WX6177));
assign II15699 = ((~_2178_))|((~II15697));
assign II22386 = ((~WX7466))|((~II22385));
assign WX6301 = (WX6299)|(WX6298);
assign WX1626 = (_2119_&WX2297);
assign II26623 = ((~WX8569))|((~II26622));
assign WX6743 = (WX8889&WX6744);
assign WX5066 = ((~WX5065));
assign II15537 = ((~WX4491))|((~II15536));
assign WX8701 = ((~WX8700));
assign WX11518 = ((~II35405))|((~II35406));
assign WX4503 = ((~WX4740));
assign WX662 = (WX174&RESET);
assign WX4168 = ((~WX4882));
assign WX4136 = ((~WX4127));
assign WX4056 = ((~WX4882));
assign WX8666 = ((~II26289))|((~II26290));
assign II30666 = ((~II30641))|((~II30665));
assign II23707 = ((~WX7102))|((~_2242_));
assign WX7407 = ((~WX7386));
assign WX9190 = ((~WX10055));
assign II26158 = ((~WX8539))|((~II26157));
assign II14630 = ((~WX4628))|((~II14622));
assign WX5884 = (WX5821&RESET);
assign II10796 = ((~II10771))|((~II10795));
assign II10299 = ((~II10275))|((~II10291));
assign WX2662 = ((~WX2661));
assign WX7447 = ((~WX7374));
assign II15316 = ((~WX4402))|((~II15314));
assign WX5420 = (WX5418)|(WX5417);
assign WX492 = (WX495&RESET);
assign II18357 = ((~WX5903))|((~II18356));
assign WX3944 = ((~WX4882));
assign WX7145 = (WX6765&RESET);
assign WX8399 = ((~WX8653));
assign II19373 = ((~WX5703))|((~II19371));
assign WX2771 = ((~WX3590));
assign II14165 = ((~WX4598))|((~II14157));
assign WX10261 = (WX10260&WX10056);
assign II26530 = ((~WX8563))|((~II26529));
assign WX3230 = (WX2634&RESET);
assign II34184 = ((~WX11345))|((~II34183));
assign WX11379 = (WX11378&WX11349);
assign II26326 = ((~II26336))|((~II26337));
assign WX6841 = (WX8938&WX6842);
assign WX8757 = ((~TM1));
assign WX10413 = ((~WX11348));
assign WX2985 = (WX2996&WX3589);
assign WX8274 = (WX8277&RESET);
assign WX2165 = (WX2102&RESET);
assign WX11098 = (WX11035&RESET);
assign WX10246 = ((~II31439))|((~II31440));
assign WX8707 = ((~WX8706));
assign II27212 = ((~WX8348))|((~WX8263));
assign WX9995 = ((~WX9973));
assign WX406 = (WX404)|(WX403);
assign II19527 = ((~_2208_))|((~II19519));
assign WX2372 = ((~WX2298));
assign II26119 = ((~WX8473))|((~II26118));
assign WX3788 = ((~II11427))|((~II11428));
assign WX5405 = ((~WX6175));
assign WX4128 = (_2189_&WX4883);
assign WX5584 = ((~WX5583));
assign WX9717 = (WX9253&RESET);
assign II18387 = ((~WX5905))|((~II18379));
assign II2299 = ((~WX1001))|((~II2298));
assign WX7079 = ((~WX7306));
assign WX10131 = (WX10129)|(WX10128);
assign II34889 = ((~II34879))|((~II34887));
assign WX9449 = ((~WX9448));
assign WX4179 = ((~WX4178));
assign II27502 = ((~_2300_))|((~II27500));
assign WX8642 = (WX8579&RESET);
assign WX9516 = ((~WX10055));
assign II2190 = ((~WX785))|((~II2189));
assign WX5720 = ((~WX6137));
assign II26569 = ((~II26559))|((~II26567));
assign WX1608 = (WX1619&WX2296);
assign II22232 = ((~WX7124))|((~II22230));
assign II18816 = ((~WX5869))|((~II18814));
assign WX9901 = (WX9838&RESET);
assign WX6865 = (WX6871&WX6866);
assign II22067 = ((~II22042))|((~II22066));
assign WX4437 = ((~WX4864));
assign II34944 = ((~WX11239))|((~II34942));
assign II22927 = ((~WX7296))|((~WX7360));
assign II18294 = ((~WX5899))|((~II18286));
assign II10751 = ((~II10741))|((~II10749));
assign WX9149 = (WX9147)|(WX9146);
assign WX365 = (WX531&WX1004);
assign II26562 = ((~WX8629))|((~II26560));
assign WX10307 = ((~II31704))|((~II31705));
assign WX11433 = ((~WX11432));
assign WX5828 = (WX5304&RESET);
assign WX3374 = (WX3311&RESET);
assign II22828 = ((~II22818))|((~II22826));
assign II14430 = ((~II14420))|((~II14428));
assign II35248 = ((~WX10936))|((~WX10853));
assign WX9469 = (WX11545&WX9470);
assign II31628 = ((~_2321_))|((~II31626));
assign II14607 = ((~WX4690))|((~WX4754));
assign II34888 = ((~II34863))|((~II34887));
assign II31321 = ((~WX9649))|((~WX9572));
assign II19242 = ((~WX5765))|((~II19241));
assign II11309 = ((~WX3185))|((~WX3109));
assign WX9285 = (WX9283)|(WX9282);
assign II30844 = ((~WX9876))|((~WX9940));
assign II27622 = ((~WX8380))|((~II27621));
assign II26344 = ((~WX8551))|((~II26343));
assign WX2953 = ((~WX3590));
assign WX9297 = (WX9303&WX9298);
assign WX3560 = ((~WX3491));
assign II34727 = ((~WX11225))|((~II34725));
assign II6109 = ((~II6084))|((~II6108));
assign WX7109 = (WX6513&RESET);
assign WX7927 = (WX8261&WX8762);
assign II35430 = ((~WX10950))|((~WX10881));
assign WX3757 = (WX3755)|(WX3754);
assign WX1024 = (WX1022)|(WX1021);
assign II30056 = ((~WX9698))|((~II30054));
assign II3197 = ((~WX507))|((~II3195));
assign WX11382 = (WX11380)|(WX11379);
assign II22910 = ((~II22920))|((~II22921));
assign WX2382 = ((~WX2381));
assign WX3102 = (WX3105&RESET);
assign II10510 = ((~WX3391))|((~II10509));
assign WX3324 = (WX3261&RESET);
assign II19137 = ((~WX5757))|((~WX5667));
assign WX7613 = (WX7065&WX7614);
assign WX2740 = (WX2738)|(WX2737);
assign II26585 = ((~II26575))|((~II26583));
assign II10447 = ((~WX3387))|((~WX3451));
assign WX8791 = ((~WX8790));
assign WX2432 = ((~II7305))|((~II7306));
assign II26810 = ((~WX8645))|((~II26808));
assign II27721 = ((~_2273_))|((~II27719));
assign II30355 = ((~II30331))|((~II30347));
assign WX5458 = ((~WX5457));
assign WX11523 = ((~WX11522));
assign II30552 = ((~WX9730))|((~II30550));
assign II26450 = ((~II26460))|((~II26461));
assign II11140 = ((~WX3172))|((~WX3083));
assign WX350 = (WX348)|(WX347);
assign II31703 = ((~WX9686))|((~_2308_));
assign II7646 = ((~WX1923))|((~II7645));
assign WX10562 = (WX10568&WX10563);
assign WX3210 = ((~WX3447));
assign WX2827 = ((~WX3590));
assign WX1655 = (WX3759&WX1656);
assign II31612 = ((~WX9671))|((~_2323_));
assign II6387 = ((~II6363))|((~II6379));
assign WX9817 = (WX9754&RESET);
assign WX3779 = ((~WX3778));
assign WX2878 = (WX5017&WX2879);
assign II19541 = ((~WX5784))|((~_2235_));
assign WX92 = (WX98&WX93);
assign WX7763 = (WX7714&WX7728);
assign II22269 = ((~WX7190))|((~II22268));
assign II14652 = ((~II14662))|((~II14663));
assign WX2499 = (WX2497)|(WX2496);
assign II15341 = ((~WX4480))|((~II15340));
assign WX6900 = (WX7006&WX7469);
assign WX3651 = ((~WX3591));
assign II22618 = ((~WX7276))|((~II22617));
assign WX3139 = ((~WX3561));
assign II22611 = ((~II22601))|((~II22609));
assign WX1949 = (WX1425&RESET);
assign WX3923 = (WX4891&WX3924);
assign II34640 = ((~II34615))|((~II34639));
assign WX4496 = ((~WX4726));
assign II6466 = ((~WX2032))|((~II6465));
assign WX6836 = (WX6847&WX7468);
assign WX3692 = (WX3180&WX3693);
assign II10774 = ((~WX3588))|((~II10773));
assign WX7589 = ((~WX7588));
assign WX5789 = ((~WX6019));
assign WX9799 = (WX9736&RESET);
assign II27226 = ((~WX8349))|((~II27225));
assign WX1046 = ((~WX1045));
assign WX86 = (DATA_9_28&WX87);
assign WX8763 = ((~WX8754));
assign WX10944 = ((~WX10912));
assign WX2440 = (WX2439&WX2298);
assign II19702 = ((~WX5809))|((~_2210_));
assign II22858 = ((~WX7228))|((~II22857));
assign II2904 = ((~WX895))|((~II2902));
assign II23617 = ((~WX7087))|((~II23616));
assign WX275 = ((~WX1003));
assign WX2468 = (WX2467&WX2298);
assign II18828 = ((~II18830))|((~II18831));
assign WX63 = (WX74&WX1003);
assign II10114 = ((~II10089))|((~II10113));
assign WX11442 = (WX11441&WX11349);
assign WX5664 = (WX5667&RESET);
assign WX5386 = (WX5384)|(WX5383);
assign II27509 = ((~II27499))|((~II27507));
assign WX7438 = ((~WX7437));
assign II26678 = ((~II26668))|((~II26676));
assign WX9203 = (WX11412&WX9204);
assign WX582 = ((~WX550));
assign WX9977 = ((~II30852))|((~II30853));
assign WX5398 = (WX6275&WX5399);
assign II26722 = ((~II26698))|((~II26714));
assign II2973 = ((~II2963))|((~II2971));
assign II23527 = ((~_2268_))|((~II23525));
assign WX5782 = ((~WX5750));
assign WX4125 = (WX4131&WX4126);
assign II2632 = ((~II2622))|((~II2630));
assign WX11437 = ((~WX11349));
assign II34615 = ((~II34625))|((~II34626));
assign II18164 = ((~WX6173))|((~II18163));
assign II10663 = ((~II10665))|((~II10666));
assign WX5220 = ((~WX5219));
assign WX7432 = ((~WX7431));
assign II2965 = ((~WX835))|((~II2964));
assign WX1200 = ((~WX1199));
assign WX194 = (WX2382&WX195);
assign II23352 = ((~WX6992))|((~II23350));
assign II19177 = ((~WX5760))|((~II19176));
assign WX5415 = ((~WX5406));
assign WX352 = (DATA_9_9&WX353);
assign WX7534 = ((~II23195))|((~II23196));
assign II6172 = ((~II6162))|((~II6170));
assign WX10582 = (WX10580)|(WX10579);
assign WX5177 = (WX5128&WX5142);
assign WX4078 = ((~WX4883));
assign WX7567 = ((~WX7566));
assign II22262 = ((~WX7466))|((~II22261));
assign WX10823 = ((~WX11348));
assign WX10607 = (_2348_&WX11348);
assign II34322 = ((~WX11135))|((~WX11199));
assign II3500 = ((~WX639))|((~_2108_));
assign WX11341 = ((~TM0));
assign WX11134 = (WX11071&RESET);
assign II22414 = ((~II22424))|((~II22425));
assign WX10933 = ((~WX10901));
assign II22020 = ((~WX7174))|((~II22012));
assign WX3517 = ((~II10982))|((~II10983));
assign WX960 = ((~WX930));
assign II2701 = ((~WX1002))|((~WX691));
assign WX7094 = ((~WX7336));
assign WX9769 = (WX9706&RESET);
assign WX6398 = ((~WX6177));
assign WX7366 = ((~II22067))|((~II22068));
assign WX1154 = (WX1153&WX1005);
assign WX5131 = ((~II15656))|((~II15657));
assign WX573 = ((~WX951));
assign II14188 = ((~II14190))|((~II14191));
assign WX4948 = ((~II15185))|((~II15186));
assign II22167 = ((~II22169))|((~II22170));
assign WX8880 = (WX8878)|(WX8877);
assign II22456 = ((~II22446))|((~II22454));
assign WX6808 = (WX6819&WX7468);
assign II22835 = ((~WX7290))|((~II22834));
assign II6759 = ((~II6735))|((~II6751));
assign WX2871 = ((~WX2862));
assign WX1971 = (WX1579&RESET);
assign WX4419 = (WX4422&RESET);
assign WX6180 = (WX5752&WX6181);
assign II31413 = ((~WX9656))|((~II31412));
assign WX10637 = ((~WX11348));
assign WX10717 = ((~WX11347));
assign WX8874 = ((~WX8873));
assign WX5532 = (WX5530)|(WX5529);
assign II35235 = ((~WX10935))|((~WX10851));
assign II6760 = ((~II6735))|((~II6759));
assign II6503 = ((~II6505))|((~II6506));
assign WX8658 = ((~II26041))|((~II26042));
assign WX2605 = (WX2535&WX2556);
assign WX6278 = (WX5766&WX6279);
assign II6844 = ((~II6846))|((~II6847));
assign WX3709 = ((~WX3708));
assign WX10375 = (WX10287&WX10314);
assign II6100 = ((~II6102))|((~II6103));
assign WX1742 = (WX1836&WX2297);
assign II22997 = ((~II22972))|((~II22996));
assign II31656 = ((~_2317_))|((~II31654));
assign WX55 = ((~WX1004));
assign WX299 = ((~WX290));
assign WX10024 = ((~WX10023));
assign II7591 = ((~_2130_))|((~II7589));
assign WX188 = ((~WX187));
assign II23105 = ((~WX6954))|((~II23103));
assign WX10710 = (WX11517&WX10711);
assign WX6220 = ((~II19151))|((~II19152));
assign WX9725 = (WX9309&RESET);
assign WX9247 = (WX9245)|(WX9244);
assign WX2065 = (WX2002&RESET);
assign II34277 = ((~WX11345))|((~II34276));
assign WX5730 = ((~WX6157));
assign II7175 = ((~WX1882))|((~II7174));
assign II10595 = ((~WX3333))|((~II10594));
assign WX223 = ((~WX1004));
assign WX1721 = (WX1727&WX1722);
assign WX9151 = (WX10091&WX9152);
assign II22974 = ((~WX7467))|((~WX7172));
assign II23416 = ((~WX7071))|((~II23415));
assign II14811 = ((~WX4576))|((~II14809));
assign WX11238 = (WX11175&RESET);
assign WX181 = ((~WX1004));
assign II19499 = ((~II19489))|((~II19497));
assign WX2047 = (WX1984&RESET);
assign WX3698 = (WX3697&WX3591);
assign WX8125 = ((~WX8762));
assign II30132 = ((~WX9830))|((~II30131));
assign WX9253 = ((~WX9252));
assign WX2475 = (WX2474&WX2298);
assign II34329 = ((~II34305))|((~II34321));
assign WX11602 = ((~II35723))|((~II35724));
assign WX3250 = (WX2774&RESET);
assign WX9175 = (WX11398&WX9176);
assign WX5126 = ((~II15621))|((~II15622));
assign WX3766 = ((~WX3765));
assign WX8013 = ((~WX8762));
assign WX1755 = (WX1753)|(WX1752);
assign II15119 = ((~WX4463))|((~WX4372));
assign WX8952 = ((~WX8951));
assign WX72 = (DATA_9_29&WX73);
assign WX6501 = (WX6507&WX6502);
assign WX4163 = (WX4161)|(WX4160);
assign WX7287 = (WX7224&RESET);
assign II6831 = ((~WX2295))|((~II6830));
assign II34331 = ((~II34321))|((~II34329));
assign II30403 = ((~WX9784))|((~II30402));
assign WX2483 = (WX1899&WX2484);
assign WX4083 = (WX4089&WX4084);
assign WX8959 = ((~WX8958));
assign WX9244 = (_2321_&WX10055);
assign WX5539 = ((~WX6176));
assign WX494 = (WX497&RESET);
assign WX3898 = (WX3828&WX3849);
assign II2878 = ((~II2854))|((~II2870));
assign WX1292 = (WX1251&WX1263);
assign WX5221 = (WX5232&WX6175);
assign II2723 = ((~II2699))|((~II2715));
assign WX993 = ((~WX992));
assign WX6239 = ((~WX6238));
assign II22409 = ((~II22399))|((~II22407));
assign II6721 = ((~WX2112))|((~WX2176));
assign WX6548 = ((~WX7469));
assign WX8173 = ((~WX8761));
assign II6026 = ((~WX1940))|((~II6024));
assign WX10626 = (WX11475&WX10627);
assign WX8492 = (WX8429&RESET);
assign WX1937 = (WX1341&RESET);
assign II22779 = ((~II22755))|((~II22771));
assign II10937 = ((~II10927))|((~II10935));
assign WX2396 = ((~WX2395));
assign WX7644 = ((~WX7643));
assign WX4958 = ((~WX4884));
assign II23391 = ((~WX6998))|((~II23389));
assign WX3503 = ((~II10548))|((~II10549));
assign II18041 = ((~WX5819))|((~II18039));
assign WX6458 = (WX6404&WX6435);
assign WX7916 = (WX7914)|(WX7913);
assign WX10353 = (WX10298&WX10314);
assign II15366 = ((~WX4482))|((~WX4410));
assign WX151 = (_2100_&WX1004);
assign II31627 = ((~WX9673))|((~II31626));
assign WX8117 = ((~WX8761));
assign WX4790 = ((~II14367))|((~II14368));
assign II3210 = ((~WX509))|((~II3208));
assign WX10468 = (DATA_0_25&WX10469);
assign WX4337 = (WX4335)|(WX4334);
assign WX5444 = ((~WX5443));
assign WX269 = ((~WX1004));
assign WX5762 = ((~WX5730));
assign WX7297 = (WX7234&RESET);
assign II6332 = ((~II6342))|((~II6343));
assign WX3646 = ((~WX3645));
assign II7645 = ((~WX1923))|((~_2121_));
assign II34262 = ((~WX11195))|((~II34260));
assign WX10617 = (WX10628&WX11347);
assign II3536 = ((~WX614))|((~II3535));
assign WX10768 = (WX10766)|(WX10765);
assign WX8164 = (WX8162)|(WX8161);
assign WX6132 = ((~WX6102));
assign WX8746 = ((~WX8670));
assign WX1511 = (WX1517&WX1512);
assign II30838 = ((~II30828))|((~II30836));
assign II34075 = ((~WX11119))|((~II34074));
assign WX3168 = ((~WX3136));
assign WX7426 = ((~WX7425));
assign WX6676 = (WX6974&WX7469);
assign WX9787 = (WX9724&RESET);
assign WX7049 = ((~WX7017));
assign II26661 = ((~II26636))|((~II26660));
assign II6239 = ((~II6249))|((~II6250));
assign WX1127 = (WX597&WX1128);
assign WX1356 = (WX1367&WX2296);
assign II22035 = ((~II22011))|((~II22027));
assign WX8857 = (WX8351&WX8858);
assign WX2325 = ((~WX2324));
assign WX5137 = ((~II15698))|((~II15699));
assign WX9749 = (WX9477&RESET);
assign II22603 = ((~WX7467))|((~II22602));
assign WX4645 = (WX4582&RESET);
assign WX1239 = ((~II3550))|((~II3551));
assign WX2225 = ((~WX2209));
assign WX7557 = (WX7057&WX7558);
assign WX9338 = (WX9349&WX10054);
assign II31231 = ((~WX9642))|((~II31230));
assign II35365 = ((~WX10945))|((~WX10871));
assign II26360 = ((~WX8759))|((~II26359));
assign II26514 = ((~WX8760))|((~WX8435));
assign II26095 = ((~WX8535))|((~WX8599));
assign II34702 = ((~II34677))|((~II34701));
assign WX8454 = (WX8170&RESET);
assign WX798 = (WX735&RESET);
assign II26567 = ((~II26543))|((~II26559));
assign WX10694 = (WX10692)|(WX10691);
assign II34657 = ((~II34647))|((~II34655));
assign II11192 = ((~WX3176))|((~WX3091));
assign II2568 = ((~II2544))|((~II2560));
assign WX1306 = (WX1245&WX1263);
assign WX11530 = ((~WX11529));
assign WX4862 = ((~WX4861));
assign WX6171 = ((~TM1));
assign WX5218 = (WX5216)|(WX5215);
assign II11374 = ((~WX3190))|((~WX3119));
assign II6024 = ((~WX2294))|((~WX1940));
assign WX10719 = (_2340_&WX11348);
assign II11310 = ((~WX3185))|((~II11309));
assign WX11082 = (WX11019&RESET);
assign WX1926 = ((~WX2172));
assign II2251 = ((~WX789))|((~WX853));
assign WX3118 = (WX3121&RESET);
assign WX8262 = (WX8265&RESET);
assign WX9295 = ((~WX9294));
assign II15594 = ((~_2195_))|((~II15592));
assign WX8989 = ((~II27508))|((~II27509));
assign WX6556 = (WX6567&WX7468);
assign WX2851 = ((~WX3590));
assign WX10664 = (DATA_0_11&WX10665);
assign WX11024 = (WX10644&RESET);
assign WX4090 = (WX4388&WX4883);
assign II30720 = ((~WX9868))|((~WX9932));
assign WX6372 = ((~WX6371));
assign WX5936 = (WX5873&RESET);
assign II26414 = ((~II26404))|((~II26412));
assign WX4699 = (WX4636&RESET);
assign WX11373 = (WX10927&WX11374);
assign WX7666 = ((~WX7665));
assign II14454 = ((~WX4744))|((~II14452));
assign WX2554 = ((~II7709))|((~II7710));
assign WX866 = (WX803&RESET);
assign WX9275 = (WX9273)|(WX9272);
assign WX217 = (WX228&WX1003);
assign II35646 = ((~WX10968))|((~II35645));
assign WX11466 = (WX11464)|(WX11463);
assign WX4045 = (WX6247&WX4046);
assign II26949 = ((~WX8760))|((~II26948));
assign II2848 = ((~II2823))|((~II2847));
assign WX11363 = ((~WX11362));
assign II26652 = ((~II26654))|((~II26655));
assign II18937 = ((~II18939))|((~II18940));
assign WX11537 = ((~WX11536));
assign WX8051 = ((~WX8762));
assign WX11505 = (WX11504&WX11349);
assign II3144 = ((~WX587))|((~II3143));
assign WX9777 = (WX9714&RESET);
assign WX1412 = (WX1423&WX2296);
assign WX2789 = (WX2800&WX3589);
assign II10781 = ((~WX3345))|((~II10780));
assign WX7419 = ((~WX7392));
assign II18466 = ((~II18456))|((~II18464));
assign WX8227 = (WX8238&WX8761);
assign II34711 = ((~WX11346))|((~II34710));
assign II26964 = ((~WX8591))|((~II26963));
assign DATA_9_11 = ((~WX1151));
assign WX9767 = (WX9704&RESET);
assign WX10395 = ((~WX11347));
assign II26188 = ((~WX8541))|((~WX8605));
assign WX10712 = (WX10710)|(WX10709);
assign WX9318 = (WX9568&WX10055);
assign WX1546 = (WX1808&WX2297);
assign WX5391 = ((~WX6175));
assign WX2532 = ((~II7555))|((~II7556));
assign WX10982 = ((~WX11233));
assign II14218 = ((~II14228))|((~II14229));
assign WX8947 = (WX8946&WX8763);
assign WX9551 = (WX9554&RESET);
assign WX4474 = ((~WX4442));
assign WX11368 = (WX11366)|(WX11365);
assign WX6283 = ((~II19268))|((~II19269));
assign II11062 = ((~WX3166))|((~WX3071));
assign II6071 = ((~WX2070))|((~II6070));
assign WX4353 = (WX6401&WX4354);
assign II18899 = ((~II18874))|((~II18898));
assign WX6806 = ((~WX6797));
assign II3429 = ((~WX609))|((~WX543));
assign WX2313 = ((~II7084))|((~II7085));
assign II34910 = ((~II34912))|((~II34913));
assign II10362 = ((~II10337))|((~II10361));
assign WX11393 = (WX11392&WX11349);
assign II26730 = ((~II26732))|((~II26733));
assign WX9657 = ((~WX9625));
assign II14056 = ((~II14032))|((~II14048));
assign II34361 = ((~II34336))|((~II34360));
assign II18991 = ((~II18967))|((~II18983));
assign II18022 = ((~II18024))|((~II18025));
assign II3079 = ((~WX582))|((~II3078));
assign II22418 = ((~WX7136))|((~II22416));
assign II2289 = ((~II2265))|((~II2281));
assign WX4020 = (WX4378&WX4883);
assign WX2842 = (WX2840)|(WX2839);
assign II15494 = ((~II15484))|((~II15492));
assign II3543 = ((~WX615))|((~II3542));
assign WX4851 = ((~WX4783));
assign WX10481 = (_2357_&WX11348);
assign WX8137 = (WX8291&WX8762);
assign WX9387 = (WX9385)|(WX9384);
assign WX1429 = (WX1427)|(WX1426);
assign WX7084 = ((~WX7316));
assign WX4161 = (WX5010&WX4162);
assign WX5567 = ((~WX6176));
assign II6084 = ((~II6094))|((~II6095));
assign II31361 = ((~WX9652))|((~II31360));
assign II18985 = ((~WX6007))|((~II18984));
assign WX6794 = (WX6805&WX7468);
assign WX7918 = ((~WX7917));
assign II30171 = ((~II30161))|((~II30169));
assign II22425 = ((~II22415))|((~II22423));
assign WX4225 = (WX4223)|(WX4222);
assign WX6308 = (WX6306)|(WX6305);
assign WX8004 = (WX8010&WX8005);
assign II10688 = ((~WX3339))|((~II10687));
assign WX4615 = (WX4552&RESET);
assign II2010 = ((~II1986))|((~II2002));
assign WX5490 = (WX5488)|(WX5487);
assign WX7047 = ((~WX7015));
assign WX1247 = ((~II3606))|((~II3607));
assign II15068 = ((~WX4459))|((~II15067));
assign WX5051 = ((~WX5050));
assign II3156 = ((~WX588))|((~WX501));
assign WX1561 = (WX2417&WX1562);
assign II15121 = ((~WX4372))|((~II15119));
assign WX7860 = (WX7858)|(WX7857);
assign WX7121 = (WX6597&RESET);
assign WX3809 = ((~II11466))|((~II11467));
assign WX3590 = ((~WX3583));
assign II18347 = ((~II18357))|((~II18358));
assign II2258 = ((~II2234))|((~II2250));
assign WX1660 = ((~WX2297));
assign WX678 = (WX286&RESET);
assign WX10160 = ((~WX10159));
assign WX2351 = ((~WX2298));
assign WX10262 = (WX9660&WX10263);
assign WX5432 = (WX5438&WX5433);
assign II23709 = ((~_2242_))|((~II23707));
assign WX4931 = (WX4929)|(WX4928);
assign WX4520 = ((~WX4774));
assign WX5712 = (WX5715&RESET);
assign II26846 = ((~II26822))|((~II26838));
assign WX2763 = ((~WX3589));
assign WX5716 = (WX5719&RESET);
assign II10641 = ((~II10616))|((~II10640));
assign WX1552 = (WX1563&WX2296);
assign II14718 = ((~WX4570))|((~II14716));
assign WX5948 = (WX5885&RESET);
assign WX2269 = ((~WX2199));
assign WX2210 = ((~II6543))|((~II6544));
assign II14205 = ((~WX4664))|((~II14204));
assign WX3644 = ((~WX3591));
assign II27474 = ((~WX8303))|((~II27472));
assign II27305 = ((~WX8277))|((~II27303));
assign WX1991 = (WX1719&RESET);
assign WX11042 = (WX10770&RESET);
assign II26919 = ((~WX8461))|((~II26917));
assign II15649 = ((~WX4508))|((~II15648));
assign II14191 = ((~WX4536))|((~II14189));
assign II27658 = ((~_2283_))|((~II27656));
assign WX1674 = ((~WX2297));
assign II18210 = ((~WX5957))|((~II18209));
assign II18178 = ((~WX5955))|((~WX6019));
assign II31661 = ((~WX9679))|((~_2315_));
assign II11680 = ((~_2148_))|((~II11678));
assign WX7410 = ((~WX7409));
assign WX8115 = (WX8126&WX8761);
assign WX10017 = ((~WX9952));
assign II30366 = ((~WX9718))|((~II30364));
assign WX3794 = ((~WX3793));
assign WX7385 = ((~II22656))|((~II22657));
assign II10260 = ((~II10262))|((~II10263));
assign WX4119 = (WX4989&WX4120);
assign WX5852 = (WX5472&RESET);
assign WX5023 = ((~WX5022));
assign II7202 = ((~WX1800))|((~II7200));
assign WX3232 = (WX2648&RESET);
assign WX8740 = ((~WX8667));
assign II2445 = ((~II2420))|((~II2444));
assign WX2009 = (WX1946&RESET);
assign WX8100 = ((~WX8099));
assign II30224 = ((~WX9836))|((~WX9900));
assign II15515 = ((~WX4518))|((~_2204_));
assign WX8329 = ((~WX8705));
assign WX3048 = (WX3046)|(WX3045);
assign II6597 = ((~WX2104))|((~WX2168));
assign II6150 = ((~WX1948))|((~II6148));
assign WX7953 = ((~WX8762));
assign II23287 = ((~WX6982))|((~II23285));
assign WX4559 = (WX4179&RESET);
assign WX5379 = (_2224_&WX6176);
assign II14477 = ((~II14467))|((~II14475));
assign WX682 = (WX314&RESET);
assign WX9502 = ((~WX10055));
assign II35482 = ((~WX10954))|((~WX10889));
assign WX9002 = ((~II27615))|((~II27616));
assign WX609 = ((~WX577));
assign WX10791 = ((~WX11348));
assign WX10236 = (WX10234)|(WX10233);
assign II35668 = ((~_2347_))|((~II35666));
assign WX5201 = (WX5116&WX5142);
assign WX1218 = (WX610&WX1219);
assign WX5748 = ((~WX6129));
assign WX10174 = ((~WX10173));
assign II10517 = ((~II10492))|((~II10516));
assign WX641 = ((~WX895));
assign WX5354 = (WX5352)|(WX5351);
assign WX8534 = (WX8471&RESET);
assign WX6572 = ((~WX7468));
assign II18434 = ((~II18409))|((~II18433));
assign WX9380 = (WX9391&WX10054);
assign WX1684 = ((~WX2297));
assign II26515 = ((~WX8760))|((~II26514));
assign WX10900 = ((~WX11325));
assign WX7793 = (WX7804&WX8761);
assign WX9048 = (WX9010&WX9021);
assign II2506 = ((~II2482))|((~II2498));
assign II14746 = ((~II14748))|((~II14749));
assign WX4719 = (WX4656&RESET);
assign WX3501 = ((~II10486))|((~II10487));
assign II3171 = ((~WX503))|((~II3169));
assign WX1304 = (WX1246&WX1263);
assign WX8739 = ((~WX8738));
assign WX6898 = ((~WX7469));
assign II34315 = ((~WX11071))|((~II34314));
assign II26748 = ((~WX8641))|((~II26746));
assign II7694 = ((~WX1931))|((~_2113_));
assign WX8972 = ((~WX8971));
assign WX3933 = (WX6191&WX3934);
assign II34107 = ((~WX11185))|((~II34105));
assign WX6085 = ((~II18434))|((~II18435));
assign WX7552 = (WX7550)|(WX7549);
assign II15210 = ((~WX4470))|((~WX4386));
assign WX9092 = ((~WX10055));
assign II19718 = ((~_2207_))|((~II19716));
assign WX5666 = (WX5669&RESET);
assign WX3174 = ((~WX3142));
assign WX1595 = (WX1601&WX1596);
assign WX11411 = ((~WX11410));
assign WX3398 = (WX3335&RESET);
assign WX1268 = (WX1261&WX1263);
assign WX8343 = ((~WX8311));
assign WX480 = (WX478)|(WX477);
assign II10378 = ((~WX3319))|((~II10377));
assign WX10107 = (WX10106&WX10056);
assign II6847 = ((~WX2184))|((~II6845));
assign WX7705 = ((~II23582))|((~II23583));
assign WX4320 = (WX4331&WX4882);
assign WX10630 = ((~WX10629));
assign WX4183 = (WX4181)|(WX4180);
assign II10837 = ((~WX3285))|((~II10835));
assign II7343 = ((~WX1895))|((~WX1822));
assign WX7658 = ((~WX7657));
assign WX4027 = (WX4033&WX4028);
assign WX8802 = ((~WX8763));
assign WX94 = (WX92)|(WX91);
assign WX4073 = (WX6261&WX4074);
assign WX2219 = ((~II6822))|((~II6823));
assign WX9881 = (WX9818&RESET);
assign II30195 = ((~WX9898))|((~II30193));
assign II2172 = ((~II2182))|((~II2183));
assign WX7058 = ((~WX7026));
assign II6916 = ((~II6906))|((~II6914));
assign WX457 = ((~WX1003));
assign II6394 = ((~II6404))|((~II6405));
assign WX8416 = (WX7904&RESET);
assign WX8181 = ((~WX8762));
assign WX2343 = (WX1879&WX2344);
assign II31621 = ((~_2322_))|((~II31619));
assign WX6088 = ((~II18527))|((~II18528));
assign WX7384 = ((~II22625))|((~II22626));
assign WX70 = (WX68)|(WX67);
assign WX2684 = (WX2682)|(WX2681);
assign WX127 = (WX497&WX1004);
assign WX79 = ((~WX1003));
assign WX9376 = ((~WX10055));
assign WX376 = (WX2473&WX377);
assign WX5807 = ((~WX6055));
assign WX10501 = ((~WX11348));
assign WX6588 = (_2262_&WX7469);
assign II15093 = ((~WX4461))|((~WX4368));
assign WX9167 = (WX9165)|(WX9164);
assign II18722 = ((~WX6174))|((~II18721));
assign WX1606 = ((~WX1597));
assign WX5304 = ((~WX5303));
assign WX3490 = ((~II10145))|((~II10146));
assign WX8646 = (WX8583&RESET);
assign WX4184 = (_2185_&WX4883);
assign II26202 = ((~II26212))|((~II26213));
assign II2420 = ((~II2430))|((~II2431));
assign WX2481 = ((~II7396))|((~II7397));
assign II19711 = ((~_2209_))|((~II19709));
assign WX7471 = ((~II23078))|((~II23079));
assign WX4938 = (WX4936)|(WX4935);
assign WX898 = (WX835&RESET);
assign WX4355 = (WX4353)|(WX4352);
assign WX5128 = ((~II15635))|((~II15636));
assign WX1181 = ((~II3378))|((~II3379));
assign WX3994 = ((~WX4883));
assign II22803 = ((~WX7288))|((~WX7352));
assign II3654 = ((~WX633))|((~_2086_));
assign WX9619 = ((~WX9992));
assign WX8689 = ((~II27002))|((~II27003));
assign II6411 = ((~WX2092))|((~WX2156));
assign WX2890 = (WX2888)|(WX2887);
assign WX2838 = (WX2836)|(WX2835);
assign II22198 = ((~II22200))|((~II22201));
assign WX6211 = ((~WX6210));
assign II14158 = ((~WX4880))|((~WX4534));
assign WX5611 = ((~WX5602));
assign II10712 = ((~WX3588))|((~II10711));
assign WX10653 = (WX10867&WX11348);
assign WX4298 = ((~WX4883));
assign WX7977 = ((~WX8761));
assign WX10006 = ((~WX10005));
assign WX2033 = (WX1970&RESET);
assign WX3244 = (WX2732&RESET);
assign WX6754 = ((~WX7468));
assign II2491 = ((~WX741))|((~II2483));
assign WX7085 = ((~WX7318));
assign II34903 = ((~WX11109))|((~II34895));
assign II34432 = ((~WX11345))|((~II34431));
assign WX9009 = ((~II27664))|((~II27665));
assign WX3707 = ((~WX3591));
assign WX10002 = ((~WX10001));
assign WX8254 = (WX8257&RESET);
assign WX5548 = (WX7645&WX5549);
assign WX3686 = ((~WX3591));
assign WX3624 = (WX3622)|(WX3621);
assign WX6357 = (WX6355)|(WX6354);
assign II14358 = ((~II14360))|((~II14361));
assign II3053 = ((~WX580))|((~II3052));
assign WX167 = ((~WX1004));
assign WX5060 = ((~II15393))|((~II15394));
assign WX7493 = (WX7492&WX7470);
assign WX4304 = ((~WX4295));
assign WX3926 = ((~WX3917));
assign II18023 = ((~WX5945))|((~WX6009));
assign II18573 = ((~WX5917))|((~II18565));
assign WX5767 = ((~WX5735));
assign WX10971 = ((~WX11211));
assign WX5519 = (_2214_&WX6176);
assign II35525 = ((~WX10976))|((~_2364_));
assign WX4458 = ((~WX4842));
assign WX3497 = ((~II10362))|((~II10363));
assign II19627 = ((~_2223_))|((~II19625));
assign WX2077 = (WX2014&RESET);
assign WX11314 = ((~WX11247));
assign WX3976 = ((~WX4883));
assign WX2323 = ((~WX2298));
assign WX9663 = ((~WX9888));
assign II10043 = ((~II10045))|((~II10046));
assign WX1079 = ((~WX1005));
assign WX7833 = ((~WX7824));
assign II34445 = ((~II34447))|((~II34448));
assign II23674 = ((~_2248_))|((~II23672));
assign WX4490 = ((~WX4458));
assign WX7649 = ((~WX7470));
assign WX10744 = (WX10750&WX10745);
assign II31335 = ((~WX9650))|((~II31334));
assign II10059 = ((~II10061))|((~II10062));
assign WX6319 = (WX6318&WX6177);
assign II30303 = ((~WX10052))|((~II30302));
assign II14399 = ((~II14389))|((~II14397));
assign WX8088 = (WX8094&WX8089);
assign WX6861 = (WX6859)|(WX6858);
assign II15080 = ((~WX4460))|((~WX4366));
assign II18286 = ((~II18288))|((~II18289));
assign II7527 = ((~WX1905))|((~II7526));
assign WX157 = ((~WX1004));
assign WX6178 = ((~II19073))|((~II19074));
assign WX4327 = (WX4325)|(WX4324);
assign WX478 = (DATA_9_0&WX479);
assign WX3204 = ((~WX3435));
assign II2121 = ((~II2111))|((~II2119));
assign WX10022 = ((~WX10021));
assign II6813 = ((~II6815))|((~II6816));
assign WX7321 = (WX7258&RESET);
assign II30448 = ((~II30424))|((~II30440));
assign II18909 = ((~WX5875))|((~II18907));
assign WX11307 = ((~WX11306));
assign II6289 = ((~WX2148))|((~II6287));
assign II18822 = ((~WX5933))|((~II18821));
assign WX10570 = (WX11447&WX10571);
assign WX6139 = ((~WX6138));
assign II19308 = ((~WX5693))|((~II19306));
assign II35417 = ((~WX10949))|((~WX10879));
assign II26864 = ((~II26854))|((~II26862));
assign II35605 = ((~_2357_))|((~II35603));
assign WX7726 = ((~II23729))|((~II23730));
assign WX1112 = (WX1111&WX1005);
assign WX8016 = ((~WX8015));
assign II31606 = ((~WX9670))|((~II31605));
assign WX7807 = (WX7818&WX8761);
assign WX9447 = (WX9445)|(WX9444);
assign WX6250 = (WX5762&WX6251);
assign WX6311 = ((~II19320))|((~II19321));
assign WX7205 = (WX7142&RESET);
assign WX9329 = (WX11475&WX9330);
assign WX1447 = (WX1445)|(WX1444);
assign WX6008 = (WX5945&RESET);
assign WX8478 = (WX8415&RESET);
assign WX6382 = (WX6381&WX6177);
assign WX47 = ((~WX38));
assign WX11249 = ((~II34206))|((~II34207));
assign WX5976 = (WX5913&RESET);
assign WX9509 = (WX9507)|(WX9506);
assign II18582 = ((~WX5981))|((~II18581));
assign II30683 = ((~II30673))|((~II30681));
assign WX9123 = (WX10077&WX9124);
assign II14126 = ((~II14128))|((~II14129));
assign WX4100 = (_2191_&WX4883);
assign WX3523 = ((~WX3522));
assign WX9417 = (WX10224&WX9418);
assign WX6435 = ((~WX6402));
assign WX10579 = (_2350_&WX11348);
assign WX10488 = (WX10486)|(WX10485);
assign II34517 = ((~II34507))|((~II34515));
assign II10006 = ((~WX3295))|((~II10005));
assign WX4916 = ((~WX4884));
assign II31270 = ((~WX9645))|((~II31269));
assign WX10284 = ((~II31543))|((~II31544));
assign II27422 = ((~WX8295))|((~II27420));
assign WX10474 = (WX10472)|(WX10471);
assign WX6811 = (WX6809)|(WX6808);
assign II27523 = ((~_2279_))|((~II27522));
assign WX10243 = (WX10241)|(WX10240);
assign WX2509 = ((~II7448))|((~II7449));
assign WX6076 = ((~II18155))|((~II18156));
assign WX1580 = (WX1591&WX2296);
assign II30651 = ((~WX9800))|((~II30650));
assign WX3653 = ((~WX3652));
assign WX8040 = (WX8889&WX8041);
assign WX5402 = ((~WX5401));
assign II6627 = ((~II6629))|((~II6630));
assign WX6259 = (WX6257)|(WX6256);
assign WX4883 = ((~WX4876));
assign WX4741 = (WX4678&RESET);
assign WX10182 = ((~WX10181));
assign WX2749 = ((~WX3589));
assign II34564 = ((~II34554))|((~II34562));
assign WX10029 = ((~WX9958));
assign WX11058 = (WX10995&RESET);
assign WX253 = (WX515&WX1004);
assign WX9111 = (WX9109)|(WX9108);
assign WX8750 = ((~WX8672));
assign WX6903 = (WX6901)|(WX6900);
assign WX6143 = ((~WX6142));
assign WX4248 = ((~WX4239));
assign WX9116 = ((~WX10054));
assign WX8464 = (WX8240&RESET);
assign II35744 = ((~WX10985))|((~II35743));
assign II23653 = ((~_2251_))|((~II23651));
assign WX118 = ((~WX117));
assign II6000 = ((~WX2002))|((~II5992));
assign WX5674 = (WX5677&RESET);
assign WX8385 = ((~WX8625));
assign II18472 = ((~II18474))|((~II18475));
assign II26376 = ((~WX8617))|((~II26374));
assign WX2634 = ((~WX2633));
assign II10480 = ((~WX3453))|((~II10478));
assign II7189 = ((~WX1798))|((~II7187));
assign WX5036 = (WX5034)|(WX5033);
assign WX1869 = ((~WX2250));
assign WX11074 = (WX11011&RESET);
assign WX3402 = (WX3339&RESET);
assign II22244 = ((~II22246))|((~II22247));
assign WX10950 = ((~WX10918));
assign II23402 = ((~WX7070))|((~WX7000));
assign WX11198 = (WX11135&RESET);
assign WX937 = ((~WX936));
assign II22717 = ((~II22693))|((~II22709));
assign II22710 = ((~WX7282))|((~WX7346));
assign WX6070 = (WX6007&RESET);
assign WX2167 = (WX2104&RESET);
assign WX8570 = (WX8507&RESET);
assign II3607 = ((~_2095_))|((~II3605));
assign II23554 = ((~WX7078))|((~II23553));
assign II14251 = ((~WX4880))|((~WX4540));
assign II18110 = ((~II18100))|((~II18108));
assign WX5046 = ((~II15367))|((~II15368));
assign II31375 = ((~WX9580))|((~II31373));
assign WX3137 = ((~WX3557));
assign WX9815 = (WX9752&RESET);
assign WX1589 = (WX2431&WX1590);
assign WX3713 = (WX3183&WX3714);
assign II15613 = ((~WX4502))|((~_2192_));
assign WX2304 = ((~WX2303));
assign WX9676 = ((~WX9914));
assign II26498 = ((~WX8561))|((~WX8625));
assign II18418 = ((~WX5907))|((~II18410));
assign WX3721 = ((~WX3591));
assign WX1914 = ((~WX2148));
assign WX10335 = (WX10305&WX10314);
assign II26051 = ((~WX8405))|((~II26049));
assign WX11402 = ((~WX11349));
assign WX10150 = (WX9644&WX10151);
assign II2041 = ((~II2017))|((~II2033));
assign WX4037 = (WX4035)|(WX4034);
assign WX10969 = ((~WX11207));
assign II22433 = ((~WX7328))|((~II22431));
assign WX11568 = (WX11567&WX11349);
assign WX4581 = (WX4333&RESET);
assign II15718 = ((~WX4520))|((~_2174_));
assign WX8818 = ((~WX8817));
assign II11167 = ((~WX3174))|((~II11166));
assign WX7541 = ((~II23208))|((~II23209));
assign II10928 = ((~WX3588))|((~WX3291));
assign II18015 = ((~WX5881))|((~II18007));
assign II14576 = ((~WX4688))|((~WX4752));
assign II11363 = ((~WX3117))|((~II11361));
assign WX4064 = ((~WX4883));
assign II30487 = ((~II30489))|((~II30490));
assign II10356 = ((~WX3445))|((~II10354));
assign WX1706 = (WX1717&WX2296);
assign II35519 = ((~II35509))|((~II35517));
assign WX5363 = ((~WX6175));
assign II18149 = ((~WX6017))|((~II18147));
assign WX9684 = ((~WX9930));
assign WX178 = (WX176)|(WX175);
assign II6704 = ((~II6714))|((~II6715));
assign II10588 = ((~WX3588))|((~II10587));
assign WX907 = ((~II2228))|((~II2229));
assign WX5115 = ((~II15544))|((~II15545));
assign II14483 = ((~WX4682))|((~WX4746));
assign II23574 = ((~WX7081))|((~_2263_));
assign WX10192 = (WX9650&WX10193);
assign II30480 = ((~II30455))|((~II30479));
assign WX6581 = (WX6579)|(WX6578);
assign II30412 = ((~WX9912))|((~II30410));
assign II31126 = ((~WX9634))|((~WX9542));
assign WX8081 = (WX8283&WX8762);
assign WX7902 = (WX7900)|(WX7899);
assign II22632 = ((~II22634))|((~II22635));
assign WX1658 = (WX1824&WX2297);
assign WX5607 = (WX5713&WX6176);
assign WX3428 = (WX3365&RESET);
assign WX8608 = (WX8545&RESET);
assign II34988 = ((~II34990))|((~II34991));
assign II10213 = ((~II10223))|((~II10224));
assign II22221 = ((~II22197))|((~II22213));
assign WX2332 = ((~WX2331));
assign II34485 = ((~II34460))|((~II34484));
assign II14283 = ((~WX4880))|((~II14282));
assign WX208 = (WX2389&WX209);
assign II11103 = ((~WX3077))|((~II11101));
assign II2173 = ((~II2175))|((~II2176));
assign II26110 = ((~II26112))|((~II26113));
assign II15238 = ((~WX4390))|((~II15236));
assign II7421 = ((~WX1901))|((~WX1834));
assign WX8830 = ((~WX8763));
assign II10478 = ((~WX3389))|((~WX3453));
assign II31400 = ((~WX9655))|((~II31399));
assign II10957 = ((~II10967))|((~II10968));
assign II26802 = ((~II26792))|((~II26800));
assign II10564 = ((~WX3331))|((~II10563));
assign II10177 = ((~II10167))|((~II10175));
assign II22339 = ((~WX7258))|((~II22338));
assign WX2708 = (WX2706)|(WX2705);
assign II11658 = ((~WX3217))|((~II11657));
assign WX5700 = (WX5703&RESET);
assign WX9487 = (WX10259&WX9488);
assign WX11607 = ((~WX11574));
assign WX4980 = (WX4978)|(WX4977);
assign WX8699 = ((~WX8698));
assign WX6657 = (WX6655)|(WX6654);
assign II3697 = ((~WX640))|((~II3696));
assign WX7167 = (WX6919&RESET);
assign WX11332 = ((~WX11256));
assign WX4271 = (WX4269)|(WX4268);
assign WX3364 = (WX3301&RESET);
assign WX173 = ((~WX164));
assign II15224 = ((~WX4471))|((~II15223));
assign II6775 = ((~WX2052))|((~II6767));
assign II23562 = ((~_2265_))|((~II23560));
assign II26491 = ((~WX8497))|((~II26490));
assign WX6707 = (WX6705)|(WX6704);
assign II19724 = ((~WX5813))|((~II19723));
assign WX2818 = (WX2824&WX2819);
assign WX8865 = ((~WX8763));
assign II30063 = ((~II30053))|((~II30061));
assign II10105 = ((~II10107))|((~II10108));
assign II18751 = ((~II18753))|((~II18754));
assign WX2955 = ((~WX2946));
assign II14609 = ((~WX4754))|((~II14607));
assign WX3845 = ((~II11700))|((~II11701));
assign II27147 = ((~WX8343))|((~WX8253));
assign WX2777 = ((~WX3589));
assign WX3551 = ((~WX3550));
assign WX2151 = (WX2088&RESET);
assign WX10012 = ((~WX10011));
assign WX4995 = ((~WX4994));
assign WX4849 = ((~WX4782));
assign II14701 = ((~WX4696))|((~II14700));
assign WX1199 = (WX1197)|(WX1196);
assign WX10294 = ((~II31613))|((~II31614));
assign WX2988 = (WX2986)|(WX2985);
assign II34967 = ((~II34957))|((~II34965));
assign II18272 = ((~WX5961))|((~II18271));
assign WX4151 = ((~WX4150));
assign WX3544 = ((~WX3515));
assign II19634 = ((~_2222_))|((~II19632));
assign WX3817 = ((~II11488))|((~II11489));
assign WX919 = ((~II2600))|((~II2601));
assign WX8544 = (WX8481&RESET);
assign WX9933 = (WX9870&RESET);
assign II26809 = ((~WX8581))|((~II26808));
assign II26800 = ((~WX8517))|((~II26792));
assign II18565 = ((~II18567))|((~II18568));
assign II35603 = ((~WX10962))|((~_2357_));
assign II10185 = ((~WX3587))|((~II10184));
assign II2322 = ((~II2312))|((~II2320));
assign WX8310 = ((~WX8731));
assign II34610 = ((~II34600))|((~II34608));
assign II15212 = ((~WX4386))|((~II15210));
assign WX9877 = (WX9814&RESET);
assign II11707 = ((~WX3226))|((~II11706));
assign II6341 = ((~WX2024))|((~II6333));
assign WX2994 = (WX3780&WX2995);
assign II6302 = ((~II6304))|((~II6305));
assign WX7947 = (WX7958&WX8761);
assign WX914 = ((~II2445))|((~II2446));
assign WX9105 = (WX11363&WX9106);
assign II34074 = ((~WX11119))|((~WX11183));
assign II22812 = ((~II22802))|((~II22810));
assign WX3761 = (WX3760&WX3591);
assign WX6392 = (WX6390)|(WX6389);
assign WX5344 = (WX5342)|(WX5341);
assign II6348 = ((~II6350))|((~II6351));
assign II35484 = ((~WX10889))|((~II35482));
assign WX40 = (WX2305&WX41);
assign WX3830 = ((~II11595))|((~II11596));
assign WX7932 = ((~WX7931));
assign WX1858 = ((~WX2228));
assign WX2027 = (WX1964&RESET);
assign WX7211 = (WX7148&RESET);
assign II31534 = ((~II31536))|((~II31537));
assign II15134 = ((~WX4374))|((~II15132));
assign II3578 = ((~WX620))|((~II3577));
assign WX6600 = ((~WX7468));
assign WX3813 = (WX3811)|(WX3810);
assign WX3781 = ((~II11414))|((~II11415));
assign II19620 = ((~_2224_))|((~II19618));
assign WX738 = (WX675&RESET);
assign WX8684 = ((~II26847))|((~II26848));
assign WX5359 = ((~WX5350));
assign WX4907 = (WX4906&WX4884);
assign WX5076 = (WX4486&WX5077);
assign WX7820 = ((~WX7819));
assign WX5314 = (WX6233&WX5315);
assign WX3565 = ((~WX3564));
assign II10038 = ((~II10028))|((~II10036));
assign WX2701 = ((~WX3590));
assign II14671 = ((~WX4758))|((~II14669));
assign II6906 = ((~II6908))|((~II6909));
assign WX1568 = ((~WX2296));
assign WX3882 = (WX3817&WX3849);
assign WX10686 = ((~WX10685));
assign WX2770 = (WX3668&WX2771);
assign II30140 = ((~II30130))|((~II30138));
assign II6039 = ((~WX2068))|((~WX2132));
assign II34848 = ((~II34850))|((~II34851));
assign WX3468 = (WX3405&RESET);
assign WX11295 = ((~WX11294));
assign II18037 = ((~II18047))|((~II18048));
assign II23299 = ((~WX7062))|((~II23298));
assign II30636 = ((~II30626))|((~II30634));
assign WX8319 = ((~WX8749));
assign WX4264 = (WX4275&WX4882);
assign II14406 = ((~WX4880))|((~WX4550));
assign II19204 = ((~WX5677))|((~II19202));
assign II10632 = ((~II10634))|((~II10635));
assign WX1559 = (WX1557)|(WX1556);
assign II7395 = ((~WX1899))|((~WX1830));
assign II10502 = ((~WX3327))|((~II10501));
assign WX10818 = (DATA_0_0&WX10819);
assign WX3225 = ((~WX3477));
assign WX7983 = (WX8269&WX8762);
assign II22903 = ((~II22879))|((~II22895));
assign WX902 = ((~II2073))|((~II2074));
assign II6822 = ((~II6797))|((~II6821));
assign II27679 = ((~_2280_))|((~II27677));
assign II22321 = ((~II22331))|((~II22332));
assign II22177 = ((~II22167))|((~II22175));
assign WX6551 = (WX7498&WX6552);
assign WX35 = (WX46&WX1003);
assign WX10271 = (WX10269)|(WX10268);
assign II7084 = ((~WX1875))|((~II7083));
assign WX1339 = (WX1337)|(WX1336);
assign II31572 = ((~_2329_))|((~II31570));
assign WX6329 = (WX6327)|(WX6326);
assign II23722 = ((~WX7105))|((~II23721));
assign II22332 = ((~II22322))|((~II22330));
assign II6909 = ((~WX2188))|((~II6907));
assign WX5467 = (WX5693&WX6176);
assign WX9050 = (WX9009&WX9021);
assign WX567 = ((~WX939));
assign II11554 = ((~_2168_))|((~II11552));
assign II22276 = ((~WX7254))|((~WX7318));
assign WX7715 = ((~II23652))|((~II23653));
assign WX8917 = ((~WX8916));
assign WX1617 = (WX2445&WX1618);
assign WX4252 = ((~WX4882));
assign WX7067 = ((~WX7035));
assign WX594 = ((~WX562));
assign WX5626 = ((~WX5625));
assign WX1775 = ((~WX1774));
assign WX8781 = ((~WX8763));
assign II2569 = ((~II2544))|((~II2568));
assign WX11462 = ((~II35301))|((~II35302));
assign WX4067 = ((~WX4066));
assign WX8335 = ((~WX8717));
assign II26275 = ((~II26265))|((~II26273));
assign WX1472 = (_2130_&WX2297);
assign II35456 = ((~WX10952))|((~WX10885));
assign II18568 = ((~WX5853))|((~II18566));
assign WX4340 = ((~WX4883));
assign WX9495 = (WX9493)|(WX9492);
assign II22665 = ((~WX7467))|((~II22664));
assign WX6350 = (WX6348)|(WX6347);
assign II2935 = ((~WX897))|((~II2933));
assign II30372 = ((~WX9782))|((~II30371));
assign II11672 = ((~WX3220))|((~II11671));
assign WX6058 = (WX5995&RESET);
assign II35717 = ((~_2339_))|((~II35715));
assign II26437 = ((~WX8557))|((~II26436));
assign WX8360 = ((~WX8328));
assign II6684 = ((~II6674))|((~II6682));
assign WX9604 = ((~WX10026));
assign WX9423 = (WX9429&WX9424);
assign II27581 = ((~_2295_))|((~II27579));
assign WX1402 = (_2135_&WX2297);
assign II34539 = ((~WX11149))|((~WX11213));
assign WX10188 = ((~WX10187));
assign WX3068 = ((~WX3067));
assign II27594 = ((~WX8376))|((~II27593));
assign WX9923 = (WX9860&RESET);
assign WX7620 = (WX7066&WX7621);
assign II34495 = ((~WX11019))|((~II34493));
assign II14839 = ((~II14841))|((~II14842));
assign II10534 = ((~II10524))|((~II10532));
assign WX1282 = (WX1255&WX1263);
assign WX8522 = (WX8459&RESET);
assign WX3888 = (WX3833&WX3849);
assign WX2730 = (WX2728)|(WX2727);
assign II14956 = ((~II14931))|((~II14955));
assign WX8780 = (WX8340&WX8781);
assign WX4432 = ((~WX4854));
assign II27517 = ((~_2300_))|((~II27515));
assign II10819 = ((~WX3411))|((~WX3475));
assign II30915 = ((~II30905))|((~II30913));
assign WX10169 = ((~II31296))|((~II31297));
assign II6746 = ((~II6736))|((~II6744));
assign WX9170 = (WX9181&WX10054);
assign WX6362 = (WX5778&WX6363);
assign WX548 = ((~WX965));
assign WX4808 = ((~II14925))|((~II14926));
assign II10248 = ((~WX3247))|((~II10246));
assign WX11546 = ((~II35457))|((~II35458));
assign WX824 = (WX761&RESET);
assign WX722 = (WX659&RESET);
assign II31710 = ((~WX9687))|((~_2307_));
assign WX9525 = (WX11573&WX9526);
assign II18301 = ((~II18303))|((~II18304));
assign WX7060 = ((~WX7028));
assign II14229 = ((~II14219))|((~II14227));
assign WX1363 = (WX1361)|(WX1360);
assign II30952 = ((~II30954))|((~II30955));
assign II15184 = ((~WX4468))|((~WX4382));
assign II7549 = ((~_2136_))|((~II7547));
assign WX3514 = ((~II10889))|((~II10890));
assign WX5656 = (WX5659&RESET);
assign WX11112 = (WX11049&RESET);
assign WX11357 = ((~II35106))|((~II35107));
assign WX9072 = (WX8999&WX9021);
assign WX10082 = (WX10080)|(WX10079);
assign II11687 = ((~_2147_))|((~II11685));
assign II18503 = ((~II18505))|((~II18506));
assign WX7486 = (WX7485&WX7470);
assign DATA_9_9 = ((~WX1165));
assign WX8324 = ((~WX8695));
assign II27434 = ((~WX8365))|((~II27433));
assign II2749 = ((~WX885))|((~II2747));
assign WX5441 = ((~WX6176));
assign WX454 = ((~WX453));
assign II19451 = ((~WX5715))|((~II19449));
assign II6157 = ((~II6147))|((~II6155));
assign WX8358 = ((~WX8326));
assign II34880 = ((~WX11171))|((~WX11235));
assign WX4968 = ((~WX4967));
assign WX604 = ((~WX572));
assign II2467 = ((~II2469))|((~II2470));
assign II2438 = ((~WX801))|((~II2437));
assign WX10238 = ((~WX10237));
assign WX3947 = (WX6198&WX3948);
assign WX10118 = ((~WX10117));
assign WX1647 = (WX1645)|(WX1644);
assign II26087 = ((~WX8471))|((~II26079));
assign WX4208 = (WX4219&WX4882);
assign II19548 = ((~WX5785))|((~_2234_));
assign WX6650 = ((~WX7469));
assign WX532 = (WX535&RESET);
assign II2337 = ((~WX731))|((~II2336));
assign WX258 = ((~WX257));
assign WX692 = (WX384&RESET);
assign WX556 = ((~WX981));
assign II14523 = ((~II14513))|((~II14521));
assign II23364 = ((~WX7067))|((~II23363));
assign II6613 = ((~WX2295))|((~WX1978));
assign WX3561 = ((~WX3560));
assign WX201 = ((~WX192));
assign WX3488 = ((~II10083))|((~II10084));
assign II22146 = ((~II22136))|((~II22144));
assign WX187 = ((~WX178));
assign WX5383 = (WX5681&WX6176);
assign WX2366 = (WX2364)|(WX2363);
assign WX7147 = (WX6779&RESET);
assign II34934 = ((~WX11111))|((~II34926));
assign WX5698 = (WX5701&RESET);
assign WX6918 = ((~WX6909));
assign II18101 = ((~WX6173))|((~WX5823));
assign II26080 = ((~WX8759))|((~WX8407));
assign WX510 = (WX513&RESET);
assign WX3063 = (WX3133&WX3590);
assign WX5739 = ((~WX6111));
assign II6164 = ((~WX2076))|((~II6163));
assign WX4453 = ((~WX4832));
assign WX3268 = (WX2900&RESET);
assign II7533 = ((~WX1906))|((~_2138_));
assign WX1709 = (WX1707)|(WX1706);
assign WX10479 = ((~WX11347));
assign WX3549 = ((~WX3548));
assign WX5175 = (WX5110&WX5142);
assign II30604 = ((~II30579))|((~II30603));
assign II30031 = ((~WX9760))|((~II30030));
assign II3456 = ((~WX611))|((~II3455));
assign WX7277 = (WX7214&RESET);
assign WX7027 = ((~WX7458));
assign II23103 = ((~WX7047))|((~WX6954));
assign WX1088 = ((~WX1087));
assign II23274 = ((~WX6980))|((~II23272));
assign WX973 = ((~WX972));
assign WX8148 = (WX10238&WX8149);
assign WX11128 = (WX11065&RESET);
assign WX10597 = (WX10859&WX11348);
assign II26126 = ((~WX8537))|((~WX8601));
assign II10253 = ((~WX3311))|((~II10245));
assign WX8556 = (WX8493&RESET);
assign WX381 = ((~WX1004));
assign WX11579 = ((~II35562))|((~II35563));
assign II10540 = ((~WX3393))|((~WX3457));
assign WX6669 = (WX6675&WX6670);
assign II6798 = ((~II6800))|((~II6801));
assign II6301 = ((~II6311))|((~II6312));
assign WX4837 = ((~WX4808));
assign WX10371 = (WX10289&WX10314);
assign WX5812 = ((~WX6065));
assign II30216 = ((~WX9772))|((~II30208));
assign WX1093 = ((~WX1005));
assign WX560 = ((~WX989));
assign II2771 = ((~WX759))|((~II2770));
assign WX9226 = (WX9237&WX10054);
assign WX1332 = (_2140_&WX2297);
assign WX6342 = ((~WX6177));
assign WX8304 = (WX8241&RESET);
assign WX9645 = ((~WX9613));
assign WX2690 = ((~WX2689));
assign II14986 = ((~II14962))|((~II14978));
assign WX7319 = (WX7256&RESET);
assign II14738 = ((~II14714))|((~II14730));
assign WX11483 = ((~II35340))|((~II35341));
assign WX2907 = ((~WX3590));
assign II7410 = ((~WX1832))|((~II7408));
assign WX3084 = (WX3087&RESET);
assign WX3967 = (WX3965)|(WX3964);
assign WX2731 = ((~WX2722));
assign WX1541 = (WX1539)|(WX1538);
assign II19695 = ((~WX5808))|((~_2211_));
assign II11692 = ((~WX3223))|((~_2146_));
assign II14614 = ((~II14590))|((~II14606));
assign II18224 = ((~II18226))|((~II18227));
assign II18209 = ((~WX5957))|((~WX6021));
assign WX5455 = ((~WX6176));
assign WX1508 = ((~WX1499));
assign II26399 = ((~II26389))|((~II26397));
assign II31512 = ((~_2316_))|((~II31504));
assign II14445 = ((~WX4616))|((~II14444));
assign WX6052 = (WX5989&RESET);
assign WX8824 = (WX8822)|(WX8821);
assign WX3032 = (WX5094&WX3033);
assign WX7051 = ((~WX7019));
assign II34144 = ((~II34119))|((~II34143));
assign II14299 = ((~WX4734))|((~II14297));
assign WX5014 = ((~WX4884));
assign II34802 = ((~II34804))|((~II34805));
assign WX2883 = ((~WX3590));
assign WX7616 = ((~WX7615));
assign WX1438 = ((~WX1429));
assign WX5525 = ((~WX6176));
assign WX4977 = (WX4976&WX4884);
assign II34787 = ((~WX11165))|((~WX11229));
assign WX925 = ((~II2786))|((~II2787));
assign II34244 = ((~II34246))|((~II34247));
assign II26755 = ((~II26745))|((~II26753));
assign II6583 = ((~WX2295))|((~II6582));
assign WX193 = (_2097_&WX1004);
assign II18201 = ((~WX5893))|((~II18193));
assign II14067 = ((~WX4528))|((~II14065));
assign WX6166 = ((~WX6087));
assign WX11555 = (WX10953&WX11556);
assign II6133 = ((~WX2074))|((~II6132));
assign WX10256 = ((~WX10056));
assign WX7341 = (WX7278&RESET);
assign II11573 = ((~WX3204))|((~_2165_));
assign WX7461 = ((~TM0));
assign II14453 = ((~WX4680))|((~II14452));
assign WX4005 = (WX4003)|(WX4002);
assign WX10936 = ((~WX10904));
assign II15552 = ((~_2201_))|((~II15550));
assign WX2298 = ((~WX2289));
assign WX8873 = (WX8871)|(WX8870);
assign II22509 = ((~WX7467))|((~WX7142));
assign II18318 = ((~WX6173))|((~WX5837));
assign WX8769 = ((~WX8768));
assign II22011 = ((~II22021))|((~II22022));
assign WX4286 = (WX4416&WX4883);
assign WX7891 = (WX7902&WX8761);
assign WX7827 = ((~WX8762));
assign II31579 = ((~_2328_))|((~II31577));
assign WX9697 = (WX9113&RESET);
assign WX1575 = (WX2424&WX1576);
assign WX7531 = (WX7529)|(WX7528);
assign WX2587 = (WX2543&WX2556);
assign WX3189 = ((~WX3157));
assign II14942 = ((~II14932))|((~II14940));
assign WX11166 = (WX11103&RESET);
assign II23157 = ((~WX6962))|((~II23155));
assign WX2196 = ((~II6109))|((~II6110));
assign WX2420 = (WX1890&WX2421);
assign II11624 = ((~_2158_))|((~II11622));
assign WX9286 = (_2318_&WX10055);
assign WX3959 = (WX3957)|(WX3956);
assign II14864 = ((~II14854))|((~II14862));
assign WX3576 = ((~WX3499));
assign WX1460 = ((~WX2297));
assign WX7185 = (WX7122&RESET);
assign II30768 = ((~WX10053))|((~II30767));
assign WX3822 = ((~II11539))|((~II11540));
assign II10865 = ((~II10867))|((~II10868));
assign II34129 = ((~WX11059))|((~II34128));
assign WX10588 = ((~WX10587));
assign II19151 = ((~WX5758))|((~II19150));
assign II18311 = ((~II18301))|((~II18309));
assign II26017 = ((~II26019))|((~II26020));
assign II2739 = ((~WX757))|((~II2731));
assign WX724 = (WX661&RESET);
assign WX1035 = (WX1034&WX1005);
assign WX2359 = (WX2357)|(WX2356);
assign WX10068 = (WX10066)|(WX10065);
assign II31717 = ((~WX9688))|((~_2306_));
assign WX11566 = ((~WX11565));
assign II11631 = ((~_2157_))|((~II11629));
assign WX7687 = ((~WX7686));
assign II10122 = ((~WX3587))|((~WX3239));
assign WX8981 = ((~II27486))|((~II27487));
assign WX1899 = ((~WX1867));
assign WX161 = (WX172&WX1003);
assign WX10341 = (WX10303&WX10314);
assign II11679 = ((~WX3221))|((~II11678));
assign II22106 = ((~WX7466))|((~WX7116));
assign II2498 = ((~II2500))|((~II2501));
assign WX2526 = ((~II7513))|((~II7514));
assign WX8927 = (WX8361&WX8928);
assign WX7680 = ((~WX7679));
assign II23623 = ((~WX7088))|((~_2256_));
assign WX2053 = (WX1990&RESET);
assign WX1455 = (WX1461&WX1456);
assign II11153 = ((~WX3173))|((~WX3085));
assign II15198 = ((~WX4469))|((~II15197));
assign II15457 = ((~WX4489))|((~WX4424));
assign WX10516 = (WX10514)|(WX10513);
assign WX6723 = ((~WX6722));
assign WX5372 = (WX5370)|(WX5369);
assign WX5082 = (WX5081&WX4884);
assign II30109 = ((~II30099))|((~II30107));
assign II22635 = ((~WX7150))|((~II22633));
assign WX7882 = (WX10105&WX7883);
assign II3571 = ((~WX619))|((~II3570));
assign II26885 = ((~II26887))|((~II26888));
assign WX3700 = ((~WX3591));
assign WX3182 = ((~WX3150));
assign II18782 = ((~II18784))|((~II18785));
assign II3614 = ((~_2094_))|((~II3612));
assign WX5477 = (_2217_&WX6176);
assign WX3053 = ((~WX3044));
assign II26900 = ((~II26902))|((~II26903));
assign WX10772 = (WX10778&WX10773);
assign WX10773 = ((~WX11347));
assign WX4978 = (WX4472&WX4979);
endmodule
