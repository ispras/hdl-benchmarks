//NOTE: no-implementation module stub

module GtCLK_NAND2 (
    output Z,
    input A,
    input B
);

endmodule
