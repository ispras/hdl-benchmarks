module bitwise_and_4_1(a, b, c);
  input [3:0] a;
  input b;
  output [3:0] c;
  assign c = a & b;
endmodule
