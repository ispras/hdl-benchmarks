module logical_not_3_1(a, b);
  input [2:0] a;
  output b;
  assign b = !a;
endmodule
