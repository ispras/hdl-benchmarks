module logical_not_3_3(a, b);
  input [2:0] a;
  output [2:0] b;
  assign b = !a;
endmodule
