//NOTE: no-implementation module stub

module SU208010 (
    input wire A0,
    input wire A1,
    input wire A2,
    input wire A3,
    input wire A4,
    input wire A5,
    input wire A6,
    input wire A7,
    input wire A8,
    input wire A9,
    input wire A10,
    input wire A11,
    `ifdef FD_PM8K
    input wire A12,
    `endif
    output wire DO0,
    output wire DO1,
    output wire DO2,
    output wire DO3,
    output wire DO4,
    output wire DO5,
    output wire DO6,
    output wire DO7,
    output wire DO8,
    output wire DO9,
    output wire DO10,
    output wire DO11,
    output wire DO12,
    output wire DO13,
    output wire DO14,
    output wire DO15,
    input wire DI0,
    input wire DI1,
    input wire DI2,
    input wire DI3,
    input wire DI4,
    input wire DI5,
    input wire DI6,
    input wire DI7,
    input wire DI8,
    input wire DI9,
    input wire DI10,
    input wire DI11,
    input wire DI12,
    input wire DI13,
    input wire DI14,
    input wire DI15,
    input wire CK,
    input wire WEB,
    input wire CS,
    input wire OE
);
endmodule

module SU210018 (
    input wire A0,
    input wire A1,
    input wire A2,
    input wire A3,
    input wire A4,
    input wire A5,
    input wire A6,
    input wire A7,
    input wire A8,
    input wire A9,
    input wire A10,
    input wire A11,
    `ifdef FD_PM8K
    // No A12 input if FD_PM8K is defined
    `else
    input wire A12,
    `endif
    output wire DO0,
    output wire DO1,
    output wire DO2,
    output wire DO3,
    output wire DO4,
    output wire DO5,
    output wire DO6,
    output wire DO7,
    output wire DO8,
    output wire DO9,
    output wire DO10,
    output wire DO11,
    output wire DO12,
    output wire DO13,
    output wire DO14,
    output wire DO15,
    output wire DO16,
    output wire DO17,
    output wire DO18,
    output wire DO19,
    output wire DO20,
    output wire DO21,
    output wire DO22,
    output wire DO23,
    input wire DI0,
    input wire DI1,
    input wire DI2,
    input wire DI3,
    input wire DI4,
    input wire DI5,
    input wire DI6,
    input wire DI7,
    input wire DI8,
    input wire DI9,
    input wire DI10,
    input wire DI11,
    input wire DI12,
    input wire DI13,
    input wire DI14,
    input wire DI15,
    input wire DI16,
    input wire DI17,
    input wire DI18,
    input wire DI19,
    input wire DI20,
    input wire DI21,
    input wire DI22,
    input wire DI23,
    input wire CK,
    input wire WEB,
    input wire CS,
    input wire OE
);
endmodule

module SU208018 (
    input wire A0,
    input wire A1,
    input wire A2,
    input wire A3,
    input wire A4,
    input wire A5,
    input wire A6,
    input wire A7,
    input wire A8,
    input wire A9,
    input wire A10,
    input wire A11,
    output wire DO0,
    output wire DO1,
    output wire DO2,
    output wire DO3,
    output wire DO4,
    output wire DO5,
    output wire DO6,
    output wire DO7,
    output wire DO8,
    output wire DO9,
    output wire DO10,
    output wire DO11,
    output wire DO12,
    output wire DO13,
    output wire DO14,
    output wire DO15,
    output wire DO16,
    output wire DO17,
    output wire DO18,
    output wire DO19,
    output wire DO20,
    output wire DO21,
    output wire DO22,
    output wire DO23,
    input wire DI0,
    input wire DI1,
    input wire DI2,
    input wire DI3,
    input wire DI4,
    input wire DI5,
    input wire DI6,
    input wire DI7,
    input wire DI8,
    input wire DI9,
    input wire DI10,
    input wire DI11,
    input wire DI12,
    input wire DI13,
    input wire DI14,
    input wire DI15,
    input wire DI16,
    input wire DI17,
    input wire DI18,
    input wire DI19,
    input wire DI20,
    input wire DI21,
    input wire DI22,
    input wire DI23,
    input wire CK,
    input wire WEB,
    input wire CS,
    input wire OE
);
endmodule

module SU20E010 (
    input wire A0,
    input wire A1,
    input wire A2,
    input wire A3,
    input wire A4,
    input wire A5,
    input wire A6,
    input wire A7,
    input wire A8,
    input wire A9,
    input wire A10,
    input wire A11,
    input wire A12,
    output wire DO0,
    output wire DO1,
    output wire DO2,
    output wire DO3,
    output wire DO4,
    output wire DO5,
    output wire DO6,
    output wire DO7,
    output wire DO8,
    output wire DO9,
    output wire DO10,
    output wire DO11,
    output wire DO12,
    output wire DO13,
    output wire DO14,
    output wire DO15,
    input wire DI0,
    input wire DI1,
    input wire DI2,
    input wire DI3,
    input wire DI4,
    input wire DI5,
    input wire DI6,
    input wire DI7,
    input wire DI8,
    input wire DI9,
    input wire DI10,
    input wire DI11,
    input wire DI12,
    input wire DI13,
    input wire DI14,
    input wire DI15,
    input wire CK,
    input wire WEB,
    input wire CS,
    input wire OE
);
endmodule

module SU210010 (
    input wire A0,
    input wire A1,
    input wire A2,
    input wire A3,
    input wire A4,
    input wire A5,
    input wire A6,
    input wire A7,
    input wire A8,
    input wire A9,
    input wire A10,
    input wire A11,
    input wire A12,
    output wire DO0,
    output wire DO1,
    output wire DO2,
    output wire DO3,
    output wire DO4,
    output wire DO5,
    output wire DO6,
    output wire DO7,
    output wire DO8,
    output wire DO9,
    output wire DO10,
    output wire DO11,
    output wire DO12,
    output wire DO13,
    output wire DO14,
    output wire DO15,
    input wire DI0,
    input wire DI1,
    input wire DI2,
    input wire DI3,
    input wire DI4,
    input wire DI5,
    input wire DI6,
    input wire DI7,
    input wire DI8,
    input wire DI9,
    input wire DI10,
    input wire DI11,
    input wire DI12,
    input wire DI13,
    input wire DI14,
    input wire DI15,
    input wire CK,
    input wire WEB,
    input wire CS,
    input wire OE
);
endmodule
