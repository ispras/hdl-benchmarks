//
// Conformal-LEC Version 15.10-d003 ( 23-Apr-2015) ( 64 bit executable)
//
module top ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 , 
    n5008 , 
    n5009 , 
    n5010 , 
    n5011 , 
    n5012 , 
    n5013 , 
    n5014 , 
    n5015 , 
    n5016 , 
    n5017 , 
    n5018 , 
    n5019 , 
    n5020 , 
    n5021 , 
    n5022 , 
    n5023 , 
    n5024 , 
    n5025 , 
    n5026 , 
    n5027 , 
    n5028 , 
    n5029 , 
    n5030 , 
    n5031 , 
    n5032 , 
    n5033 , 
    n5034 , 
    n5035 , 
    n5036 , 
    n5037 , 
    n5038 , 
    n5039 , 
    n5040 , 
    n5041 , 
    n5042 , 
    n5043 , 
    n5044 , 
    n5045 , 
    n5046 , 
    n5047 , 
    n5048 , 
    n5049 , 
    n5050 , 
    n5051 , 
    n5052 , 
    n5053 , 
    n5054 , 
    n5055 , 
    n5056 , 
    n5057 , 
    n5058 , 
    n5059 , 
    n5060 , 
    n5061 , 
    n5062 , 
    n5063 , 
    n5064 , 
    n5065 , 
    n5066 , 
    n5067 , 
    n5068 , 
    n5069 , 
    n5070 , 
    n5071 , 
    n5072 , 
    n5073 , 
    n5074 , 
    n5075 , 
    n5076 , 
    n5077 , 
    n5078 , 
    n5079 , 
    n5080 , 
    n5081 , 
    n5082 , 
    n5083 , 
    n5084 , 
    n5085 , 
    n5086 , 
    n5087 , 
    n5088 , 
    n5089 , 
    n5090 , 
    n5091 , 
    n5092 , 
    n5093 , 
    n5094 , 
    n5095 , 
    n5096 , 
    n5097 , 
    n5098 , 
    n5099 , 
    n5100 , 
    n5101 , 
    n5102 , 
    n5103 , 
    n5104 , 
    n5105 , 
    n5106 , 
    n5107 , 
    n5108 , 
    n5109 , 
    n5110 , 
    n5111 , 
    n5112 , 
    n5113 , 
    n5114 , 
    n5115 , 
    n5116 , 
    n5117 , 
    n5118 , 
    n5119 , 
    n5120 , 
    n5121 , 
    n5122 , 
    n5123 , 
    n5124 , 
    n5125 , 
    n5126 , 
    n5127 , 
    n5128 , 
    n5129 , 
    n5130 , 
    n5131 , 
    n5132 , 
    n5133 , 
    n5134 , 
    n5135 , 
    n5136 , 
    n5137 , 
    n5138 , 
    n5139 , 
    n5140 , 
    n5141 , 
    n5142 , 
    n5143 , 
    n5144 , 
    n5145 , 
    n5146 , 
    n5147 , 
    n5148 , 
    n5149 , 
    n5150 , 
    n5151 , 
    n5152 , 
    n5153 , 
    n5154 , 
    n5155 , 
    n5156 , 
    n5157 , 
    n5158 , 
    n5159 , 
    n5160 , 
    n5161 , 
    n5162 , 
    n5163 , 
    n5164 , 
    n5165 , 
    n5166 , 
    n5167 , 
    n5168 , 
    n5169 , 
    n5170 , 
    n5171 , 
    n5172 , 
    n5173 , 
    n5174 , 
    n5175 , 
    n5176 , 
    n5177 , 
    n5178 , 
    n5179 , 
    n5180 , 
    n5181 , 
    n5182 , 
    n5183 , 
    n5184 , 
    n5185 , 
    n5186 , 
    n5187 , 
    n5188 , 
    n5189 , 
    n5190 , 
    n5191 , 
    n5192 , 
    n5193 , 
    n5194 , 
    n5195 , 
    n5196 , 
    n5197 , 
    n5198 , 
    n5199 , 
    n5200 , 
    n5201 , 
    n5202 , 
    n5203 , 
    n5204 , 
    n5205 , 
    n5206 , 
    n5207 , 
    n5208 , 
    n5209 , 
    n5210 , 
    n5211 , 
    n5212 , 
    n5213 , 
    n5214 , 
    n5215 , 
    n5216 , 
    n5217 , 
    n5218 , 
    n5219 , 
    n5220 , 
    n5221 , 
    n5222 , 
    n5223 , 
    n5224 , 
    n5225 , 
    n5226 , 
    n5227 , 
    n5228 , 
    n5229 , 
    n5230 , 
    n5231 , 
    n5232 , 
    n5233 , 
    n5234 , 
    n5235 , 
    n5236 , 
    n5237 , 
    n5238 , 
    n5239 , 
    n5240 , 
    n5241 , 
    n5242 , 
    n5243 , 
    n5244 , 
    n5245 , 
    n5246 , 
    n5247 , 
    n5248 , 
    n5249 , 
    n5250 , 
    n5251 , 
    n5252 , 
    n5253 , 
    n5254 , 
    n5255 , 
    n5256 , 
    n5257 , 
    n5258 , 
    n5259 , 
    n5260 , 
    n5261 , 
    n5262 , 
    n5263 , 
    n5264 , 
    n5265 , 
    n5266 , 
    n5267 , 
    n5268 , 
    n5269 , 
    n5270 , 
    n5271 , 
    n5272 , 
    n5273 , 
    n5274 , 
    n5275 , 
    n5276 , 
    n5277 , 
    n5278 , 
    n5279 , 
    n5280 , 
    n5281 , 
    n5282 , 
    n5283 , 
    n5284 , 
    n5285 , 
    n5286 , 
    n5287 , 
    n5288 , 
    n5289 , 
    n5290 , 
    n5291 , 
    n5292 , 
    n5293 , 
    n5294 , 
    n5295 , 
    n5296 , 
    n5297 , 
    n5298 , 
    n5299 , 
    n5300 , 
    n5301 , 
    n5302 , 
    n5303 , 
    n5304 , 
    n5305 , 
    n5306 , 
    n5307 , 
    n5308 , 
    n5309 , 
    n5310 , 
    n5311 , 
    n5312 , 
    n5313 , 
    n5314 , 
    n5315 , 
    n5316 , 
    n5317 , 
    n5318 , 
    n5319 , 
    n5320 , 
    n5321 , 
    n5322 , 
    n5323 , 
    n5324 , 
    n5325 , 
    n5326 , 
    n5327 , 
    n5328 , 
    n5329 , 
    n5330 , 
    n5331 , 
    n5332 , 
    n5333 , 
    n5334 , 
    n5335 , 
    n5336 , 
    n5337 , 
    n5338 , 
    n5339 , 
    n5340 , 
    n5341 , 
    n5342 , 
    n5343 , 
    n5344 , 
    n5345 , 
    n5346 , 
    n5347 , 
    n5348 , 
    n5349 , 
    n5350 , 
    n5351 , 
    n5352 , 
    n5353 , 
    n5354 , 
    n5355 , 
    n5356 , 
    n5357 , 
    n5358 , 
    n5359 , 
    n5360 , 
    n5361 , 
    n5362 , 
    n5363 , 
    n5364 , 
    n5365 , 
    n5366 , 
    n5367 , 
    n5368 , 
    n5369 , 
    n5370 , 
    n5371 , 
    n5372 , 
    n5373 , 
    n5374 , 
    n5375 , 
    n5376 , 
    n5377 , 
    n5378 , 
    n5379 , 
    n5380 , 
    n5381 , 
    n5382 , 
    n5383 , 
    n5384 , 
    n5385 , 
    n5386 , 
    n5387 , 
    n5388 , 
    n5389 , 
    n5390 , 
    n5391 , 
    n5392 , 
    n5393 , 
    n5394 , 
    n5395 , 
    n5396 , 
    n5397 , 
    n5398 , 
    n5399 , 
    n5400 , 
    n5401 , 
    n5402 , 
    n5403 , 
    n5404 , 
    n5405 , 
    n5406 , 
    n5407 , 
    n5408 , 
    n5409 , 
    n5410 , 
    n5411 , 
    n5412 , 
    n5413 , 
    n5414 , 
    n5415 , 
    n5416 , 
    n5417 , 
    n5418 , 
    n5419 , 
    n5420 , 
    n5421 , 
    n5422 , 
    n5423 , 
    n5424 , 
    n5425 , 
    n5426 , 
    n5427 , 
    n5428 , 
    n5429 , 
    n5430 , 
    n5431 , 
    n5432 , 
    n5433 , 
    n5434 , 
    n5435 , 
    n5436 , 
    n5437 , 
    n5438 , 
    n5439 , 
    n5440 , 
    n5441 , 
    n5442 , 
    n5443 , 
    n5444 , 
    n5445 , 
    n5446 , 
    n5447 , 
    n5448 , 
    n5449 , 
    n5450 , 
    n5451 , 
    n5452 , 
    n5453 , 
    n5454 , 
    n5455 , 
    n5456 , 
    n5457 , 
    n5458 , 
    n5459 , 
    n5460 , 
    n5461 , 
    n5462 , 
    n5463 , 
    n5464 , 
    n5465 , 
    n5466 , 
    n5467 , 
    n5468 , 
    n5469 , 
    n5470 , 
    n5471 , 
    n5472 , 
    n5473 , 
    n5474 , 
    n5475 , 
    n5476 , 
    n5477 , 
    n5478 , 
    n5479 , 
    n5480 , 
    n5481 , 
    n5482 , 
    n5483 , 
    n5484 , 
    n5485 , 
    n5486 , 
    n5487 , 
    n5488 , 
    n5489 , 
    n5490 , 
    n5491 , 
    n5492 , 
    n5493 , 
    n5494 , 
    n5495 , 
    n5496 , 
    n5497 , 
    n5498 , 
    n5499 , 
    n5500 , 
    n5501 , 
    n5502 , 
    n5503 , 
    n5504 , 
    n5505 , 
    n5506 , 
    n5507 , 
    n5508 , 
    n5509 , 
    n5510 , 
    n5511 , 
    n5512 , 
    n5513 , 
    n5514 , 
    n5515 , 
    n5516 , 
    n5517 , 
    n5518 , 
    n5519 , 
    n5520 , 
    n5521 , 
    n5522 , 
    n5523 , 
    n5524 , 
    n5525 , 
    n5526 , 
    n5527 , 
    n5528 , 
    n5529 , 
    n5530 , 
    n5531 , 
    n5532 , 
    n5533 , 
    n5534 , 
    n5535 , 
    n5536 , 
    n5537 , 
    n5538 , 
    n5539 , 
    n5540 , 
    n5541 , 
    n5542 , 
    n5543 , 
    n5544 , 
    n5545 , 
    n5546 , 
    n5547 , 
    n5548 , 
    n5549 , 
    n5550 , 
    n5551 , 
    n5552 , 
    n5553 , 
    n5554 , 
    n5555 , 
    n5556 , 
    n5557 , 
    n5558 , 
    n5559 , 
    n5560 , 
    n5561 , 
    n5562 , 
    n5563 , 
    n5564 , 
    n5565 , 
    n5566 , 
    n5567 , 
    n5568 , 
    n5569 , 
    n5570 , 
    n5571 , 
    n5572 , 
    n5573 , 
    n5574 , 
    n5575 , 
    n5576 , 
    n5577 , 
    n5578 , 
    n5579 , 
    n5580 , 
    n5581 , 
    n5582 , 
    n5583 , 
    n5584 , 
    n5585 , 
    n5586 , 
    n5587 , 
    n5588 , 
    n5589 , 
    n5590 , 
    n5591 , 
    n5592 , 
    n5593 , 
    n5594 , 
    n5595 , 
    n5596 , 
    n5597 , 
    n5598 , 
    n5599 , 
    n5600 , 
    n5601 , 
    n5602 , 
    n5603 , 
    n5604 , 
    n5605 , 
    n5606 , 
    n5607 , 
    n5608 , 
    n5609 , 
    n5610 , 
    n5611 , 
    n5612 , 
    n5613 , 
    n5614 , 
    n5615 , 
    n5616 , 
    n5617 , 
    n5618 , 
    n5619 , 
    n5620 , 
    n5621 , 
    n5622 , 
    n5623 , 
    n5624 , 
    n5625 , 
    n5626 , 
    n5627 , 
    n5628 , 
    n5629 , 
    n5630 , 
    n5631 , 
    n5632 , 
    n5633 , 
    n5634 , 
    n5635 , 
    n5636 , 
    n5637 , 
    n5638 , 
    n5639 , 
    n5640 , 
    n5641 , 
    n5642 , 
    n5643 , 
    n5644 , 
    n5645 , 
    n5646 , 
    n5647 , 
    n5648 , 
    n5649 , 
    n5650 , 
    n5651 , 
    n5652 , 
    n5653 , 
    n5654 , 
    n5655 , 
    n5656 , 
    n5657 , 
    n5658 , 
    n5659 , 
    n5660 , 
    n5661 , 
    n5662 , 
    n5663 , 
    n5664 , 
    n5665 , 
    n5666 , 
    n5667 , 
    n5668 , 
    n5669 , 
    n5670 , 
    n5671 , 
    n5672 , 
    n5673 , 
    n5674 , 
    n5675 , 
    n5676 , 
    n5677 , 
    n5678 , 
    n5679 , 
    n5680 , 
    n5681 , 
    n5682 , 
    n5683 , 
    n5684 , 
    n5685 , 
    n5686 , 
    n5687 , 
    n5688 , 
    n5689 , 
    n5690 , 
    n5691 , 
    n5692 , 
    n5693 , 
    n5694 , 
    n5695 , 
    n5696 , 
    n5697 , 
    n5698 , 
    n5699 , 
    n5700 , 
    n5701 , 
    n5702 , 
    n5703 , 
    n5704 , 
    n5705 , 
    n5706 , 
    n5707 , 
    n5708 , 
    n5709 , 
    n5710 , 
    n5711 , 
    n5712 , 
    n5713 , 
    n5714 , 
    n5715 , 
    n5716 , 
    n5717 , 
    n5718 , 
    n5719 , 
    n5720 , 
    n5721 , 
    n5722 , 
    n5723 , 
    n5724 , 
    n5725 , 
    n5726 , 
    n5727 , 
    n5728 , 
    n5729 , 
    n5730 , 
    n5731 , 
    n5732 , 
    n5733 , 
    n5734 , 
    n5735 , 
    n5736 , 
    n5737 , 
    n5738 , 
    n5739 , 
    n5740 , 
    n5741 , 
    n5742 , 
    n5743 , 
    n5744 , 
    n5745 , 
    n5746 , 
    n5747 , 
    n5748 , 
    n5749 , 
    n5750 , 
    n5751 , 
    n5752 , 
    n5753 , 
    n5754 , 
    n5755 , 
    n5756 , 
    n5757 , 
    n5758 , 
    n5759 , 
    n5760 , 
    n5761 , 
    n5762 , 
    n5763 , 
    n5764 , 
    n5765 , 
    n5766 , 
    n5767 , 
    n5768 , 
    n5769 , 
    n5770 , 
    n5771 , 
    n5772 , 
    n5773 , 
    n5774 , 
    n5775 , 
    n5776 , 
    n5777 , 
    n5778 , 
    n5779 , 
    n5780 , 
    n5781 , 
    n5782 , 
    n5783 , 
    n5784 , 
    n5785 , 
    n5786 , 
    n5787 , 
    n5788 , 
    n5789 , 
    n5790 , 
    n5791 , 
    n5792 , 
    n5793 , 
    n5794 , 
    n5795 , 
    n5796 , 
    n5797 , 
    n5798 , 
    n5799 , 
    n5800 , 
    n5801 , 
    n5802 , 
    n5803 , 
    n5804 , 
    n5805 , 
    n5806 , 
    n5807 , 
    n5808 , 
    n5809 , 
    n5810 , 
    n5811 , 
    n5812 , 
    n5813 , 
    n5814 , 
    n5815 , 
    n5816 , 
    n5817 , 
    n5818 , 
    n5819 , 
    n5820 , 
    n5821 , 
    n5822 , 
    n5823 , 
    n5824 , 
    n5825 , 
    n5826 , 
    n5827 , 
    n5828 , 
    n5829 , 
    n5830 , 
    n5831 , 
    n5832 , 
    n5833 , 
    n5834 , 
    n5835 , 
    n5836 , 
    n5837 , 
    n5838 , 
    n5839 , 
    n5840 , 
    n5841 , 
    n5842 , 
    n5843 , 
    n5844 , 
    n5845 , 
    n5846 , 
    n5847 , 
    n5848 , 
    n5849 , 
    n5850 , 
    n5851 , 
    n5852 , 
    n5853 , 
    n5854 , 
    n5855 , 
    n5856 , 
    n5857 , 
    n5858 , 
    n5859 , 
    n5860 , 
    n5861 , 
    n5862 , 
    n5863 , 
    n5864 , 
    n5865 , 
    n5866 , 
    n5867 , 
    n5868 , 
    n5869 , 
    n5870 , 
    n5871 , 
    n5872 , 
    n5873 , 
    n5874 , 
    n5875 , 
    n5876 , 
    n5877 , 
    n5878 , 
    n5879 , 
    n5880 , 
    n5881 , 
    n5882 , 
    n5883 , 
    n5884 , 
    n5885 , 
    n5886 , 
    n5887 , 
    n5888 , 
    n5889 , 
    n5890 , 
    n5891 , 
    n5892 , 
    n5893 , 
    n5894 , 
    n5895 , 
    n5896 , 
    n5897 , 
    n5898 , 
    n5899 , 
    n5900 , 
    n5901 , 
    n5902 , 
    n5903 , 
    n5904 , 
    n5905 , 
    n5906 , 
    n5907 , 
    n5908 , 
    n5909 , 
    n5910 , 
    n5911 , 
    n5912 , 
    n5913 , 
    n5914 , 
    n5915 , 
    n5916 , 
    n5917 , 
    n5918 , 
    n5919 , 
    n5920 , 
    n5921 , 
    n5922 , 
    n5923 , 
    n5924 , 
    n5925 , 
    n5926 , 
    n5927 , 
    n5928 , 
    n5929 , 
    n5930 , 
    n5931 , 
    n5932 , 
    n5933 , 
    n5934 , 
    n5935 , 
    n5936 , 
    n5937 , 
    n5938 , 
    n5939 , 
    n5940 , 
    n5941 , 
    n5942 , 
    n5943 , 
    n5944 , 
    n5945 , 
    n5946 , 
    n5947 , 
    n5948 , 
    n5949 , 
    n5950 , 
    n5951 , 
    n5952 , 
    n5953 , 
    n5954 , 
    n5955 , 
    n5956 , 
    n5957 , 
    n5958 , 
    n5959 , 
    n5960 , 
    n5961 , 
    n5962 , 
    n5963 , 
    n5964 , 
    n5965 , 
    n5966 , 
    n5967 , 
    n5968 , 
    n5969 , 
    n5970 , 
    n5971 , 
    n5972 , 
    n5973 , 
    n5974 , 
    n5975 , 
    n5976 , 
    n5977 , 
    n5978 , 
    n5979 , 
    n5980 , 
    n5981 , 
    n5982 , 
    n5983 , 
    n5984 , 
    n5985 , 
    n5986 , 
    n5987 , 
    n5988 , 
    n5989 , 
    n5990 , 
    n5991 , 
    n5992 , 
    n5993 , 
    n5994 , 
    n5995 , 
    n5996 , 
    n5997 , 
    n5998 , 
    n5999 , 
    n6000 , 
    n6001 , 
    n6002 , 
    n6003 , 
    n6004 , 
    n6005 , 
    n6006 , 
    n6007 , 
    n6008 , 
    n6009 , 
    n6010 , 
    n6011 , 
    n6012 , 
    n6013 , 
    n6014 , 
    n6015 , 
    n6016 , 
    n6017 , 
    n6018 , 
    n6019 , 
    n6020 , 
    n6021 , 
    n6022 , 
    n6023 , 
    n6024 , 
    n6025 , 
    n6026 , 
    n6027 , 
    n6028 , 
    n6029 , 
    n6030 , 
    n6031 , 
    n6032 , 
    n6033 , 
    n6034 , 
    n6035 , 
    n6036 , 
    n6037 , 
    n6038 , 
    n6039 , 
    n6040 , 
    n6041 , 
    n6042 , 
    n6043 , 
    n6044 , 
    n6045 , 
    n6046 , 
    n6047 , 
    n6048 , 
    n6049 , 
    n6050 , 
    n6051 , 
    n6052 , 
    n6053 , 
    n6054 , 
    n6055 , 
    n6056 , 
    n6057 , 
    n6058 , 
    n6059 , 
    n6060 , 
    n6061 , 
    n6062 , 
    n6063 , 
    n6064 , 
    n6065 , 
    n6066 , 
    n6067 , 
    n6068 , 
    n6069 , 
    n6070 , 
    n6071 , 
    n6072 , 
    n6073 , 
    n6074 , 
    n6075 , 
    n6076 , 
    n6077 , 
    n6078 , 
    n6079 , 
    n6080 , 
    n6081 , 
    n6082 , 
    n6083 , 
    n6084 , 
    n6085 , 
    n6086 , 
    n6087 , 
    n6088 , 
    n6089 , 
    n6090 , 
    n6091 , 
    n6092 , 
    n6093 , 
    n6094 , 
    n6095 , 
    n6096 , 
    n6097 , 
    n6098 , 
    n6099 , 
    n6100 , 
    n6101 , 
    n6102 , 
    n6103 , 
    n6104 , 
    n6105 , 
    n6106 , 
    n6107 , 
    n6108 , 
    n6109 , 
    n6110 , 
    n6111 , 
    n6112 , 
    n6113 , 
    n6114 , 
    n6115 , 
    n6116 , 
    n6117 , 
    n6118 , 
    n6119 , 
    n6120 , 
    n6121 , 
    n6122 , 
    n6123 , 
    n6124 , 
    n6125 , 
    n6126 , 
    n6127 , 
    n6128 , 
    n6129 , 
    n6130 , 
    n6131 , 
    n6132 , 
    n6133 , 
    n6134 , 
    n6135 , 
    n6136 , 
    n6137 , 
    n6138 , 
    n6139 , 
    n6140 , 
    n6141 , 
    n6142 , 
    n6143 , 
    n6144 , 
    n6145 , 
    n6146 , 
    n6147 , 
    n6148 , 
    n6149 , 
    n6150 , 
    n6151 , 
    n6152 , 
    n6153 , 
    n6154 , 
    n6155 , 
    n6156 , 
    n6157 , 
    n6158 , 
    n6159 , 
    n6160 , 
    n6161 , 
    n6162 , 
    n6163 , 
    n6164 , 
    n6165 , 
    n6166 , 
    n6167 , 
    n6168 , 
    n6169 , 
    n6170 , 
    n6171 , 
    n6172 , 
    n6173 , 
    n6174 , 
    n6175 , 
    n6176 , 
    n6177 , 
    n6178 , 
    n6179 , 
    n6180 , 
    n6181 , 
    n6182 , 
    n6183 , 
    n6184 , 
    n6185 , 
    n6186 , 
    n6187 , 
    n6188 , 
    n6189 , 
    n6190 , 
    n6191 , 
    n6192 , 
    n6193 , 
    n6194 , 
    n6195 , 
    n6196 , 
    n6197 , 
    n6198 , 
    n6199 , 
    n6200 , 
    n6201 , 
    n6202 , 
    n6203 , 
    n6204 , 
    n6205 , 
    n6206 , 
    n6207 , 
    n6208 , 
    n6209 , 
    n6210 , 
    n6211 , 
    n6212 , 
    n6213 , 
    n6214 , 
    n6215 , 
    n6216 , 
    n6217 , 
    n6218 , 
    n6219 , 
    n6220 , 
    n6221 , 
    n6222 , 
    n6223 , 
    n6224 , 
    n6225 , 
    n6226 , 
    n6227 , 
    n6228 , 
    n6229 , 
    n6230 , 
    n6231 , 
    n6232 , 
    n6233 , 
    n6234 , 
    n6235 , 
    n6236 , 
    n6237 , 
    n6238 , 
    n6239 , 
    n6240 , 
    n6241 , 
    n6242 , 
    n6243 , 
    n6244 , 
    n6245 , 
    n6246 , 
    n6247 , 
    n6248 , 
    n6249 , 
    n6250 , 
    n6251 , 
    n6252 , 
    n6253 , 
    n6254 , 
    n6255 , 
    n6256 , 
    n6257 , 
    n6258 , 
    n6259 , 
    n6260 , 
    n6261 , 
    n6262 , 
    n6263 , 
    n6264 , 
    n6265 , 
    n6266 , 
    n6267 , 
    n6268 , 
    n6269 , 
    n6270 , 
    n6271 , 
    n6272 , 
    n6273 , 
    n6274 , 
    n6275 , 
    n6276 , 
    n6277 , 
    n6278 , 
    n6279 , 
    n6280 , 
    n6281 , 
    n6282 , 
    n6283 , 
    n6284 , 
    n6285 , 
    n6286 , 
    n6287 , 
    n6288 , 
    n6289 , 
    n6290 , 
    n6291 , 
    n6292 , 
    n6293 , 
    n6294 , 
    n6295 , 
    n6296 , 
    n6297 , 
    n6298 , 
    n6299 , 
    n6300 , 
    n6301 , 
    n6302 , 
    n6303 , 
    n6304 , 
    n6305 , 
    n6306 , 
    n6307 , 
    n6308 , 
    n6309 , 
    n6310 , 
    n6311 , 
    n6312 , 
    n6313 , 
    n6314 , 
    n6315 , 
    n6316 , 
    n6317 , 
    n6318 , 
    n6319 , 
    n6320 , 
    n6321 , 
    n6322 , 
    n6323 , 
    n6324 , 
    n6325 , 
    n6326 , 
    n6327 , 
    n6328 , 
    n6329 , 
    n6330 , 
    n6331 , 
    n6332 , 
    n6333 , 
    n6334 , 
    n6335 , 
    n6336 , 
    n6337 , 
    n6338 , 
    n6339 , 
    n6340 , 
    n6341 , 
    n6342 , 
    n6343 , 
    n6344 , 
    n6345 , 
    n6346 , 
    n6347 , 
    n6348 , 
    n6349 , 
    n6350 , 
    n6351 , 
    n6352 , 
    n6353 , 
    n6354 , 
    n6355 , 
    n6356 , 
    n6357 , 
    n6358 , 
    n6359 , 
    n6360 , 
    n6361 , 
    n6362 , 
    n6363 , 
    n6364 , 
    n6365 , 
    n6366 , 
    n6367 , 
    n6368 , 
    n6369 , 
    n6370 , 
    n6371 , 
    n6372 , 
    n6373 , 
    n6374 , 
    n6375 , 
    n6376 , 
    n6377 , 
    n6378 , 
    n6379 , 
    n6380 , 
    n6381 , 
    n6382 , 
    n6383 , 
    n6384 , 
    n6385 , 
    n6386 , 
    n6387 , 
    n6388 , 
    n6389 , 
    n6390 , 
    n6391 , 
    n6392 , 
    n6393 , 
    n6394 , 
    n6395 , 
    n6396 , 
    n6397 , 
    n6398 , 
    n6399 , 
    n6400 , 
    n6401 , 
    n6402 , 
    n6403 , 
    n6404 , 
    n6405 , 
    n6406 , 
    n6407 , 
    n6408 , 
    n6409 , 
    n6410 , 
    n6411 , 
    n6412 , 
    n6413 , 
    n6414 , 
    n6415 , 
    n6416 , 
    n6417 , 
    n6418 , 
    n6419 , 
    n6420 , 
    n6421 , 
    n6422 , 
    n6423 , 
    n6424 , 
    n6425 , 
    n6426 , 
    n6427 , 
    n6428 , 
    n6429 , 
    n6430 , 
    n6431 , 
    n6432 , 
    n6433 , 
    n6434 , 
    n6435 , 
    n6436 , 
    n6437 , 
    n6438 , 
    n6439 , 
    n6440 , 
    n6441 , 
    n6442 , 
    n6443 , 
    n6444 , 
    n6445 , 
    n6446 , 
    n6447 , 
    n6448 , 
    n6449 , 
    n6450 , 
    n6451 , 
    n6452 , 
    n6453 , 
    n6454 , 
    n6455 , 
    n6456 , 
    n6457 , 
    n6458 , 
    n6459 , 
    n6460 , 
    n6461 , 
    n6462 , 
    n6463 , 
    n6464 , 
    n6465 , 
    n6466 , 
    n6467 , 
    n6468 , 
    n6469 , 
    n6470 , 
    n6471 , 
    n6472 , 
    n6473 , 
    n6474 , 
    n6475 , 
    n6476 , 
    n6477 , 
    n6478 , 
    n6479 , 
    n6480 , 
    n6481 , 
    n6482 , 
    n6483 , 
    n6484 , 
    n6485 , 
    n6486 , 
    n6487 , 
    n6488 , 
    n6489 , 
    n6490 , 
    n6491 , 
    n6492 , 
    n6493 , 
    n6494 , 
    n6495 , 
    n6496 , 
    n6497 , 
    n6498 , 
    n6499 , 
    n6500 , 
    n6501 , 
    n6502 , 
    n6503 , 
    n6504 , 
    n6505 , 
    n6506 , 
    n6507 , 
    n6508 , 
    n6509 , 
    n6510 , 
    n6511 , 
    n6512 , 
    n6513 , 
    n6514 , 
    n6515 , 
    n6516 , 
    n6517 , 
    n6518 , 
    n6519 , 
    n6520 , 
    n6521 , 
    n6522 , 
    n6523 , 
    n6524 , 
    n6525 , 
    n6526 , 
    n6527 , 
    n6528 , 
    n6529 , 
    n6530 , 
    n6531 , 
    n6532 , 
    n6533 , 
    n6534 , 
    n6535 , 
    n6536 , 
    n6537 , 
    n6538 , 
    n6539 , 
    n6540 , 
    n6541 , 
    n6542 , 
    n6543 , 
    n6544 , 
    n6545 , 
    n6546 , 
    n6547 , 
    n6548 , 
    n6549 , 
    n6550 , 
    n6551 , 
    n6552 , 
    n6553 , 
    n6554 , 
    n6555 , 
    n6556 , 
    n6557 , 
    n6558 , 
    n6559 , 
    n6560 , 
    n6561 , 
    n6562 , 
    n6563 , 
    n6564 , 
    n6565 , 
    n6566 , 
    n6567 , 
    n6568 , 
    n6569 , 
    n6570 , 
    n6571 , 
    n6572 , 
    n6573 , 
    n6574 , 
    n6575 , 
    n6576 , 
    n6577 , 
    n6578 , 
    n6579 , 
    n6580 , 
    n6581 , 
    n6582 , 
    n6583 , 
    n6584 , 
    n6585 , 
    n6586 , 
    n6587 , 
    n6588 , 
    n6589 , 
    n6590 , 
    n6591 , 
    n6592 , 
    n6593 , 
    n6594 , 
    n6595 , 
    n6596 , 
    n6597 , 
    n6598 , 
    n6599 , 
    n6600 , 
    n6601 , 
    n6602 , 
    n6603 , 
    n6604 , 
    n6605 , 
    n6606 , 
    n6607 , 
    n6608 , 
    n6609 , 
    n6610 , 
    n6611 , 
    n6612 , 
    n6613 , 
    n6614 , 
    n6615 , 
    n6616 , 
    n6617 , 
    n6618 , 
    n6619 , 
    n6620 , 
    n6621 , 
    n6622 , 
    n6623 , 
    n6624 , 
    n6625 , 
    n6626 , 
    n6627 , 
    n6628 , 
    n6629 , 
    n6630 , 
    n6631 , 
    n6632 , 
    n6633 , 
    n6634 , 
    n6635 , 
    n6636 , 
    n6637 , 
    n6638 , 
    n6639 , 
    n6640 , 
    n6641 , 
    n6642 , 
    n6643 , 
    n6644 , 
    n6645 , 
    n6646 , 
    n6647 , 
    n6648 , 
    n6649 , 
    n6650 , 
    n6651 , 
    n6652 , 
    n6653 , 
    n6654 , 
    n6655 , 
    n6656 , 
    n6657 , 
    n6658 , 
    n6659 , 
    n6660 , 
    n6661 , 
    n6662 , 
    n6663 , 
    n6664 , 
    n6665 , 
    n6666 , 
    n6667 , 
    n6668 , 
    n6669 , 
    n6670 , 
    n6671 , 
    n6672 , 
    n6673 , 
    n6674 , 
    n6675 , 
    n6676 , 
    n6677 , 
    n6678 , 
    n6679 , 
    n6680 , 
    n6681 , 
    n6682 , 
    n6683 , 
    n6684 , 
    n6685 , 
    n6686 , 
    n6687 , 
    n6688 , 
    n6689 , 
    n6690 , 
    n6691 , 
    n6692 , 
    n6693 , 
    n6694 , 
    n6695 , 
    n6696 , 
    n6697 , 
    n6698 , 
    n6699 , 
    n6700 , 
    n6701 , 
    n6702 , 
    n6703 , 
    n6704 , 
    n6705 , 
    n6706 , 
    n6707 , 
    n6708 , 
    n6709 , 
    n6710 , 
    n6711 , 
    n6712 , 
    n6713 , 
    n6714 , 
    n6715 , 
    n6716 , 
    n6717 , 
    n6718 , 
    n6719 , 
    n6720 , 
    n6721 , 
    n6722 , 
    n6723 , 
    n6724 , 
    n6725 , 
    n6726 , 
    n6727 , 
    n6728 , 
    n6729 , 
    n6730 , 
    n6731 , 
    n6732 , 
    n6733 , 
    n6734 , 
    n6735 , 
    n6736 , 
    n6737 , 
    n6738 , 
    n6739 , 
    n6740 , 
    n6741 , 
    n6742 , 
    n6743 , 
    n6744 , 
    n6745 , 
    n6746 , 
    n6747 , 
    n6748 , 
    n6749 , 
    n6750 , 
    n6751 , 
    n6752 , 
    n6753 , 
    n6754 , 
    n6755 , 
    n6756 , 
    n6757 , 
    n6758 , 
    n6759 , 
    n6760 );
input 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 ;
output 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 , 
    n5008 , 
    n5009 , 
    n5010 , 
    n5011 , 
    n5012 , 
    n5013 , 
    n5014 , 
    n5015 , 
    n5016 , 
    n5017 , 
    n5018 , 
    n5019 , 
    n5020 , 
    n5021 , 
    n5022 , 
    n5023 , 
    n5024 , 
    n5025 , 
    n5026 , 
    n5027 , 
    n5028 , 
    n5029 , 
    n5030 , 
    n5031 , 
    n5032 , 
    n5033 , 
    n5034 , 
    n5035 , 
    n5036 , 
    n5037 , 
    n5038 , 
    n5039 , 
    n5040 , 
    n5041 , 
    n5042 , 
    n5043 , 
    n5044 , 
    n5045 , 
    n5046 , 
    n5047 , 
    n5048 , 
    n5049 , 
    n5050 , 
    n5051 , 
    n5052 , 
    n5053 , 
    n5054 , 
    n5055 , 
    n5056 , 
    n5057 , 
    n5058 , 
    n5059 , 
    n5060 , 
    n5061 , 
    n5062 , 
    n5063 , 
    n5064 , 
    n5065 , 
    n5066 , 
    n5067 , 
    n5068 , 
    n5069 , 
    n5070 , 
    n5071 , 
    n5072 , 
    n5073 , 
    n5074 , 
    n5075 , 
    n5076 , 
    n5077 , 
    n5078 , 
    n5079 , 
    n5080 , 
    n5081 , 
    n5082 , 
    n5083 , 
    n5084 , 
    n5085 , 
    n5086 , 
    n5087 , 
    n5088 , 
    n5089 , 
    n5090 , 
    n5091 , 
    n5092 , 
    n5093 , 
    n5094 , 
    n5095 , 
    n5096 , 
    n5097 , 
    n5098 , 
    n5099 , 
    n5100 , 
    n5101 , 
    n5102 , 
    n5103 , 
    n5104 , 
    n5105 , 
    n5106 , 
    n5107 , 
    n5108 , 
    n5109 , 
    n5110 , 
    n5111 , 
    n5112 , 
    n5113 , 
    n5114 , 
    n5115 , 
    n5116 , 
    n5117 , 
    n5118 , 
    n5119 , 
    n5120 , 
    n5121 , 
    n5122 , 
    n5123 , 
    n5124 , 
    n5125 , 
    n5126 , 
    n5127 , 
    n5128 , 
    n5129 , 
    n5130 , 
    n5131 , 
    n5132 , 
    n5133 , 
    n5134 , 
    n5135 , 
    n5136 , 
    n5137 , 
    n5138 , 
    n5139 , 
    n5140 , 
    n5141 , 
    n5142 , 
    n5143 , 
    n5144 , 
    n5145 , 
    n5146 , 
    n5147 , 
    n5148 , 
    n5149 , 
    n5150 , 
    n5151 , 
    n5152 , 
    n5153 , 
    n5154 , 
    n5155 , 
    n5156 , 
    n5157 , 
    n5158 , 
    n5159 , 
    n5160 , 
    n5161 , 
    n5162 , 
    n5163 , 
    n5164 , 
    n5165 , 
    n5166 , 
    n5167 , 
    n5168 , 
    n5169 , 
    n5170 , 
    n5171 , 
    n5172 , 
    n5173 , 
    n5174 , 
    n5175 , 
    n5176 , 
    n5177 , 
    n5178 , 
    n5179 , 
    n5180 , 
    n5181 , 
    n5182 , 
    n5183 , 
    n5184 , 
    n5185 , 
    n5186 , 
    n5187 , 
    n5188 , 
    n5189 , 
    n5190 , 
    n5191 , 
    n5192 , 
    n5193 , 
    n5194 , 
    n5195 , 
    n5196 , 
    n5197 , 
    n5198 , 
    n5199 , 
    n5200 , 
    n5201 , 
    n5202 , 
    n5203 , 
    n5204 , 
    n5205 , 
    n5206 , 
    n5207 , 
    n5208 , 
    n5209 , 
    n5210 , 
    n5211 , 
    n5212 , 
    n5213 , 
    n5214 , 
    n5215 , 
    n5216 , 
    n5217 , 
    n5218 , 
    n5219 , 
    n5220 , 
    n5221 , 
    n5222 , 
    n5223 , 
    n5224 , 
    n5225 , 
    n5226 , 
    n5227 , 
    n5228 , 
    n5229 , 
    n5230 , 
    n5231 , 
    n5232 , 
    n5233 , 
    n5234 , 
    n5235 , 
    n5236 , 
    n5237 , 
    n5238 , 
    n5239 , 
    n5240 , 
    n5241 , 
    n5242 , 
    n5243 , 
    n5244 , 
    n5245 , 
    n5246 , 
    n5247 , 
    n5248 , 
    n5249 , 
    n5250 , 
    n5251 , 
    n5252 , 
    n5253 , 
    n5254 , 
    n5255 , 
    n5256 , 
    n5257 , 
    n5258 , 
    n5259 , 
    n5260 , 
    n5261 , 
    n5262 , 
    n5263 , 
    n5264 , 
    n5265 , 
    n5266 , 
    n5267 , 
    n5268 , 
    n5269 , 
    n5270 , 
    n5271 , 
    n5272 , 
    n5273 , 
    n5274 , 
    n5275 , 
    n5276 , 
    n5277 , 
    n5278 , 
    n5279 , 
    n5280 , 
    n5281 , 
    n5282 , 
    n5283 , 
    n5284 , 
    n5285 , 
    n5286 , 
    n5287 , 
    n5288 , 
    n5289 , 
    n5290 , 
    n5291 , 
    n5292 , 
    n5293 , 
    n5294 , 
    n5295 , 
    n5296 , 
    n5297 , 
    n5298 , 
    n5299 , 
    n5300 , 
    n5301 , 
    n5302 , 
    n5303 , 
    n5304 , 
    n5305 , 
    n5306 , 
    n5307 , 
    n5308 , 
    n5309 , 
    n5310 , 
    n5311 , 
    n5312 , 
    n5313 , 
    n5314 , 
    n5315 , 
    n5316 , 
    n5317 , 
    n5318 , 
    n5319 , 
    n5320 , 
    n5321 , 
    n5322 , 
    n5323 , 
    n5324 , 
    n5325 , 
    n5326 , 
    n5327 , 
    n5328 , 
    n5329 , 
    n5330 , 
    n5331 , 
    n5332 , 
    n5333 , 
    n5334 , 
    n5335 , 
    n5336 , 
    n5337 , 
    n5338 , 
    n5339 , 
    n5340 , 
    n5341 , 
    n5342 , 
    n5343 , 
    n5344 , 
    n5345 , 
    n5346 , 
    n5347 , 
    n5348 , 
    n5349 , 
    n5350 , 
    n5351 , 
    n5352 , 
    n5353 , 
    n5354 , 
    n5355 , 
    n5356 , 
    n5357 , 
    n5358 , 
    n5359 , 
    n5360 , 
    n5361 , 
    n5362 , 
    n5363 , 
    n5364 , 
    n5365 , 
    n5366 , 
    n5367 , 
    n5368 , 
    n5369 , 
    n5370 , 
    n5371 , 
    n5372 , 
    n5373 , 
    n5374 , 
    n5375 , 
    n5376 , 
    n5377 , 
    n5378 , 
    n5379 , 
    n5380 , 
    n5381 , 
    n5382 , 
    n5383 , 
    n5384 , 
    n5385 , 
    n5386 , 
    n5387 , 
    n5388 , 
    n5389 , 
    n5390 , 
    n5391 , 
    n5392 , 
    n5393 , 
    n5394 , 
    n5395 , 
    n5396 , 
    n5397 , 
    n5398 , 
    n5399 , 
    n5400 , 
    n5401 , 
    n5402 , 
    n5403 , 
    n5404 , 
    n5405 , 
    n5406 , 
    n5407 , 
    n5408 , 
    n5409 , 
    n5410 , 
    n5411 , 
    n5412 , 
    n5413 , 
    n5414 , 
    n5415 , 
    n5416 , 
    n5417 , 
    n5418 , 
    n5419 , 
    n5420 , 
    n5421 , 
    n5422 , 
    n5423 , 
    n5424 , 
    n5425 , 
    n5426 , 
    n5427 , 
    n5428 , 
    n5429 , 
    n5430 , 
    n5431 , 
    n5432 , 
    n5433 , 
    n5434 , 
    n5435 , 
    n5436 , 
    n5437 , 
    n5438 , 
    n5439 , 
    n5440 , 
    n5441 , 
    n5442 , 
    n5443 , 
    n5444 , 
    n5445 , 
    n5446 , 
    n5447 , 
    n5448 , 
    n5449 , 
    n5450 , 
    n5451 , 
    n5452 , 
    n5453 , 
    n5454 , 
    n5455 , 
    n5456 , 
    n5457 , 
    n5458 , 
    n5459 , 
    n5460 , 
    n5461 , 
    n5462 , 
    n5463 , 
    n5464 , 
    n5465 , 
    n5466 , 
    n5467 , 
    n5468 , 
    n5469 , 
    n5470 , 
    n5471 , 
    n5472 , 
    n5473 , 
    n5474 , 
    n5475 , 
    n5476 , 
    n5477 , 
    n5478 , 
    n5479 , 
    n5480 , 
    n5481 , 
    n5482 , 
    n5483 , 
    n5484 , 
    n5485 , 
    n5486 , 
    n5487 , 
    n5488 , 
    n5489 , 
    n5490 , 
    n5491 , 
    n5492 , 
    n5493 , 
    n5494 , 
    n5495 , 
    n5496 , 
    n5497 , 
    n5498 , 
    n5499 , 
    n5500 , 
    n5501 , 
    n5502 , 
    n5503 , 
    n5504 , 
    n5505 , 
    n5506 , 
    n5507 , 
    n5508 , 
    n5509 , 
    n5510 , 
    n5511 , 
    n5512 , 
    n5513 , 
    n5514 , 
    n5515 , 
    n5516 , 
    n5517 , 
    n5518 , 
    n5519 , 
    n5520 , 
    n5521 , 
    n5522 , 
    n5523 , 
    n5524 , 
    n5525 , 
    n5526 , 
    n5527 , 
    n5528 , 
    n5529 , 
    n5530 , 
    n5531 , 
    n5532 , 
    n5533 , 
    n5534 , 
    n5535 , 
    n5536 , 
    n5537 , 
    n5538 , 
    n5539 , 
    n5540 , 
    n5541 , 
    n5542 , 
    n5543 , 
    n5544 , 
    n5545 , 
    n5546 , 
    n5547 , 
    n5548 , 
    n5549 , 
    n5550 , 
    n5551 , 
    n5552 , 
    n5553 , 
    n5554 , 
    n5555 , 
    n5556 , 
    n5557 , 
    n5558 , 
    n5559 , 
    n5560 , 
    n5561 , 
    n5562 , 
    n5563 , 
    n5564 , 
    n5565 , 
    n5566 , 
    n5567 , 
    n5568 , 
    n5569 , 
    n5570 , 
    n5571 , 
    n5572 , 
    n5573 , 
    n5574 , 
    n5575 , 
    n5576 , 
    n5577 , 
    n5578 , 
    n5579 , 
    n5580 , 
    n5581 , 
    n5582 , 
    n5583 , 
    n5584 , 
    n5585 , 
    n5586 , 
    n5587 , 
    n5588 , 
    n5589 , 
    n5590 , 
    n5591 , 
    n5592 , 
    n5593 , 
    n5594 , 
    n5595 , 
    n5596 , 
    n5597 , 
    n5598 , 
    n5599 , 
    n5600 , 
    n5601 , 
    n5602 , 
    n5603 , 
    n5604 , 
    n5605 , 
    n5606 , 
    n5607 , 
    n5608 , 
    n5609 , 
    n5610 , 
    n5611 , 
    n5612 , 
    n5613 , 
    n5614 , 
    n5615 , 
    n5616 , 
    n5617 , 
    n5618 , 
    n5619 , 
    n5620 , 
    n5621 , 
    n5622 , 
    n5623 , 
    n5624 , 
    n5625 , 
    n5626 , 
    n5627 , 
    n5628 , 
    n5629 , 
    n5630 , 
    n5631 , 
    n5632 , 
    n5633 , 
    n5634 , 
    n5635 , 
    n5636 , 
    n5637 , 
    n5638 , 
    n5639 , 
    n5640 , 
    n5641 , 
    n5642 , 
    n5643 , 
    n5644 , 
    n5645 , 
    n5646 , 
    n5647 , 
    n5648 , 
    n5649 , 
    n5650 , 
    n5651 , 
    n5652 , 
    n5653 , 
    n5654 , 
    n5655 , 
    n5656 , 
    n5657 , 
    n5658 , 
    n5659 , 
    n5660 , 
    n5661 , 
    n5662 , 
    n5663 , 
    n5664 , 
    n5665 , 
    n5666 , 
    n5667 , 
    n5668 , 
    n5669 , 
    n5670 , 
    n5671 , 
    n5672 , 
    n5673 , 
    n5674 , 
    n5675 , 
    n5676 , 
    n5677 , 
    n5678 , 
    n5679 , 
    n5680 , 
    n5681 , 
    n5682 , 
    n5683 , 
    n5684 , 
    n5685 , 
    n5686 , 
    n5687 , 
    n5688 , 
    n5689 , 
    n5690 , 
    n5691 , 
    n5692 , 
    n5693 , 
    n5694 , 
    n5695 , 
    n5696 , 
    n5697 , 
    n5698 , 
    n5699 , 
    n5700 , 
    n5701 , 
    n5702 , 
    n5703 , 
    n5704 , 
    n5705 , 
    n5706 , 
    n5707 , 
    n5708 , 
    n5709 , 
    n5710 , 
    n5711 , 
    n5712 , 
    n5713 , 
    n5714 , 
    n5715 , 
    n5716 , 
    n5717 , 
    n5718 , 
    n5719 , 
    n5720 , 
    n5721 , 
    n5722 , 
    n5723 , 
    n5724 , 
    n5725 , 
    n5726 , 
    n5727 , 
    n5728 , 
    n5729 , 
    n5730 , 
    n5731 , 
    n5732 , 
    n5733 , 
    n5734 , 
    n5735 , 
    n5736 , 
    n5737 , 
    n5738 , 
    n5739 , 
    n5740 , 
    n5741 , 
    n5742 , 
    n5743 , 
    n5744 , 
    n5745 , 
    n5746 , 
    n5747 , 
    n5748 , 
    n5749 , 
    n5750 , 
    n5751 , 
    n5752 , 
    n5753 , 
    n5754 , 
    n5755 , 
    n5756 , 
    n5757 , 
    n5758 , 
    n5759 , 
    n5760 , 
    n5761 , 
    n5762 , 
    n5763 , 
    n5764 , 
    n5765 , 
    n5766 , 
    n5767 , 
    n5768 , 
    n5769 , 
    n5770 , 
    n5771 , 
    n5772 , 
    n5773 , 
    n5774 , 
    n5775 , 
    n5776 , 
    n5777 , 
    n5778 , 
    n5779 , 
    n5780 , 
    n5781 , 
    n5782 , 
    n5783 , 
    n5784 , 
    n5785 , 
    n5786 , 
    n5787 , 
    n5788 , 
    n5789 , 
    n5790 , 
    n5791 , 
    n5792 , 
    n5793 , 
    n5794 , 
    n5795 , 
    n5796 , 
    n5797 , 
    n5798 , 
    n5799 , 
    n5800 , 
    n5801 , 
    n5802 , 
    n5803 , 
    n5804 , 
    n5805 , 
    n5806 , 
    n5807 , 
    n5808 , 
    n5809 , 
    n5810 , 
    n5811 , 
    n5812 , 
    n5813 , 
    n5814 , 
    n5815 , 
    n5816 , 
    n5817 , 
    n5818 , 
    n5819 , 
    n5820 , 
    n5821 , 
    n5822 , 
    n5823 , 
    n5824 , 
    n5825 , 
    n5826 , 
    n5827 , 
    n5828 , 
    n5829 , 
    n5830 , 
    n5831 , 
    n5832 , 
    n5833 , 
    n5834 , 
    n5835 , 
    n5836 , 
    n5837 , 
    n5838 , 
    n5839 , 
    n5840 , 
    n5841 , 
    n5842 , 
    n5843 , 
    n5844 , 
    n5845 , 
    n5846 , 
    n5847 , 
    n5848 , 
    n5849 , 
    n5850 , 
    n5851 , 
    n5852 , 
    n5853 , 
    n5854 , 
    n5855 , 
    n5856 , 
    n5857 , 
    n5858 , 
    n5859 , 
    n5860 , 
    n5861 , 
    n5862 , 
    n5863 , 
    n5864 , 
    n5865 , 
    n5866 , 
    n5867 , 
    n5868 , 
    n5869 , 
    n5870 , 
    n5871 , 
    n5872 , 
    n5873 , 
    n5874 , 
    n5875 , 
    n5876 , 
    n5877 , 
    n5878 , 
    n5879 , 
    n5880 , 
    n5881 , 
    n5882 , 
    n5883 , 
    n5884 , 
    n5885 , 
    n5886 , 
    n5887 , 
    n5888 , 
    n5889 , 
    n5890 , 
    n5891 , 
    n5892 , 
    n5893 , 
    n5894 , 
    n5895 , 
    n5896 , 
    n5897 , 
    n5898 , 
    n5899 , 
    n5900 , 
    n5901 , 
    n5902 , 
    n5903 , 
    n5904 , 
    n5905 , 
    n5906 , 
    n5907 , 
    n5908 , 
    n5909 , 
    n5910 , 
    n5911 , 
    n5912 , 
    n5913 , 
    n5914 , 
    n5915 , 
    n5916 , 
    n5917 , 
    n5918 , 
    n5919 , 
    n5920 , 
    n5921 , 
    n5922 , 
    n5923 , 
    n5924 , 
    n5925 , 
    n5926 , 
    n5927 , 
    n5928 , 
    n5929 , 
    n5930 , 
    n5931 , 
    n5932 , 
    n5933 , 
    n5934 , 
    n5935 , 
    n5936 , 
    n5937 , 
    n5938 , 
    n5939 , 
    n5940 , 
    n5941 , 
    n5942 , 
    n5943 , 
    n5944 , 
    n5945 , 
    n5946 , 
    n5947 , 
    n5948 , 
    n5949 , 
    n5950 , 
    n5951 , 
    n5952 , 
    n5953 , 
    n5954 , 
    n5955 , 
    n5956 , 
    n5957 , 
    n5958 , 
    n5959 , 
    n5960 , 
    n5961 , 
    n5962 , 
    n5963 , 
    n5964 , 
    n5965 , 
    n5966 , 
    n5967 , 
    n5968 , 
    n5969 , 
    n5970 , 
    n5971 , 
    n5972 , 
    n5973 , 
    n5974 , 
    n5975 , 
    n5976 , 
    n5977 , 
    n5978 , 
    n5979 , 
    n5980 , 
    n5981 , 
    n5982 , 
    n5983 , 
    n5984 , 
    n5985 , 
    n5986 , 
    n5987 , 
    n5988 , 
    n5989 , 
    n5990 , 
    n5991 , 
    n5992 , 
    n5993 , 
    n5994 , 
    n5995 , 
    n5996 , 
    n5997 , 
    n5998 , 
    n5999 , 
    n6000 , 
    n6001 , 
    n6002 , 
    n6003 , 
    n6004 , 
    n6005 , 
    n6006 , 
    n6007 , 
    n6008 , 
    n6009 , 
    n6010 , 
    n6011 , 
    n6012 , 
    n6013 , 
    n6014 , 
    n6015 , 
    n6016 , 
    n6017 , 
    n6018 , 
    n6019 , 
    n6020 , 
    n6021 , 
    n6022 , 
    n6023 , 
    n6024 , 
    n6025 , 
    n6026 , 
    n6027 , 
    n6028 , 
    n6029 , 
    n6030 , 
    n6031 , 
    n6032 , 
    n6033 , 
    n6034 , 
    n6035 , 
    n6036 , 
    n6037 , 
    n6038 , 
    n6039 , 
    n6040 , 
    n6041 , 
    n6042 , 
    n6043 , 
    n6044 , 
    n6045 , 
    n6046 , 
    n6047 , 
    n6048 , 
    n6049 , 
    n6050 , 
    n6051 , 
    n6052 , 
    n6053 , 
    n6054 , 
    n6055 , 
    n6056 , 
    n6057 , 
    n6058 , 
    n6059 , 
    n6060 , 
    n6061 , 
    n6062 , 
    n6063 , 
    n6064 , 
    n6065 , 
    n6066 , 
    n6067 , 
    n6068 , 
    n6069 , 
    n6070 , 
    n6071 , 
    n6072 , 
    n6073 , 
    n6074 , 
    n6075 , 
    n6076 , 
    n6077 , 
    n6078 , 
    n6079 , 
    n6080 , 
    n6081 , 
    n6082 , 
    n6083 , 
    n6084 , 
    n6085 , 
    n6086 , 
    n6087 , 
    n6088 , 
    n6089 , 
    n6090 , 
    n6091 , 
    n6092 , 
    n6093 , 
    n6094 , 
    n6095 , 
    n6096 , 
    n6097 , 
    n6098 , 
    n6099 , 
    n6100 , 
    n6101 , 
    n6102 , 
    n6103 , 
    n6104 , 
    n6105 , 
    n6106 , 
    n6107 , 
    n6108 , 
    n6109 , 
    n6110 , 
    n6111 , 
    n6112 , 
    n6113 , 
    n6114 , 
    n6115 , 
    n6116 , 
    n6117 , 
    n6118 , 
    n6119 , 
    n6120 , 
    n6121 , 
    n6122 , 
    n6123 , 
    n6124 , 
    n6125 , 
    n6126 , 
    n6127 , 
    n6128 , 
    n6129 , 
    n6130 , 
    n6131 , 
    n6132 , 
    n6133 , 
    n6134 , 
    n6135 , 
    n6136 , 
    n6137 , 
    n6138 , 
    n6139 , 
    n6140 , 
    n6141 , 
    n6142 , 
    n6143 , 
    n6144 , 
    n6145 , 
    n6146 , 
    n6147 , 
    n6148 , 
    n6149 , 
    n6150 , 
    n6151 , 
    n6152 , 
    n6153 , 
    n6154 , 
    n6155 , 
    n6156 , 
    n6157 , 
    n6158 , 
    n6159 , 
    n6160 , 
    n6161 , 
    n6162 , 
    n6163 , 
    n6164 , 
    n6165 , 
    n6166 , 
    n6167 , 
    n6168 , 
    n6169 , 
    n6170 , 
    n6171 , 
    n6172 , 
    n6173 , 
    n6174 , 
    n6175 , 
    n6176 , 
    n6177 , 
    n6178 , 
    n6179 , 
    n6180 , 
    n6181 , 
    n6182 , 
    n6183 , 
    n6184 , 
    n6185 , 
    n6186 , 
    n6187 , 
    n6188 , 
    n6189 , 
    n6190 , 
    n6191 , 
    n6192 , 
    n6193 , 
    n6194 , 
    n6195 , 
    n6196 , 
    n6197 , 
    n6198 , 
    n6199 , 
    n6200 , 
    n6201 , 
    n6202 , 
    n6203 , 
    n6204 , 
    n6205 , 
    n6206 , 
    n6207 , 
    n6208 , 
    n6209 , 
    n6210 , 
    n6211 , 
    n6212 , 
    n6213 , 
    n6214 , 
    n6215 , 
    n6216 , 
    n6217 , 
    n6218 , 
    n6219 , 
    n6220 , 
    n6221 , 
    n6222 , 
    n6223 , 
    n6224 , 
    n6225 , 
    n6226 , 
    n6227 , 
    n6228 , 
    n6229 , 
    n6230 , 
    n6231 , 
    n6232 , 
    n6233 , 
    n6234 , 
    n6235 , 
    n6236 , 
    n6237 , 
    n6238 , 
    n6239 , 
    n6240 , 
    n6241 , 
    n6242 , 
    n6243 , 
    n6244 , 
    n6245 , 
    n6246 , 
    n6247 , 
    n6248 , 
    n6249 , 
    n6250 , 
    n6251 , 
    n6252 , 
    n6253 , 
    n6254 , 
    n6255 , 
    n6256 , 
    n6257 , 
    n6258 , 
    n6259 , 
    n6260 , 
    n6261 , 
    n6262 , 
    n6263 , 
    n6264 , 
    n6265 , 
    n6266 , 
    n6267 , 
    n6268 , 
    n6269 , 
    n6270 , 
    n6271 , 
    n6272 , 
    n6273 , 
    n6274 , 
    n6275 , 
    n6276 , 
    n6277 , 
    n6278 , 
    n6279 , 
    n6280 , 
    n6281 , 
    n6282 , 
    n6283 , 
    n6284 , 
    n6285 , 
    n6286 , 
    n6287 , 
    n6288 , 
    n6289 , 
    n6290 , 
    n6291 , 
    n6292 , 
    n6293 , 
    n6294 , 
    n6295 , 
    n6296 , 
    n6297 , 
    n6298 , 
    n6299 , 
    n6300 , 
    n6301 , 
    n6302 , 
    n6303 , 
    n6304 , 
    n6305 , 
    n6306 , 
    n6307 , 
    n6308 , 
    n6309 , 
    n6310 , 
    n6311 , 
    n6312 , 
    n6313 , 
    n6314 , 
    n6315 , 
    n6316 , 
    n6317 , 
    n6318 , 
    n6319 , 
    n6320 , 
    n6321 , 
    n6322 , 
    n6323 , 
    n6324 , 
    n6325 , 
    n6326 , 
    n6327 , 
    n6328 , 
    n6329 , 
    n6330 , 
    n6331 , 
    n6332 , 
    n6333 , 
    n6334 , 
    n6335 , 
    n6336 , 
    n6337 , 
    n6338 , 
    n6339 , 
    n6340 , 
    n6341 , 
    n6342 , 
    n6343 , 
    n6344 , 
    n6345 , 
    n6346 , 
    n6347 , 
    n6348 , 
    n6349 , 
    n6350 , 
    n6351 , 
    n6352 , 
    n6353 , 
    n6354 , 
    n6355 , 
    n6356 , 
    n6357 , 
    n6358 , 
    n6359 , 
    n6360 , 
    n6361 , 
    n6362 , 
    n6363 , 
    n6364 , 
    n6365 , 
    n6366 , 
    n6367 , 
    n6368 , 
    n6369 , 
    n6370 , 
    n6371 , 
    n6372 , 
    n6373 , 
    n6374 , 
    n6375 , 
    n6376 , 
    n6377 , 
    n6378 , 
    n6379 , 
    n6380 , 
    n6381 , 
    n6382 , 
    n6383 , 
    n6384 , 
    n6385 , 
    n6386 , 
    n6387 , 
    n6388 , 
    n6389 , 
    n6390 , 
    n6391 , 
    n6392 , 
    n6393 , 
    n6394 , 
    n6395 , 
    n6396 , 
    n6397 , 
    n6398 , 
    n6399 , 
    n6400 , 
    n6401 , 
    n6402 , 
    n6403 , 
    n6404 , 
    n6405 , 
    n6406 , 
    n6407 , 
    n6408 , 
    n6409 , 
    n6410 , 
    n6411 , 
    n6412 , 
    n6413 , 
    n6414 , 
    n6415 , 
    n6416 , 
    n6417 , 
    n6418 , 
    n6419 , 
    n6420 , 
    n6421 , 
    n6422 , 
    n6423 , 
    n6424 , 
    n6425 , 
    n6426 , 
    n6427 , 
    n6428 , 
    n6429 , 
    n6430 , 
    n6431 , 
    n6432 , 
    n6433 , 
    n6434 , 
    n6435 , 
    n6436 , 
    n6437 , 
    n6438 , 
    n6439 , 
    n6440 , 
    n6441 , 
    n6442 , 
    n6443 , 
    n6444 , 
    n6445 , 
    n6446 , 
    n6447 , 
    n6448 , 
    n6449 , 
    n6450 , 
    n6451 , 
    n6452 , 
    n6453 , 
    n6454 , 
    n6455 , 
    n6456 , 
    n6457 , 
    n6458 , 
    n6459 , 
    n6460 , 
    n6461 , 
    n6462 , 
    n6463 , 
    n6464 , 
    n6465 , 
    n6466 , 
    n6467 , 
    n6468 , 
    n6469 , 
    n6470 , 
    n6471 , 
    n6472 , 
    n6473 , 
    n6474 , 
    n6475 , 
    n6476 , 
    n6477 , 
    n6478 , 
    n6479 , 
    n6480 , 
    n6481 , 
    n6482 , 
    n6483 , 
    n6484 , 
    n6485 , 
    n6486 , 
    n6487 , 
    n6488 , 
    n6489 , 
    n6490 , 
    n6491 , 
    n6492 , 
    n6493 , 
    n6494 , 
    n6495 , 
    n6496 , 
    n6497 , 
    n6498 , 
    n6499 , 
    n6500 , 
    n6501 , 
    n6502 , 
    n6503 , 
    n6504 , 
    n6505 , 
    n6506 , 
    n6507 , 
    n6508 , 
    n6509 , 
    n6510 , 
    n6511 , 
    n6512 , 
    n6513 , 
    n6514 , 
    n6515 , 
    n6516 , 
    n6517 , 
    n6518 , 
    n6519 , 
    n6520 , 
    n6521 , 
    n6522 , 
    n6523 , 
    n6524 , 
    n6525 , 
    n6526 , 
    n6527 , 
    n6528 , 
    n6529 , 
    n6530 , 
    n6531 , 
    n6532 , 
    n6533 , 
    n6534 , 
    n6535 , 
    n6536 , 
    n6537 , 
    n6538 , 
    n6539 , 
    n6540 , 
    n6541 , 
    n6542 , 
    n6543 , 
    n6544 , 
    n6545 , 
    n6546 , 
    n6547 , 
    n6548 , 
    n6549 , 
    n6550 , 
    n6551 , 
    n6552 , 
    n6553 , 
    n6554 , 
    n6555 , 
    n6556 , 
    n6557 , 
    n6558 , 
    n6559 , 
    n6560 , 
    n6561 , 
    n6562 , 
    n6563 , 
    n6564 , 
    n6565 , 
    n6566 , 
    n6567 , 
    n6568 , 
    n6569 , 
    n6570 , 
    n6571 , 
    n6572 , 
    n6573 , 
    n6574 , 
    n6575 , 
    n6576 , 
    n6577 , 
    n6578 , 
    n6579 , 
    n6580 , 
    n6581 , 
    n6582 , 
    n6583 , 
    n6584 , 
    n6585 , 
    n6586 , 
    n6587 , 
    n6588 , 
    n6589 , 
    n6590 , 
    n6591 , 
    n6592 , 
    n6593 , 
    n6594 , 
    n6595 , 
    n6596 , 
    n6597 , 
    n6598 , 
    n6599 , 
    n6600 , 
    n6601 , 
    n6602 , 
    n6603 , 
    n6604 , 
    n6605 , 
    n6606 , 
    n6607 , 
    n6608 , 
    n6609 , 
    n6610 , 
    n6611 , 
    n6612 , 
    n6613 , 
    n6614 , 
    n6615 , 
    n6616 , 
    n6617 , 
    n6618 , 
    n6619 , 
    n6620 , 
    n6621 , 
    n6622 , 
    n6623 , 
    n6624 , 
    n6625 , 
    n6626 , 
    n6627 , 
    n6628 , 
    n6629 , 
    n6630 , 
    n6631 , 
    n6632 , 
    n6633 , 
    n6634 , 
    n6635 , 
    n6636 , 
    n6637 , 
    n6638 , 
    n6639 , 
    n6640 , 
    n6641 , 
    n6642 , 
    n6643 , 
    n6644 , 
    n6645 , 
    n6646 , 
    n6647 , 
    n6648 , 
    n6649 , 
    n6650 , 
    n6651 , 
    n6652 , 
    n6653 , 
    n6654 , 
    n6655 , 
    n6656 , 
    n6657 , 
    n6658 , 
    n6659 , 
    n6660 , 
    n6661 , 
    n6662 , 
    n6663 , 
    n6664 , 
    n6665 , 
    n6666 , 
    n6667 , 
    n6668 , 
    n6669 , 
    n6670 , 
    n6671 , 
    n6672 , 
    n6673 , 
    n6674 , 
    n6675 , 
    n6676 , 
    n6677 , 
    n6678 , 
    n6679 , 
    n6680 , 
    n6681 , 
    n6682 , 
    n6683 , 
    n6684 , 
    n6685 , 
    n6686 , 
    n6687 , 
    n6688 , 
    n6689 , 
    n6690 , 
    n6691 , 
    n6692 , 
    n6693 , 
    n6694 , 
    n6695 , 
    n6696 , 
    n6697 , 
    n6698 , 
    n6699 , 
    n6700 , 
    n6701 , 
    n6702 , 
    n6703 , 
    n6704 , 
    n6705 , 
    n6706 , 
    n6707 , 
    n6708 , 
    n6709 , 
    n6710 , 
    n6711 , 
    n6712 , 
    n6713 , 
    n6714 , 
    n6715 , 
    n6716 , 
    n6717 , 
    n6718 , 
    n6719 , 
    n6720 , 
    n6721 , 
    n6722 , 
    n6723 , 
    n6724 , 
    n6725 , 
    n6726 , 
    n6727 , 
    n6728 , 
    n6729 , 
    n6730 , 
    n6731 , 
    n6732 , 
    n6733 , 
    n6734 , 
    n6735 , 
    n6736 , 
    n6737 , 
    n6738 , 
    n6739 , 
    n6740 , 
    n6741 , 
    n6742 , 
    n6743 , 
    n6744 , 
    n6745 , 
    n6746 , 
    n6747 , 
    n6748 , 
    n6749 , 
    n6750 , 
    n6751 , 
    n6752 , 
    n6753 , 
    n6754 , 
    n6755 , 
    n6756 , 
    n6757 , 
    n6758 , 
    n6759 , 
    n6760 ;

wire  C0 , C1 , 
    RI15b3e9d0_1 , 
    RI15b56850_817 , 
    RI15b51120_631 , 
    RI15b51288_634 , 
    RI15b51198_632 , 
    RI15b51210_633 , 
    RI15b4c2d8_464 , 
    RI15b51030_629 , 
    RI15b4c260_463 , 
    RI15b50fb8_628 , 
    RI15b4c1e8_462 , 
    RI15b50f40_627 , 
    RI15b4c170_461 , 
    RI15b50ec8_626 , 
    RI15b4c0f8_460 , 
    RI15b50e50_625 , 
    RI15b57750_849 , 
    RI15b4fb90_585 , 
    RI15b4f7d0_577 , 
    RI15b4f410_569 , 
    RI15b4f050_561 , 
    RI15b4ec90_553 , 
    RI15b4e8d0_545 , 
    RI15b4e510_537 , 
    RI15b4e150_529 , 
    RI15b4dd90_521 , 
    RI15b4d9d0_513 , 
    RI15b4d610_505 , 
    RI15b4d250_497 , 
    RI15b4ce90_489 , 
    RI15b4cad0_481 , 
    RI15b4c710_473 , 
    RI15b4c350_465 , 
    RI15b4fc08_586 , 
    RI15b4f848_578 , 
    RI15b4f488_570 , 
    RI15b4f0c8_562 , 
    RI15b4ed08_554 , 
    RI15b4e948_546 , 
    RI15b4e588_538 , 
    RI15b4e1c8_530 , 
    RI15b4de08_522 , 
    RI15b4da48_514 , 
    RI15b4d688_506 , 
    RI15b4d2c8_498 , 
    RI15b4cf08_490 , 
    RI15b4cb48_482 , 
    RI15b4c788_474 , 
    RI15b4c3c8_466 , 
    RI15b4fc80_587 , 
    RI15b4f8c0_579 , 
    RI15b4f500_571 , 
    RI15b4f140_563 , 
    RI15b4ed80_555 , 
    RI15b4e9c0_547 , 
    RI15b4e600_539 , 
    RI15b4e240_531 , 
    RI15b4de80_523 , 
    RI15b4dac0_515 , 
    RI15b4d700_507 , 
    RI15b4d340_499 , 
    RI15b4cf80_491 , 
    RI15b4cbc0_483 , 
    RI15b4c800_475 , 
    RI15b4c440_467 , 
    RI15b4fcf8_588 , 
    RI15b4f938_580 , 
    RI15b4f578_572 , 
    RI15b4f1b8_564 , 
    RI15b4edf8_556 , 
    RI15b4ea38_548 , 
    RI15b4e678_540 , 
    RI15b4e2b8_532 , 
    RI15b4def8_524 , 
    RI15b4db38_516 , 
    RI15b4d778_508 , 
    RI15b4d3b8_500 , 
    RI15b4cff8_492 , 
    RI15b4cc38_484 , 
    RI15b4c878_476 , 
    RI15b4c4b8_468 , 
    RI15b4fd70_589 , 
    RI15b4f9b0_581 , 
    RI15b4f5f0_573 , 
    RI15b4f230_565 , 
    RI15b4ee70_557 , 
    RI15b4eab0_549 , 
    RI15b4e6f0_541 , 
    RI15b4e330_533 , 
    RI15b4df70_525 , 
    RI15b4dbb0_517 , 
    RI15b4d7f0_509 , 
    RI15b4d430_501 , 
    RI15b4d070_493 , 
    RI15b4ccb0_485 , 
    RI15b4c8f0_477 , 
    RI15b4c530_469 , 
    RI15b4fde8_590 , 
    RI15b4fa28_582 , 
    RI15b4f668_574 , 
    RI15b4f2a8_566 , 
    RI15b4eee8_558 , 
    RI15b4eb28_550 , 
    RI15b4e768_542 , 
    RI15b4e3a8_534 , 
    RI15b4dfe8_526 , 
    RI15b4dc28_518 , 
    RI15b4d868_510 , 
    RI15b4d4a8_502 , 
    RI15b4d0e8_494 , 
    RI15b4cd28_486 , 
    RI15b4c968_478 , 
    RI15b4c5a8_470 , 
    RI15b4fe60_591 , 
    RI15b4faa0_583 , 
    RI15b4f6e0_575 , 
    RI15b4f320_567 , 
    RI15b4ef60_559 , 
    RI15b4eba0_551 , 
    RI15b4e7e0_543 , 
    RI15b4e420_535 , 
    RI15b4e060_527 , 
    RI15b4dca0_519 , 
    RI15b4d8e0_511 , 
    RI15b4d520_503 , 
    RI15b4d160_495 , 
    RI15b4cda0_487 , 
    RI15b4c9e0_479 , 
    RI15b4c620_471 , 
    RI15b4fed8_592 , 
    RI15b4fb18_584 , 
    RI15b4f758_576 , 
    RI15b4f398_568 , 
    RI15b4efd8_560 , 
    RI15b4ec18_552 , 
    RI15b4e858_544 , 
    RI15b4e498_536 , 
    RI15b4e0d8_528 , 
    RI15b4dd18_520 , 
    RI15b4d958_512 , 
    RI15b4d598_504 , 
    RI15b4d1d8_496 , 
    RI15b4ce18_488 , 
    RI15b4ca58_480 , 
    RI15b4c698_472 , 
    RI15b54780_747 , 
    RI15b547f8_748 , 
    RI15b54870_749 , 
    RI15b667c8_1362 , 
    RI15b66840_1363 , 
    RI15b54690_745 , 
    RI15b55950_785 , 
    RI15b576d8_848 , 
    RI15b57660_847 , 
    RI15b56670_813 , 
    RI15b558d8_784 , 
    RI15b55860_783 , 
    RI15b557e8_782 , 
    RI15b57570_845 , 
    RI15b574f8_844 , 
    RI15b57480_843 , 
    RI15b57408_842 , 
    RI15b57390_841 , 
    RI15b57318_840 , 
    RI15b572a0_839 , 
    RI15b57228_838 , 
    RI15b571b0_837 , 
    RI15b57138_836 , 
    RI15b570c0_835 , 
    RI15b57048_834 , 
    RI15b56fd0_833 , 
    RI15b56f58_832 , 
    RI15b56ee0_831 , 
    RI15b56e68_830 , 
    RI15b56df0_829 , 
    RI15b56d78_828 , 
    RI15b56d00_827 , 
    RI15b56c88_826 , 
    RI15b56c10_825 , 
    RI15b56b98_824 , 
    RI15b56b20_823 , 
    RI15b56aa8_822 , 
    RI15b56a30_821 , 
    RI15b569b8_820 , 
    RI15b56940_819 , 
    RI15b568c8_818 , 
    RI15b567d8_816 , 
    RI15b56760_815 , 
    RI15b566e8_814 , 
    RI15b3ea48_2 , 
    RI15b58740_883 , 
    RI15b5d498_1048 , 
    RI15b586c8_882 , 
    RI15b5d420_1047 , 
    RI15b58650_881 , 
    RI15b5d3a8_1046 , 
    RI15b585d8_880 , 
    RI15b5d330_1045 , 
    RI15b58560_879 , 
    RI15b5d2b8_1044 , 
    RI15b62f10_1241 , 
    RI15b5c778_1020 , 
    RI15b5c700_1019 , 
    RI15b5c688_1018 , 
    RI15b5c610_1017 , 
    RI15b5c598_1016 , 
    RI15b5c520_1015 , 
    RI15b5c4a8_1014 , 
    RI15b5c430_1013 , 
    RI15b5c3b8_1012 , 
    RI15b5c340_1011 , 
    RI15b5bf80_1003 , 
    RI15b5bbc0_995 , 
    RI15b5b800_987 , 
    RI15b5b440_979 , 
    RI15b5b080_971 , 
    RI15b5acc0_963 , 
    RI15b5a900_955 , 
    RI15b5a540_947 , 
    RI15b5a180_939 , 
    RI15b59dc0_931 , 
    RI15b59a00_923 , 
    RI15b59640_915 , 
    RI15b59280_907 , 
    RI15b58ec0_899 , 
    RI15b58b00_891 , 
    RI15b5c2c8_1010 , 
    RI15b5bf08_1002 , 
    RI15b5bb48_994 , 
    RI15b5b788_986 , 
    RI15b5b3c8_978 , 
    RI15b5b008_970 , 
    RI15b5ac48_962 , 
    RI15b5a888_954 , 
    RI15b5a4c8_946 , 
    RI15b5a108_938 , 
    RI15b59d48_930 , 
    RI15b59988_922 , 
    RI15b595c8_914 , 
    RI15b59208_906 , 
    RI15b58e48_898 , 
    RI15b58a88_890 , 
    RI15b5c250_1009 , 
    RI15b5be90_1001 , 
    RI15b5bad0_993 , 
    RI15b5b710_985 , 
    RI15b5b350_977 , 
    RI15b5af90_969 , 
    RI15b5abd0_961 , 
    RI15b5a810_953 , 
    RI15b5a450_945 , 
    RI15b5a090_937 , 
    RI15b59cd0_929 , 
    RI15b59910_921 , 
    RI15b59550_913 , 
    RI15b59190_905 , 
    RI15b58dd0_897 , 
    RI15b58a10_889 , 
    RI15b5c1d8_1008 , 
    RI15b5be18_1000 , 
    RI15b5ba58_992 , 
    RI15b5b698_984 , 
    RI15b5b2d8_976 , 
    RI15b5af18_968 , 
    RI15b5ab58_960 , 
    RI15b5a798_952 , 
    RI15b5a3d8_944 , 
    RI15b5a018_936 , 
    RI15b59c58_928 , 
    RI15b59898_920 , 
    RI15b594d8_912 , 
    RI15b59118_904 , 
    RI15b58d58_896 , 
    RI15b58998_888 , 
    RI15b5c160_1007 , 
    RI15b5bda0_999 , 
    RI15b5b9e0_991 , 
    RI15b5b620_983 , 
    RI15b5b260_975 , 
    RI15b5aea0_967 , 
    RI15b5aae0_959 , 
    RI15b5a720_951 , 
    RI15b5a360_943 , 
    RI15b59fa0_935 , 
    RI15b59be0_927 , 
    RI15b59820_919 , 
    RI15b59460_911 , 
    RI15b590a0_903 , 
    RI15b58ce0_895 , 
    RI15b58920_887 , 
    RI15b5c0e8_1006 , 
    RI15b5bd28_998 , 
    RI15b5b968_990 , 
    RI15b5b5a8_982 , 
    RI15b5b1e8_974 , 
    RI15b5ae28_966 , 
    RI15b5aa68_958 , 
    RI15b5a6a8_950 , 
    RI15b5a2e8_942 , 
    RI15b59f28_934 , 
    RI15b59b68_926 , 
    RI15b597a8_918 , 
    RI15b593e8_910 , 
    RI15b59028_902 , 
    RI15b58c68_894 , 
    RI15b588a8_886 , 
    RI15b5c070_1005 , 
    RI15b5bcb0_997 , 
    RI15b5b8f0_989 , 
    RI15b5b530_981 , 
    RI15b5b170_973 , 
    RI15b5adb0_965 , 
    RI15b5a9f0_957 , 
    RI15b5a630_949 , 
    RI15b5a270_941 , 
    RI15b59eb0_933 , 
    RI15b59af0_925 , 
    RI15b59730_917 , 
    RI15b59370_909 , 
    RI15b58fb0_901 , 
    RI15b58bf0_893 , 
    RI15b58830_885 , 
    RI15b5bff8_1004 , 
    RI15b5bc38_996 , 
    RI15b5b878_988 , 
    RI15b5b4b8_980 , 
    RI15b5b0f8_972 , 
    RI15b5ad38_964 , 
    RI15b5a978_956 , 
    RI15b5a5b8_948 , 
    RI15b5a1f8_940 , 
    RI15b59e38_932 , 
    RI15b59a78_924 , 
    RI15b596b8_916 , 
    RI15b592f8_908 , 
    RI15b58f38_900 , 
    RI15b58b78_892 , 
    RI15b587b8_884 , 
    RI15b5d588_1050 , 
    RI15b5d6f0_1053 , 
    RI15b5d600_1051 , 
    RI15b5d678_1052 , 
    RI15b62e98_1240 , 
    RI15b62e20_1239 , 
    RI15b62da8_1238 , 
    RI15b62d30_1237 , 
    RI15b62cb8_1236 , 
    RI15b62c40_1235 , 
    RI15b62bc8_1234 , 
    RI15b606c0_1155 , 
    RI15b63e10_1273 , 
    RI15b4b090_425 , 
    RI15b44cb8_212 , 
    RI15b44e20_215 , 
    RI15b44d30_213 , 
    RI15b44da8_214 , 
    RI15b3fe70_45 , 
    RI15b44bc8_210 , 
    RI15b3fdf8_44 , 
    RI15b44b50_209 , 
    RI15b3fd80_43 , 
    RI15b44ad8_208 , 
    RI15b3fd08_42 , 
    RI15b44a60_207 , 
    RI15b3fc90_41 , 
    RI15b449e8_206 , 
    RI15b4bf90_457 , 
    RI15b43728_166 , 
    RI15b43368_158 , 
    RI15b42fa8_150 , 
    RI15b42be8_142 , 
    RI15b42828_134 , 
    RI15b42468_126 , 
    RI15b420a8_118 , 
    RI15b41ce8_110 , 
    RI15b41928_102 , 
    RI15b41568_94 , 
    RI15b411a8_86 , 
    RI15b40de8_78 , 
    RI15b40a28_70 , 
    RI15b40668_62 , 
    RI15b402a8_54 , 
    RI15b3fee8_46 , 
    RI15b437a0_167 , 
    RI15b433e0_159 , 
    RI15b43020_151 , 
    RI15b42c60_143 , 
    RI15b428a0_135 , 
    RI15b424e0_127 , 
    RI15b42120_119 , 
    RI15b41d60_111 , 
    RI15b419a0_103 , 
    RI15b415e0_95 , 
    RI15b41220_87 , 
    RI15b40e60_79 , 
    RI15b40aa0_71 , 
    RI15b406e0_63 , 
    RI15b40320_55 , 
    RI15b3ff60_47 , 
    RI15b43818_168 , 
    RI15b43458_160 , 
    RI15b43098_152 , 
    RI15b42cd8_144 , 
    RI15b42918_136 , 
    RI15b42558_128 , 
    RI15b42198_120 , 
    RI15b41dd8_112 , 
    RI15b41a18_104 , 
    RI15b41658_96 , 
    RI15b41298_88 , 
    RI15b40ed8_80 , 
    RI15b40b18_72 , 
    RI15b40758_64 , 
    RI15b40398_56 , 
    RI15b3ffd8_48 , 
    RI15b43890_169 , 
    RI15b434d0_161 , 
    RI15b43110_153 , 
    RI15b42d50_145 , 
    RI15b42990_137 , 
    RI15b425d0_129 , 
    RI15b42210_121 , 
    RI15b41e50_113 , 
    RI15b41a90_105 , 
    RI15b416d0_97 , 
    RI15b41310_89 , 
    RI15b40f50_81 , 
    RI15b40b90_73 , 
    RI15b407d0_65 , 
    RI15b40410_57 , 
    RI15b40050_49 , 
    RI15b43908_170 , 
    RI15b43548_162 , 
    RI15b43188_154 , 
    RI15b42dc8_146 , 
    RI15b42a08_138 , 
    RI15b42648_130 , 
    RI15b42288_122 , 
    RI15b41ec8_114 , 
    RI15b41b08_106 , 
    RI15b41748_98 , 
    RI15b41388_90 , 
    RI15b40fc8_82 , 
    RI15b40c08_74 , 
    RI15b40848_66 , 
    RI15b40488_58 , 
    RI15b400c8_50 , 
    RI15b43980_171 , 
    RI15b435c0_163 , 
    RI15b43200_155 , 
    RI15b42e40_147 , 
    RI15b42a80_139 , 
    RI15b426c0_131 , 
    RI15b42300_123 , 
    RI15b41f40_115 , 
    RI15b41b80_107 , 
    RI15b417c0_99 , 
    RI15b41400_91 , 
    RI15b41040_83 , 
    RI15b40c80_75 , 
    RI15b408c0_67 , 
    RI15b40500_59 , 
    RI15b40140_51 , 
    RI15b439f8_172 , 
    RI15b43638_164 , 
    RI15b43278_156 , 
    RI15b42eb8_148 , 
    RI15b42af8_140 , 
    RI15b42738_132 , 
    RI15b42378_124 , 
    RI15b41fb8_116 , 
    RI15b41bf8_108 , 
    RI15b41838_100 , 
    RI15b41478_92 , 
    RI15b410b8_84 , 
    RI15b40cf8_76 , 
    RI15b40938_68 , 
    RI15b40578_60 , 
    RI15b401b8_52 , 
    RI15b43a70_173 , 
    RI15b436b0_165 , 
    RI15b432f0_157 , 
    RI15b42f30_149 , 
    RI15b42b70_141 , 
    RI15b427b0_133 , 
    RI15b423f0_125 , 
    RI15b42030_117 , 
    RI15b41c70_109 , 
    RI15b418b0_101 , 
    RI15b414f0_93 , 
    RI15b41130_85 , 
    RI15b40d70_77 , 
    RI15b409b0_69 , 
    RI15b405f0_61 , 
    RI15b40230_53 , 
    RI15b48318_328 , 
    RI15b48390_329 , 
    RI15b48408_330 , 
    RI15b668b8_1364 , 
    RI15b3fba0_39 , 
    RI15b47df0_317 , 
    RI15b4a190_393 , 
    RI15b4bf18_456 , 
    RI15b4bea0_455 , 
    RI15b4be28_454 , 
    RI15b4bdb0_453 , 
    RI15b4bd38_452 , 
    RI15b4bcc0_451 , 
    RI15b4bc48_450 , 
    RI15b4bbd0_449 , 
    RI15b4bb58_448 , 
    RI15b4bae0_447 , 
    RI15b4ba68_446 , 
    RI15b4b9f0_445 , 
    RI15b4b978_444 , 
    RI15b4b900_443 , 
    RI15b4b888_442 , 
    RI15b4b810_441 , 
    RI15b4b798_440 , 
    RI15b4b720_439 , 
    RI15b4b6a8_438 , 
    RI15b4b630_437 , 
    RI15b4b5b8_436 , 
    RI15b4b540_435 , 
    RI15b4b4c8_434 , 
    RI15b4b450_433 , 
    RI15b4b3d8_432 , 
    RI15b4b360_431 , 
    RI15b4b2e8_430 , 
    RI15b4b270_429 , 
    RI15b4b1f8_428 , 
    RI15b4a208_394 , 
    RI15b4a118_392 , 
    RI15b4a0a0_391 , 
    RI15b4a028_390 , 
    RI15b49fb0_389 , 
    RI15b49f38_388 , 
    RI15b49ec0_387 , 
    RI15b49e48_386 , 
    RI15b49dd0_385 , 
    RI15b49d58_384 , 
    RI15b49ce0_383 , 
    RI15b49c68_382 , 
    RI15b49bf0_381 , 
    RI15b49b78_380 , 
    RI15b49b00_379 , 
    RI15b49a88_378 , 
    RI15b49a10_377 , 
    RI15b49998_376 , 
    RI15b49920_375 , 
    RI15b498a8_374 , 
    RI15b49830_373 , 
    RI15b497b8_372 , 
    RI15b49740_371 , 
    RI15b496c8_370 , 
    RI15b49650_369 , 
    RI15b495d8_368 , 
    RI15b49560_367 , 
    RI15b494e8_366 , 
    RI15b49470_365 , 
    RI15b493f8_364 , 
    RI15b49380_363 , 
    RI15b4b108_426 , 
    RI15b4b018_424 , 
    RI15b4afa0_423 , 
    RI15b4af28_422 , 
    RI15b4aeb0_421 , 
    RI15b4ae38_420 , 
    RI15b4adc0_419 , 
    RI15b4ad48_418 , 
    RI15b4acd0_417 , 
    RI15b4ac58_416 , 
    RI15b4abe0_415 , 
    RI15b4ab68_414 , 
    RI15b4aaf0_413 , 
    RI15b4aa78_412 , 
    RI15b4aa00_411 , 
    RI15b4a988_410 , 
    RI15b4a910_409 , 
    RI15b4a898_408 , 
    RI15b4a820_407 , 
    RI15b4a7a8_406 , 
    RI15b4a730_405 , 
    RI15b4a6b8_404 , 
    RI15b4a640_403 , 
    RI15b4a5c8_402 , 
    RI15b4a550_401 , 
    RI15b4a4d8_400 , 
    RI15b4a460_399 , 
    RI15b4a3e8_398 , 
    RI15b4a370_397 , 
    RI15b4a2f8_396 , 
    RI15b4a280_395 , 
    RI15b50928_614 , 
    RI15b508b0_613 , 
    RI15b50838_612 , 
    RI15b507c0_611 , 
    RI15b50748_610 , 
    RI15b506d0_609 , 
    RI15b50658_608 , 
    RI15b505e0_607 , 
    RI15b50568_606 , 
    RI15b504f0_605 , 
    RI15b50478_604 , 
    RI15b50400_603 , 
    RI15b50388_602 , 
    RI15b50310_601 , 
    RI15b50298_600 , 
    RI15b50220_599 , 
    RI15b501a8_598 , 
    RI15b50130_597 , 
    RI15b500b8_596 , 
    RI15b50040_595 , 
    RI15b4ffc8_594 , 
    RI15b4ff50_593 , 
    RI15b57fc0_867 , 
    RI15b57de0_863 , 
    RI15b55fe0_799 , 
    RI15b57d68_862 , 
    RI15b57cf0_861 , 
    RI15b57c78_860 , 
    RI15b57c00_859 , 
    RI15b57b88_858 , 
    RI15b57b10_857 , 
    RI15b57a98_856 , 
    RI15b57a20_855 , 
    RI15b579a8_854 , 
    RI15b57930_853 , 
    RI15b578b8_852 , 
    RI15b57840_851 , 
    RI15b577c8_850 , 
    RI15b55f68_798 , 
    RI15b55ef0_797 , 
    RI15b55e78_796 , 
    RI15b55e00_795 , 
    RI15b55d88_794 , 
    RI15b55d10_793 , 
    RI15b55c98_792 , 
    RI15b55c20_791 , 
    RI15b55ba8_790 , 
    RI15b55b30_789 , 
    RI15b55ab8_788 , 
    RI15b55a40_787 , 
    RI15b559c8_786 , 
    RI15b65850_1329 , 
    RI15b666d8_1360 , 
    RI15b658c8_1330 , 
    RI15b65940_1331 , 
    RI15b659b8_1332 , 
    RI15b65a30_1333 , 
    RI15b65aa8_1334 , 
    RI15b65b20_1335 , 
    RI15b65b98_1336 , 
    RI15b65fd0_1345 , 
    RI15b65f58_1344 , 
    RI15b65ee0_1343 , 
    RI15b65e68_1342 , 
    RI15b65df0_1341 , 
    RI15b65d78_1340 , 
    RI15b65d00_1339 , 
    RI15b65c88_1338 , 
    RI15b65c10_1337 , 
    RI15b66660_1359 , 
    RI15b665e8_1358 , 
    RI15b66570_1357 , 
    RI15b664f8_1356 , 
    RI15b66480_1355 , 
    RI15b66408_1354 , 
    RI15b66390_1353 , 
    RI15b66318_1352 , 
    RI15b662a0_1351 , 
    RI15b66228_1350 , 
    RI15b661b0_1349 , 
    RI15b66138_1348 , 
    RI15b660c0_1347 , 
    RI15b66048_1346 , 
    RI15b62b50_1233 , 
    RI15b63a50_1265 , 
    RI15b60be8_1166 , 
    RI15b60c60_1167 , 
    RI15b60cd8_1168 , 
    RI15b66750_1361 , 
    RI15b3fb28_38 , 
    RI15b61c50_1201 , 
    RI15b58470_877 , 
    RI15b583f8_876 , 
    RI15b58380_875 , 
    RI15b58308_874 , 
    RI15b58290_873 , 
    RI15b58218_872 , 
    RI15b581a0_871 , 
    RI15b58128_870 , 
    RI15b580b0_869 , 
    RI15b58038_868 , 
    RI15b57f48_866 , 
    RI15b57ed0_865 , 
    RI15b57e58_864 , 
    RI15b565f8_812 , 
    RI15b56580_811 , 
    RI15b56508_810 , 
    RI15b56490_809 , 
    RI15b56418_808 , 
    RI15b563a0_807 , 
    RI15b56328_806 , 
    RI15b562b0_805 , 
    RI15b56238_804 , 
    RI15b561c0_803 , 
    RI15b56148_802 , 
    RI15b560d0_801 , 
    RI15b56058_800 , 
    RI15b605d0_1153 , 
    RI15b60648_1154 , 
    RI15b54168_734 , 
    RI15b541e0_735 , 
    RI15b47d00_315 , 
    RI15b47d78_316 , 
    RI15b51558_640 , 
    RI15b450f0_221 , 
    RI15b4c008_458 , 
    RI15b63d98_1272 , 
    RI15b575e8_846 , 
    RI15b648d8_1296 , 
    RI15b63ac8_1266 , 
    RI15b64860_1295 , 
    RI15b647e8_1294 , 
    RI15b64770_1293 , 
    RI15b646f8_1292 , 
    RI15b64680_1291 , 
    RI15b64608_1290 , 
    RI15b64590_1289 , 
    RI15b64518_1288 , 
    RI15b644a0_1287 , 
    RI15b64428_1286 , 
    RI15b643b0_1285 , 
    RI15b64338_1284 , 
    RI15b642c0_1283 , 
    RI15b64248_1282 , 
    RI15b641d0_1281 , 
    RI15b64158_1280 , 
    RI15b640e0_1279 , 
    RI15b64068_1278 , 
    RI15b63ff0_1277 , 
    RI15b63f78_1276 , 
    RI15b63f00_1275 , 
    RI15b63e88_1274 , 
    RI15b63d20_1271 , 
    RI15b63ca8_1270 , 
    RI15b63c30_1269 , 
    RI15b63bb8_1268 , 
    RI15b63b40_1267 , 
    RI15b5d948_1058 , 
    RI15b467e8_270 , 
    RI15b48480_331 , 
    RI15b49308_362 , 
    RI15b484f8_332 , 
    RI15b48570_333 , 
    RI15b485e8_334 , 
    RI15b48660_335 , 
    RI15b486d8_336 , 
    RI15b48750_337 , 
    RI15b487c8_338 , 
    RI15b48840_339 , 
    RI15b488b8_340 , 
    RI15b48930_341 , 
    RI15b489a8_342 , 
    RI15b48a20_343 , 
    RI15b48a98_344 , 
    RI15b48b10_345 , 
    RI15b48b88_346 , 
    RI15b5e5f0_1085 , 
    RI15b5e6e0_1087 , 
    RI15b5d9c0_1059 , 
    RI15b5da38_1060 , 
    RI15b5dab0_1061 , 
    RI15b5db28_1062 , 
    RI15b5dba0_1063 , 
    RI15b5dc18_1064 , 
    RI15b5dc90_1065 , 
    RI15b5dd08_1066 , 
    RI15b5dd80_1067 , 
    RI15b5ddf8_1068 , 
    RI15b5de70_1069 , 
    RI15b5dee8_1070 , 
    RI15b5df60_1071 , 
    RI15b5dfd8_1072 , 
    RI15b5e050_1073 , 
    RI15b5e0c8_1074 , 
    RI15b5e140_1075 , 
    RI15b5e1b8_1076 , 
    RI15b5e230_1077 , 
    RI15b5e2a8_1078 , 
    RI15b5e320_1079 , 
    RI15b5e398_1080 , 
    RI15b5e410_1081 , 
    RI15b5e488_1082 , 
    RI15b5e500_1083 , 
    RI15b5e578_1084 , 
    RI15b5e668_1086 , 
    RI15b3f948_34 , 
    RI15b64950_1297 , 
    RI15b3eac0_3 , 
    RI15b657d8_1328 , 
    RI15b3f8d0_33 , 
    RI15b649c8_1298 , 
    RI15b3f858_32 , 
    RI15b64a40_1299 , 
    RI15b3f7e0_31 , 
    RI15b64ab8_1300 , 
    RI15b3f768_30 , 
    RI15b64b30_1301 , 
    RI15b3f6f0_29 , 
    RI15b64ba8_1302 , 
    RI15b3f678_28 , 
    RI15b64c20_1303 , 
    RI15b3f600_27 , 
    RI15b64c98_1304 , 
    RI15b3f1c8_18 , 
    RI15b650d0_1313 , 
    RI15b3f240_19 , 
    RI15b65058_1312 , 
    RI15b3f2b8_20 , 
    RI15b64fe0_1311 , 
    RI15b3f330_21 , 
    RI15b64f68_1310 , 
    RI15b3f3a8_22 , 
    RI15b64ef0_1309 , 
    RI15b3f420_23 , 
    RI15b64e78_1308 , 
    RI15b3f498_24 , 
    RI15b64e00_1307 , 
    RI15b3f510_25 , 
    RI15b64d88_1306 , 
    RI15b3f588_26 , 
    RI15b64d10_1305 , 
    RI15b3eb38_4 , 
    RI15b65760_1327 , 
    RI15b3ebb0_5 , 
    RI15b656e8_1326 , 
    RI15b3ec28_6 , 
    RI15b65670_1325 , 
    RI15b3eca0_7 , 
    RI15b655f8_1324 , 
    RI15b3ed18_8 , 
    RI15b65580_1323 , 
    RI15b3ed90_9 , 
    RI15b65508_1322 , 
    RI15b3ee08_10 , 
    RI15b65490_1321 , 
    RI15b3ee80_11 , 
    RI15b65418_1320 , 
    RI15b3eef8_12 , 
    RI15b653a0_1319 , 
    RI15b3ef70_13 , 
    RI15b65328_1318 , 
    RI15b3efe8_14 , 
    RI15b652b0_1317 , 
    RI15b3f060_15 , 
    RI15b65238_1316 , 
    RI15b3f0d8_16 , 
    RI15b651c0_1315 , 
    RI15b3f150_17 , 
    RI15b65148_1314 , 
    RI15b62f88_1242 , 
    RI15b5c7f0_1021 , 
    RI15b479b8_308 , 
    RI15b47b98_312 , 
    RI15b52278_668 , 
    RI15b52458_672 , 
    RI15b523e0_671 , 
    RI15b52368_670 , 
    RI15b522f0_669 , 
    RI15b51300_635 , 
    RI15b51378_636 , 
    RI15b513f0_637 , 
    RI15b51468_638 , 
    RI15b534c0_707 , 
    RI15b52f98_696 , 
    RI15b548e8_750 , 
    RI15b55770_781 , 
    RI15b54960_751 , 
    RI15b549d8_752 , 
    RI15b54a50_753 , 
    RI15b54ac8_754 , 
    RI15b54b40_755 , 
    RI15b54bb8_756 , 
    RI15b54c30_757 , 
    RI15b54ca8_758 , 
    RI15b54d20_759 , 
    RI15b54d98_760 , 
    RI15b54e10_761 , 
    RI15b54e88_762 , 
    RI15b54f00_763 , 
    RI15b54f78_764 , 
    RI15b54ff0_765 , 
    RI15b514e0_639 , 
    RI15b515d0_641 , 
    RI15b51648_642 , 
    RI15b516c0_643 , 
    RI15b51738_644 , 
    RI15b517b0_645 , 
    RI15b51828_646 , 
    RI15b518a0_647 , 
    RI15b51918_648 , 
    RI15b51990_649 , 
    RI15b51a08_650 , 
    RI15b51a80_651 , 
    RI15b51af8_652 , 
    RI15b51b70_653 , 
    RI15b51be8_654 , 
    RI15b51c60_655 , 
    RI15b51cd8_656 , 
    RI15b51d50_657 , 
    RI15b51dc8_658 , 
    RI15b51e40_659 , 
    RI15b51eb8_660 , 
    RI15b51f30_661 , 
    RI15b51fa8_662 , 
    RI15b52020_663 , 
    RI15b52098_664 , 
    RI15b52110_665 , 
    RI15b52188_666 , 
    RI15b52200_667 , 
    RI15b50b08_618 , 
    RI15b50a90_617 , 
    RI15b50a18_616 , 
    RI15b509a0_615 , 
    RI15b46e00_283 , 
    RI15b4b180_427 , 
    RI15b48228_326 , 
    RI15b482a0_327 , 
    RI15b45348_226 , 
    RI15b4c080_459 , 
    RI15b55680_779 , 
    RI15b55608_778 , 
    RI15b55590_777 , 
    RI15b55518_776 , 
    RI15b554a0_775 , 
    RI15b55428_774 , 
    RI15b553b0_773 , 
    RI15b55338_772 , 
    RI15b552c0_771 , 
    RI15b55248_770 , 
    RI15b551d0_769 , 
    RI15b55158_768 , 
    RI15b550e0_767 , 
    RI15b55068_766 , 
    RI15b52908_682 , 
    RI15b53f10_729 , 
    RI15b556f8_780 , 
    RI15b52b60_687 , 
    RI15b61d40_1203 , 
    RI15b62ad8_1232 , 
    RI15b61cc8_1202 , 
    RI15b639d8_1264 , 
    RI15b63960_1263 , 
    RI15b638e8_1262 , 
    RI15b63870_1261 , 
    RI15b637f8_1260 , 
    RI15b63780_1259 , 
    RI15b63708_1258 , 
    RI15b63690_1257 , 
    RI15b63618_1256 , 
    RI15b635a0_1255 , 
    RI15b63528_1254 , 
    RI15b634b0_1253 , 
    RI15b63438_1252 , 
    RI15b633c0_1251 , 
    RI15b63348_1250 , 
    RI15b632d0_1249 , 
    RI15b63258_1248 , 
    RI15b631e0_1247 , 
    RI15b63168_1246 , 
    RI15b630f0_1245 , 
    RI15b63078_1244 , 
    RI15b63000_1243 , 
    RI15b5f658_1120 , 
    RI15b5fdd8_1136 , 
    RI15b60d50_1169 , 
    RI15b61bd8_1200 , 
    RI15b60dc8_1170 , 
    RI15b60e40_1171 , 
    RI15b60eb8_1172 , 
    RI15b60f30_1173 , 
    RI15b60fa8_1174 , 
    RI15b61020_1175 , 
    RI15b61098_1176 , 
    RI15b61110_1177 , 
    RI15b61188_1178 , 
    RI15b61200_1179 , 
    RI15b61278_1180 , 
    RI15b612f0_1181 , 
    RI15b61368_1182 , 
    RI15b613e0_1183 , 
    RI15b61458_1184 , 
    RI15b62100_1211 , 
    RI15b62088_1210 , 
    RI15b62010_1209 , 
    RI15b61f98_1208 , 
    RI15b61f20_1207 , 
    RI15b61ea8_1206 , 
    RI15b61e30_1205 , 
    RI15b61db8_1204 , 
    RI15b45438_228 , 
    RI15b477d8_304 , 
    RI15b5cf70_1037 , 
    RI15b5cef8_1036 , 
    RI15b5ce80_1035 , 
    RI15b5ce08_1034 , 
    RI15b5cd90_1033 , 
    RI15b5cd18_1032 , 
    RI15b5cca0_1031 , 
    RI15b5cc28_1030 , 
    RI15b5cbb0_1029 , 
    RI15b5cb38_1028 , 
    RI15b5cac0_1027 , 
    RI15b5ca48_1026 , 
    RI15b5c9d0_1025 , 
    RI15b5c958_1024 , 
    RI15b5c8e0_1023 , 
    RI15b5c868_1022 , 
    RI15b5f388_1114 , 
    RI15b60738_1156 , 
    RI15b3f9c0_35 , 
    RI15b3fa38_36 , 
    RI15b60828_1158 , 
    RI15b5e848_1090 , 
    RI15b46950_273 , 
    RI15b470d0_289 , 
    RI15b44880_203 , 
    RI15b44808_202 , 
    RI15b44790_201 , 
    RI15b44718_200 , 
    RI15b446a0_199 , 
    RI15b44628_198 , 
    RI15b445b0_197 , 
    RI15b44538_196 , 
    RI15b444c0_195 , 
    RI15b44448_194 , 
    RI15b443d0_193 , 
    RI15b44358_192 , 
    RI15b442e0_191 , 
    RI15b44268_190 , 
    RI15b441f0_189 , 
    RI15b44178_188 , 
    RI15b44100_187 , 
    RI15b44088_186 , 
    RI15b44010_185 , 
    RI15b43f98_184 , 
    RI15b43f20_183 , 
    RI15b43ea8_182 , 
    RI15b43e30_181 , 
    RI15b43db8_180 , 
    RI15b43d40_179 , 
    RI15b43cc8_178 , 
    RI15b43c50_177 , 
    RI15b43bd8_176 , 
    RI15b43b60_175 , 
    RI15b43ae8_174 , 
    RI15b532e0_703 , 
    RI15b62a60_1231 , 
    RI15b629e8_1230 , 
    RI15b62970_1229 , 
    RI15b628f8_1228 , 
    RI15b62880_1227 , 
    RI15b62808_1226 , 
    RI15b62790_1225 , 
    RI15b62718_1224 , 
    RI15b626a0_1223 , 
    RI15b62628_1222 , 
    RI15b625b0_1221 , 
    RI15b62538_1220 , 
    RI15b624c0_1219 , 
    RI15b62448_1218 , 
    RI15b623d0_1217 , 
    RI15b62358_1216 , 
    RI15b622e0_1215 , 
    RI15b62268_1214 , 
    RI15b621f0_1213 , 
    RI15b62178_1212 , 
    RI15b5f6d0_1121 , 
    RI15b5d1c8_1042 , 
    RI15b5d150_1041 , 
    RI15b5d0d8_1040 , 
    RI15b5d060_1039 , 
    RI15b5cfe8_1038 , 
    RI15b45618_232 , 
    RI15b52c50_689 , 
    RI15b5e8c0_1091 , 
    RI15b5e7d0_1089 , 
    RI15b5e758_1088 , 
    RI15b5d768_1054 , 
    RI15b5d7e0_1055 , 
    RI15b5d858_1056 , 
    RI15b5d8d0_1057 , 
    RI15b53538_708 , 
    RI15b5f9a0_1127 , 
    RI15b5ec08_1098 , 
    RI15b614d0_1185 , 
    RI15b61b60_1199 , 
    RI15b61ae8_1198 , 
    RI15b61a70_1197 , 
    RI15b619f8_1196 , 
    RI15b61980_1195 , 
    RI15b61908_1194 , 
    RI15b61890_1193 , 
    RI15b61818_1192 , 
    RI15b617a0_1191 , 
    RI15b61728_1190 , 
    RI15b616b0_1189 , 
    RI15b61638_1188 , 
    RI15b615c0_1187 , 
    RI15b61548_1186 , 
    RI15b526b0_677 , 
    RI15b53100_699 , 
    RI15b52cc8_690 , 
    RI15b46ba8_278 , 
    RI15b52bd8_688 , 
    RI15b53f88_730 , 
    RI15b603f0_1149 , 
    RI15b45d98_248 , 
    RI15b50dd8_624 , 
    RI15b50d60_623 , 
    RI15b50ce8_622 , 
    RI15b50c70_621 , 
    RI15b50bf8_620 , 
    RI15b50b80_619 , 
    RI15b475f8_300 , 
    RI15b3fab0_37 , 
    RI15b45168_222 , 
    RI15b542d0_737 , 
    RI15b45ac8_242 , 
    RI15b527a0_679 , 
    RI15b53088_698 , 
    RI15b53808_714 , 
    RI15b5ee60_1103 , 
    RI15b60468_1150 , 
    RI15b54618_744 , 
    RI15b54708_746 , 
    RI15b46fe0_287 , 
    RI15b60918_1160 , 
    RI15b52d40_691 , 
    RI15b460e0_255 , 
    RI15b476e8_302 , 
    RI15b48c00_347 , 
    RI15b49290_361 , 
    RI15b49218_360 , 
    RI15b491a0_359 , 
    RI15b49128_358 , 
    RI15b490b0_357 , 
    RI15b49038_356 , 
    RI15b48fc0_355 , 
    RI15b48f48_354 , 
    RI15b48ed0_353 , 
    RI15b48e58_352 , 
    RI15b48de0_351 , 
    RI15b48d68_350 , 
    RI15b48cf0_349 , 
    RI15b48c78_348 , 
    RI15b52638_676 , 
    RI15b53c40_723 , 
    RI15b468d8_272 , 
    RI15b45ff0_253 , 
    RI15b45f78_252 , 
    RI15b45f00_251 , 
    RI15b45e88_250 , 
    RI15b44e98_216 , 
    RI15b44f10_217 , 
    RI15b44f88_218 , 
    RI15b45000_219 , 
    RI15b54258_736 , 
    RI15b53b50_721 , 
    RI15b5f0b8_1108 , 
    RI15b53da8_726 , 
    RI15b469c8_274 , 
    RI15b5f220_1111 , 
    RI15b47328_294 , 
    RI15b45a50_241 , 
    RI15b584e8_878 , 
    RI15b5d240_1043 , 
    RI15b52e30_693 , 
    RI15b535b0_709 , 
    RI15b53e20_727 , 
    RI15b60288_1146 , 
    RI15b3fc18_40 , 
    RI15b44970_205 , 
    RI15b448f8_204 , 
    RI15b608a0_1159 , 
    RI15b45780_235 , 
    RI15b525c0_675 , 
    RI15b47418_296 , 
    RI15b5f310_1113 , 
    RI15b44c40_211 , 
    RI15b46a40_275 , 
    RI15b60af8_1164 , 
    RI15b47f58_320 , 
    RI15b53718_712 , 
    RI15b5fb80_1131 , 
    RI15b52db8_692 , 
    RI15b45d20_247 , 
    RI15b52f20_695 , 
    RI15b47ee0_319 , 
    RI15b543c0_739 , 
    RI15b5ef50_1105 , 
    RI15b5ec80_1099 , 
    RI15b53448_706 , 
    RI15b529f8_684 , 
    RI15b54000_731 , 
    RI15b5f838_1124 , 
    RI15b53880_715 , 
    RI15b5fce8_1134 , 
    RI15b46d10_281 , 
    RI15b52890_681 , 
    RI15b5f5e0_1119 , 
    RI15b5fd60_1135 , 
    RI15b454b0_229 , 
    RI15b46860_271 , 
    RI15b46ab8_276 , 
    RI15b5f478_1116 , 
    RI15b540f0_733 , 
    RI15b60558_1152 , 
    RI15b47490_297 , 
    RI15b471c0_291 , 
    RI15b47238_292 , 
    RI15b53268_702 , 
    RI15b539e8_718 , 
    RI15b5f130_1109 , 
    RI15b5fb08_1130 , 
    RI15b607b0_1157 , 
    RI15b544b0_741 , 
    RI15b5eed8_1104 , 
    RI15b604e0_1151 , 
    RI15b510a8_630 , 
    RI15b463b0_261 , 
    RI15b46428_262 , 
    RI15b5f298_1112 , 
    RI15b5f1a8_1110 , 
    RI15b47a30_309 , 
    RI15b53bc8_722 , 
    RI15b46338_260 , 
    RI15b47c10_313 , 
    RI15b48048_322 , 
    RI15b464a0_263 , 
    RI15b5ecf8_1100 , 
    RI15b52ea8_694 , 
    RI15b53628_710 , 
    RI15b47850_305 , 
    RI15b46068_254 , 
    RI15b47670_301 , 
    RI15b524d0_673 , 
    RI15b53178_700 , 
    RI15b52ae8_686 , 
    RI15b451e0_223 , 
    RI15b52548_674 , 
    RI15b60030_1141 , 
    RI15b457f8_236 , 
    RI15b60990_1161 , 
    RI15b53ad8_720 , 
    RI15b5ff40_1139 , 
    RI15b45528_230 , 
    RI15b5fa18_1128 , 
    RI15b53358_704 , 
    RI15b5f7c0_1123 , 
    RI15b462c0_259 , 
    RI15b453c0_227 , 
    RI15b45870_237 , 
    RI15b46518_264 , 
    RI15b47058_288 , 
    RI15b60b70_1165 , 
    RI15b45bb8_244 , 
    RI15b533d0_705 , 
    RI15b47e68_318 , 
    RI15b47fd0_321 , 
    RI15b5f568_1118 , 
    RI15b480c0_323 , 
    RI15b45960_239 , 
    RI15b52980_683 , 
    RI15b53cb8_724 , 
    RI15b60120_1143 , 
    RI15b5f4f0_1117 , 
    RI15b46248_258 , 
    RI15b46e78_284 , 
    RI15b46590_265 , 
    RI15b5fe50_1137 , 
    RI15b47aa8_310 , 
    RI15b47b20_311 , 
    RI15b5efc8_1106 , 
    RI15b60378_1148 , 
    RI15b5ed70_1101 , 
    RI15b46c20_279 , 
    RI15b5d510_1049 , 
    RI15b45258_224 , 
    RI15b46f68_286 , 
    RI15b461d0_257 , 
    RI15b472b0_293 , 
    RI15b5f928_1126 , 
    RI15b536a0_711 , 
    RI15b45b40_243 , 
    RI15b48138_324 , 
    RI15b5f400_1115 , 
    RI15b46b30_277 , 
    RI15b46608_266 , 
    RI15b45690_233 , 
    RI15b53790_713 , 
    RI15b5fbf8_1132 , 
    RI15b54078_732 , 
    RI15b46c98_280 , 
    RI15b53e98_728 , 
    RI15b455a0_231 , 
    RI15b47940_307 , 
    RI15b45e10_249 , 
    RI15b5fa90_1129 , 
    RI15b54348_738 , 
    RI15b60a08_1162 , 
    RI15b531f0_701 , 
    RI15b60210_1145 , 
    RI15b478c8_306 , 
    RI15b47c88_314 , 
    RI15b46680_267 , 
    RI15b46158_256 , 
    RI15b5fc70_1133 , 
    RI15b53a60_719 , 
    RI15b538f8_716 , 
    RI15b5eb18_1096 , 
    RI15b5f040_1107 , 
    RI15b52728_678 , 
    RI15b5eaa0_1095 , 
    RI15b600a8_1142 , 
    RI15b5ede8_1102 , 
    RI15b5eb90_1097 , 
    RI15b60198_1144 , 
    RI15b481b0_325 , 
    RI15b545a0_743 , 
    RI15b452d0_225 , 
    RI15b46d88_282 , 
    RI15b5ea28_1094 , 
    RI15b54438_740 , 
    RI15b47508_298 , 
    RI15b466f8_268 , 
    RI15b47148_290 , 
    RI15b458e8_238 , 
    RI15b52a70_685 , 
    RI15b52818_680 , 
    RI15b5e9b0_1093 , 
    RI15b5ffb8_1140 , 
    RI15b5f8b0_1125 , 
    RI15b46ef0_285 , 
    RI15b45ca8_246 , 
    RI15b53970_717 , 
    RI15b47580_299 , 
    RI15b53010_697 , 
    RI15b5e938_1092 , 
    RI15b45078_220 , 
    RI15b60300_1147 , 
    RI15b46770_269 , 
    RI15b60a80_1163 , 
    RI15b473a0_295 , 
    RI15b47760_303 , 
    RI15b5f748_1122 , 
    RI15b5fec8_1138 , 
    RI15b45c30_245 , 
    RI15b53d30_725 , 
    RI15b45708_234 , 
    RI15b54528_742 , 
    RI15b459d8_240 , 
    R_187c_13cca558 , 
    R_125d_156aaaf8 , 
    R_c3e_13d2c178 , 
    R_61f_117eb278 , 
    R_187d_117f5b38 , 
    R_125e_13b8fe18 , 
    R_c3f_123b4358 , 
    R_187b_13ccb278 , 
    R_620_13dfb518 , 
    R_125c_15816b78 , 
    R_c3d_13c22918 , 
    R_61e_14a0c538 , 
    R_5e7_10080958 , 
    R_c06_170189e8 , 
    R_18b4_1162f978 , 
    R_1225_13c08298 , 
    R_1844_117ef378 , 
    R_1295_123bcf58 , 
    R_c76_15ff42e8 , 
    R_657_13bf5c78 , 
    R_187e_140ac0d8 , 
    R_125f_13c0f638 , 
    R_c40_1580a9b8 , 
    R_621_11c70318 , 
    R_187a_13ddd2d8 , 
    R_61d_123b84f8 , 
    R_125b_1162bf58 , 
    R_c3c_15ff9928 , 
    R_12be_13ccf378 , 
    R_5be_11c6a738 , 
    R_bdd_17016508 , 
    R_c9f_11636598 , 
    R_11fc_13ddf7b8 , 
    R_680_10085638 , 
    R_181b_13d430d8 , 
    R_18dd_13c062b8 , 
    R_180c_156b4eb8 , 
    R_12cd_13d535d8 , 
    R_5af_1700c3c8 , 
    R_cae_14a14ff8 , 
    R_bce_15ff4608 , 
    R_68f_13befcd8 , 
    R_18ec_13d204b8 , 
    R_11ed_116361d8 , 
    R_187f_15811038 , 
    R_1260_13d3b6f8 , 
    R_c41_14a0bef8 , 
    R_622_123b3bd8 , 
    R_61c_13d56378 , 
    R_c3b_150e7c58 , 
    R_1879_15ff5c88 , 
    R_125a_13bf58b8 , 
    R_f82_13c1cd38 , 
    R_963_13c209d8 , 
    R_8fa_117ec678 , 
    R_f19_15ff0648 , 
    R_1538_13d29bf8 , 
    R_15a1_150e22f8 , 
    R_158f_13cd9058 , 
    R_f70_17015608 , 
    R_951_156b2578 , 
    R_90c_13c0e0f8 , 
    R_f2b_140b8838 , 
    R_154a_1587f278 , 
    R_1880_13c22738 , 
    R_1261_13ccc0d8 , 
    R_c42_117eb818 , 
    R_623_140b3158 , 
    R_61b_11c70458 , 
    R_c3a_13b96218 , 
    R_1259_13d23578 , 
    R_1878_1162da38 , 
    R_ce6_14875d78 , 
    R_1924_13d1df38 , 
    R_11b5_13d56f58 , 
    R_577_1162c818 , 
    R_6c7_10082438 , 
    R_17d4_13cda278 , 
    R_1305_10081fd8 , 
    R_b96_15812b18 , 
    R_1881_156b0638 , 
    R_1262_12fc1698 , 
    R_c43_140b0138 , 
    R_624_13d421d8 , 
    R_61a_14b2a318 , 
    R_c39_117eaeb8 , 
    R_1258_117e8618 , 
    R_1877_1162cdb8 , 
    R_119b_15ffa3c8 , 
    R_55d_13b8e5b8 , 
    R_131f_158106d8 , 
    R_6e1_13c0fb38 , 
    R_17ba_15fed6c8 , 
    R_b7c_13b96e98 , 
    R_193e_123b6018 , 
    R_d00_117ec358 , 
    R_1323_13d5b878 , 
    R_6e5_15ff5328 , 
    R_559_13c024d8 , 
    R_1197_13bf4918 , 
    R_1942_11c6dd98 , 
    R_d04_14a16df8 , 
    R_17b6_13dec158 , 
    R_b78_13c10c18 , 
    R_13ca_13d2c718 , 
    R_19e9_13bf62b8 , 
    R_170f_150defb8 , 
    R_10f0_140b1ad8 , 
    R_ad1_11c6ac38 , 
    R_78c_13d5d3f8 , 
    R_dab_140b3dd8 , 
    R_883_13b936f8 , 
    R_ff9_11631958 , 
    R_ea2_150dd758 , 
    R_9da_13cd8018 , 
    R_1618_117f3658 , 
    R_14c1_123ba4d8 , 
    R_b5e_14a0f918 , 
    R_179c_123bb018 , 
    R_133d_13cd4e18 , 
    R_6ff_14a0a918 , 
    R_195c_150ddf78 , 
    R_117d_123b8c78 , 
    R_d1e_124c2cd8 , 
    R_5f7_12fbf758 , 
    R_c16_13df9858 , 
    R_1235_15880cb8 , 
    R_1854_1580fd78 , 
    R_18a4_13bf2d98 , 
    R_1285_100890f8 , 
    R_c66_13bed2f8 , 
    R_647_13d51af8 , 
    R_1882_13d1fbf8 , 
    R_1263_123be498 , 
    R_c44_13c229b8 , 
    R_625_13c1e638 , 
    R_619_156b6718 , 
    R_c38_117efd78 , 
    R_1257_14a0f0f8 , 
    R_1876_15ffcb28 , 
    R_985_1587c4d8 , 
    R_1516_12fc1eb8 , 
    R_15c3_13c02078 , 
    R_8d8_13d22fd8 , 
    R_fa4_13d1e898 , 
    R_ef7_1162bd78 , 
    R_1663_124c2698 , 
    R_838_1580b8b8 , 
    R_a25_13bf4ff8 , 
    R_1476_1486bd78 , 
    R_1044_13d57818 , 
    R_e57_13b8f738 , 
    R_15fa_13c0bb78 , 
    R_ec0_13c1bf78 , 
    R_fdb_15ff7308 , 
    R_14df_14a0cdf8 , 
    R_9bc_15812758 , 
    R_8a1_13d21818 , 
    R_1883_13d41058 , 
    R_1264_13c02758 , 
    R_c45_13d24c98 , 
    R_626_123b86d8 , 
    R_618_1587ea58 , 
    R_c37_13c0bfd8 , 
    R_1256_13d54258 , 
    R_1875_158179d8 , 
    R_1145_13b98658 , 
    R_737_116313b8 , 
    R_b26_1486a518 , 
    R_d56_117e9d38 , 
    R_1764_13ccf7d8 , 
    R_1375_13c275f8 , 
    R_1994_123bac58 , 
    R_143d_13bf2258 , 
    R_a5e_1587ed78 , 
    R_e1e_13c1bbb8 , 
    R_107d_15888418 , 
    R_7ff_13cd45f8 , 
    R_169c_15885fd8 , 
    R_1a5c_13de04d8 , 
    R_1a48_13c1ff38 , 
    R_a72_1486d358 , 
    R_1429_13d23438 , 
    R_1091_14a11d58 , 
    R_e0a_13bfa3b8 , 
    R_16b0_140aae18 , 
    R_7eb_123b8278 , 
    R_12c6_13cd49b8 , 
    R_5b6_117f1f38 , 
    R_ca7_140b4418 , 
    R_bd5_13d51698 , 
    R_688_13b99af8 , 
    R_11f4_13d1e6b8 , 
    R_18e5_13d45658 , 
    R_1813_13d29c98 , 
    R_16d9_14a17cf8 , 
    R_1a1f_11c70958 , 
    R_1400_14b29b98 , 
    R_de1_13cd0638 , 
    R_7c2_15ffa508 , 
    R_a9b_100865d8 , 
    R_10ba_15881938 , 
    R_1805_14b271b8 , 
    R_5a8_123b8318 , 
    R_cb5_170107e8 , 
    R_bc7_13c2a758 , 
    R_696_10082ed8 , 
    R_18f3_15ffc628 , 
    R_11e6_14b222f8 , 
    R_12d4_11634d38 , 
    R_119f_156b4738 , 
    R_561_1162a658 , 
    R_6dd_117f36f8 , 
    R_131b_15ff76c8 , 
    R_17be_15816538 , 
    R_b80_13cd8338 , 
    R_cfc_1700d2c8 , 
    R_193a_15885718 , 
    R_5da_13df70f8 , 
    R_18c1_11c6f738 , 
    R_bf9_13d28ed8 , 
    R_12a2_13bf2578 , 
    R_1218_13d28078 , 
    R_c83_13d59f78 , 
    R_1837_13deb9d8 , 
    R_664_123b47b8 , 
    R_e39_156b3518 , 
    R_a43_14b1feb8 , 
    R_81a_13cceb58 , 
    R_1062_117eedd8 , 
    R_1458_13df07f8 , 
    R_1681_140b99b8 , 
    R_1327_124c2b98 , 
    R_6e9_156b3158 , 
    R_555_13d59b18 , 
    R_1193_13b97438 , 
    R_1946_14a16858 , 
    R_d08_13d59938 , 
    R_b74_123c0478 , 
    R_17b2_13cd6498 , 
    R_113a_117eb458 , 
    R_742_14a129d8 , 
    R_b1b_11629758 , 
    R_d61_11633618 , 
    R_1380_15887338 , 
    R_1759_14874518 , 
    R_199f_13d3c9b8 , 
    R_1884_13cd1c18 , 
    R_1265_156b0818 , 
    R_c46_1580b598 , 
    R_627_117efb98 , 
    R_617_158807b8 , 
    R_c36_156b63f8 , 
    R_1255_1580dbb8 , 
    R_1874_13df9c18 , 
    R_87a_13c286d8 , 
    R_1002_14a17938 , 
    R_e99_123ba258 , 
    R_9e3_170110a8 , 
    R_1621_117eacd8 , 
    R_14b8_123b31d8 , 
    R_edf_117f5bd8 , 
    R_14fe_13d55518 , 
    R_15db_117f7258 , 
    R_fbc_13beb9f8 , 
    R_8c0_11631ef8 , 
    R_99d_13cd4d78 , 
    R_845_15888918 , 
    R_1656_117f4af8 , 
    R_1483_13d53d58 , 
    R_a18_12fbdef8 , 
    R_e64_14875058 , 
    R_1037_15815098 , 
    R_d8e_11630878 , 
    R_172c_13d39d58 , 
    R_13ad_14a12618 , 
    R_19cc_13cda1d8 , 
    R_110d_13dd5cb8 , 
    R_aee_117e9478 , 
    R_76f_117f4378 , 
    R_ccd_13b8c8f8 , 
    R_590_13dd64d8 , 
    R_17ed_156b36f8 , 
    R_190b_14872038 , 
    R_6ae_156ab958 , 
    R_baf_1700cd28 , 
    R_12ec_124c3778 , 
    R_11ce_11c6cad8 , 
    R_17a3_150e7398 , 
    R_1336_148754b8 , 
    R_6f8_13c1c018 , 
    R_1184_150e6498 , 
    R_1955_14b235b8 , 
    R_d17_14b27398 , 
    R_b65_13dde318 , 
    R_1885_1486cdb8 , 
    R_1266_14a12438 , 
    R_c47_100803b8 , 
    R_628_117eb098 , 
    R_616_170152e8 , 
    R_c35_123b88b8 , 
    R_1254_150e59f8 , 
    R_1873_12fc2278 , 
    R_74a_1008cb18 , 
    R_1132_15880e98 , 
    R_d69_14b23158 , 
    R_b13_140b3d38 , 
    R_1388_140aaf58 , 
    R_19a7_140b9b98 , 
    R_1751_1007feb8 , 
    R_b57_13ccd6b8 , 
    R_1344_117f3018 , 
    R_1795_1008b678 , 
    R_706_1580bd18 , 
    R_1963_13d1f478 , 
    R_1176_17015b08 , 
    R_d25_15882298 , 
    R_1590_150e4b98 , 
    R_f71_124c4998 , 
    R_952_14b26e98 , 
    R_90b_13d41af8 , 
    R_f2a_1162a158 , 
    R_1549_1587ff98 , 
    R_5c6_15816218 , 
    R_12b6_1587db58 , 
    R_be5_140b5818 , 
    R_c97_156b09f8 , 
    R_1204_13c23b38 , 
    R_678_15884ef8 , 
    R_1823_13d53df8 , 
    R_18d5_11636098 , 
    R_ed8_117e9c98 , 
    R_15e2_14a140f8 , 
    R_14f7_13b965d8 , 
    R_fc3_14b27e38 , 
    R_8b9_14875e18 , 
    R_9a4_117ee018 , 
    R_1a04_13c22b98 , 
    R_13e5_13de07f8 , 
    R_16f4_123b9fd8 , 
    R_dc6_14873f78 , 
    R_10d5_13b94a58 , 
    R_7a7_116355f8 , 
    R_ab6_15814e18 , 
    R_1886_11638c58 , 
    R_1267_14b23f18 , 
    R_c48_13bf5e58 , 
    R_629_150e7e38 , 
    R_615_13c1d7d8 , 
    R_c34_15ff1228 , 
    R_1253_13d222b8 , 
    R_1872_13ccb4f8 , 
    R_16f6_116389d8 , 
    R_10d7_156b5778 , 
    R_ab8_156ac8f8 , 
    R_1a02_13cd8298 , 
    R_13e3_14a0a7d8 , 
    R_7a5_13d456f8 , 
    R_dc4_11634b58 , 
    R_b4d_1700f208 , 
    R_710_156ac718 , 
    R_178b_1580ca38 , 
    R_196d_117eb8b8 , 
    R_d2f_13dedf58 , 
    R_116c_140b8338 , 
    R_134e_13d282f8 , 
    R_1a06_1486e1b8 , 
    R_13e7_116377b8 , 
    R_dc8_1162b058 , 
    R_7a9_123bd458 , 
    R_16f2_158857b8 , 
    R_ab4_12fbed58 , 
    R_10d3_158899f8 , 
    R_85a_156b1a38 , 
    R_1498_15811c18 , 
    R_1641_150db8b8 , 
    R_a03_123bd818 , 
    R_e79_13cd8658 , 
    R_1022_11c6cf38 , 
    R_150d_14b21678 , 
    R_15cc_14a0ba98 , 
    R_8cf_13ded9b8 , 
    R_fad_140ac038 , 
    R_eee_11632e98 , 
    R_98e_12fbecb8 , 
    R_13bd_13df6c98 , 
    R_19dc_156b6858 , 
    R_171c_117ecb78 , 
    R_10fd_117eef18 , 
    R_ade_13dd7658 , 
    R_77f_117f4558 , 
    R_d9e_13ddc3d8 , 
    R_16f8_14a0e018 , 
    R_10d9_123b9538 , 
    R_aba_13c29678 , 
    R_7a3_13ccb138 , 
    R_dc2_158108b8 , 
    R_13e1_156b8478 , 
    R_1a00_123b7f58 , 
    R_971_13df5618 , 
    R_8ec_123bbd38 , 
    R_15af_14866eb8 , 
    R_f0b_13cd72f8 , 
    R_f90_15812438 , 
    R_152a_13df8818 , 
    R_c15_15fee528 , 
    R_1234_15ff9e28 , 
    R_1853_13dd8738 , 
    R_18a5_170177c8 , 
    R_1286_124c4858 , 
    R_c67_13ccba98 , 
    R_648_15814058 , 
    R_5f6_13cce018 , 
    R_c05_14866d78 , 
    R_18b5_10087cf8 , 
    R_1224_13ccff58 , 
    R_1296_13dda7b8 , 
    R_1843_1580a878 , 
    R_c77_13d523b8 , 
    R_658_140ae1f8 , 
    R_5e6_13d46698 , 
    R_1a08_14b1b958 , 
    R_13e9_13d22358 , 
    R_dca_14b297d8 , 
    R_7ab_15887ab8 , 
    R_ab2_13df75f8 , 
    R_10d1_13d55d38 , 
    R_16f0_14b1e978 , 
    R_d87_123bae38 , 
    R_1733_15ff79e8 , 
    R_13a6_156b1718 , 
    R_1114_13d46ff8 , 
    R_19c5_13bf6ad8 , 
    R_af5_13c1b6b8 , 
    R_768_158896d8 , 
    R_964_123c1f58 , 
    R_8f9_117ee658 , 
    R_f18_14a19d78 , 
    R_1537_117e9b58 , 
    R_15a2_13ccce98 , 
    R_f83_14a0e978 , 
    R_1887_17018da8 , 
    R_1268_13d38278 , 
    R_c49_123b36d8 , 
    R_62a_13d42278 , 
    R_614_13c2a258 , 
    R_c33_150e7bb8 , 
    R_1252_116378f8 , 
    R_1871_13defad8 , 
    R_11a3_13c1be38 , 
    R_565_13ddbb18 , 
    R_6d9_11636818 , 
    R_1317_1580c5d8 , 
    R_17c2_13c03518 , 
    R_b84_156b5278 , 
    R_cf8_15881a78 , 
    R_1936_13d2a558 , 
    R_13b4_156abb38 , 
    R_19d3_13bf92d8 , 
    R_1725_13cd9a58 , 
    R_1106_14b1c718 , 
    R_ae7_13cd22f8 , 
    R_776_14873bb8 , 
    R_d95_15815778 , 
    R_feb_1486c818 , 
    R_eb0_13d53498 , 
    R_14cf_14b1bd18 , 
    R_9cc_158172f8 , 
    R_160a_17010ce8 , 
    R_891_13b8ab98 , 
    R_132b_1007f7d8 , 
    R_6ed_140b6538 , 
    R_118f_14b1ee78 , 
    R_194a_13d2ae18 , 
    R_d0c_13dee8b8 , 
    R_b70_13d20f58 , 
    R_17ae_13d29a18 , 
    R_1a3c_13b95278 , 
    R_109d_10084878 , 
    R_141d_13d441b8 , 
    R_16bc_14a0bdb8 , 
    R_dfe_15ff38e8 , 
    R_7df_1587d338 , 
    R_a7e_14a0bb38 , 
    R_151f_12fbe998 , 
    R_97c_13d528b8 , 
    R_15ba_1008b0d8 , 
    R_8e1_15889818 , 
    R_f00_17017ae8 , 
    R_f9b_13b974d8 , 
    R_16fa_14b299b8 , 
    R_10db_13cd6cb8 , 
    R_abc_15882b58 , 
    R_7a1_15ffcd08 , 
    R_dc0_117f53b8 , 
    R_13df_156b9238 , 
    R_19fe_13c01fd8 , 
    R_5cf_124c4678 , 
    R_12ad_13cca878 , 
    R_bee_156ac498 , 
    R_c8e_156b6cb8 , 
    R_120d_123be218 , 
    R_66f_13df8d18 , 
    R_182c_13b90598 , 
    R_18cc_170190c8 , 
    R_1505_13d27858 , 
    R_15d4_13d3a078 , 
    R_fb5_13c265b8 , 
    R_8c7_13ccf738 , 
    R_996_13cd1498 , 
    R_ee6_156ae158 , 
    R_1a0a_140b9238 , 
    R_13eb_150e7438 , 
    R_dcc_15815c78 , 
    R_7ad_1008c078 , 
    R_ab0_11629618 , 
    R_10cf_1580df78 , 
    R_16ee_123bf758 , 
    R_1660_13dd6258 , 
    R_83b_117f03b8 , 
    R_a22_156b92d8 , 
    R_1479_13ddc518 , 
    R_1041_14a0db18 , 
    R_e5a_11633118 , 
    R_1711_11c69d38 , 
    R_10f2_1486ad38 , 
    R_ad3_13d5a5b8 , 
    R_78a_13dfa2f8 , 
    R_da9_123bc9b8 , 
    R_13c8_11628e98 , 
    R_19e7_14a10098 , 
    R_eb5_13cd9cd8 , 
    R_fe6_13df1d38 , 
    R_14d4_13c27a58 , 
    R_9c7_140af5f8 , 
    R_896_123b6658 , 
    R_1605_156b1b78 , 
    R_1888_1580c858 , 
    R_1269_13b99c38 , 
    R_c4a_14a0cb78 , 
    R_62b_1162a1f8 , 
    R_613_124c47b8 , 
    R_c32_14b23518 , 
    R_1251_13d3fed8 , 
    R_1870_13b92bb8 , 
    R_16cc_156ba318 , 
    R_1a2c_156b08b8 , 
    R_140d_11638258 , 
    R_dee_13c0e058 , 
    R_7cf_123bbe78 , 
    R_a8e_170160a8 , 
    R_10ad_10082618 , 
    R_11b0_13b99f58 , 
    R_572_140ab458 , 
    R_6cc_117e8a78 , 
    R_130a_13dda498 , 
    R_17cf_13d389f8 , 
    R_b91_14b1f418 , 
    R_ceb_13d56d78 , 
    R_1929_13cd4af8 , 
    R_f72_13c2a1b8 , 
    R_953_14b20a98 , 
    R_90a_156ae658 , 
    R_f29_11630698 , 
    R_1548_140ac538 , 
    R_1591_13c25618 , 
    R_16fc_156b9a58 , 
    R_10dd_13d551f8 , 
    R_abe_14a15958 , 
    R_79f_140af7d8 , 
    R_dbe_13cd4c38 , 
    R_13dd_15884b38 , 
    R_19fc_13b96fd8 , 
    R_ff0_123b3b38 , 
    R_eab_11634518 , 
    R_9d1_13d4ed58 , 
    R_14ca_11631e58 , 
    R_160f_170102e8 , 
    R_88c_116319f8 , 
    R_e36_13c05b38 , 
    R_a46_11637e98 , 
    R_817_116294d8 , 
    R_1065_13c0b218 , 
    R_1455_117ef238 , 
    R_1684_13dd5ad8 , 
    R_e2b_13d28578 , 
    R_a51_11630ff8 , 
    R_80c_13d2acd8 , 
    R_1070_150e2d98 , 
    R_1a69_11c6fe18 , 
    R_168f_13d295b8 , 
    R_144a_1580c678 , 
    R_1a0c_13ccacd8 , 
    R_13ed_13cd4ff8 , 
    R_dce_14871f98 , 
    R_7af_11633578 , 
    R_aae_15814238 , 
    R_10cd_13d20878 , 
    R_16ec_13df6a18 , 
    R_1889_13bf9c38 , 
    R_126a_15886a78 , 
    R_c4b_13cd76b8 , 
    R_62c_10086038 , 
    R_612_10088dd8 , 
    R_c31_13b90778 , 
    R_1250_13d58c18 , 
    R_186f_1162dcb8 , 
    R_1a21_150e5598 , 
    R_1402_140b1cb8 , 
    R_de3_140b0778 , 
    R_7c4_13cd5138 , 
    R_a99_13cd0a98 , 
    R_10b8_13bea7d8 , 
    R_16d7_15888a58 , 
    R_b23_1587bc18 , 
    R_d59_14868cb8 , 
    R_1378_14b28158 , 
    R_1761_11631f98 , 
    R_1997_13d45158 , 
    R_1142_117f06d8 , 
    R_73a_13de1158 , 
    R_1a35_1486d7b8 , 
    R_16c3_13c01498 , 
    R_1416_1162ee38 , 
    R_df7_117f35b8 , 
    R_7d8_156abc78 , 
    R_a85_17014168 , 
    R_10a4_1486b0f8 , 
    R_a59_14a1a1d8 , 
    R_e23_13df5f78 , 
    R_1078_1580f558 , 
    R_804_156b6f38 , 
    R_1697_13d59d98 , 
    R_1a61_14a195f8 , 
    R_1442_14a18c98 , 
    R_1096_13dd6f78 , 
    R_1424_13b906d8 , 
    R_16b5_13c045f8 , 
    R_e05_140ad938 , 
    R_7e6_1486dd58 , 
    R_a77_100895f8 , 
    R_1a43_170104c8 , 
    R_15ef_15889318 , 
    R_ecb_13df7198 , 
    R_14ea_13cd2078 , 
    R_fd0_13cd59f8 , 
    R_8ac_15889278 , 
    R_9b1_1008a3b8 , 
    R_cc2_14a11218 , 
    R_17f8_13c28d18 , 
    R_59b_15812bb8 , 
    R_1900_1486c318 , 
    R_6a3_11c69658 , 
    R_bba_13deb7f8 , 
    R_12e1_123bbf18 , 
    R_11d9_14a18518 , 
    R_1125_124c3e58 , 
    R_d76_156b6218 , 
    R_b06_14b24af8 , 
    R_1395_13c0d978 , 
    R_19b4_14a10598 , 
    R_1744_11c6e3d8 , 
    R_757_13d3ceb8 , 
    R_16fe_123b51b8 , 
    R_10df_156b31f8 , 
    R_ac0_123c19b8 , 
    R_79d_13ddd698 , 
    R_dbc_13d207d8 , 
    R_13db_13d412d8 , 
    R_19fa_140afeb8 , 
    R_188a_14a0dd98 , 
    R_126b_170193e8 , 
    R_c4c_14874a18 , 
    R_62d_123c23b8 , 
    R_611_156aa558 , 
    R_c30_13cd8158 , 
    R_124f_13cd9418 , 
    R_186e_1162cb38 , 
    R_1233_13d5c318 , 
    R_1852_11635698 , 
    R_18a6_15885218 , 
    R_1287_13c29e98 , 
    R_c68_12fc1cd8 , 
    R_649_150e1f38 , 
    R_5f5_13bf7398 , 
    R_c14_13defe98 , 
    R_18c2_13d5d998 , 
    R_bf8_13bf77f8 , 
    R_12a3_14b20278 , 
    R_1217_123bdd18 , 
    R_c84_123bee98 , 
    R_1836_14a16038 , 
    R_665_117eefb8 , 
    R_5d9_15fed588 , 
    R_84f_1587bdf8 , 
    R_148d_156b2d98 , 
    R_164c_156b65d8 , 
    R_a0e_13cd5098 , 
    R_e6e_13c1e818 , 
    R_102d_14a14878 , 
    R_d7b_1007dbb8 , 
    R_1120_13cd3158 , 
    R_139a_12fbf398 , 
    R_b01_1587af98 , 
    R_19b9_116327b8 , 
    R_75c_13d54b18 , 
    R_173f_14a0d1b8 , 
    R_ca0_117f3978 , 
    R_bdc_14867a98 , 
    R_11fb_13d26638 , 
    R_681_13c02c58 , 
    R_18de_1162c638 , 
    R_181a_15887fb8 , 
    R_12bf_12fbe3f8 , 
    R_5bd_123b9678 , 
    R_1a0e_1486b698 , 
    R_13ef_156ba1d8 , 
    R_dd0_12fc0798 , 
    R_7b1_14a13478 , 
    R_aac_116311d8 , 
    R_10cb_150dccb8 , 
    R_16ea_140b6cb8 , 
    R_ffe_13ccf198 , 
    R_e9d_13d27038 , 
    R_9df_14a17398 , 
    R_161d_13b962b8 , 
    R_14bc_117f0598 , 
    R_87e_140b08b8 , 
    R_5a1_13d446b8 , 
    R_cbc_12fc1b98 , 
    R_bc0_13dfb338 , 
    R_69d_11c69798 , 
    R_18fa_140b5098 , 
    R_11df_15880998 , 
    R_12db_156b4af8 , 
    R_17fe_1580f5f8 , 
    R_191b_13c25f78 , 
    R_580_1162b4b8 , 
    R_6be_158101d8 , 
    R_17dd_14872358 , 
    R_12fc_15813dd8 , 
    R_b9f_140b49b8 , 
    R_cdd_13bf42d8 , 
    R_11be_150e4378 , 
    R_eba_13d29158 , 
    R_fe1_13d2bef8 , 
    R_14d9_13c21338 , 
    R_9c2_116297f8 , 
    R_89b_117ed118 , 
    R_1600_117e96f8 , 
    R_585_14a19b98 , 
    R_1916_150e99b8 , 
    R_17e2_123c1d78 , 
    R_6b9_150dc998 , 
    R_ba4_13c04d78 , 
    R_12f7_117f4ff8 , 
    R_11c3_117ee158 , 
    R_cd8_150deab8 , 
    R_15c4_13d46e18 , 
    R_8d7_13de10b8 , 
    R_fa5_13df4858 , 
    R_ef6_13c1f358 , 
    R_986_11631278 , 
    R_1515_13ccb8b8 , 
    R_11a7_123b9b78 , 
    R_569_12fbfd98 , 
    R_6d5_14b25958 , 
    R_1313_1587dab8 , 
    R_17c6_13d290b8 , 
    R_b88_14a0d9d8 , 
    R_cf4_13bea558 , 
    R_1932_13cd1538 , 
    R_1778_11631598 , 
    R_d42_1580f918 , 
    R_1159_148722b8 , 
    R_1361_14a18658 , 
    R_b3a_11637678 , 
    R_1980_15883a58 , 
    R_723_14a0aeb8 , 
    R_ec5_123c1eb8 , 
    R_fd6_15ff7448 , 
    R_14e4_14a121b8 , 
    R_9b7_117eaaf8 , 
    R_8a6_156b3018 , 
    R_15f5_140ade38 , 
    R_d45_117f4418 , 
    R_1775_140b5d18 , 
    R_1364_13c1d918 , 
    R_1156_15ff6fe8 , 
    R_1983_100863f8 , 
    R_726_13d39498 , 
    R_b37_10089b98 , 
    R_15e9_11636db8 , 
    R_14f0_13b92398 , 
    R_fca_156b44b8 , 
    R_8b2_11629078 , 
    R_9ab_14866698 , 
    R_ed1_158870b8 , 
    R_1632_117f1178 , 
    R_9f4_1486d2b8 , 
    R_e88_124c4498 , 
    R_1013_14a135b8 , 
    R_14a7_15814af8 , 
    R_869_14a19e18 , 
    R_132f_13c0b8f8 , 
    R_6f1_150df878 , 
    R_118b_14b27618 , 
    R_194e_14b236f8 , 
    R_d10_123b2d78 , 
    R_b6c_123b8138 , 
    R_17aa_13dfac58 , 
    R_188b_117e9978 , 
    R_126c_1580edd8 , 
    R_c4d_13d24b58 , 
    R_62e_13bf7438 , 
    R_610_14a186f8 , 
    R_c2f_14a0c038 , 
    R_124e_117ee338 , 
    R_186d_15fee348 , 
    R_e8c_1587e738 , 
    R_162e_123b25f8 , 
    R_9f0_140abe58 , 
    R_14ab_13dd50d8 , 
    R_86d_14a18dd8 , 
    R_100f_13d5dad8 , 
    R_8f8_15ff8668 , 
    R_f17_14a18e78 , 
    R_1536_14a0dc58 , 
    R_15a3_12fc08d8 , 
    R_f84_117e8d98 , 
    R_965_140b2578 , 
    R_d71_14b23018 , 
    R_b0b_13c21e78 , 
    R_1390_17016a08 , 
    R_19af_11636458 , 
    R_1749_117ec178 , 
    R_752_15ff64a8 , 
    R_112a_1587e0f8 , 
    R_18b6_13bf3018 , 
    R_1223_13dd8418 , 
    R_1297_13b99738 , 
    R_1842_123b43f8 , 
    R_c78_15887018 , 
    R_659_123b34f8 , 
    R_5e5_13df0578 , 
    R_c04_13cd6f38 , 
    R_954_17014988 , 
    R_909_13d3efd8 , 
    R_f28_13bf6fd8 , 
    R_1547_13df7b98 , 
    R_1592_156b9918 , 
    R_f73_13d22a38 , 
    R_70d_13beb098 , 
    R_178e_13c1cb58 , 
    R_196a_156b6d58 , 
    R_d2c_14a0ec98 , 
    R_116f_13d3e7b8 , 
    R_134b_15ff6cc8 , 
    R_b50_15815598 , 
    R_caf_156adc58 , 
    R_bcd_1162baf8 , 
    R_690_13c1e098 , 
    R_18ed_124c3278 , 
    R_11ec_1008d0b8 , 
    R_12ce_13c071b8 , 
    R_180b_1008abd8 , 
    R_5ae_13cd7ed8 , 
    R_177b_1007d6b8 , 
    R_d3f_13cd10d8 , 
    R_115c_150e8f18 , 
    R_135e_11c696f8 , 
    R_b3d_13dddeb8 , 
    R_720_13d395d8 , 
    R_197d_14a15458 , 
    R_1700_140ae8d8 , 
    R_10e1_13c07758 , 
    R_ac2_156ad2f8 , 
    R_79b_15886398 , 
    R_dba_116373f8 , 
    R_13d9_14a14378 , 
    R_19f8_117ef558 , 
    R_595_13def178 , 
    R_17f2_1580c998 , 
    R_1906_13ccad78 , 
    R_6a9_15ff4ba8 , 
    R_bb4_117f4d78 , 
    R_12e7_13cd42d8 , 
    R_11d3_1162b0f8 , 
    R_cc8_123b7738 , 
    R_d48_13c21c98 , 
    R_1772_14a16998 , 
    R_1367_15880858 , 
    R_1153_117f1678 , 
    R_1986_11c6c038 , 
    R_729_117f72f8 , 
    R_b34_158825b8 , 
    R_ff5_13c2a618 , 
    R_ea6_150dd7f8 , 
    R_9d6_13c01f38 , 
    R_14c5_14a0e518 , 
    R_1614_156b2b18 , 
    R_887_14a18298 , 
    R_848_13ddf218 , 
    R_1653_14869438 , 
    R_1486_156afe18 , 
    R_a15_1700ed08 , 
    R_e67_117f4e18 , 
    R_1034_156ac5d8 , 
    R_8eb_150db1d8 , 
    R_15b0_1580bdb8 , 
    R_f0a_14a0ce98 , 
    R_f91_117f6f38 , 
    R_1529_123bca58 , 
    R_972_13ccc038 , 
    R_1a10_123b4718 , 
    R_13f1_13d24298 , 
    R_dd2_14a19198 , 
    R_7b3_13c07938 , 
    R_aaa_13b8cfd8 , 
    R_10c9_15812a78 , 
    R_16e8_13cd8d38 , 
    R_d64_15ff5968 , 
    R_b18_117f40f8 , 
    R_1383_13c2a438 , 
    R_19a2_117f01d8 , 
    R_1756_123c0f18 , 
    R_1137_13d20ff8 , 
    R_745_13c1d5f8 , 
    R_1636_14b22618 , 
    R_9f8_13decdd8 , 
    R_e84_14875b98 , 
    R_1017_13d3bbf8 , 
    R_865_13d4e7b8 , 
    R_14a3_11c6d078 , 
    R_83e_13d43ad8 , 
    R_a1f_13d22d58 , 
    R_147c_1580d398 , 
    R_103e_13d57958 , 
    R_e5d_1486ddf8 , 
    R_165d_13bec038 , 
    R_1494_117f6718 , 
    R_1645_11c6c178 , 
    R_a07_14b251d8 , 
    R_e75_1580a5f8 , 
    R_1026_158103b8 , 
    R_856_13cd2a78 , 
    R_188c_13d39ad8 , 
    R_126d_11636638 , 
    R_c4e_13c0fe58 , 
    R_62f_116305f8 , 
    R_60f_13bf44b8 , 
    R_c2e_156b6c18 , 
    R_124d_123b5438 , 
    R_186c_15817758 , 
    R_57b_12fc1f58 , 
    R_6c3_14a11718 , 
    R_17d8_13bf24d8 , 
    R_1301_13ccee78 , 
    R_b9a_140b40f8 , 
    R_ce2_156b49b8 , 
    R_11b9_13d5d5d8 , 
    R_1920_117ea198 , 
    R_1713_14a0f878 , 
    R_10f4_13de4c18 , 
    R_ad5_117ed1b8 , 
    R_788_117e8ed8 , 
    R_da7_11635ff8 , 
    R_13c6_123c10f8 , 
    R_19e5_1580eb58 , 
    R_e90_11637038 , 
    R_9ec_117eb958 , 
    R_162a_117ec0d8 , 
    R_14af_156abdb8 , 
    R_871_1587f138 , 
    R_100b_11631d18 , 
    R_111b_1580faf8 , 
    R_139f_150df058 , 
    R_afc_117f8158 , 
    R_19be_13ccfff8 , 
    R_761_12fbf078 , 
    R_173a_156b5a98 , 
    R_d80_13c1d418 , 
    R_58a_13ddaf38 , 
    R_1911_124c4038 , 
    R_17e7_15883198 , 
    R_6b4_15881bb8 , 
    R_ba9_13d5c958 , 
    R_12f2_17013c68 , 
    R_11c8_11634fb8 , 
    R_cd3_13c06178 , 
    R_6fc_13de34f8 , 
    R_1180_13ddc298 , 
    R_1959_14a14698 , 
    R_d1b_13cd9558 , 
    R_b61_13d22538 , 
    R_179f_150e5818 , 
    R_133a_13d57138 , 
    R_be4_15817bb8 , 
    R_c98_13dec298 , 
    R_1203_1587d978 , 
    R_679_123b7918 , 
    R_1822_117e9018 , 
    R_18d6_13c2ad98 , 
    R_5c5_1162b5f8 , 
    R_12b7_117f83d8 , 
    R_ca8_14a11038 , 
    R_bd4_11637ad8 , 
    R_689_158869d8 , 
    R_11f3_116300f8 , 
    R_18e6_156b1678 , 
    R_1812_11c6f558 , 
    R_12c7_13b97c58 , 
    R_5b5_11637fd8 , 
    R_177e_14b1a738 , 
    R_d3c_13b8b278 , 
    R_115f_156ac7b8 , 
    R_135b_13d38b38 , 
    R_b40_158142d8 , 
    R_71d_13c1ea98 , 
    R_197a_13c0a318 , 
    R_e16_17018088 , 
    R_1085_13c03e78 , 
    R_7f7_15888b98 , 
    R_16a4_158821f8 , 
    R_1a54_13de0438 , 
    R_1435_10082258 , 
    R_a66_15882838 , 
    R_703_14867bd8 , 
    R_1960_1162c958 , 
    R_1179_13d3c7d8 , 
    R_d22_13d599d8 , 
    R_b5a_13bf68f8 , 
    R_1341_13d458d8 , 
    R_1798_1700e9e8 , 
    R_171e_13df60b8 , 
    R_10ff_13ddcab8 , 
    R_ae0_14a11f38 , 
    R_77d_13d27df8 , 
    R_d9c_13ccd4d8 , 
    R_13bb_1587d478 , 
    R_19da_13dd5a38 , 
    R_108a_1486e938 , 
    R_e11_13cd8c98 , 
    R_16a9_14a130b8 , 
    R_7f2_156b2938 , 
    R_1a4f_13d3a618 , 
    R_a6b_13b8e1f8 , 
    R_1430_13dd84b8 , 
    R_d4b_117f6178 , 
    R_176f_13d447f8 , 
    R_136a_13c26838 , 
    R_1150_15ff71c8 , 
    R_1989_13ccbc78 , 
    R_72c_10083c98 , 
    R_b31_13d44c58 , 
    R_814_13d51eb8 , 
    R_1068_1580ea18 , 
    R_1687_123b81d8 , 
    R_1452_13df0938 , 
    R_e33_14a0c3f8 , 
    R_a49_14a0eb58 , 
    R_1851_13d5b058 , 
    R_18a7_13b96858 , 
    R_1288_13c1daf8 , 
    R_c69_156af738 , 
    R_64a_11629438 , 
    R_5f4_140b13f8 , 
    R_c13_1162db78 , 
    R_1232_156aaa58 , 
    R_15bb_117f3338 , 
    R_8e0_14a0f698 , 
    R_f9c_14a104f8 , 
    R_eff_13d381d8 , 
    R_151e_15883af8 , 
    R_97d_14a16178 , 
    R_1702_13cd9198 , 
    R_10e3_117f2f78 , 
    R_ac4_1700f028 , 
    R_799_13d5a018 , 
    R_db8_150e6998 , 
    R_13d7_14b1d1b8 , 
    R_19f6_1580aa58 , 
    R_14fd_156b56d8 , 
    R_15dc_123bfd98 , 
    R_fbd_14a0b098 , 
    R_8bf_14875f58 , 
    R_99e_15ff9388 , 
    R_ede_11634338 , 
    R_188d_17018e48 , 
    R_126e_150e04f8 , 
    R_c4f_15814918 , 
    R_630_13d25558 , 
    R_60e_13cd3d38 , 
    R_c2d_1580aaf8 , 
    R_124c_13d40018 , 
    R_186b_13d42bd8 , 
    R_1a23_13d52458 , 
    R_1404_1486a8d8 , 
    R_de5_11633a78 , 
    R_7c6_156b9738 , 
    R_a97_13c05e58 , 
    R_10b6_124c3638 , 
    R_16d5_123bc4b8 , 
    R_bed_13b90db8 , 
    R_c8f_117ef4b8 , 
    R_120c_13ddcd38 , 
    R_670_13ccfaf8 , 
    R_182b_13cd80b8 , 
    R_18cd_13c1ca18 , 
    R_5ce_14b1ded8 , 
    R_12ae_13c1f178 , 
    R_bc6_13cd7bb8 , 
    R_697_13bf83d8 , 
    R_18f4_15881cf8 , 
    R_11e5_1162add8 , 
    R_12d5_17015928 , 
    R_1804_150e44b8 , 
    R_5a7_12fbe178 , 
    R_cb6_1162e398 , 
    R_110f_15887518 , 
    R_19ca_156b8a18 , 
    R_af0_17012a48 , 
    R_76d_156b1df8 , 
    R_d8c_15814b98 , 
    R_172e_117ed438 , 
    R_13ab_13b99878 , 
    R_1a12_13d52ef8 , 
    R_13f3_156b74d8 , 
    R_dd4_140ac5d8 , 
    R_7b5_13c1f718 , 
    R_aa8_14a0ea18 , 
    R_10c7_13df2c38 , 
    R_16e6_156b9eb8 , 
    R_15cd_13cd86f8 , 
    R_8ce_13d1e2f8 , 
    R_fae_13bf6df8 , 
    R_eed_15812578 , 
    R_98f_117f62b8 , 
    R_150c_15ff3848 , 
    R_908_123c0658 , 
    R_f27_13cd08b8 , 
    R_1546_14a18f18 , 
    R_1593_13d58e98 , 
    R_f74_158805d8 , 
    R_955_1580f0f8 , 
    R_d5c_1580ed38 , 
    R_137b_13d5cc78 , 
    R_175e_15813478 , 
    R_199a_117e8b18 , 
    R_113f_123b3098 , 
    R_73d_13c220f8 , 
    R_b20_13c06c18 , 
    R_163a_13d3ddb8 , 
    R_9fc_14a0b818 , 
    R_e80_11633ed8 , 
    R_101b_123b6518 , 
    R_861_124c3bd8 , 
    R_149f_123b5e38 , 
    R_1080_14a149b8 , 
    R_7fc_13d3f258 , 
    R_169f_124c2d78 , 
    R_1a59_117eded8 , 
    R_143a_14a0edd8 , 
    R_a61_1700dd68 , 
    R_e1b_13cd1178 , 
    R_140f_117f1cb8 , 
    R_df0_13c09cd8 , 
    R_7d1_14b28978 , 
    R_a8c_123c0338 , 
    R_10ab_13df0398 , 
    R_16ca_13d52f98 , 
    R_1a2e_13c22698 , 
    R_b10_14b21fd8 , 
    R_138b_156b0318 , 
    R_19aa_14a194b8 , 
    R_174e_15811a38 , 
    R_74d_117f0e58 , 
    R_112f_156aac38 , 
    R_d6c_156b62b8 , 
    R_1781_1162d5d8 , 
    R_d39_15811b78 , 
    R_1162_124c2558 , 
    R_1358_156b8e78 , 
    R_b43_13c06858 , 
    R_71a_117ee798 , 
    R_1977_15880b78 , 
    R_1108_13ccfb98 , 
    R_ae9_1580cd58 , 
    R_774_1700a7a8 , 
    R_d93_13cce0b8 , 
    R_13b2_15886898 , 
    R_1727_14870e18 , 
    R_19d1_123b5b18 , 
    R_188e_11c6a698 , 
    R_126f_14b23c98 , 
    R_c50_13d471d8 , 
    R_631_13ddd7d8 , 
    R_60d_117f3a18 , 
    R_c2c_13d2c498 , 
    R_124b_156b97d8 , 
    R_186a_13ddb118 , 
    R_fdc_1162ca98 , 
    R_14de_13c202f8 , 
    R_9bd_11632cb8 , 
    R_8a0_13bf81f8 , 
    R_15fb_123ba078 , 
    R_ebf_13b91678 , 
    R_e94_148719f8 , 
    R_9e8_15ff97e8 , 
    R_1626_13de2918 , 
    R_14b3_13dde9f8 , 
    R_875_156aea18 , 
    R_1007_15881578 , 
    R_14f6_11638938 , 
    R_fc4_1580d578 , 
    R_8b8_123ba2f8 , 
    R_9a5_117ecc18 , 
    R_ed7_14a0da78 , 
    R_15e3_123c0158 , 
    R_e0c_1700d0e8 , 
    R_16ae_123b38b8 , 
    R_7ed_117ef738 , 
    R_1a4a_12fc1c38 , 
    R_a70_150dbc78 , 
    R_142b_15889bd8 , 
    R_108f_13de36d8 , 
    R_d4e_11c6b6d8 , 
    R_176c_13ddfcb8 , 
    R_136d_11634dd8 , 
    R_114d_158861b8 , 
    R_198c_13d53a38 , 
    R_72f_11637498 , 
    R_b2e_170098a8 , 
    R_8f7_13b8e298 , 
    R_f16_1587d838 , 
    R_1535_13ded2d8 , 
    R_15a4_1162bcd8 , 
    R_f85_170174a8 , 
    R_966_156acd58 , 
    R_12a4_13cd0db8 , 
    R_1216_13c26518 , 
    R_c85_13d505b8 , 
    R_1835_13b8eb58 , 
    R_666_13cd8798 , 
    R_5d8_14a11fd8 , 
    R_18c3_156b8c98 , 
    R_bf7_156b4418 , 
    R_15d5_117ed898 , 
    R_fb6_14b24558 , 
    R_8c6_13d442f8 , 
    R_997_123bb478 , 
    R_ee5_14a14af8 , 
    R_1504_13d553d8 , 
    R_6d1_158167b8 , 
    R_130f_156ab4f8 , 
    R_17ca_150df9b8 , 
    R_b8c_124c3ef8 , 
    R_cf0_11c6a878 , 
    R_192e_150e8a18 , 
    R_11ab_13d29d38 , 
    R_56d_156b76b8 , 
    R_1704_13bf4238 , 
    R_10e5_14871778 , 
    R_ac6_1587bcb8 , 
    R_797_14b1c178 , 
    R_db6_13ddd058 , 
    R_13d5_1587c618 , 
    R_19f4_150e3ab8 , 
    R_1298_156b1d58 , 
    R_1841_13d2c538 , 
    R_c79_156b5598 , 
    R_65a_14874ab8 , 
    R_5e4_13bf0278 , 
    R_c03_14a0d2f8 , 
    R_18b7_13ccd1b8 , 
    R_1222_14b1acd8 , 
    R_1073_14b20f98 , 
    R_809_13d3e678 , 
    R_1a66_123b6158 , 
    R_1692_117f31f8 , 
    R_1447_13b93338 , 
    R_e28_156abbd8 , 
    R_a54_13cce838 , 
    R_1054_13bf8ab8 , 
    R_1466_13d5abf8 , 
    R_1673_1580e798 , 
    R_e47_1587b178 , 
    R_a35_117f5db8 , 
    R_828_10081f38 , 
    R_1469_1587ee18 , 
    R_1051_11635c38 , 
    R_e4a_11629118 , 
    R_1670_1007f238 , 
    R_82b_13cd7258 , 
    R_a32_1486afb8 , 
    R_1187_117f4198 , 
    R_1952_14a0c0d8 , 
    R_d14_13dee778 , 
    R_b68_10089d78 , 
    R_17a6_15811f38 , 
    R_1333_117f21b8 , 
    R_6f5_13d43678 , 
    R_6c8_1580d758 , 
    R_1306_1580d938 , 
    R_17d3_13d3a578 , 
    R_b95_117f7618 , 
    R_ce7_13d27218 , 
    R_1925_15ff0328 , 
    R_11b4_13b8ec98 , 
    R_576_13d2bf98 , 
    R_e00_13cd8bf8 , 
    R_7e1_150e4058 , 
    R_a7c_156b7118 , 
    R_1a3e_14a0b278 , 
    R_109b_123bd4f8 , 
    R_141f_1008c578 , 
    R_16ba_156b6e98 , 
    R_188f_156b5458 , 
    R_1270_14a103b8 , 
    R_c51_11630af8 , 
    R_632_13ccde38 , 
    R_60c_13dd9c78 , 
    R_c2b_14b23478 , 
    R_124a_140b7898 , 
    R_1869_14b29cd8 , 
    R_1a14_117ebbd8 , 
    R_13f5_13cd8a18 , 
    R_dd6_13de0d98 , 
    R_7b7_15816a38 , 
    R_aa6_13d28c58 , 
    R_10c5_11632998 , 
    R_16e4_10087078 , 
    R_190c_13d1d998 , 
    R_6af_124c33b8 , 
    R_bae_1587b5d8 , 
    R_12ed_14a176b8 , 
    R_11cd_13cd27f8 , 
    R_cce_116331b8 , 
    R_58f_156b9558 , 
    R_17ec_13dd7fb8 , 
    R_1057_123bd278 , 
    R_1463_124c4b78 , 
    R_1676_140ae6f8 , 
    R_e44_148741f8 , 
    R_a38_150dc3f8 , 
    R_825_123b3278 , 
    R_18a8_1580c8f8 , 
    R_1289_13c09738 , 
    R_c6a_15811fd8 , 
    R_64b_1007d938 , 
    R_5f3_116307d8 , 
    R_c12_1162cc78 , 
    R_1231_13dee9f8 , 
    R_1850_1587f778 , 
    R_146c_14872f38 , 
    R_104e_1580f7d8 , 
    R_e4d_14b20d18 , 
    R_166d_13d20058 , 
    R_82e_1580f2d8 , 
    R_a2f_123b3db8 , 
    R_19c3_116340b8 , 
    R_af7_13cd2d98 , 
    R_766_13c07618 , 
    R_1735_13bf9f58 , 
    R_d85_13dd7518 , 
    R_13a4_150ea138 , 
    R_1116_13c02438 , 
    R_df9_13dd9458 , 
    R_7da_14a16fd8 , 
    R_a83_13b9a278 , 
    R_10a2_123b3d18 , 
    R_1a37_1587f958 , 
    R_16c1_13d3d458 , 
    R_1418_13d2b1d8 , 
    R_ea1_156b5c78 , 
    R_9db_13c05bd8 , 
    R_1619_15888d78 , 
    R_14c0_17012fe8 , 
    R_882_13dee458 , 
    R_ffa_11c68f78 , 
    R_1967_15ff9608 , 
    R_1172_170122c8 , 
    R_d29_13bed898 , 
    R_1348_156b1178 , 
    R_b53_1162fe78 , 
    R_1791_15ff73a8 , 
    R_70a_13dee818 , 
    R_8ea_13b91c18 , 
    R_15b1_140b0d18 , 
    R_f09_13d4f9d8 , 
    R_f92_13b99238 , 
    R_1528_13cca918 , 
    R_973_12fc1738 , 
    R_907_13d1cef8 , 
    R_f26_13d51378 , 
    R_1545_13ddab78 , 
    R_1594_123b52f8 , 
    R_f75_1587ec38 , 
    R_956_117f3bf8 , 
    R_a1c_13d42098 , 
    R_147f_15ffd208 , 
    R_103b_12fbfbb8 , 
    R_e60_13b98dd8 , 
    R_165a_156b9418 , 
    R_841_13de1e78 , 
    R_1715_13c03ab8 , 
    R_10f6_1587fc78 , 
    R_ad7_11c6aaf8 , 
    R_786_13bf7938 , 
    R_da5_13c24c18 , 
    R_13c4_156adbb8 , 
    R_19e3_13b8b4f8 , 
    R_15c5_13cce478 , 
    R_8d6_14a156d8 , 
    R_fa6_13ccd7f8 , 
    R_ef5_13c0f8b8 , 
    R_987_148737f8 , 
    R_1514_13d4ea38 , 
    R_d36_13cd2938 , 
    R_1165_1700dae8 , 
    R_1355_13c0e2d8 , 
    R_b46_12fbedf8 , 
    R_717_13c1ebd8 , 
    R_1974_13b938d8 , 
    R_1784_14b1b3b8 , 
    R_156d_13b91d58 , 
    R_f4e_13d2bb38 , 
    R_156c_1486f8d8 , 
    R_92f_1587e418 , 
    R_f4d_158174d8 , 
    R_92e_15880df8 , 
    R_156e_13bee0b8 , 
    R_f4f_13d1f298 , 
    R_930_117f5818 , 
    R_156b_13cd6a38 , 
    R_f4c_13d4edf8 , 
    R_92d_13b93838 , 
    R_156f_1700c828 , 
    R_f50_13d5d038 , 
    R_931_1007f198 , 
    R_92c_13bef238 , 
    R_156a_14a0d7f8 , 
    R_f4b_1162df38 , 
    R_682_13dd6a78 , 
    R_11fa_12fbfe38 , 
    R_18df_1162e1b8 , 
    R_1819_117f44b8 , 
    R_12c0_156b3478 , 
    R_5bc_150db098 , 
    R_ca1_15888af8 , 
    R_bdb_123b9178 , 
    R_1890_13c0a4f8 , 
    R_1271_13cd3e78 , 
    R_c52_11629cf8 , 
    R_633_1587c6b8 , 
    R_60b_17014c08 , 
    R_c2a_13c01d58 , 
    R_1249_150de798 , 
    R_1868_13cd62b8 , 
    R_105a_14a112b8 , 
    R_1460_158862f8 , 
    R_1679_13cd44b8 , 
    R_e41_14a14e18 , 
    R_a3b_13cd1998 , 
    R_822_117e9158 , 
    R_1570_13d44118 , 
    R_f51_13ccb778 , 
    R_932_15810d18 , 
    R_92b_14a180b8 , 
    R_f4a_1162c8b8 , 
    R_1569_13bede38 , 
    R_163e_12fc0338 , 
    R_a00_13df4df8 , 
    R_e7c_13c08798 , 
    R_101f_117ed9d8 , 
    R_85d_117f4738 , 
    R_149b_13cd1038 , 
    R_146f_117f47d8 , 
    R_104b_158885f8 , 
    R_e50_12fbe858 , 
    R_166a_1587c938 , 
    R_831_156b2398 , 
    R_a2c_11c701d8 , 
    R_801_150e6e98 , 
    R_169a_13b94878 , 
    R_1a5e_1162d3f8 , 
    R_143f_13b8c218 , 
    R_a5c_13b8c178 , 
    R_e20_13ddd0f8 , 
    R_107b_156b2118 , 
    R_d51_13df3b38 , 
    R_1769_14b21038 , 
    R_1370_13cd2618 , 
    R_114a_13c218d8 , 
    R_198f_13d28bb8 , 
    R_732_13d55fb8 , 
    R_b2b_13ccd2f8 , 
    R_1571_1580af58 , 
    R_f52_12fc1ff8 , 
    R_933_14868718 , 
    R_92a_13c01a38 , 
    R_f49_13d4f4d8 , 
    R_1568_1580c218 , 
    R_1706_15814eb8 , 
    R_10e7_14a160d8 , 
    R_ac8_156afa58 , 
    R_795_14a12b18 , 
    R_db4_117edd98 , 
    R_13d3_13b90f98 , 
    R_19f2_12fbf258 , 
    R_17b9_156b0b38 , 
    R_193f_13d3aa78 , 
    R_b7b_13befeb8 , 
    R_d01_140ab318 , 
    R_119a_13b8a5f8 , 
    R_1320_14b27f78 , 
    R_55c_11630e18 , 
    R_6e2_158149b8 , 
    R_106b_117f3518 , 
    R_168a_117eb598 , 
    R_144f_14b26718 , 
    R_e30_123b3e58 , 
    R_a4c_170172c8 , 
    R_811_15882478 , 
    R_1406_148665f8 , 
    R_de7_1007fcd8 , 
    R_7c8_156b7f78 , 
    R_a95_117f6cb8 , 
    R_10b4_13d3d598 , 
    R_16d3_1700be28 , 
    R_1a25_13b9a318 , 
    R_1572_156b67b8 , 
    R_f53_123c01f8 , 
    R_934_156b0958 , 
    R_929_13d5bf58 , 
    R_f48_13c256b8 , 
    R_1567_13b91e98 , 
    R_1943_11c70598 , 
    R_d05_13c0cd98 , 
    R_b77_13d415f8 , 
    R_17b5_14a12118 , 
    R_1324_15887298 , 
    R_6e6_13becb78 , 
    R_558_116299d8 , 
    R_1196_13d4f398 , 
    R_e98_13d433f8 , 
    R_9e4_13cccdf8 , 
    R_1622_13c044b8 , 
    R_14b7_13d21318 , 
    R_879_15884c78 , 
    R_1003_124c39f8 , 
    R_1a16_1486b418 , 
    R_13f7_13d24338 , 
    R_dd8_1587fd18 , 
    R_7b9_13c0f458 , 
    R_aa4_13c1d0f8 , 
    R_10c3_13ccbef8 , 
    R_16e2_140b6df8 , 
    R_1573_14a0c498 , 
    R_f54_11632858 , 
    R_935_150e5318 , 
    R_928_156aab98 , 
    R_f47_13cd9238 , 
    R_1566_123b2a58 , 
    R_a0b_11637858 , 
    R_e71_14b21a38 , 
    R_102a_11c6ccb8 , 
    R_852_14b1d938 , 
    R_1490_13bf8158 , 
    R_1649_13dd4f98 , 
    R_a12_1008b358 , 
    R_e6a_156b7a78 , 
    R_1031_14b25778 , 
    R_84b_156ad1b8 , 
    R_1650_13dd4e58 , 
    R_1489_13c21978 , 
    R_7e8_1486a0b8 , 
    R_1a45_1162e2f8 , 
    R_a75_156b0778 , 
    R_1426_11637718 , 
    R_1094_13d28398 , 
    R_16b3_117efeb8 , 
    R_e07_13d453d8 , 
    R_17bd_1162b918 , 
    R_b7f_14a0be58 , 
    R_cfd_13d1d038 , 
    R_193b_13d39f38 , 
    R_119e_13c1bcf8 , 
    R_560_12fbf118 , 
    R_6de_13cd4058 , 
    R_131c_13c245d8 , 
    R_1891_123b9858 , 
    R_1272_13dd9ef8 , 
    R_c53_15ff5148 , 
    R_634_11631818 , 
    R_60a_156b2758 , 
    R_c29_13cd0598 , 
    R_1248_12fbfcf8 , 
    R_1867_14a0ded8 , 
    R_9cd_13d1f518 , 
    R_14ce_1008b5d8 , 
    R_160b_14b24cd8 , 
    R_890_11628df8 , 
    R_fec_13ccc5d8 , 
    R_eaf_13d5baf8 , 
    R_15bc_15889138 , 
    R_8df_11637358 , 
    R_f9d_158889b8 , 
    R_efe_11632b78 , 
    R_97e_13c29718 , 
    R_151d_1700bc48 , 
    R_ae2_123bdef8 , 
    R_77b_17011828 , 
    R_d9a_13c047d8 , 
    R_13b9_15ffc948 , 
    R_19d8_14870b98 , 
    R_1720_156b9198 , 
    R_1101_140b7398 , 
    R_1202_15881898 , 
    R_67a_13de2878 , 
    R_1821_117f1c18 , 
    R_18d7_1580f378 , 
    R_5c4_14868fd8 , 
    R_12b8_11631b38 , 
    R_be3_13de2198 , 
    R_c99_13c029d8 , 
    R_fd1_13c1d058 , 
    R_14e9_14868538 , 
    R_9b2_1580b6d8 , 
    R_8ab_14a0fc38 , 
    R_15f0_140ae3d8 , 
    R_eca_14a11df8 , 
    R_1574_13cd7cf8 , 
    R_f55_14b1ac38 , 
    R_936_140acf38 , 
    R_927_124c4178 , 
    R_f46_14a0af58 , 
    R_1565_1700e808 , 
    R_14d3_1580e5b8 , 
    R_9c8_15fef248 , 
    R_895_13d532b8 , 
    R_1606_1007ef18 , 
    R_eb4_117eda78 , 
    R_fe7_1162ba58 , 
    R_8f6_156b7b18 , 
    R_f15_158819d8 , 
    R_15a5_158168f8 , 
    R_1534_123b9c18 , 
    R_f86_13c1ce78 , 
    R_967_11c68938 , 
    R_1901_15817ed8 , 
    R_6a4_1162c1d8 , 
    R_bb9_156ab1d8 , 
    R_12e2_11636a98 , 
    R_11d8_156aa738 , 
    R_cc3_15887c98 , 
    R_59a_117f76b8 , 
    R_17f7_117e9838 , 
    R_105d_123b4998 , 
    R_145d_123bec18 , 
    R_167c_140b6178 , 
    R_e3e_150da7d8 , 
    R_a3e_11635cd8 , 
    R_81f_156b45f8 , 
    R_120b_13def358 , 
    R_671_140b4058 , 
    R_182a_117ef698 , 
    R_18ce_156b4e18 , 
    R_5cd_14a185b8 , 
    R_12af_15ff69a8 , 
    R_bec_124c2878 , 
    R_c90_117eb778 , 
    R_1386_14a0c7b8 , 
    R_19a5_1008a598 , 
    R_1753_13cd1218 , 
    R_748_13d3b518 , 
    R_1134_1580ad78 , 
    R_d67_13d3caf8 , 
    R_b15_156b2078 , 
    R_128a_15880718 , 
    R_c6b_14a13518 , 
    R_64c_148739d8 , 
    R_5f2_13dd5538 , 
    R_c11_15ff5aa8 , 
    R_1230_124c42b8 , 
    R_184f_1587fa98 , 
    R_18a9_11c6f918 , 
    R_bbf_1587ddd8 , 
    R_69e_123b5bb8 , 
    R_18fb_13df16f8 , 
    R_11de_10089058 , 
    R_12dc_13c0bc18 , 
    R_17fd_13d408d8 , 
    R_5a0_11631db8 , 
    R_cbd_14872df8 , 
    R_691_15883378 , 
    R_18ee_14a171b8 , 
    R_11eb_13d4f078 , 
    R_12cf_158850d8 , 
    R_180a_13d3fc58 , 
    R_5ad_14a0c2b8 , 
    R_cb0_13de1658 , 
    R_bcc_13df1f18 , 
    R_1472_13d3c698 , 
    R_1048_13df8bd8 , 
    R_e53_10087b18 , 
    R_1667_13beaf58 , 
    R_834_15888698 , 
    R_a29_13de0618 , 
    R_1575_13d42598 , 
    R_f56_13c0c578 , 
    R_937_15886c58 , 
    R_926_158846d8 , 
    R_f45_13d4f438 , 
    R_1564_1587b038 , 
    R_906_14a145f8 , 
    R_f25_13d24e78 , 
    R_1544_124c4fd8 , 
    R_1595_14b1f698 , 
    R_f76_117f6fd8 , 
    R_957_15888878 , 
    R_c7a_140ac998 , 
    R_65b_1580b778 , 
    R_5e3_117eba98 , 
    R_c02_123b2f58 , 
    R_18b8_12fc05b8 , 
    R_1221_15812cf8 , 
    R_1299_14b1fc38 , 
    R_1840_13d549d8 , 
    R_1947_156ac3f8 , 
    R_d09_150dd438 , 
    R_b73_117f7938 , 
    R_17b1_14a0dcf8 , 
    R_1328_13d2aeb8 , 
    R_6ea_123bbb58 , 
    R_1192_1587dbf8 , 
    R_137e_13c27738 , 
    R_175b_15883ff8 , 
    R_199d_1008a6d8 , 
    R_113c_13d20eb8 , 
    R_740_13bf6b78 , 
    R_b1d_123c1918 , 
    R_d5f_15888c38 , 
    R_fcb_13def8f8 , 
    R_8b1_170124a8 , 
    R_9ac_14a190f8 , 
    R_ed0_13d23d98 , 
    R_15ea_1580e658 , 
    R_14ef_123bead8 , 
    R_d33_123bd8b8 , 
    R_1168_156b6fd8 , 
    R_1352_13c10b78 , 
    R_b49_14a158b8 , 
    R_714_1587c898 , 
    R_1971_13ddfe98 , 
    R_1787_1486e2f8 , 
    R_68a_14a15b38 , 
    R_11f2_1162a6f8 , 
    R_18e7_13c08c98 , 
    R_1811_117e9a18 , 
    R_12c8_140aa878 , 
    R_5b4_140b2a78 , 
    R_ca9_15887e78 , 
    R_bd3_13c0e9b8 , 
    R_195d_15884818 , 
    R_117c_14874838 , 
    R_d1f_1007f698 , 
    R_b5d_123bb8d8 , 
    R_133e_13d55dd8 , 
    R_179b_12fbde58 , 
    R_700_13cd9878 , 
    R_1576_1700c6e8 , 
    R_f57_14a14198 , 
    R_938_13bedc58 , 
    R_925_13df1338 , 
    R_f44_156b99b8 , 
    R_1563_158841d8 , 
    R_c86_14a12e38 , 
    R_1834_13cd3f18 , 
    R_667_1486b558 , 
    R_5d7_156b0c78 , 
    R_18c4_11c709f8 , 
    R_bf6_11c6f378 , 
    R_12a5_1162d718 , 
    R_1215_117f51d8 , 
    R_1892_13d3b1f8 , 
    R_1273_13dd5c18 , 
    R_c54_13becd58 , 
    R_635_13d2c678 , 
    R_609_1580ef18 , 
    R_c28_140ba098 , 
    R_1247_13ccda78 , 
    R_1866_13bf9eb8 , 
    R_9d2_13ccb958 , 
    R_14c9_117f80b8 , 
    R_1610_1700a988 , 
    R_88b_1587e5f8 , 
    R_ff1_13b8bd18 , 
    R_eaa_13dd6618 , 
    R_1708_11630558 , 
    R_10e9_123c2138 , 
    R_aca_14a131f8 , 
    R_793_12fc2138 , 
    R_db2_123b68d8 , 
    R_13d1_156ac998 , 
    R_19f0_13d47138 , 
    R_7d3_13dd99f8 , 
    R_a8a_150e0ef8 , 
    R_10a9_1486ae78 , 
    R_16c8_13dfaed8 , 
    R_1a30_14a19698 , 
    R_1411_13dfa438 , 
    R_df2_150e09f8 , 
    R_14e3_11634838 , 
    R_9b8_13d43b78 , 
    R_8a5_13bee798 , 
    R_15f6_117f0458 , 
    R_ec4_11c68a78 , 
    R_fd7_116387f8 , 
    R_17c1_13d57d18 , 
    R_b83_13bedd98 , 
    R_cf9_1587d798 , 
    R_1937_150e3c98 , 
    R_11a2_13c05138 , 
    R_564_15815278 , 
    R_6da_13c00f98 , 
    R_1318_1008a9f8 , 
    R_faf_158866b8 , 
    R_8cd_15ff2ee8 , 
    R_eec_117f7078 , 
    R_990_11633c58 , 
    R_150b_13cd8dd8 , 
    R_15ce_13df0898 , 
    R_1766_116318b8 , 
    R_1373_15810598 , 
    R_1147_13b8d438 , 
    R_1992_13b8d1b8 , 
    R_735_13cd4cd8 , 
    R_b28_1162fab8 , 
    R_d54_150e15d8 , 
    R_1577_13d44ed8 , 
    R_f58_13d3e178 , 
    R_939_123b2878 , 
    R_924_140b7118 , 
    R_f43_140aeab8 , 
    R_1562_100874d8 , 
    R_17ce_13d50b58 , 
    R_b90_14a17e38 , 
    R_cec_156b8fb8 , 
    R_192a_13df93f8 , 
    R_11af_156b2a78 , 
    R_571_13b96ad8 , 
    R_6cd_150dc5d8 , 
    R_130b_14b1eab8 , 
    R_19b7_117f7758 , 
    R_75a_150de5b8 , 
    R_1741_100824d8 , 
    R_d79_1008a638 , 
    R_1122_150e9a58 , 
    R_1398_10083978 , 
    R_b03_158129d8 , 
    R_14d8_13cd4698 , 
    R_9c3_13befa58 , 
    R_89a_117edb18 , 
    R_1601_13d272b8 , 
    R_eb9_11638438 , 
    R_fe2_13defdf8 , 
    R_13f9_1580cb78 , 
    R_dda_117f7118 , 
    R_7bb_13bf54f8 , 
    R_aa2_12fc1a58 , 
    R_10c1_13b901d8 , 
    R_16e0_158811b8 , 
    R_1a18_156b8bf8 , 
    R_fbe_13cd90f8 , 
    R_8be_13df3278 , 
    R_99f_123b6b58 , 
    R_edd_13b99cd8 , 
    R_15dd_156aef18 , 
    R_14fc_140b09f8 , 
    R_19b2_150e0318 , 
    R_1746_123b75f8 , 
    R_755_14a13338 , 
    R_1127_13de3318 , 
    R_d74_17011d28 , 
    R_b08_150dce98 , 
    R_1393_11c68c58 , 
    R_1956_15813158 , 
    R_d18_156b9698 , 
    R_b64_156b3a18 , 
    R_17a2_117e8758 , 
    R_1337_13d20af8 , 
    R_6f9_17012b88 , 
    R_1183_1580f698 , 
    R_bb3_17013d08 , 
    R_12e8_14b1e158 , 
    R_11d2_124c3318 , 
    R_cc9_11c6e018 , 
    R_594_13cd9698 , 
    R_17f1_13c0bdf8 , 
    R_1907_13ccaa58 , 
    R_6aa_13de4038 , 
    R_ba3_13cd5bd8 , 
    R_12f8_13cd2758 , 
    R_11c2_13c1fc18 , 
    R_cd9_14b1f878 , 
    R_584_12fc0bf8 , 
    R_1917_13d21f98 , 
    R_17e1_13d37878 , 
    R_6ba_11637b78 , 
    R_8e9_13cd6b78 , 
    R_15b2_117f08b8 , 
    R_f08_156b5db8 , 
    R_f93_13b92758 , 
    R_1527_13ccaeb8 , 
    R_974_13c0c2f8 , 
    R_ad9_150e2a78 , 
    R_784_13dfa4d8 , 
    R_da3_14a0cd58 , 
    R_13c2_13d2a4b8 , 
    R_19e1_1700c5a8 , 
    R_1717_13df61f8 , 
    R_10f8_156b7258 , 
    R_1578_123bab18 , 
    R_f59_13c10358 , 
    R_93a_1486f978 , 
    R_923_11632178 , 
    R_f42_14b1f9b8 , 
    R_1561_13bf4a58 , 
    R_1060_13c0b358 , 
    R_145a_14a12bb8 , 
    R_167f_14a19378 , 
    R_e3b_13dd7f18 , 
    R_a41_14a10d18 , 
    R_81c_13bf79d8 , 
    R_12fd_1007d9d8 , 
    R_b9e_123ba618 , 
    R_cde_13d39218 , 
    R_11bd_11c6dcf8 , 
    R_191c_1580c038 , 
    R_57f_158160d8 , 
    R_6bf_13df4e98 , 
    R_17dc_15ff5508 , 
    R_1893_117f0d18 , 
    R_1274_156b1218 , 
    R_c55_13cce338 , 
    R_636_123c1238 , 
    R_608_13d58678 , 
    R_c27_13bf2a78 , 
    R_1246_14b229d8 , 
    R_1865_156b4d78 , 
    R_772_11634a18 , 
    R_d91_13c0fdb8 , 
    R_13b0_1486d0d8 , 
    R_1729_123b6338 , 
    R_19cf_11c70c78 , 
    R_110a_156b12b8 , 
    R_aeb_11638758 , 
    R_e78_117ef0f8 , 
    R_1023_15ff3ac8 , 
    R_859_13c0f098 , 
    R_1497_116337f8 , 
    R_1642_1162e578 , 
    R_a04_13c22e18 , 
    R_76b_13ddaad8 , 
    R_d8a_10085458 , 
    R_1730_11c6fd78 , 
    R_13a9_15887978 , 
    R_1111_11629c58 , 
    R_19c8_123b61f8 , 
    R_af2_11635558 , 
    R_1045_13c2abb8 , 
    R_e56_13c1f0d8 , 
    R_1664_1700d9a8 , 
    R_837_13d43c18 , 
    R_a26_13c28c78 , 
    R_1475_123b8bd8 , 
    R_e63_156b1358 , 
    R_1038_10085f98 , 
    R_1657_13cd2c58 , 
    R_844_117f3ab8 , 
    R_1482_140b29d8 , 
    R_a19_156ad4d8 , 
    R_18f5_1587d518 , 
    R_11e4_158159f8 , 
    R_12d6_11c6c5d8 , 
    R_1803_123b54d8 , 
    R_5a6_13ccf5f8 , 
    R_cb7_1162c458 , 
    R_bc5_14a0c5d8 , 
    R_698_14a0feb8 , 
    R_194b_15882658 , 
    R_d0d_1580bef8 , 
    R_b6f_117eb638 , 
    R_17ad_156b4f58 , 
    R_132c_158823d8 , 
    R_6ee_14a0faf8 , 
    R_118e_156ab3b8 , 
    R_75f_14870918 , 
    R_173c_123b9218 , 
    R_d7e_11634018 , 
    R_111d_13beeb58 , 
    R_139d_100868f8 , 
    R_afe_15ff7ee8 , 
    R_19bc_17010248 , 
    R_1175_11634c98 , 
    R_d26_1587cf78 , 
    R_b56_13c236d8 , 
    R_1345_13cd4738 , 
    R_1794_15813338 , 
    R_707_13d580d8 , 
    R_1964_13d42b38 , 
    R_f24_13b92938 , 
    R_1543_15ff0828 , 
    R_1596_15ff8a28 , 
    R_f77_158124d8 , 
    R_958_13df5bb8 , 
    R_905_13d4f758 , 
    R_1579_13b8d078 , 
    R_f5a_15884d18 , 
    R_93b_1580c3f8 , 
    R_922_140af198 , 
    R_f41_156b7cf8 , 
    R_1560_14a14cd8 , 
    R_c6c_14b20318 , 
    R_64d_13ccebf8 , 
    R_5f1_15814c38 , 
    R_c10_15817898 , 
    R_122f_13d22038 , 
    R_184e_14b1b8b8 , 
    R_18aa_11638b18 , 
    R_128b_1587eaf8 , 
    R_1695_14a12ed8 , 
    R_1a63_1486ec58 , 
    R_1444_15ff0788 , 
    R_a57_13d5aa18 , 
    R_e25_14a17078 , 
    R_1076_1587b678 , 
    R_806_14a0bd18 , 
    R_fb7_15887158 , 
    R_8c5_1008b2b8 , 
    R_998_13d573b8 , 
    R_ee4_15ff7da8 , 
    R_1503_150daf58 , 
    R_15d6_117ed398 , 
    R_7ca_150de978 , 
    R_a93_156af4b8 , 
    R_10b2_100826b8 , 
    R_16d1_156b27f8 , 
    R_1a27_13cd2118 , 
    R_1408_1587fbd8 , 
    R_de9_13cd12b8 , 
    R_9e0_15ffc9e8 , 
    R_161e_123b8a98 , 
    R_14bb_10081cb8 , 
    R_87d_123b9498 , 
    R_fff_12fbe5d8 , 
    R_e9c_13df34f8 , 
    R_ba8_123c12d8 , 
    R_12f3_11634f18 , 
    R_11c7_17013b28 , 
    R_cd4_13c2b018 , 
    R_589_14a19058 , 
    R_1912_156aacd8 , 
    R_17e6_140b2758 , 
    R_6b5_1587d658 , 
    R_f14_13d26458 , 
    R_15a6_1162eb18 , 
    R_1533_14b268f8 , 
    R_f87_11637998 , 
    R_968_13d2b958 , 
    R_8f5_13bebe58 , 
    R_8d5_150e1c18 , 
    R_fa7_12fbff78 , 
    R_ef4_1162ea78 , 
    R_988_15814198 , 
    R_1513_13c06498 , 
    R_15c6_12fbf2f8 , 
    R_8b7_15ffa468 , 
    R_9a6_13d46058 , 
    R_ed6_13d57598 , 
    R_15e4_156aeb58 , 
    R_14f5_13c29178 , 
    R_fc5_13b8d258 , 
    R_acc_13df8638 , 
    R_791_13d42818 , 
    R_db0_13bf9418 , 
    R_13cf_123c2318 , 
    R_19ee_11630cd8 , 
    R_170a_13d25698 , 
    R_10eb_13debbb8 , 
    R_19ad_1587f9f8 , 
    R_174b_15ff3528 , 
    R_750_1008c9d8 , 
    R_112c_13c015d8 , 
    R_d6f_117eae18 , 
    R_b0d_13d41c38 , 
    R_138e_158113f8 , 
    R_168d_156b2f78 , 
    R_144c_14a0dbb8 , 
    R_e2d_1587d3d8 , 
    R_a4f_15814418 , 
    R_80e_156ac218 , 
    R_106e_14a15318 , 
    R_157a_156b4198 , 
    R_f5b_1162d7b8 , 
    R_93c_13b933d8 , 
    R_921_15813298 , 
    R_f40_13cd1fd8 , 
    R_155f_148745b8 , 
    R_1275_13d26bd8 , 
    R_c56_12fbf438 , 
    R_637_14b20db8 , 
    R_607_15886258 , 
    R_c26_13d3ac58 , 
    R_1245_13d261d8 , 
    R_1864_13ddb2f8 , 
    R_1894_13cd6998 , 
    R_9d7_1580ac38 , 
    R_1615_150e0598 , 
    R_14c4_15ffa148 , 
    R_886_156aa9b8 , 
    R_ff6_13d424f8 , 
    R_ea5_13d23b18 , 
    R_1a51_13cda098 , 
    R_a69_123b4f38 , 
    R_1432_14b1d258 , 
    R_1088_13bec3f8 , 
    R_e13_140ab1d8 , 
    R_16a7_156afb98 , 
    R_7f4_14b238d8 , 
    R_17c5_12fc1058 , 
    R_b87_140b0db8 , 
    R_cf5_156ab818 , 
    R_1933_11633258 , 
    R_11a6_13c243f8 , 
    R_568_13ccd9d8 , 
    R_6d6_13ccc498 , 
    R_1314_13b93158 , 
    R_a81_11c6b098 , 
    R_10a0_148694d8 , 
    R_1a39_150e4cd8 , 
    R_16bf_13d3e8f8 , 
    R_141a_13ccc678 , 
    R_dfb_123b4c18 , 
    R_7dc_14b22578 , 
    R_116b_13ddcb58 , 
    R_134f_14b1c7b8 , 
    R_b4c_13d41eb8 , 
    R_711_140b8798 , 
    R_178a_13b96538 , 
    R_196e_150e3658 , 
    R_d30_13df5118 , 
    R_b99_13df2ff8 , 
    R_ce3_10088b58 , 
    R_11b8_156b8798 , 
    R_1921_13b91df8 , 
    R_57a_13ccb818 , 
    R_6c4_15887798 , 
    R_17d7_11c6faf8 , 
    R_1302_12fbe8f8 , 
    R_65c_117f0278 , 
    R_5e2_117ef198 , 
    R_c01_13df0118 , 
    R_18b9_13ded058 , 
    R_1220_117f77f8 , 
    R_129a_14a10ef8 , 
    R_183f_140b7f78 , 
    R_c7b_1580c178 , 
    R_7bd_12fc1558 , 
    R_aa0_11c6be58 , 
    R_10bf_13df54d8 , 
    R_16de_13de3138 , 
    R_1a1a_156b8ab8 , 
    R_13fb_156b4b98 , 
    R_ddc_11632df8 , 
    R_a7a_11c6b1d8 , 
    R_1a40_140b6d58 , 
    R_1099_116354b8 , 
    R_1421_117ef7d8 , 
    R_16b8_13d3ea38 , 
    R_e02_15ff37a8 , 
    R_7e3_15812118 , 
    R_1a56_13bf0818 , 
    R_1437_123bad98 , 
    R_a64_13beb318 , 
    R_e18_156afc38 , 
    R_1083_123c0a18 , 
    R_7f9_156b30b8 , 
    R_16a2_150e9418 , 
    R_18e0_13c201b8 , 
    R_1818_140b47d8 , 
    R_12c1_123bb838 , 
    R_5bb_156b5638 , 
    R_ca2_13dd9d18 , 
    R_bda_13b985b8 , 
    R_683_11634478 , 
    R_11f9_13ccd938 , 
    R_157b_1486f0b8 , 
    R_f5c_13de2378 , 
    R_93d_117f0ef8 , 
    R_920_13df90d8 , 
    R_f3f_13bf1a38 , 
    R_155e_123c0d38 , 
    R_8de_13d4e0d8 , 
    R_f9e_13b8a738 , 
    R_efd_123bfed8 , 
    R_97f_123c21d8 , 
    R_151c_13d5c4f8 , 
    R_15bd_13df43f8 , 
    R_1763_13d44618 , 
    R_1995_17017548 , 
    R_1144_17018948 , 
    R_738_1700bce8 , 
    R_b25_1162ad38 , 
    R_d57_13c242b8 , 
    R_1376_117f5098 , 
    R_9be_140aaaf8 , 
    R_89f_156b2ed8 , 
    R_15fc_13c28db8 , 
    R_ebe_13cd5c78 , 
    R_fdd_1162dd58 , 
    R_14dd_123b8db8 , 
    R_14aa_13c0f9f8 , 
    R_86c_13df77d8 , 
    R_1010_15884278 , 
    R_e8b_15880ad8 , 
    R_162f_15ff7808 , 
    R_9f1_123be718 , 
    R_1457_13d54758 , 
    R_1682_1587fb38 , 
    R_e38_150debf8 , 
    R_a44_1580d618 , 
    R_819_14873898 , 
    R_1063_13cd8978 , 
    R_1a4c_156b8b58 , 
    R_a6e_117ec3f8 , 
    R_142d_14b1c998 , 
    R_108d_14a0a878 , 
    R_e0e_156b9f58 , 
    R_16ac_13bf1218 , 
    R_7ef_1700c788 , 
    R_1014_13c079d8 , 
    R_868_1587de78 , 
    R_14a6_10081998 , 
    R_1633_117e9ab8 , 
    R_9f5_13d25c38 , 
    R_e87_15ff9ce8 , 
    R_1829_123b40d8 , 
    R_18cf_13ded238 , 
    R_5cc_156aa698 , 
    R_12b0_14a177f8 , 
    R_beb_13cca738 , 
    R_c91_15ff1cc8 , 
    R_120a_13cd9738 , 
    R_672_13c06fd8 , 
    R_779_13cd2258 , 
    R_d98_13b958b8 , 
    R_13b7_1700e308 , 
    R_19d6_117ecfd8 , 
    R_1722_123b5a78 , 
    R_1103_117f7bb8 , 
    R_ae4_11634ab8 , 
    R_c57_15814f58 , 
    R_638_14a151d8 , 
    R_606_13d50838 , 
    R_c25_10083bf8 , 
    R_1244_13ddb898 , 
    R_1863_123b9f38 , 
    R_1895_13df3a98 , 
    R_1276_123bda98 , 
    R_1042_13cd6718 , 
    R_e59_1587dd38 , 
    R_1661_13de0758 , 
    R_83a_13d21598 , 
    R_a23_14869cf8 , 
    R_1478_13cd7618 , 
    R_668_11c6aff8 , 
    R_5d6_13d24158 , 
    R_18c5_123b5f78 , 
    R_bf5_123ba7f8 , 
    R_12a6_148674f8 , 
    R_1214_15886cf8 , 
    R_c87_13c21bf8 , 
    R_1833_117f3838 , 
    R_1820_14872a38 , 
    R_18d8_13b8ef18 , 
    R_5c3_10080778 , 
    R_12b9_140abb38 , 
    R_be2_13b98338 , 
    R_c9a_13cd1f38 , 
    R_1201_15ff65e8 , 
    R_67b_13c02bb8 , 
    R_1542_14a19cd8 , 
    R_1597_117ee478 , 
    R_f78_156af198 , 
    R_959_11631bd8 , 
    R_904_13bebbd8 , 
    R_f23_13c2b338 , 
    R_157c_14a0eab8 , 
    R_f5d_15817c58 , 
    R_93e_13cd6858 , 
    R_91f_117f7d98 , 
    R_f3e_1700a708 , 
    R_155d_1700fa28 , 
    R_764_150dee78 , 
    R_1737_13cd6538 , 
    R_d83_150dc678 , 
    R_1118_13cce3d8 , 
    R_13a2_13df95d8 , 
    R_af9_14b1bc78 , 
    R_19c1_15811358 , 
    R_14ae_14b22438 , 
    R_870_158800d8 , 
    R_100c_14b1bef8 , 
    R_e8f_13c27cd8 , 
    R_9ed_150e3a18 , 
    R_162b_13d24478 , 
    R_64e_12fbeb78 , 
    R_5f0_13d25738 , 
    R_c0f_1587ef58 , 
    R_122e_14a181f8 , 
    R_184d_1486ac98 , 
    R_18ab_13bf9d78 , 
    R_128c_11c6a378 , 
    R_c6d_13d3be78 , 
    R_d11_117f09f8 , 
    R_b6b_13c0e878 , 
    R_17a9_15ff62c8 , 
    R_1330_1580d6b8 , 
    R_6f2_123ba398 , 
    R_118a_13c1eef8 , 
    R_194f_13c0e738 , 
    R_1758_14a14eb8 , 
    R_19a0_13c204d8 , 
    R_1139_117ef878 , 
    R_743_13d5a478 , 
    R_b1a_13c01038 , 
    R_d62_15811df8 , 
    R_1381_123b3a98 , 
    R_e6d_123b7238 , 
    R_102e_150ddd98 , 
    R_84e_15883418 , 
    R_164d_14a0c678 , 
    R_148c_1580e8d8 , 
    R_a0f_15ffbae8 , 
    R_12ee_13d3d958 , 
    R_11cc_14a11a38 , 
    R_ccf_15812258 , 
    R_58e_150e4558 , 
    R_17eb_150e6538 , 
    R_190d_14b294b8 , 
    R_6b0_14a172f8 , 
    R_bad_15883c38 , 
    R_1018_13d2a878 , 
    R_864_13c09238 , 
    R_14a2_13cd9e18 , 
    R_1637_1162fbf8 , 
    R_9f9_156b7438 , 
    R_e83_15886438 , 
    R_1a5b_13df6158 , 
    R_143c_15ff2a88 , 
    R_a5f_13df1518 , 
    R_e1d_13c288b8 , 
    R_107e_13c1c298 , 
    R_7fe_117f30b8 , 
    R_169d_156abf98 , 
    R_15b3_13cd6e98 , 
    R_f07_13b953b8 , 
    R_f94_13d25198 , 
    R_1526_1486bf58 , 
    R_975_13d529f8 , 
    R_8e8_117f0bd8 , 
    R_78f_1162c9f8 , 
    R_dae_11c6d578 , 
    R_13cd_14a162b8 , 
    R_19ec_15814738 , 
    R_170c_13ccdd98 , 
    R_10ed_15882dd8 , 
    R_ace_15885cb8 , 
    R_157d_13cd56d8 , 
    R_f5e_140b53b8 , 
    R_93f_13d57778 , 
    R_91e_15886f78 , 
    R_f3d_11634798 , 
    R_155c_156adf78 , 
    R_782_15ffd168 , 
    R_da1_14b290f8 , 
    R_13c0_117f6b78 , 
    R_19df_117eb318 , 
    R_1719_13c1f8f8 , 
    R_10fa_13decd38 , 
    R_adb_17014708 , 
    R_a88_13cd40f8 , 
    R_10a7_117eb1d8 , 
    R_16c6_158880f8 , 
    R_1a32_15818018 , 
    R_1413_13d57ef8 , 
    R_df4_17013f88 , 
    R_7d5_15889098 , 
    R_639_13df0cf8 , 
    R_605_14b1c3f8 , 
    R_c24_11632d58 , 
    R_1243_158151d8 , 
    R_1862_140b94b8 , 
    R_1896_13c0a598 , 
    R_1277_13c27378 , 
    R_c58_13dddc38 , 
    R_15a7_17013448 , 
    R_1532_156b4ff8 , 
    R_f88_13d225d8 , 
    R_969_13cce298 , 
    R_8f4_156b9af8 , 
    R_f13_13c2b478 , 
    R_1750_14a13018 , 
    R_74b_123b9998 , 
    R_1131_13d21c78 , 
    R_d6a_13c0c118 , 
    R_b12_1587bb78 , 
    R_1389_13c2a4d8 , 
    R_19a8_124c5578 , 
    R_a9e_13de43f8 , 
    R_10bd_1162e6b8 , 
    R_16dc_14b1f058 , 
    R_1a1c_13cda138 , 
    R_13fd_14a0e0b8 , 
    R_dde_15ffc448 , 
    R_7bf_123bb0b8 , 
    R_1027_13c277d8 , 
    R_855_14a117b8 , 
    R_1493_13bee3d8 , 
    R_1646_13ccbdb8 , 
    R_a08_15ffa5a8 , 
    R_e74_123b4678 , 
    R_12d0_14a11cb8 , 
    R_1809_13d4f7f8 , 
    R_5ac_11c6e838 , 
    R_cb1_13d2c998 , 
    R_bcb_1007e3d8 , 
    R_692_1587be98 , 
    R_18ef_13d28758 , 
    R_11ea_1580f238 , 
    R_991_1007ff58 , 
    R_eeb_12fbe0d8 , 
    R_150a_14a0b3b8 , 
    R_15cf_10085958 , 
    R_fb0_117f5318 , 
    R_8cc_13bf3338 , 
    R_ce8_11c6a7d8 , 
    R_1926_116372b8 , 
    R_11b3_13cd3fb8 , 
    R_575_15817438 , 
    R_6c9_13dee318 , 
    R_1307_15ff2da8 , 
    R_17d2_156b8978 , 
    R_b94_1587e198 , 
    R_1810_117f12b8 , 
    R_12c9_17017868 , 
    R_5b3_123baa78 , 
    R_caa_15fedbc8 , 
    R_bd2_1580d9d8 , 
    R_68b_13ddf038 , 
    R_11f1_13c2a938 , 
    R_18e8_123bd638 , 
    R_157e_13dee278 , 
    R_f5f_1162d038 , 
    R_940_1486f838 , 
    R_91d_14b1cdf8 , 
    R_f3c_148682b8 , 
    R_155b_12fc0158 , 
    R_14b2_15ff2628 , 
    R_874_123c0298 , 
    R_1008_1587dc98 , 
    R_e93_13cd4878 , 
    R_9e9_123b4498 , 
    R_1627_156b7578 , 
    R_cf1_124c34f8 , 
    R_192f_14a12cf8 , 
    R_11aa_117e9bf8 , 
    R_56c_140ab598 , 
    R_6d2_1162ec58 , 
    R_1310_13ddf538 , 
    R_17c9_11638578 , 
    R_b8b_13df36d8 , 
    R_a91_13ccfeb8 , 
    R_10b0_117ea418 , 
    R_16cf_11c6b138 , 
    R_1a29_13d384f8 , 
    R_140a_140aa5f8 , 
    R_deb_140b71b8 , 
    R_7cc_13cd94b8 , 
    R_1a47_100862b8 , 
    R_a73_123be538 , 
    R_1428_13dde3b8 , 
    R_1092_15ff41a8 , 
    R_e09_15887a18 , 
    R_16b1_13c0c258 , 
    R_7ea_11c6e518 , 
    R_e66_170138a8 , 
    R_1035_1162a478 , 
    R_847_14a15a98 , 
    R_1654_1580fff8 , 
    R_1485_117f6358 , 
    R_a16_14b25638 , 
    R_b60_13b97b18 , 
    R_179e_156b3c98 , 
    R_133b_13ddde18 , 
    R_6fd_156b8338 , 
    R_117f_13cd7578 , 
    R_195a_150e1218 , 
    R_d1c_13d3fd98 , 
    R_134c_14a11ad8 , 
    R_b4f_12fbee98 , 
    R_70e_124c25f8 , 
    R_178d_11638a78 , 
    R_196b_1580a918 , 
    R_d2d_13cd54f8 , 
    R_116e_117ebb38 , 
    R_5e1_14b286f8 , 
    R_c00_150df558 , 
    R_18ba_11638bb8 , 
    R_121f_13dfa1b8 , 
    R_129b_13cd3298 , 
    R_183e_1587c398 , 
    R_c7c_11c6a558 , 
    R_65d_13cd74d8 , 
    R_9b3_13df8138 , 
    R_8aa_13dd9a98 , 
    R_15f1_156b5d18 , 
    R_ec9_1587c1b8 , 
    R_fd2_13c05098 , 
    R_14e8_1700a528 , 
    R_11dd_14875918 , 
    R_12dd_14a0e158 , 
    R_17fc_11635eb8 , 
    R_59f_14a14c38 , 
    R_cbe_116357d8 , 
    R_bbe_15881438 , 
    R_18fc_17009bc8 , 
    R_69f_13d56b98 , 
    R_1598_13cd92d8 , 
    R_f79_13bf2e38 , 
    R_95a_13d37698 , 
    R_903_117ec7b8 , 
    R_f22_14a13978 , 
    R_1541_15886758 , 
    R_12e3_17014028 , 
    R_11d7_1587d5b8 , 
    R_cc4_13bead78 , 
    R_599_150dcf38 , 
    R_17f6_117f1498 , 
    R_1902_14b1af58 , 
    R_6a5_13df56b8 , 
    R_bb8_124c3b38 , 
    R_14bf_150dd938 , 
    R_881_150db278 , 
    R_ffb_15813ab8 , 
    R_ea0_13b95778 , 
    R_9dc_15ff19a8 , 
    R_161a_14b23bf8 , 
    R_1454_123b4538 , 
    R_e35_11c70098 , 
    R_a47_1486f3d8 , 
    R_816_13c06cb8 , 
    R_1066_13bee838 , 
    R_1685_15ff1d68 , 
    R_8b0_15813c98 , 
    R_9ad_13de0bb8 , 
    R_ecf_13c26798 , 
    R_15eb_140b6498 , 
    R_14ee_13d5a298 , 
    R_fcc_150e33d8 , 
    R_101c_11c6ce98 , 
    R_860_14a17b18 , 
    R_149e_11c6edd8 , 
    R_163b_13c04b98 , 
    R_9fd_117ebf98 , 
    R_e7f_117f6038 , 
    R_604_15811718 , 
    R_c23_123bfc58 , 
    R_1242_10080c78 , 
    R_1861_12fbf7f8 , 
    R_1897_13d3d1d8 , 
    R_1278_117f4f58 , 
    R_c59_116304b8 , 
    R_63a_13c0a278 , 
    R_b59_15feff68 , 
    R_1342_148716d8 , 
    R_1797_117f7e38 , 
    R_704_123b2ff8 , 
    R_1961_1162de98 , 
    R_1178_13cd24d8 , 
    R_d23_11c68618 , 
    R_157f_13b8ce98 , 
    R_f60_140af9b8 , 
    R_941_13df8b38 , 
    R_91c_13df6d38 , 
    R_f3b_15810c78 , 
    R_155a_15882338 , 
    R_e5c_117f6df8 , 
    R_165e_117edf78 , 
    R_83d_13c24ad8 , 
    R_a20_15883738 , 
    R_147b_1700f5c8 , 
    R_103f_123b9ad8 , 
    R_5ef_1162a018 , 
    R_c0e_158802b8 , 
    R_122d_150e4eb8 , 
    R_184c_14a19418 , 
    R_18ac_117f13f8 , 
    R_128d_123b2af8 , 
    R_c6e_15ff6408 , 
    R_64f_13bf1ad8 , 
    R_9a0_13dd6078 , 
    R_edc_123be678 , 
    R_15de_15ff2268 , 
    R_14fb_13c29038 , 
    R_fbf_150e4f58 , 
    R_8bd_13cd5ef8 , 
    R_1998_14b279d8 , 
    R_1141_1580bbd8 , 
    R_73b_14a15638 , 
    R_b22_13cce8d8 , 
    R_d5a_13bf6178 , 
    R_1379_123bdbd8 , 
    R_1760_117f7f78 , 
    R_1981_1587b7b8 , 
    R_b39_15ffae68 , 
    R_724_117ec8f8 , 
    R_1777_1587ccf8 , 
    R_d43_13beedd8 , 
    R_1362_150dfcd8 , 
    R_1158_13bf0f98 , 
    R_770_15888058 , 
    R_d8f_11629f78 , 
    R_13ae_13bf3478 , 
    R_172b_156b88d8 , 
    R_19cd_117ed578 , 
    R_110c_15810458 , 
    R_aed_14a0e298 , 
    R_1449_14b26678 , 
    R_e2a_13c29858 , 
    R_a52_140af378 , 
    R_80b_158154f8 , 
    R_1071_123c1378 , 
    R_1a68_117ed618 , 
    R_1690_13c216f8 , 
    R_ef3_13cd06d8 , 
    R_989_13c068f8 , 
    R_1512_1162e078 , 
    R_15c7_13d3c4b8 , 
    R_8d4_123c1738 , 
    R_fa8_123be858 , 
    R_1984_1162e438 , 
    R_727_1700aca8 , 
    R_b36_123bb338 , 
    R_d46_13cd3338 , 
    R_1774_13c26c98 , 
    R_1365_150db818 , 
    R_1155_17012868 , 
    R_b3c_13cd4eb8 , 
    R_721_156b7d98 , 
    R_197e_13d5c8b8 , 
    R_177a_123c1418 , 
    R_d40_11635af8 , 
    R_115b_123bf2f8 , 
    R_135f_11c6da78 , 
    R_894_1587b2b8 , 
    R_1607_123bd138 , 
    R_eb3_123b5cf8 , 
    R_fe8_15816678 , 
    R_14d2_11636e58 , 
    R_9c9_13cce798 , 
    R_160c_117f74d8 , 
    R_88f_13c0d338 , 
    R_fed_12fc1198 , 
    R_eae_13cd1d58 , 
    R_9ce_1162c6d8 , 
    R_14cd_10081178 , 
    R_dac_14a109f8 , 
    R_13cb_13ccf0f8 , 
    R_19ea_11629b18 , 
    R_170e_1580e338 , 
    R_10ef_14a199b8 , 
    R_ad0_123b65b8 , 
    R_78d_15817618 , 
    R_999_1008a138 , 
    R_ee3_158135b8 , 
    R_1502_117ea238 , 
    R_15d7_11c6ab98 , 
    R_fb8_156b7bb8 , 
    R_8c4_117f8018 , 
    R_efc_12fc14b8 , 
    R_980_13d2b9f8 , 
    R_151b_14a153b8 , 
    R_15be_11629bb8 , 
    R_8dd_13d1dcb8 , 
    R_f9f_13bf1858 , 
    R_8a4_13cd4418 , 
    R_15f7_117ea878 , 
    R_ec3_14a15e58 , 
    R_fd8_117f1718 , 
    R_14e2_13ddc478 , 
    R_9b9_1008a458 , 
    R_1580_123b3958 , 
    R_f61_14867318 , 
    R_942_140b3a18 , 
    R_91b_156b0d18 , 
    R_f3a_1007f4b8 , 
    R_1559_13c234f8 , 
    R_1441_13ded378 , 
    R_a5a_13c097d8 , 
    R_e22_117eccb8 , 
    R_1079_13beb6d8 , 
    R_803_140b8158 , 
    R_1698_15811998 , 
    R_1a60_14b1b778 , 
    R_1987_140b7cf8 , 
    R_72a_158127f8 , 
    R_b33_13d2aaf8 , 
    R_d49_15811678 , 
    R_1771_17009c68 , 
    R_1368_1587e9b8 , 
    R_1152_13c0bd58 , 
    R_5d5_123be038 , 
    R_18c6_13d3a1b8 , 
    R_bf4_1587cb18 , 
    R_12a7_15817cf8 , 
    R_1213_140ad078 , 
    R_c88_17017cc8 , 
    R_1832_123bc2d8 , 
    R_669_116322b8 , 
    R_769_150da558 , 
    R_d88_117f22f8 , 
    R_1732_123b2558 , 
    R_13a7_13c08ab8 , 
    R_1113_123c1e18 , 
    R_19c6_13cd18f8 , 
    R_af4_1580feb8 , 
    R_b3f_13c22198 , 
    R_71e_140aec98 , 
    R_197b_123c14b8 , 
    R_177d_17012728 , 
    R_d3d_13c053b8 , 
    R_115e_15885c18 , 
    R_135c_13cda3b8 , 
    R_12d7_13cd2578 , 
    R_1802_13d3fbb8 , 
    R_5a5_13d375f8 , 
    R_cb8_11c6c218 , 
    R_bc4_14b2a138 , 
    R_699_15888ff8 , 
    R_18f6_124c27d8 , 
    R_11e3_1162fa18 , 
    R_b67_13cd4f58 , 
    R_17a5_116334d8 , 
    R_1334_13cd5598 , 
    R_6f6_117f1858 , 
    R_1186_11635d78 , 
    R_1953_117eb6d8 , 
    R_d15_123b5578 , 
    R_603_13ddbe38 , 
    R_c22_117f71b8 , 
    R_1241_1162a5b8 , 
    R_1860_13ccdf78 , 
    R_1898_11c6bb38 , 
    R_1279_15887478 , 
    R_c5a_14a16538 , 
    R_63b_15883cd8 , 
    R_10bb_1587d8d8 , 
    R_16da_124c3db8 , 
    R_1a1e_11c6ed38 , 
    R_13ff_17012c28 , 
    R_de0_13d3abb8 , 
    R_7c1_156b3bf8 , 
    R_a9c_1162e4d8 , 
    R_18d0_117f1358 , 
    R_5cb_12fc0d38 , 
    R_12b1_124c38b8 , 
    R_bea_13ccb098 , 
    R_c92_150e3838 , 
    R_1209_14a0aa58 , 
    R_673_14a13fb8 , 
    R_1828_1580ab98 , 
    R_14b6_1587d1f8 , 
    R_878_13c100d8 , 
    R_1004_156ab318 , 
    R_e97_14866918 , 
    R_9e5_1587d6f8 , 
    R_1623_13b96178 , 
    R_11d1_1162f6f8 , 
    R_cca_117eebf8 , 
    R_593_117ee0b8 , 
    R_17f0_100833d8 , 
    R_1908_1162f5b8 , 
    R_6ab_13ccbe58 , 
    R_bb2_15810278 , 
    R_12e9_13d26818 , 
    R_f89_13d51738 , 
    R_96a_1587c258 , 
    R_8f3_10082b18 , 
    R_f12_1162b2d8 , 
    R_15a8_14b25db8 , 
    R_1531_13c0ac78 , 
    R_12c2_13d4e2b8 , 
    R_5ba_13b94d78 , 
    R_ca3_13ddaa38 , 
    R_bd9_13d54398 , 
    R_684_117f5a98 , 
    R_11f8_13bf1538 , 
    R_18e1_17010388 , 
    R_1817_1580f9b8 , 
    R_a7f_117ebc78 , 
    R_1a3b_13d275d8 , 
    R_109e_14a11538 , 
    R_16bd_117eb9f8 , 
    R_141c_123b3f98 , 
    R_dfd_1700cf08 , 
    R_7de_15881ed8 , 
    R_f95_13d51058 , 
    R_1525_140b5598 , 
    R_976_140b2f78 , 
    R_8e7_13dd8ff8 , 
    R_15b4_13dee598 , 
    R_f06_14b29238 , 
    R_899_13d5a8d8 , 
    R_1602_13c28ef8 , 
    R_eb8_13c1c0b8 , 
    R_fe3_13ccb598 , 
    R_14d7_14a0fb98 , 
    R_9c4_123c1a58 , 
    R_1599_13bf40f8 , 
    R_f7a_13d510f8 , 
    R_95b_15813838 , 
    R_902_14a0aff8 , 
    R_f21_15812398 , 
    R_1540_14871458 , 
    R_1321_156b1038 , 
    R_1199_13cd3bf8 , 
    R_6e3_140b27f8 , 
    R_55b_13d54f78 , 
    R_1940_117ed758 , 
    R_17b8_14b1ca38 , 
    R_d02_14b21998 , 
    R_b7a_140b8298 , 
    R_ed5_123b27d8 , 
    R_15e5_13d3e0d8 , 
    R_14f4_1580cad8 , 
    R_fc6_117f2078 , 
    R_8b6_12fbe7b8 , 
    R_9a7_13dd6118 , 
    R_d96_13c23778 , 
    R_13b5_124c31d8 , 
    R_19d4_123b6798 , 
    R_1724_117edcf8 , 
    R_1105_158130b8 , 
    R_ae6_14873e38 , 
    R_777_17012228 , 
    R_1581_10080458 , 
    R_f62_13ccaff8 , 
    R_943_156b21b8 , 
    R_91a_13d23e38 , 
    R_f39_117f5778 , 
    R_1558_15ffb2c8 , 
    R_88a_15880c18 , 
    R_ff2_13d42638 , 
    R_ea9_15810ef8 , 
    R_9d3_12fc1e18 , 
    R_14c8_13d50d38 , 
    R_1611_13df2b98 , 
    R_5c2_150db138 , 
    R_12ba_158138d8 , 
    R_be1_10082898 , 
    R_c9b_13b977f8 , 
    R_1200_13d3d778 , 
    R_67c_13dec978 , 
    R_181f_156b4558 , 
    R_18d9_117f3e78 , 
    R_1743_15ff3488 , 
    R_758_13cd0ef8 , 
    R_1124_14a17d98 , 
    R_d77_14a0ca38 , 
    R_1396_156ace98 , 
    R_b05_13d37d78 , 
    R_19b5_13cd3c98 , 
    R_d9f_1580b818 , 
    R_13be_156af5f8 , 
    R_19dd_13d56238 , 
    R_171b_14a0ac38 , 
    R_10fc_13d52c78 , 
    R_add_17015ce8 , 
    R_780_13cd31f8 , 
    R_198a_12fc1af8 , 
    R_72d_13d467d8 , 
    R_b30_156ac358 , 
    R_d4c_11633d98 , 
    R_176e_12fbe678 , 
    R_136b_15810638 , 
    R_114f_123ba1b8 , 
    R_119d_123ba578 , 
    R_55f_13cce658 , 
    R_6df_13bf5ef8 , 
    R_131d_14a11c18 , 
    R_17bc_15886d98 , 
    R_b7e_123b7eb8 , 
    R_cfe_123b7418 , 
    R_193c_123b6298 , 
    R_b42_116296b8 , 
    R_71b_13cd8fb8 , 
    R_1978_1587e698 , 
    R_1780_1587b718 , 
    R_d3a_117f6678 , 
    R_1161_13beb3b8 , 
    R_1359_11c6d9d8 , 
    R_1325_156ac178 , 
    R_6e7_15882fb8 , 
    R_557_15885f38 , 
    R_1195_116363b8 , 
    R_1944_124c2918 , 
    R_d06_13dde818 , 
    R_b76_13d41b98 , 
    R_17b4_13d29ab8 , 
    R_1020_117ed258 , 
    R_85c_1580fc38 , 
    R_149a_13bf0ef8 , 
    R_163f_13de4218 , 
    R_a01_156b1498 , 
    R_e7b_1486b738 , 
    R_11c1_123b5618 , 
    R_cda_156b9878 , 
    R_1918_15880f38 , 
    R_583_13cccb78 , 
    R_17e0_14a15d18 , 
    R_6bb_117f2398 , 
    R_ba2_14a0e5b8 , 
    R_12f9_13d5c9f8 , 
    R_5ee_12fc0c98 , 
    R_c0d_13b93fb8 , 
    R_122c_14b217b8 , 
    R_18ad_13cd6358 , 
    R_184b_1486d3f8 , 
    R_128e_13b91a38 , 
    R_c6f_150e83d8 , 
    R_650_116346f8 , 
    R_5e0_13df04d8 , 
    R_bff_123b92b8 , 
    R_18bb_11c6f698 , 
    R_121e_14b1d438 , 
    R_129c_1007ebf8 , 
    R_183d_15882e78 , 
    R_c7d_13c108f8 , 
    R_65e_13d43998 , 
    R_75d_156ad118 , 
    R_173e_148678b8 , 
    R_d7c_123be998 , 
    R_111f_14a110d8 , 
    R_139b_156b35b8 , 
    R_b00_13ccf558 , 
    R_19ba_17014d48 , 
    R_a78_13cd1cb8 , 
    R_1a42_15817118 , 
    R_1097_13d240b8 , 
    R_1423_13c05a98 , 
    R_16b6_140aab98 , 
    R_e04_156b17b8 , 
    R_7e5_14b1e798 , 
    R_746_170166e8 , 
    R_1136_13d56558 , 
    R_d65_1008bb78 , 
    R_b17_123bcc38 , 
    R_1384_140b3298 , 
    R_19a3_117eaa58 , 
    R_1755_10087258 , 
    R_c21_1700d4a8 , 
    R_1240_11630238 , 
    R_185f_13bf7118 , 
    R_1899_156b1fd8 , 
    R_127a_14b28298 , 
    R_c5b_13d26278 , 
    R_63c_1587b538 , 
    R_602_156afff8 , 
    R_753_116336b8 , 
    R_1129_13ccc3f8 , 
    R_d72_13b95e58 , 
    R_b0a_156ad438 , 
    R_1391_15886578 , 
    R_19b0_17014a28 , 
    R_1748_117eeab8 , 
    R_e32_13c05c78 , 
    R_a4a_117e8bb8 , 
    R_813_11631318 , 
    R_1069_116369f8 , 
    R_1688_156b6a38 , 
    R_1451_150e6b78 , 
    R_cdf_150dfa58 , 
    R_11bc_11c6a9b8 , 
    R_191d_13c10678 , 
    R_57e_1162f338 , 
    R_6c0_13b98c98 , 
    R_17db_117f6858 , 
    R_12fe_116291b8 , 
    R_b9d_14872678 , 
    R_1349_13d26db8 , 
    R_b52_1162a978 , 
    R_1790_117e9798 , 
    R_70b_17018808 , 
    R_1968_13bf0318 , 
    R_d2a_15fef568 , 
    R_1171_117f5278 , 
    R_192b_11633cf8 , 
    R_11ae_123bc238 , 
    R_570_117ec218 , 
    R_6ce_13dee1d8 , 
    R_130c_15ff67c8 , 
    R_17cd_13b91858 , 
    R_b8f_14b25b38 , 
    R_ced_14a0a558 , 
    R_1582_150e7ed8 , 
    R_f63_13cca7d8 , 
    R_944_13d1fab8 , 
    R_919_123bdf98 , 
    R_f38_13d26958 , 
    R_1557_14a16c18 , 
    R_10ae_123b9358 , 
    R_16cd_117eee78 , 
    R_1a2b_140accb8 , 
    R_140c_11c6f058 , 
    R_ded_14a14738 , 
    R_7ce_13d45d38 , 
    R_a8f_17014de8 , 
    R_10a5_13d564b8 , 
    R_16c4_1580f878 , 
    R_1a34_14a19558 , 
    R_1415_158165d8 , 
    R_df6_156b2bb8 , 
    R_7d7_13c29998 , 
    R_a86_123bc0f8 , 
    R_165b_13de0898 , 
    R_840_156b26b8 , 
    R_a1d_14a15778 , 
    R_147e_11638078 , 
    R_103c_140b0ef8 , 
    R_e5f_150e3d38 , 
    R_11c6_13def038 , 
    R_cd5_13cd09f8 , 
    R_588_13de09d8 , 
    R_1913_13beef18 , 
    R_17e5_150de518 , 
    R_6b6_13d519b8 , 
    R_ba7_13d2ca38 , 
    R_12f4_11c6ca38 , 
    R_19e8_15888e18 , 
    R_1710_13bf6718 , 
    R_10f1_124c52f8 , 
    R_ad2_156b8658 , 
    R_78b_1162ddf8 , 
    R_daa_1008ced8 , 
    R_13c9_13de18d8 , 
    R_11a1_117e91f8 , 
    R_563_13d1ea78 , 
    R_6db_13dd91d8 , 
    R_1319_117f10d8 , 
    R_17c0_15ff4888 , 
    R_b82_13beff58 , 
    R_cfa_14b21ad8 , 
    R_1938_13df6ab8 , 
    R_82a_14a0cfd8 , 
    R_a33_11c70278 , 
    R_1468_158803f8 , 
    R_1052_117f42d8 , 
    R_1671_13dd6898 , 
    R_e49_15ff8f28 , 
    R_1329_14a16ad8 , 
    R_6eb_13d45b58 , 
    R_1191_15881618 , 
    R_1948_13c26a18 , 
    R_d0a_158820b8 , 
    R_b72_13c103f8 , 
    R_17b0_13decf18 , 
    R_a36_13b92438 , 
    R_827_123b8f98 , 
    R_1055_11635738 , 
    R_1465_14a18ab8 , 
    R_1674_11636c78 , 
    R_e46_15884098 , 
    R_851_11635238 , 
    R_148f_13df4358 , 
    R_164a_13c1e318 , 
    R_a0c_100899b8 , 
    R_e70_117ec538 , 
    R_102b_13d38d18 , 
    R_198d_156b4378 , 
    R_730_123bb518 , 
    R_b2d_124c29b8 , 
    R_d4f_13cd15d8 , 
    R_176b_150e5bd8 , 
    R_136e_15ff6b88 , 
    R_114c_140b06d8 , 
    R_16f5_13d39b78 , 
    R_1a03_14b23338 , 
    R_10d6_150df4b8 , 
    R_13e4_13cd99b8 , 
    R_ab7_1700b748 , 
    R_dc5_15ff3f28 , 
    R_7a6_150dad78 , 
    R_1a05_1162d498 , 
    R_13e6_1486e578 , 
    R_dc7_13cd2398 , 
    R_16f3_10088bf8 , 
    R_7a8_13beac38 , 
    R_10d4_13d1de98 , 
    R_ab5_13df25f8 , 
    R_82d_13c24b78 , 
    R_a30_117ef9b8 , 
    R_146b_150da9b8 , 
    R_104f_170118c8 , 
    R_e4c_13ddfd58 , 
    R_166e_123be3f8 , 
    R_73e_15883878 , 
    R_b1f_11631098 , 
    R_d5d_11636778 , 
    R_137c_11634e78 , 
    R_175d_13df13d8 , 
    R_199b_150dc8f8 , 
    R_113e_10081ad8 , 
    R_b45_13cce978 , 
    R_718_123b4fd8 , 
    R_1975_13deedb8 , 
    R_1783_15817e38 , 
    R_d37_13d26d18 , 
    R_1164_13df29b8 , 
    R_1356_15884958 , 
    R_16f7_140b9558 , 
    R_10d8_13d55158 , 
    R_ab9_14a16358 , 
    R_1a01_14a0bf98 , 
    R_7a4_13cca698 , 
    R_13e2_13d50338 , 
    R_dc3_13d5b918 , 
    R_1509_13c080b8 , 
    R_15d0_13d5d7b8 , 
    R_fb1_17011fa8 , 
    R_8cb_1162afb8 , 
    R_992_158117b8 , 
    R_eea_158843b8 , 
    R_1a07_15817f78 , 
    R_13e8_13d57458 , 
    R_dc9_13dedb98 , 
    R_7aa_14a113f8 , 
    R_ab3_13ccea18 , 
    R_16f1_13c2b298 , 
    R_10d2_14a0f4b8 , 
    R_84a_1700eee8 , 
    R_1651_100849b8 , 
    R_1488_15811858 , 
    R_a13_117f7ed8 , 
    R_e69_14b24ff8 , 
    R_1032_15884638 , 
    R_1434_15884a98 , 
    R_a67_1587c9d8 , 
    R_e15_117f6538 , 
    R_1086_158844f8 , 
    R_16a5_1587d018 , 
    R_7f6_14a10318 , 
    R_1a53_11c70b38 , 
    R_f7b_13c24f38 , 
    R_95c_13b8ad78 , 
    R_901_15ff0dc8 , 
    R_f20_11633078 , 
    R_153f_140abef8 , 
    R_159a_13d58d58 , 
    R_1a20_117f5638 , 
    R_1401_14a19918 , 
    R_de2_123bef38 , 
    R_7c3_14a0f058 , 
    R_a9a_15816f38 , 
    R_10b9_15ff6908 , 
    R_16d8_14b209f8 , 
    R_1583_13b8ba98 , 
    R_f64_123b9718 , 
    R_945_123bcaf8 , 
    R_918_13c20ed8 , 
    R_f37_158875b8 , 
    R_1556_140b5db8 , 
    R_a39_17016d28 , 
    R_824_140b4b98 , 
    R_1058_13b8c7b8 , 
    R_1462_13d228f8 , 
    R_1677_1008aef8 , 
    R_e43_140ab8b8 , 
    R_123f_12fc2458 , 
    R_185e_100815d8 , 
    R_189a_15ff14a8 , 
    R_127b_13de1a18 , 
    R_c5c_140b8518 , 
    R_63d_13df0438 , 
    R_601_14a12c58 , 
    R_c20_1486b7d8 , 
    R_15fd_156b4c38 , 
    R_ebd_117f1ad8 , 
    R_fde_13d429f8 , 
    R_14dc_13ddc5b8 , 
    R_9bf_15ff2128 , 
    R_89e_123bbdd8 , 
    R_16f9_13cd6218 , 
    R_10da_14a0d4d8 , 
    R_abb_14b262b8 , 
    R_7a2_13de1fb8 , 
    R_dc1_13c211f8 , 
    R_13e0_1486e4d8 , 
    R_19ff_123b42b8 , 
    R_1739_15ff78a8 , 
    R_d81_140ad4d8 , 
    R_111a_13d42ef8 , 
    R_13a0_117f2bb8 , 
    R_afb_13bf4af8 , 
    R_19bf_117f5e58 , 
    R_762_156b33d8 , 
    R_1a09_1162d358 , 
    R_13ea_1580dc58 , 
    R_dcb_1162f798 , 
    R_7ac_13c08838 , 
    R_ab1_150e1b78 , 
    R_10d0_150e7938 , 
    R_16ef_14a136f8 , 
    R_a6c_123b7378 , 
    R_142f_117f79d8 , 
    R_108b_156b83d8 , 
    R_e10_14a0b4f8 , 
    R_16aa_150e47d8 , 
    R_7f1_123bc378 , 
    R_1a4e_123b60b8 , 
    R_5b2_1486f018 , 
    R_cab_15fee028 , 
    R_bd1_1587dfb8 , 
    R_68c_123c1b98 , 
    R_11f0_13cd3a18 , 
    R_18e9_13b98a18 , 
    R_180f_13c1cbf8 , 
    R_12ca_14a13dd8 , 
    R_1000_13d4e858 , 
    R_e9b_13cd5f98 , 
    R_9e1_13bea878 , 
    R_161f_10080098 , 
    R_14ba_1580ba98 , 
    R_87c_13dee6d8 , 
    R_830_1008cc58 , 
    R_a2d_13d43f38 , 
    R_146e_17010ba8 , 
    R_104c_13d1f658 , 
    R_e4f_13ccef18 , 
    R_166b_116345b8 , 
    R_ff7_13c0cf78 , 
    R_ea4_117ea738 , 
    R_9d8_156b6ad8 , 
    R_1616_17009da8 , 
    R_14c3_116384d8 , 
    R_885_13de02f8 , 
    R_11b7_11c6de38 , 
    R_1922_13c26018 , 
    R_579_13d5d358 , 
    R_6c5_13d59398 , 
    R_17d6_11c6d258 , 
    R_1303_156b3d38 , 
    R_b98_14b1aeb8 , 
    R_ce4_117f17b8 , 
    R_96b_15816c18 , 
    R_8f2_158891d8 , 
    R_f11_124c3598 , 
    R_15a9_1007e0b8 , 
    R_1530_13c1c5b8 , 
    R_f8a_1580da78 , 
    R_5ab_13d20b98 , 
    R_cb2_15883eb8 , 
    R_bca_1162ecf8 , 
    R_693_1580e978 , 
    R_18f0_14868178 , 
    R_11e9_12fc0518 , 
    R_12d1_15ff4388 , 
    R_1808_117ec998 , 
    R_112e_124c40d8 , 
    R_d6d_10080278 , 
    R_b0f_150e1e98 , 
    R_138c_14a12938 , 
    R_19ab_1486d5d8 , 
    R_174d_13c05318 , 
    R_74e_117e9dd8 , 
    R_5d4_1587e918 , 
    R_18c7_117ed7f8 , 
    R_bf3_158826f8 , 
    R_12a8_140b92d8 , 
    R_1212_13debed8 , 
    R_c89_15886078 , 
    R_1831_13b99eb8 , 
    R_66a_117f7c58 , 
    R_16fb_13d39a38 , 
    R_10dc_140acad8 , 
    R_abd_12fbf938 , 
    R_7a0_1162cef8 , 
    R_dbf_13d1dd58 , 
    R_13de_13bf51d8 , 
    R_19fd_13c22cd8 , 
    R_a62_11630378 , 
    R_e1a_13d29f18 , 
    R_1081_156ae298 , 
    R_7fb_13c27c38 , 
    R_16a0_1007f9b8 , 
    R_1a58_123b6a18 , 
    R_1439_11637c18 , 
    R_1511_1162c778 , 
    R_15c8_10085a98 , 
    R_8d3_15fefba8 , 
    R_fa9_150dc218 , 
    R_ef2_13d3af78 , 
    R_98a_11629578 , 
    R_151a_15ff8d48 , 
    R_15bf_15ff4f68 , 
    R_8dc_13dd7b58 , 
    R_fa0_1162a838 , 
    R_efb_13ccc2b8 , 
    R_981_156acad8 , 
    R_133f_11636ef8 , 
    R_179a_13ccf918 , 
    R_701_13dd6438 , 
    R_195e_15817578 , 
    R_117b_156b5f98 , 
    R_d20_1162aa18 , 
    R_b5c_116370d8 , 
    R_c0c_13d3f7f8 , 
    R_122b_117ec498 , 
    R_18ae_13d39998 , 
    R_184a_124c54d8 , 
    R_128f_123b97b8 , 
    R_c70_15885998 , 
    R_651_14a122f8 , 
    R_5ed_13cccad8 , 
    R_1a0b_1486ee38 , 
    R_13ec_117f2758 , 
    R_dcd_13d1e438 , 
    R_7ae_13d3c058 , 
    R_aaf_140af698 , 
    R_10ce_11637538 , 
    R_16ed_156af558 , 
    R_a55_12fbef38 , 
    R_e27_13d405b8 , 
    R_1074_14b1a878 , 
    R_808_13c22c38 , 
    R_1693_13cd4558 , 
    R_1a65_1587f8b8 , 
    R_1446_1587eff8 , 
    R_a3c_150e6038 , 
    R_821_117f1b78 , 
    R_105b_13cd2f78 , 
    R_145f_13b8d398 , 
    R_167a_13df45d8 , 
    R_e40_13c26f18 , 
    R_1584_1580b318 , 
    R_f65_13d3b5b8 , 
    R_946_14a10a98 , 
    R_917_117f5458 , 
    R_f36_14a118f8 , 
    R_1555_15815638 , 
    R_cd0_117f6d58 , 
    R_58d_1587f3b8 , 
    R_17ea_15ffadc8 , 
    R_190e_13bf3d38 , 
    R_6b1_15ffc808 , 
    R_bac_13c0a098 , 
    R_12ef_14b277f8 , 
    R_11cb_15ff6f48 , 
    R_977_1580b1d8 , 
    R_8e6_1580c0d8 , 
    R_15b5_14866f58 , 
    R_f05_123b8ef8 , 
    R_f96_15885538 , 
    R_1524_1162d178 , 
    R_11a5_156b5138 , 
    R_567_13bf17b8 , 
    R_6d7_12fc12d8 , 
    R_1315_123b2698 , 
    R_17c4_13ccc718 , 
    R_b86_123b9a38 , 
    R_cf6_14b29738 , 
    R_1934_123bf7f8 , 
    R_1338_116375d8 , 
    R_6fa_13bec218 , 
    R_1182_13c1c658 , 
    R_1957_13d3ec18 , 
    R_d19_13def3f8 , 
    R_b63_15ffbb88 , 
    R_17a1_117f24d8 , 
    R_132d_1587ce38 , 
    R_6ef_158893b8 , 
    R_118d_124c3958 , 
    R_194c_1587cbb8 , 
    R_d0e_13c10998 , 
    R_b6e_117ef5f8 , 
    R_17ac_1486cb38 , 
    R_12b2_156ab458 , 
    R_be9_14867638 , 
    R_c93_14a12258 , 
    R_1208_13bec358 , 
    R_674_123c0018 , 
    R_1827_13c01b78 , 
    R_18d1_117e98d8 , 
    R_5ca_13ccca38 , 
    R_16fd_13bf4378 , 
    R_10de_140b68f8 , 
    R_abf_13befd78 , 
    R_79e_15817b18 , 
    R_dbd_117f2b18 , 
    R_13dc_13d1ce58 , 
    R_19fb_150e3978 , 
    R_858_150dae18 , 
    R_1496_13b8b098 , 
    R_1643_1162c278 , 
    R_a05_117f4cd8 , 
    R_e77_1486b878 , 
    R_1024_11635058 , 
    R_733_10086998 , 
    R_b2a_150dd2f8 , 
    R_d52_1580c498 , 
    R_1768_15813b58 , 
    R_1371_156b10d8 , 
    R_1149_156aff58 , 
    R_1990_117f1df8 , 
    R_185d_1162a0b8 , 
    R_189b_123bccd8 , 
    R_127c_1580f198 , 
    R_c5d_13bf88d8 , 
    R_63e_170163c8 , 
    R_600_150e8798 , 
    R_c1f_117ebdb8 , 
    R_123e_13ccb318 , 
    R_bfe_17018b28 , 
    R_18bc_123b9df8 , 
    R_121d_11632718 , 
    R_129d_117f6998 , 
    R_183c_14b21498 , 
    R_c7e_14a0d6b8 , 
    R_65f_14874978 , 
    R_5df_13c24178 , 
    R_833_117f3dd8 , 
    R_a2a_14869bb8 , 
    R_1471_140adbb8 , 
    R_1049_11636138 , 
    R_e52_13d4e498 , 
    R_1668_13b909f8 , 
    R_15df_14b24c38 , 
    R_14fa_15ff7128 , 
    R_fc0_13beba98 , 
    R_8bc_14a0e338 , 
    R_9a1_123b5758 , 
    R_edb_17017048 , 
    R_1a0d_13ccaaf8 , 
    R_13ee_13d23398 , 
    R_dcf_13cccfd8 , 
    R_7b0_123bf4d8 , 
    R_aad_14873a78 , 
    R_10cc_13cd01d8 , 
    R_16eb_150e81f8 , 
    R_172d_13cda318 , 
    R_13ac_116343d8 , 
    R_110e_14a11998 , 
    R_19cb_13d3a758 , 
    R_aef_13d50dd8 , 
    R_76e_13bf8d38 , 
    R_d8d_13dd52b8 , 
    R_715_13b94ff8 , 
    R_1972_156aa918 , 
    R_1786_140b5778 , 
    R_d34_15ff3b68 , 
    R_1167_1587c7f8 , 
    R_1353_123c05b8 , 
    R_b48_15814378 , 
    R_17fb_11c6bd18 , 
    R_59e_13cd0098 , 
    R_cbf_15fed948 , 
    R_bbd_13b8f418 , 
    R_18fd_15882798 , 
    R_6a0_117edbb8 , 
    R_11dc_150db458 , 
    R_12de_117e9658 , 
    R_19db_123b8458 , 
    R_171d_13d45e78 , 
    R_10fe_117ebd18 , 
    R_adf_13ccfcd8 , 
    R_77e_123bcff8 , 
    R_d9d_12fc0298 , 
    R_13bc_13c07cf8 , 
    R_142a_14a0f2d8 , 
    R_1090_1486e7f8 , 
    R_e0b_156b7758 , 
    R_16af_1486be18 , 
    R_7ec_123b4038 , 
    R_1a49_13ccbb38 , 
    R_a71_117f59f8 , 
    R_15f2_13d4fe38 , 
    R_ec8_15883058 , 
    R_fd3_10088798 , 
    R_14e7_14b1ce98 , 
    R_9b4_13bf5b38 , 
    R_8a9_13c21298 , 
    R_ece_11634bf8 , 
    R_15ec_13d3f4d8 , 
    R_14ed_117f5f98 , 
    R_fcd_1580d258 , 
    R_8af_13ddfb78 , 
    R_9ae_140b18f8 , 
    R_1501_117f0a98 , 
    R_15d8_11c6ea18 , 
    R_fb9_15ff0be8 , 
    R_8c3_10081498 , 
    R_99a_15ffaaa8 , 
    R_ee2_13cd1b78 , 
    R_1712_11637178 , 
    R_10f3_14a19238 , 
    R_ad4_14a0a5f8 , 
    R_789_140b2cf8 , 
    R_da8_140b3838 , 
    R_13c7_13df0ed8 , 
    R_19e6_11636958 , 
    R_95d_117f8338 , 
    R_900_140b74d8 , 
    R_f1f_1587f1d8 , 
    R_153e_13d410f8 , 
    R_159b_1162f658 , 
    R_f7c_15ffc268 , 
    R_cc5_13b8c858 , 
    R_598_17015108 , 
    R_17f5_13c1c798 , 
    R_1903_1162d2b8 , 
    R_6a6_15816df8 , 
    R_bb7_14a17a78 , 
    R_12e4_13df4678 , 
    R_11d6_13cccf38 , 
    R_a4d_14a159f8 , 
    R_810_1007f918 , 
    R_106c_13cd4238 , 
    R_168b_13d20d78 , 
    R_144e_17019028 , 
    R_e2f_123b83b8 , 
    R_f66_1700e448 , 
    R_947_13cd36f8 , 
    R_916_12fbefd8 , 
    R_f35_13dd5fd8 , 
    R_1554_13c04918 , 
    R_1585_117efe18 , 
    R_16ff_13b95318 , 
    R_10e0_1580e478 , 
    R_ac1_13d23078 , 
    R_79c_1162d8f8 , 
    R_dbb_1580e018 , 
    R_13da_123c03d8 , 
    R_19f9_13cd81f8 , 
    R_a3f_13c012b8 , 
    R_81e_140b4cd8 , 
    R_105e_156ba278 , 
    R_145c_13ddc0b8 , 
    R_167d_124c5438 , 
    R_e3d_15889778 , 
    R_be0_117ea5f8 , 
    R_c9c_13b8ed38 , 
    R_11ff_14a17618 , 
    R_67d_156b7398 , 
    R_181e_13c04e18 , 
    R_18da_13cd38d8 , 
    R_5c1_13c0a818 , 
    R_12bb_13b8a918 , 
    R_ca4_156b1c18 , 
    R_bd8_117e87f8 , 
    R_685_13bf38d8 , 
    R_11f7_10080b38 , 
    R_18e2_13becfd8 , 
    R_1816_14b1ff58 , 
    R_12c3_10083478 , 
    R_5b9_140b2bb8 , 
    R_1630_123b9cb8 , 
    R_e8a_14b1db18 , 
    R_9f2_10089418 , 
    R_14a9_156acb78 , 
    R_1011_12fbe218 , 
    R_86b_124c4e98 , 
    R_1726_14869a78 , 
    R_19d2_13d533f8 , 
    R_1107_13df9038 , 
    R_ae8_13bef5f8 , 
    R_775_158109f8 , 
    R_d94_12fbf6b8 , 
    R_13b3_13d40158 , 
    R_1658_13bf9ff8 , 
    R_843_150e0458 , 
    R_1481_117e8e38 , 
    R_a1a_15fefd88 , 
    R_1039_13ddba78 , 
    R_e62_13c23098 , 
    R_1a0f_13c24038 , 
    R_13f0_11c6e338 , 
    R_dd1_13de4a38 , 
    R_7b2_13bf2898 , 
    R_aab_13c1cfb8 , 
    R_10ca_1700ac08 , 
    R_16e9_15ff3668 , 
    R_1793_150de018 , 
    R_708_14a0d258 , 
    R_1965_13ccb6d8 , 
    R_1174_11c6c358 , 
    R_d27_13dee138 , 
    R_b55_15ffb0e8 , 
    R_1346_13d3f2f8 , 
    R_e1f_123b6ab8 , 
    R_107c_117f4058 , 
    R_800_13d219f8 , 
    R_169b_150e49b8 , 
    R_1a5d_1486e398 , 
    R_143e_14a19f58 , 
    R_a5d_15880498 , 
    R_1a22_15810b38 , 
    R_1403_124c5398 , 
    R_de4_117f6498 , 
    R_7c5_15ffbe08 , 
    R_a98_1486db78 , 
    R_10b7_14a17578 , 
    R_16d6_14a10458 , 
    R_1a2d_13b8fcd8 , 
    R_140e_13def718 , 
    R_def_13d3eb78 , 
    R_7d0_156b2e38 , 
    R_a8d_11632678 , 
    R_10ac_156b5958 , 
    R_16cb_156b72f8 , 
    R_1634_17018c68 , 
    R_9f6_158867f8 , 
    R_e86_14a183d8 , 
    R_1015_14b1e6f8 , 
    R_867_15881398 , 
    R_14a5_11629ed8 , 
    R_e8e_150da878 , 
    R_9ee_13d54618 , 
    R_162c_13b96c18 , 
    R_14ad_12fbf618 , 
    R_86f_15ff83e8 , 
    R_100d_158136f8 , 
    R_189c_14a10c78 , 
    R_127d_11636318 , 
    R_c5e_15882a18 , 
    R_63f_156b5b38 , 
    R_5ff_13d40ab8 , 
    R_c1e_14a0b958 , 
    R_123d_13ddd5f8 , 
    R_185c_11630738 , 
    R_141e_13b90818 , 
    R_16bb_123b7d78 , 
    R_dff_117eeb58 , 
    R_7e0_13dfacf8 , 
    R_a7d_123b7af8 , 
    R_1a3d_156b9cd8 , 
    R_109c_13b98d38 , 
    R_cb9_150db638 , 
    R_bc3_156b6678 , 
    R_69a_13b8b6d8 , 
    R_18f7_13b90bd8 , 
    R_11e2_13d1e4d8 , 
    R_12d8_13d43718 , 
    R_1801_13c013f8 , 
    R_5a4_15ff7d08 , 
    R_13a5_13d45338 , 
    R_1115_11630b98 , 
    R_19c4_17016fa8 , 
    R_af6_117f49b8 , 
    R_767_117f2d98 , 
    R_d86_15fef7e8 , 
    R_1734_1580c718 , 
    R_836_123b33b8 , 
    R_a27_117ede38 , 
    R_1474_13c042d8 , 
    R_1046_123bc918 , 
    R_e55_124c3a98 , 
    R_1665_156ac678 , 
    R_122a_14a0b318 , 
    R_18af_11c6f7d8 , 
    R_1849_140b6358 , 
    R_1290_13dd8b98 , 
    R_c71_14a11e98 , 
    R_652_13d386d8 , 
    R_5ec_14868df8 , 
    R_c0b_13b8c038 , 
    R_574_13d4ec18 , 
    R_6ca_156b3f18 , 
    R_1308_117f2438 , 
    R_17d1_11c6fa58 , 
    R_b93_15881078 , 
    R_ce9_156b86f8 , 
    R_1927_123bb6f8 , 
    R_11b2_14a101d8 , 
    R_8f1_14a0fcd8 , 
    R_f10_156ab778 , 
    R_15aa_13c1f498 , 
    R_152f_158884b8 , 
    R_f8b_13dda218 , 
    R_96c_15ff4e28 , 
    R_948_15ff1728 , 
    R_915_158834b8 , 
    R_f34_123bd958 , 
    R_1553_1162fdd8 , 
    R_1586_13cd7938 , 
    R_f67_156b54f8 , 
    R_1701_117ee5b8 , 
    R_10e2_13b97cf8 , 
    R_ac3_13d41ff8 , 
    R_79a_13b8d758 , 
    R_db9_13d4e358 , 
    R_13d8_13c10178 , 
    R_19f7_123b4218 , 
    R_ec2_156acdf8 , 
    R_fd9_13cd6038 , 
    R_14e1_13d4fbb8 , 
    R_9ba_13d3b018 , 
    R_8a3_117f3298 , 
    R_15f8_150dd618 , 
    R_b1c_10084238 , 
    R_d60_1700c1e8 , 
    R_137f_13d27fd8 , 
    R_175a_15fedda8 , 
    R_199e_123b8d18 , 
    R_113b_11c703b8 , 
    R_741_156b0278 , 
    R_15e6_140b4238 , 
    R_14f3_10088a18 , 
    R_fc7_117e8c58 , 
    R_8b5_13ccefb8 , 
    R_9a8_14a19af8 , 
    R_ed4_150e1998 , 
    R_d68_15885b78 , 
    R_b14_11c6b8b8 , 
    R_1387_117eaf58 , 
    R_19a6_14a19738 , 
    R_1752_150e4738 , 
    R_749_123b2918 , 
    R_1133_1587e378 , 
    R_1417_15ff4428 , 
    R_df8_15888eb8 , 
    R_7d9_124c3098 , 
    R_a84_13b8b778 , 
    R_10a3_13c1e4f8 , 
    R_1a36_14b1b318 , 
    R_16c2_156b1e98 , 
    R_1a11_123b7b98 , 
    R_13f2_13de2738 , 
    R_dd3_14a19a58 , 
    R_7b4_15885a38 , 
    R_aa9_13cd5818 , 
    R_10c8_14a14058 , 
    R_16e7_117eea18 , 
    R_b27_10087e38 , 
    R_d55_117f0f98 , 
    R_1765_12fbdf98 , 
    R_1374_17015888 , 
    R_1146_123bed58 , 
    R_1993_13d53b78 , 
    R_736_15ff9108 , 
    R_56b_123b7558 , 
    R_6d3_1007e1f8 , 
    R_1311_10087a78 , 
    R_17c8_13d50a18 , 
    R_b8a_14b26858 , 
    R_cf2_14a17438 , 
    R_1930_13c083d8 , 
    R_11a9_117f1038 , 
    R_1638_15815818 , 
    R_9fa_123b77d8 , 
    R_e82_13df3ef8 , 
    R_1019_158858f8 , 
    R_863_13d47318 , 
    R_14a1_117ed938 , 
    R_eb2_11c6d2f8 , 
    R_fe9_1162ed98 , 
    R_14d1_1587ae58 , 
    R_9ca_1587bd58 , 
    R_893_13ccf238 , 
    R_1608_117f45f8 , 
    R_6f3_17012cc8 , 
    R_1189_13de2d78 , 
    R_1950_123b8098 , 
    R_d12_13cd6d58 , 
    R_b6a_140afff8 , 
    R_17a8_13d3cf58 , 
    R_1331_148755f8 , 
    R_e9f_17016288 , 
    R_9dd_156ab8b8 , 
    R_161b_13d3ca58 , 
    R_14be_13b98478 , 
    R_880_117ea2d8 , 
    R_ffc_13b8acd8 , 
    R_1789_13cca9b8 , 
    R_196f_13bf01d8 , 
    R_d31_156b13f8 , 
    R_116a_13c23e58 , 
    R_1350_11632498 , 
    R_b4b_156ad398 , 
    R_712_13b90d18 , 
    R_e92_117f2ed8 , 
    R_9ea_123b7e18 , 
    R_1628_123b7698 , 
    R_14b1_14a16e98 , 
    R_873_14a14238 , 
    R_1009_13b980b8 , 
    R_bf2_170099e8 , 
    R_12a9_1162d0d8 , 
    R_1211_150e5278 , 
    R_c8a_150e3798 , 
    R_1830_13bf6358 , 
    R_66b_150e1498 , 
    R_5d3_158808f8 , 
    R_18c8_13cd9f58 , 
    R_a42_15888198 , 
    R_81b_12fbec18 , 
    R_1061_13d3c558 , 
    R_1459_17016aa8 , 
    R_1680_1486aab8 , 
    R_e3a_123bb798 , 
    R_17ef_15889958 , 
    R_1909_15815e58 , 
    R_6ac_12fc1918 , 
    R_bb1_14874d38 , 
    R_12ea_13ddf358 , 
    R_11d0_170096c8 , 
    R_ccb_117ec038 , 
    R_592_13c23958 , 
    R_fee_14b29f58 , 
    R_ead_13c22378 , 
    R_9cf_1162e118 , 
    R_14cc_123c0b58 , 
    R_160d_123bff78 , 
    R_88e_123c0fb8 , 
    R_8ff_156b7c58 , 
    R_f1e_15880038 , 
    R_153d_15811218 , 
    R_159c_15815db8 , 
    R_f7d_13cd0778 , 
    R_95e_13b98018 , 
    R_189d_13cd3518 , 
    R_127e_13d4f118 , 
    R_c5f_12fbfa78 , 
    R_640_140b2258 , 
    R_5fe_15888558 , 
    R_c1d_13dfb1f8 , 
    R_123c_15fee708 , 
    R_185b_14b21538 , 
    R_15d1_123b63d8 , 
    R_fb2_15810818 , 
    R_8ca_15815bd8 , 
    R_993_11c6b598 , 
    R_ee9_1700fca8 , 
    R_1508_156b7898 , 
    R_121c_158871f8 , 
    R_129e_13d3cb98 , 
    R_183b_13c20bb8 , 
    R_c7f_13cd6ad8 , 
    R_660_156ba458 , 
    R_5de_123b7cd8 , 
    R_18bd_140b9878 , 
    R_bfd_11c6f238 , 
    R_16b4_117ead78 , 
    R_e06_1580ff58 , 
    R_7e7_15885858 , 
    R_1a44_1162c4f8 , 
    R_a76_13d38638 , 
    R_1095_156b0ef8 , 
    R_1425_13d571d8 , 
    R_8e5_150db318 , 
    R_15b6_1580e838 , 
    R_f04_15885038 , 
    R_f97_1700c288 , 
    R_1523_140b8e78 , 
    R_978_156b6498 , 
    R_914_13d54c58 , 
    R_f33_13d59258 , 
    R_1552_13ccfa58 , 
    R_1587_140aacd8 , 
    R_f68_140acb78 , 
    R_949_14b26a38 , 
    R_15c0_158147d8 , 
    R_8db_1580e158 , 
    R_fa1_1162ffb8 , 
    R_efa_13bf5818 , 
    R_982_13debcf8 , 
    R_1519_15813e78 , 
    R_164e_117eb138 , 
    R_148b_15886118 , 
    R_a10_13df0f78 , 
    R_e6c_15ff0d28 , 
    R_102f_123c08d8 , 
    R_84d_15feee88 , 
    R_1703_13c254d8 , 
    R_10e4_158894f8 , 
    R_ac5_15883558 , 
    R_798_123beb78 , 
    R_db7_14869938 , 
    R_13d6_156ae8d8 , 
    R_19f5_13d2c2b8 , 
    R_eb7_11c6d1b8 , 
    R_fe4_12fc21d8 , 
    R_14d6_1008b178 , 
    R_9c5_14b21d58 , 
    R_898_123b5c58 , 
    R_1603_14872fd8 , 
    R_1714_15889638 , 
    R_10f5_140b5f98 , 
    R_ad6_14873258 , 
    R_787_14a0e838 , 
    R_da6_13ddc158 , 
    R_13c5_15fee208 , 
    R_19e4_13de3a98 , 
    R_98b_13b8dcf8 , 
    R_ef1_13b924d8 , 
    R_8d2_156ad578 , 
    R_faa_156b0458 , 
    R_1510_13d1f0b8 , 
    R_15c9_13bf0b38 , 
    R_aa7_13d451f8 , 
    R_7b6_14a18018 , 
    R_dd5_124c5258 , 
    R_10c6_1700ff28 , 
    R_13f4_14a0b778 , 
    R_16e5_13c07ed8 , 
    R_1a13_117ef058 , 
    R_839_14b28f18 , 
    R_e58_158814d8 , 
    R_a24_123b5938 , 
    R_1043_14b26538 , 
    R_1477_117f0098 , 
    R_1662_13df1978 , 
    R_854_15ff3e88 , 
    R_e73_14b288d8 , 
    R_a09_123bb158 , 
    R_1028_117f4eb8 , 
    R_1492_13cd4378 , 
    R_1647_12fc19b8 , 
    R_be8_15ffcee8 , 
    R_5c9_14b27438 , 
    R_675_156aec98 , 
    R_c94_13b8fb98 , 
    R_1207_156b81f8 , 
    R_12b3_13ddf718 , 
    R_1826_140b01d8 , 
    R_18d2_13c290d8 , 
    R_cac_123c1058 , 
    R_5b1_13d28e38 , 
    R_68d_1700f2a8 , 
    R_bd0_13ccc538 , 
    R_11ef_117f3d38 , 
    R_12cb_123bfe38 , 
    R_180e_1580c7b8 , 
    R_18ea_14a115d8 , 
    R_d75_1486bc38 , 
    R_756_13b8ae18 , 
    R_b07_140aaa58 , 
    R_1126_156aaeb8 , 
    R_1394_15814878 , 
    R_1745_123b4cb8 , 
    R_19b3_123bc558 , 
    R_d7a_13b95ef8 , 
    R_75b_15814558 , 
    R_b02_14a13f18 , 
    R_1121_150e9c38 , 
    R_1399_158830f8 , 
    R_1740_13cd6fd8 , 
    R_19b8_15812c58 , 
    R_c0a_14a19ff8 , 
    R_5eb_15feeac8 , 
    R_653_123be358 , 
    R_c72_13df6fb8 , 
    R_1229_156b7938 , 
    R_1291_14a0d758 , 
    R_1848_14a197d8 , 
    R_18b0_15815a98 , 
    R_a96_150e8478 , 
    R_7c7_13d45c98 , 
    R_de6_13c05778 , 
    R_10b5_156ab6d8 , 
    R_1405_14a192d8 , 
    R_16d4_14868c18 , 
    R_1a24_116348d8 , 
    R_85f_13dd89b8 , 
    R_e7e_140ad6b8 , 
    R_9fe_13c02d98 , 
    R_101d_123b5d98 , 
    R_149d_156b8dd8 , 
    R_163c_1486a6f8 , 
    R_d9b_13d3dbd8 , 
    R_77c_116359b8 , 
    R_ae1_15fed768 , 
    R_1100_10085818 , 
    R_13ba_15881d98 , 
    R_171f_13bf08b8 , 
    R_19d9_1700c508 , 
    R_889_15ff9b08 , 
    R_9d4_11c6e6f8 , 
    R_ea8_13d1fe78 , 
    R_ff3_117efc38 , 
    R_14c7_140b4918 , 
    R_1612_13cd0278 , 
    R_582_14869118 , 
    R_cdb_14a0ae18 , 
    R_ba1_13d29338 , 
    R_6bc_13cd53b8 , 
    R_11c0_13deef98 , 
    R_12fa_11631638 , 
    R_17df_13cd0e58 , 
    R_1919_1587e2d8 , 
    R_e24_13ddcfb8 , 
    R_a58_14a18a18 , 
    R_805_1580a7d8 , 
    R_1077_11c6d898 , 
    R_1443_13d3f9d8 , 
    R_1696_156afd78 , 
    R_1a62_14b1b138 , 
    R_94a_156b24d8 , 
    R_f32_116350f8 , 
    R_913_100840f8 , 
    R_f69_117f0c78 , 
    R_1551_150dde38 , 
    R_1588_150e7d98 , 
    R_a50_13df7698 , 
    R_e2c_15881e38 , 
    R_80d_14a16a38 , 
    R_106f_156ad938 , 
    R_144b_1486ce58 , 
    R_168e_123bbc98 , 
    R_6fe_13bf5318 , 
    R_b5f_13cd4918 , 
    R_d1d_13def2b8 , 
    R_117e_14a0ccb8 , 
    R_133c_117f2938 , 
    R_179d_10085138 , 
    R_195b_14b1c8f8 , 
    R_cb3_1587b358 , 
    R_5aa_13dd5678 , 
    R_694_11636b38 , 
    R_bc9_124c3d18 , 
    R_11e8_13ccd258 , 
    R_12d2_123bdc78 , 
    R_1807_117ee298 , 
    R_18f1_156aba98 , 
    R_c1c_156ba3b8 , 
    R_5fd_14a10958 , 
    R_641_123b90d8 , 
    R_c60_158171b8 , 
    R_123b_1162cd18 , 
    R_127f_13b8a558 , 
    R_185a_15814cd8 , 
    R_189e_13bf8e78 , 
    R_877_13d3e498 , 
    R_9e6_14b28838 , 
    R_e96_156b4a58 , 
    R_1005_13c1edb8 , 
    R_14b5_15882018 , 
    R_1624_10086cb8 , 
    R_db5_117ece98 , 
    R_796_156b0138 , 
    R_ac7_148725d8 , 
    R_10e6_11630918 , 
    R_13d4_15882bf8 , 
    R_1705_10085db8 , 
    R_19f3_1008c618 , 
    R_96d_1162e7f8 , 
    R_f0f_13d3d9f8 , 
    R_8f0_13d29838 , 
    R_f8c_117f2578 , 
    R_152e_117f3f18 , 
    R_15ab_13ccc358 , 
    R_587_124c5118 , 
    R_cd6_13d39178 , 
    R_ba6_156ad9d8 , 
    R_6b7_13c0b718 , 
    R_11c5_13d39538 , 
    R_12f5_158104f8 , 
    R_17e4_156acf38 , 
    R_1914_10084f58 , 
    R_846_100885b8 , 
    R_e65_15810318 , 
    R_a17_13ccf878 , 
    R_1036_140b5278 , 
    R_1484_11c6b778 , 
    R_1655_1700cdc8 , 
    R_a45_17017188 , 
    R_e37_10083018 , 
    R_818_13b8dbb8 , 
    R_1064_1700d5e8 , 
    R_1456_13cd8518 , 
    R_1683_1587f6d8 , 
    R_57d_14b1ef18 , 
    R_ce0_1580ccb8 , 
    R_b9c_15884e58 , 
    R_6c1_156b1538 , 
    R_11bb_117ed2f8 , 
    R_12ff_17012408 , 
    R_17da_123bf398 , 
    R_191e_140b0c78 , 
    R_d58_13df39f8 , 
    R_b24_15815958 , 
    R_739_123c1698 , 
    R_1143_13cd7078 , 
    R_1377_158873d8 , 
    R_1762_140aef18 , 
    R_1996_156b4058 , 
    R_95f_13bf9918 , 
    R_f1d_15ff80c8 , 
    R_8fe_13d4f898 , 
    R_f7e_156b42d8 , 
    R_153c_13c1d698 , 
    R_159d_1162b198 , 
    R_aa5_156b4238 , 
    R_7b8_1162e9d8 , 
    R_dd7_140b62b8 , 
    R_10c4_12fc1878 , 
    R_13f6_1700d728 , 
    R_16e3_123b4d58 , 
    R_1a15_13d3e998 , 
    R_b0c_123c1878 , 
    R_d70_13b96038 , 
    R_751_13bf12b8 , 
    R_112b_13d5c3b8 , 
    R_138f_13df66f8 , 
    R_174a_13d24658 , 
    R_19ae_1587f818 , 
    R_a8b_117f7898 , 
    R_7d2_10082a78 , 
    R_df1_15884778 , 
    R_10aa_13c28458 , 
    R_1410_13cd5a98 , 
    R_16c9_13c03018 , 
    R_1a2f_15886b18 , 
    R_d7f_117f5ef8 , 
    R_760_13cce6f8 , 
    R_afd_156ae018 , 
    R_111c_13c0f138 , 
    R_139e_15ff9428 , 
    R_173b_13d23758 , 
    R_19bd_150e0c78 , 
    R_70f_14b26038 , 
    R_b4e_158835f8 , 
    R_d2e_15ff2d08 , 
    R_116d_14a0bc78 , 
    R_134d_13cd26b8 , 
    R_178c_13d39718 , 
    R_196c_117ef418 , 
    R_705_17018768 , 
    R_b58_12fc00b8 , 
    R_d24_13c0ca78 , 
    R_1177_13d5b558 , 
    R_1343_13d298d8 , 
    R_1796_156ae338 , 
    R_1962_13d5d218 , 
    R_c9d_13c00ef8 , 
    R_bdf_117f0638 , 
    R_5c0_117ea0f8 , 
    R_67e_14a0b8b8 , 
    R_11fe_124c36d8 , 
    R_12bc_13b981f8 , 
    R_181d_123ba758 , 
    R_18db_11c6d7f8 , 
    R_ebc_1580cfd8 , 
    R_89d_11c693d8 , 
    R_9c0_13d46b98 , 
    R_fdf_158176b8 , 
    R_14db_156b5e58 , 
    R_15fe_140b97d8 , 
    R_ee1_13d40c98 , 
    R_99b_156b3838 , 
    R_8c2_15813518 , 
    R_fba_140aebf8 , 
    R_1500_1700e8a8 , 
    R_15d9_13d53538 , 
    R_eda_13d57638 , 
    R_9a2_13c28bd8 , 
    R_8bb_13d43498 , 
    R_fc1_156b40f8 , 
    R_14f9_13cd6178 , 
    R_15e0_13cd0458 , 
    R_d8b_150dc7b8 , 
    R_76c_150e63f8 , 
    R_af1_13b8c3f8 , 
    R_1110_13d5cdb8 , 
    R_13aa_14b1d898 , 
    R_172f_11c6dbb8 , 
    R_19c9_1509b4f8 , 
    R_55a_158145f8 , 
    R_6e4_11630a58 , 
    R_b79_13ccfd78 , 
    R_d03_124c2eb8 , 
    R_1198_117f3b58 , 
    R_1322_15ff6ea8 , 
    R_17b7_15810bd8 , 
    R_1941_117ed4d8 , 
    R_6cf_1486c6d8 , 
    R_56f_14a0b598 , 
    R_cee_13cd9c38 , 
    R_b8e_150e97d8 , 
    R_11ad_13d569b8 , 
    R_130d_124c3818 , 
    R_17cc_117e9298 , 
    R_192c_13b94918 , 
    R_94b_100881f8 , 
    R_f31_13c231d8 , 
    R_912_11630f58 , 
    R_f6a_117ea058 , 
    R_1550_17014668 , 
    R_1589_123b7198 , 
    R_bd7_14a0ef18 , 
    R_ca5_1007eb58 , 
    R_5b8_170170e8 , 
    R_686_15810f98 , 
    R_11f6_14b22bb8 , 
    R_12c4_15ff0008 , 
    R_1815_156b1cb8 , 
    R_18e3_13ccb9f8 , 
    R_6e0_14a15f98 , 
    R_55e_148707d8 , 
    R_cff_14a0b458 , 
    R_b7d_156b6df8 , 
    R_119c_14872ad8 , 
    R_131e_13dd6e38 , 
    R_17bb_13bf1d58 , 
    R_193d_11c70638 , 
    R_d92_14b21358 , 
    R_773_117f54f8 , 
    R_aea_17012908 , 
    R_1109_15ff3de8 , 
    R_13b1_150dc358 , 
    R_1728_13d5beb8 , 
    R_19d0_14870af8 , 
    R_e12_13b8cc18 , 
    R_a6a_13d1d218 , 
    R_7f3_148688f8 , 
    R_1089_123b6838 , 
    R_1431_15812ed8 , 
    R_16a8_123bf118 , 
    R_1a50_117ed6b8 , 
    R_6f7_117e93d8 , 
    R_b66_14a0f238 , 
    R_d16_13c1b7f8 , 
    R_1185_13d1ecf8 , 
    R_1335_13bf1f38 , 
    R_17a4_14b1ea18 , 
    R_1954_15ff1ae8 , 
    R_e17_13df86d8 , 
    R_a65_14b22b18 , 
    R_7f8_1700bec8 , 
    R_1084_13d39038 , 
    R_1436_15fef608 , 
    R_16a3_15ff2768 , 
    R_1a55_123b5898 , 
    R_a21_1587bad8 , 
    R_83c_13cd7398 , 
    R_e5b_123bf898 , 
    R_1040_1008ac78 , 
    R_147a_13c04378 , 
    R_165f_13cd97d8 , 
    R_bfc_13d53cb8 , 
    R_5dd_123b45d8 , 
    R_661_13d3c2d8 , 
    R_c80_1008ca78 , 
    R_121b_14b24698 , 
    R_129f_1008b7b8 , 
    R_183a_156acc18 , 
    R_18be_14a0de38 , 
    R_c1b_123b48f8 , 
    R_5fc_140b3518 , 
    R_642_14a0d118 , 
    R_c61_13c06718 , 
    R_123a_15ffcf88 , 
    R_1280_14a106d8 , 
    R_1859_13d25378 , 
    R_189f_14a13c98 , 
    R_556_13d2a2d8 , 
    R_6e8_12fbf4d8 , 
    R_b75_156ae838 , 
    R_d07_156abe58 , 
    R_1194_1580f058 , 
    R_1326_11c684d8 , 
    R_17b3_13ddb4d8 , 
    R_1945_14b22898 , 
    R_bf1_13df18d8 , 
    R_5d2_10088f18 , 
    R_66c_123c06f8 , 
    R_c8b_13c0e5f8 , 
    R_1210_117f56d8 , 
    R_12aa_140afb98 , 
    R_182f_13d58998 , 
    R_18c9_11c6eb58 , 
    R_cc0_1580fcd8 , 
    R_59d_13df9d58 , 
    R_6a1_13cd9b98 , 
    R_bbc_13d4e678 , 
    R_11db_124c45d8 , 
    R_12df_13d27178 , 
    R_17fa_13beb8b8 , 
    R_18fe_1587ca78 , 
    R_d63_117f68f8 , 
    R_b19_158882d8 , 
    R_744_123bea38 , 
    R_1138_14869ed8 , 
    R_1382_13b8b958 , 
    R_1757_13de1978 , 
    R_19a1_123b3598 , 
    R_db3_14869898 , 
    R_794_17016788 , 
    R_ac9_15811cb8 , 
    R_10e8_140b1538 , 
    R_13d2_13c292b8 , 
    R_1707_13ddd9b8 , 
    R_19f1_13cce518 , 
    R_ecd_13d5b5f8 , 
    R_9af_1587fdb8 , 
    R_8ae_11631778 , 
    R_fce_13c051d8 , 
    R_14ec_156b01d8 , 
    R_15ed_1008af98 , 
    R_da4_13cd7438 , 
    R_785_116381b8 , 
    R_ad8_117f7a78 , 
    R_10f7_1587f598 , 
    R_13c3_13cd0b38 , 
    R_1716_123b6bf8 , 
    R_19e2_13d567d8 , 
    R_58c_1587fe58 , 
    R_cd1_1486dc18 , 
    R_bab_13df0e38 , 
    R_6b2_14867ef8 , 
    R_11ca_123bd9f8 , 
    R_12f0_158817f8 , 
    R_17e9_123bb5b8 , 
    R_190f_15881b18 , 
    R_979_117efcd8 , 
    R_f03_13c06f38 , 
    R_8e4_123b2b98 , 
    R_f98_13d588f8 , 
    R_1522_15817d98 , 
    R_15b7_11636bd8 , 
    R_c09_14a18bf8 , 
    R_5ea_1162b558 , 
    R_654_150e54f8 , 
    R_c73_15810958 , 
    R_1228_150e4ff8 , 
    R_1292_117e9fb8 , 
    R_1847_13d54898 , 
    R_18b1_1162ae78 , 
    R_ec7_10083838 , 
    R_8a8_140b6858 , 
    R_9b5_156b6038 , 
    R_fd4_13bef878 , 
    R_14e6_123be178 , 
    R_15f3_1580b958 , 
    R_6dc_13d56738 , 
    R_562_11630198 , 
    R_cfb_156b77f8 , 
    R_b81_14b23658 , 
    R_11a0_117f1a38 , 
    R_131a_13cd6678 , 
    R_17bf_1162eed8 , 
    R_1939_13b99198 , 
    R_85b_150e9ff8 , 
    R_e7a_13df06b8 , 
    R_a02_13d20378 , 
    R_1021_14873438 , 
    R_1499_13c056d8 , 
    R_1640_15816e98 , 
    R_6c6_14b27a78 , 
    R_578_13c06678 , 
    R_ce5_117e9518 , 
    R_b97_116328f8 , 
    R_11b6_123b6478 , 
    R_1304_150e5a98 , 
    R_17d5_13cd9eb8 , 
    R_1923_10086ad8 , 
    R_aa3_123ba9d8 , 
    R_7ba_17013308 , 
    R_dd9_1587f4f8 , 
    R_10c2_13de4358 , 
    R_13f8_14866c38 , 
    R_16e1_1587e058 , 
    R_1a17_13d3a398 , 
    R_ea3_117f04f8 , 
    R_884_124c4358 , 
    R_9d9_14a0c178 , 
    R_ff8_14a15098 , 
    R_14c2_13d50e78 , 
    R_1617_13de3e58 , 
    R_e0d_13c081f8 , 
    R_a6f_140ab4f8 , 
    R_7ee_117eb4f8 , 
    R_108e_117ecf38 , 
    R_142c_13d55f18 , 
    R_16ad_15885df8 , 
    R_1a4b_13d3a118 , 
    R_e01_13b8ca38 , 
    R_a7b_150e6f38 , 
    R_7e2_116332f8 , 
    R_109a_140adc58 , 
    R_1420_1580acd8 , 
    R_16b9_13b972f8 , 
    R_1a3f_13cd8f18 , 
    R_597_156aeab8 , 
    R_cc6_1486fd38 , 
    R_bb6_13d58fd8 , 
    R_6a7_140b7938 , 
    R_11d5_14871bd8 , 
    R_12e5_14b28bf8 , 
    R_17f4_156b4cd8 , 
    R_1904_140b9058 , 
    R_dfa_1486ff18 , 
    R_a82_116368b8 , 
    R_7db_150dd1b8 , 
    R_10a1_123b8598 , 
    R_1419_13df1b58 , 
    R_16c0_13b994b8 , 
    R_1a38_13ccab98 , 
    R_911_14b22078 , 
    R_94c_123bc7d8 , 
    R_f30_12fbf898 , 
    R_f6b_13c0a6d8 , 
    R_154f_1700ea88 , 
    R_158a_13c25758 , 
    R_d44_13b99418 , 
    R_b38_13d23618 , 
    R_725_13d4f618 , 
    R_1157_14a13298 , 
    R_1363_124c4718 , 
    R_1776_15882518 , 
    R_1982_15816fd8 , 
    R_983_1700b4c8 , 
    R_ef9_1007e338 , 
    R_8da_1587ba38 , 
    R_fa2_15ffaf08 , 
    R_1518_13c09ff8 , 
    R_15c1_13c1e138 , 
    R_d41_13bf8f18 , 
    R_722_14b26fd8 , 
    R_b3b_14a0f378 , 
    R_115a_156af9b8 , 
    R_1360_156aa5f8 , 
    R_1779_13dec3d8 , 
    R_197f_1700ba68 , 
    R_7fd_13d29658 , 
    R_e1c_156b8158 , 
    R_a60_124c2738 , 
    R_107f_13d55ab8 , 
    R_143b_13cd5458 , 
    R_169e_13d59618 , 
    R_1a5a_117ecd58 , 
    R_a94_158121b8 , 
    R_7c9_13c1bb18 , 
    R_de8_13df22d8 , 
    R_10b3_17011328 , 
    R_1407_140b9cd8 , 
    R_16d2_150e0098 , 
    R_1a26_14868678 , 
    R_e9a_14a0e1f8 , 
    R_87b_123b2e18 , 
    R_9e2_148680d8 , 
    R_1001_100877f8 , 
    R_14b9_150dda78 , 
    R_1620_117efff8 , 
    R_bc2_1580b098 , 
    R_cba_13c20118 , 
    R_5a3_13b98298 , 
    R_69b_13bf94b8 , 
    R_11e1_1486a798 , 
    R_12d9_123ba118 , 
    R_1800_15888378 , 
    R_18f8_156ac538 , 
    R_960_13ccf418 , 
    R_f1c_13df79b8 , 
    R_8fd_123b6fb8 , 
    R_f7f_140aa558 , 
    R_153b_117f5d18 , 
    R_159e_14871db8 , 
    R_d47_13d27998 , 
    R_b35_1587cc58 , 
    R_728_140ba318 , 
    R_1154_117e95b8 , 
    R_1366_17015568 , 
    R_1773_156ac2b8 , 
    R_1985_1162c3b8 , 
    R_b11_15883698 , 
    R_d6b_123b8958 , 
    R_74c_150e17b8 , 
    R_1130_13bef0f8 , 
    R_138a_13d25cd8 , 
    R_174f_13df2058 , 
    R_19a9_1486eed8 , 
    R_6ec_13c03b58 , 
    R_b71_140afd78 , 
    R_d0b_1587d158 , 
    R_1190_13c09198 , 
    R_132a_13d44bb8 , 
    R_17af_123b9d58 , 
    R_1949_140b51d8 , 
    R_815_158140f8 , 
    R_a48_13bed6b8 , 
    R_e34_13cd7e38 , 
    R_1067_13b93ab8 , 
    R_1453_15ff99c8 , 
    R_1686_1008c258 , 
    R_af8_148696b8 , 
    R_d84_156b3e78 , 
    R_765_13df9678 , 
    R_1117_140b2398 , 
    R_13a3_123bd598 , 
    R_1736_117f1218 , 
    R_19c2_14871098 , 
    R_d3e_14870198 , 
    R_71f_123b6e78 , 
    R_b3e_11631138 , 
    R_115d_1008bd58 , 
    R_135d_13cd9d78 , 
    R_177c_11629258 , 
    R_197c_13bec8f8 , 
    R_96e_1162bff8 , 
    R_f0e_17010f68 , 
    R_8ef_13dd96d8 , 
    R_f8d_13cd51d8 , 
    R_152d_13d1f8d8 , 
    R_15ac_12fc1418 , 
    R_ee8_13d55658 , 
    R_994_13c086f8 , 
    R_8c9_1162f838 , 
    R_fb3_11c6c7b8 , 
    R_1507_14b218f8 , 
    R_15d2_11c6e978 , 
    R_ed3_13b93018 , 
    R_9a9_140ac3f8 , 
    R_8b4_150e2e38 , 
    R_fc8_14875238 , 
    R_14f2_13cd1718 , 
    R_15e7_150e0e58 , 
    R_c1a_13d3c198 , 
    R_5fb_156b22f8 , 
    R_643_117ea698 , 
    R_c62_1162c598 , 
    R_1239_15817938 , 
    R_1281_158887d8 , 
    R_1858_13bea9b8 , 
    R_18a0_123bfcf8 , 
    R_98c_13c21f18 , 
    R_ef0_13d51418 , 
    R_8d1_12fc06f8 , 
    R_fab_14a127f8 , 
    R_150f_15817398 , 
    R_15ca_156b71b8 , 
    R_c95_123be2b8 , 
    R_be7_1162d858 , 
    R_5c8_15feeca8 , 
    R_676_13d37e18 , 
    R_1206_13ddcc98 , 
    R_12b4_10087938 , 
    R_1825_1486a298 , 
    R_18d3_17018f88 , 
    R_d5b_150e0958 , 
    R_b21_14b21e98 , 
    R_73c_13bec858 , 
    R_1140_13b98798 , 
    R_137a_13dd7018 , 
    R_175f_15ff7f88 , 
    R_1999_117f2118 , 
    R_d4a_13df40d8 , 
    R_b32_13c268d8 , 
    R_72b_11632c18 , 
    R_1151_11638898 , 
    R_1369_117f5138 , 
    R_1770_124c2a58 , 
    R_1988_150dfaf8 , 
    R_db1_13bf06d8 , 
    R_792_13ccb638 , 
    R_acb_13d2a378 , 
    R_10ea_13d2b598 , 
    R_13d0_1700b388 , 
    R_1709_1162a298 , 
    R_19ef_150de1f8 , 
    R_ae3_14b24738 , 
    R_d99_156abef8 , 
    R_77a_13c0f3b8 , 
    R_1102_11632358 , 
    R_13b8_13c29c18 , 
    R_1721_14870f58 , 
    R_19d7_13de38b8 , 
    R_6d8_1580ebf8 , 
    R_566_140b4f58 , 
    R_cf7_13d26778 , 
    R_b85_13df3958 , 
    R_11a4_140b1178 , 
    R_1316_13c24718 , 
    R_17c3_13df1e78 , 
    R_1935_14a13798 , 
    R_a0d_14a0f198 , 
    R_850_1700cbe8 , 
    R_e6f_117ee6f8 , 
    R_102c_156ae3d8 , 
    R_148e_17014208 , 
    R_164b_123b8638 , 
    R_f2f_13ccded8 , 
    R_910_158144b8 , 
    R_94d_13de1dd8 , 
    R_f6c_140aca38 , 
    R_154e_158131f8 , 
    R_158b_123b5078 , 
    R_70c_1162a338 , 
    R_b51_13df4c18 , 
    R_d2b_123bacf8 , 
    R_1170_13ddca18 , 
    R_134a_123bdb38 , 
    R_178f_14a0df78 , 
    R_1969_13c0e918 , 
    R_ec1_13c0ddd8 , 
    R_8a2_13dd9638 , 
    R_9bb_14a13d38 , 
    R_fda_14876098 , 
    R_14e0_117ea9b8 , 
    R_15f9_13d4fcf8 , 
    R_d3b_150e4a58 , 
    R_71c_150dba98 , 
    R_b41_100844b8 , 
    R_1160_14a16498 , 
    R_135a_156b8838 , 
    R_177f_13ccedd8 , 
    R_1979_156ad7f8 , 
    R_80a_11c686b8 , 
    R_a53_13d54ed8 , 
    R_e29_124c3138 , 
    R_1072_13d5c598 , 
    R_1448_156b5098 , 
    R_1691_13bf8478 , 
    R_1a67_13d3a898 , 
    R_aa1_13ccbd18 , 
    R_7bc_13ccc218 , 
    R_ddb_15812618 , 
    R_10c0_15816d58 , 
    R_13fa_14b29a58 , 
    R_16df_10084eb8 , 
    R_1a19_11c70a98 , 
    R_a1e_13de1338 , 
    R_83f_123bc5f8 , 
    R_e5e_13c25258 , 
    R_103d_123b2738 , 
    R_147d_13d53e98 , 
    R_165c_123b57f8 , 
    R_c74_14b242d8 , 
    R_c08_13ded7d8 , 
    R_5e9_15816178 , 
    R_655_13c026b8 , 
    R_1227_123b72d8 , 
    R_1293_1008c6b8 , 
    R_1846_13c22af8 , 
    R_18b2_150dd4d8 , 
    R_a14_11632038 , 
    R_849_123c1af8 , 
    R_e68_15887658 , 
    R_1033_13bf8518 , 
    R_1487_1007fc38 , 
    R_1652_11635418 , 
    R_68e_11630eb8 , 
    R_bcf_1486c4f8 , 
    R_cad_150e5c78 , 
    R_5b0_13d20c38 , 
    R_11ee_13df5938 , 
    R_12cc_156aee78 , 
    R_180d_13d29dd8 , 
    R_18eb_13cd2bb8 , 
    R_7e9_13b903b8 , 
    R_e08_14a11498 , 
    R_a74_13c02a78 , 
    R_1093_123bddb8 , 
    R_1427_1580dd98 , 
    R_16b2_123b89f8 , 
    R_1a46_150dff58 , 
    R_c81_140ac718 , 
    R_bfb_117e8f78 , 
    R_5dc_13cd21b8 , 
    R_662_11c6af58 , 
    R_121a_13dd6bb8 , 
    R_12a0_156af7d8 , 
    R_1839_10083a18 , 
    R_18bf_13cd63f8 , 
    R_d4d_14b1c218 , 
    R_b2f_14a168f8 , 
    R_72e_15885178 , 
    R_114e_14866878 , 
    R_136c_13d5ce58 , 
    R_176d_15883e18 , 
    R_198b_123ba938 , 
    R_bb0_11635198 , 
    R_6ad_14b295f8 , 
    R_591_123b56b8 , 
    R_ccc_13c02f78 , 
    R_11cf_13dedd78 , 
    R_12eb_156ab598 , 
    R_17ee_117f2a78 , 
    R_190a_1162b238 , 
    R_7d4_14a0fe18 , 
    R_df3_14b1e478 , 
    R_a89_13dd9278 , 
    R_10a8_13d52958 , 
    R_1412_11c6f198 , 
    R_16c7_13d27d58 , 
    R_1a31_140b9d78 , 
    R_c19_1700d408 , 
    R_5fa_13df88b8 , 
    R_644_13d23938 , 
    R_c63_1162e258 , 
    R_1238_13df9a38 , 
    R_1282_13c2acf8 , 
    R_1857_13cd2ed8 , 
    R_18a1_156aefb8 , 
    R_6f0_140ae658 , 
    R_b6d_123b4178 , 
    R_d0f_150df0f8 , 
    R_118c_14a17898 , 
    R_132e_13bed758 , 
    R_17ab_13cd0d18 , 
    R_194d_1008c438 , 
    R_802_13d3e5d8 , 
    R_e21_14a0aaf8 , 
    R_a5b_13bf7e38 , 
    R_107a_13d1ed98 , 
    R_1440_124c4d58 , 
    R_1699_140b0318 , 
    R_1a5f_124c5618 , 
    R_8fc_13bebd18 , 
    R_961_12fbe358 , 
    R_f1b_13ddafd8 , 
    R_f80_1486f478 , 
    R_153a_116341f8 , 
    R_159f_1008d338 , 
    R_ada_15812f78 , 
    R_da2_156b5ef8 , 
    R_783_123ba898 , 
    R_10f9_123b7a58 , 
    R_13c1_13d3bfb8 , 
    R_1718_156b8018 , 
    R_19e0_13dd4ef8 , 
    R_6cb_117f2258 , 
    R_573_1162dfd8 , 
    R_cea_13d5be18 , 
    R_b92_13c01998 , 
    R_11b1_1700a208 , 
    R_1309_117e8898 , 
    R_17d0_156b8d38 , 
    R_1928_14a0f738 , 
    R_eb1_156b8f18 , 
    R_892_11c69018 , 
    R_9cb_13bed1b8 , 
    R_fea_13d2b3b8 , 
    R_14d0_13ccf698 , 
    R_1609_13cd30b8 , 
    R_67f_13cd88d8 , 
    R_c9e_1580ee78 , 
    R_bde_123b3138 , 
    R_5bf_117f0b38 , 
    R_11fd_1162f3d8 , 
    R_12bd_13bf9698 , 
    R_181c_13bf7758 , 
    R_18dc_15817258 , 
    R_c8c_13b97258 , 
    R_bf0_13c26d38 , 
    R_5d1_14875af8 , 
    R_66d_1700eda8 , 
    R_120f_156b0a98 , 
    R_12ab_1486c278 , 
    R_182e_116366d8 , 
    R_18ca_11c708b8 , 
    R_f2e_13dddb98 , 
    R_90f_13b8e3d8 , 
    R_94e_117f3c98 , 
    R_f6d_13bf7a78 , 
    R_154d_13df8c78 , 
    R_158c_13d278f8 , 
    R_702_13de3598 , 
    R_b5b_13d45bf8 , 
    R_d21_156ac038 , 
    R_117a_14b292d8 , 
    R_1340_123bbab8 , 
    R_1799_13df1018 , 
    R_195f_13b92e38 , 
    R_d38_156afaf8 , 
    R_719_13d1d498 , 
    R_b44_13df7238 , 
    R_1163_13b91358 , 
    R_1357_13d5bcd8 , 
    R_1782_1486c138 , 
    R_1976_14b1de38 , 
    R_695_13b93b58 , 
    R_bc8_13dfb3d8 , 
    R_cb4_15817078 , 
    R_5a9_156b6998 , 
    R_11e7_13bf3298 , 
    R_12d3_14b28338 , 
    R_1806_123b6dd8 , 
    R_18f2_13d40338 , 
    R_a06_158876f8 , 
    R_857_14874dd8 , 
    R_e76_13bf0958 , 
    R_1025_13d59438 , 
    R_1495_14870238 , 
    R_1644_15ff4d88 , 
    R_6fb_156b9378 , 
    R_b62_123bb298 , 
    R_d1a_117ee1f8 , 
    R_1181_148748d8 , 
    R_1339_1580de38 , 
    R_17a0_13dd7478 , 
    R_1958_156ae5b8 , 
    R_97a_117eaff8 , 
    R_f02_13d538f8 , 
    R_8e3_13c107b8 , 
    R_f99_1580efb8 , 
    R_1521_148676d8 , 
    R_15b8_13b93e78 , 
    R_829_13b954f8 , 
    R_a34_156b03b8 , 
    R_e48_15813d38 , 
    R_1053_13cd3478 , 
    R_1467_13b8be58 , 
    R_1672_13cd1df8 , 
    R_e89_13de0078 , 
    R_9f3_156b0598 , 
    R_86a_13b94378 , 
    R_1012_123bf618 , 
    R_14a8_13becdf8 , 
    R_1631_1486c9f8 , 
    R_acd_1008bfd8 , 
    R_daf_123b59d8 , 
    R_790_13d2bd18 , 
    R_10ec_1700b6a8 , 
    R_13ce_13df2a58 , 
    R_170b_14b26178 , 
    R_19ed_148709b8 , 
    R_a31_13cd7d98 , 
    R_82c_140b1e98 , 
    R_e4b_116316d8 , 
    R_1050_13d3d138 , 
    R_146a_123bd318 , 
    R_166f_140ad118 , 
    R_eac_1007f418 , 
    R_88d_13bf99b8 , 
    R_9d0_17010748 , 
    R_fef_1580b138 , 
    R_14cb_13d44258 , 
    R_160e_11632a38 , 
    R_826_13c24cb8 , 
    R_a37_158112b8 , 
    R_e45_15fee168 , 
    R_1056_15fedc68 , 
    R_1464_13d3fa78 , 
    R_1675_14b28dd8 , 
    R_eb6_11c69518 , 
    R_897_11c69338 , 
    R_9c6_156ad258 , 
    R_fe5_14b1f4b8 , 
    R_14d5_14871a98 , 
    R_1604_13beed38 , 
    R_9ef_14a126b8 , 
    R_e8d_13c07578 , 
    R_86e_13ded738 , 
    R_100e_100810d8 , 
    R_14ac_13cce158 , 
    R_162d_13c0adb8 , 
    R_7cb_14a0acd8 , 
    R_dea_123c0798 , 
    R_a92_13d25238 , 
    R_10b1_13d55478 , 
    R_1409_1587f638 , 
    R_16d0_13c02ed8 , 
    R_1a28_14a12398 , 
    R_ee0_13d1ffb8 , 
    R_99c_14a0f418 , 
    R_8c1_14b25818 , 
    R_fbb_123b70f8 , 
    R_14ff_1580bf98 , 
    R_15da_140ba138 , 
    R_687_14b23fb8 , 
    R_bd6_13dd71f8 , 
    R_ca6_123bd098 , 
    R_5b7_117e8cf8 , 
    R_11f5_15815318 , 
    R_12c5_14a0f7d8 , 
    R_1814_170116e8 , 
    R_18e4_12fc1d78 , 
    R_812_12fc0018 , 
    R_a4b_13bf22f8 , 
    R_e31_13bee338 , 
    R_106a_13d56a58 , 
    R_1450_1580a738 , 
    R_1689_14a0c218 , 
    R_e85_156aa878 , 
    R_9f7_13d246f8 , 
    R_866_15ffb868 , 
    R_1016_156af698 , 
    R_14a4_11c6ec98 , 
    R_1635_15ff7588 , 
    R_8ee_140ae338 , 
    R_96f_13d3b8d8 , 
    R_f0d_13d4fa78 , 
    R_f8e_13d541b8 , 
    R_152c_156b2258 , 
    R_15ad_13d58218 , 
    R_9de_124c3458 , 
    R_e9e_123b9038 , 
    R_87f_117f0958 , 
    R_ffd_13c27f58 , 
    R_14bd_13cd71b8 , 
    R_161c_156b6178 , 
    R_aec_14866b98 , 
    R_d90_10081718 , 
    R_771_1007ee78 , 
    R_110b_14b24f58 , 
    R_13af_158110d8 , 
    R_172a_11c6feb8 , 
    R_19ce_11c6fc38 , 
    R_6d4_15ff47e8 , 
    R_56a_17018268 , 
    R_cf3_150e21b8 , 
    R_b89_13cd67b8 , 
    R_11a8_13c0ab38 , 
    R_1312_15881758 , 
    R_17c7_1580cf38 , 
    R_1931_11c6b4f8 , 
    R_7be_13d51918 , 
    R_ddd_10083fb8 , 
    R_a9f_140b7b18 , 
    R_10be_1162c138 , 
    R_13fc_13b967b8 , 
    R_16dd_15ffb728 , 
    R_1a1b_13d3ab18 , 
    R_a2e_1580aeb8 , 
    R_82f_14b26cb8 , 
    R_e4e_13dec798 , 
    R_104d_13de2af8 , 
    R_146d_156b1998 , 
    R_166c_117f5958 , 
    R_d50_156b51d8 , 
    R_b2c_12fc0478 , 
    R_731_15ffaa08 , 
    R_114b_13ddbed8 , 
    R_136f_11c6c718 , 
    R_176a_11628f38 , 
    R_198e_150e3518 , 
    R_ed9_15ff7948 , 
    R_9a3_13c1fad8 , 
    R_8ba_116386b8 , 
    R_fc2_1700f7a8 , 
    R_14f8_117f15d8 , 
    R_15e1_150dcd58 , 
    R_b16_13c1c1f8 , 
    R_d66_13b8b1d8 , 
    R_747_158864d8 , 
    R_1135_156b68f8 , 
    R_1385_1580b278 , 
    R_1754_156add98 , 
    R_19a4_13d4fd98 , 
    R_823_11c6f2d8 , 
    R_a3a_14871318 , 
    R_e42_156ade38 , 
    R_1059_13c0f318 , 
    R_1461_14a1a138 , 
    R_1678_14a0fd78 , 
    R_8d9_158837d8 , 
    R_984_15882d38 , 
    R_ef8_15816998 , 
    R_fa3_15815458 , 
    R_1517_156ad898 , 
    R_15c2_11630c38 , 
    R_af3_13beae18 , 
    R_d89_117e8938 , 
    R_76a_123bceb8 , 
    R_1112_13c20c58 , 
    R_13a8_117f4a58 , 
    R_1731_1008a818 , 
    R_19c7_13d38bd8 , 
    R_b04_156aed38 , 
    R_d78_13cd7758 , 
    R_759_11629938 , 
    R_1123_15ffb908 , 
    R_1397_13d37a58 , 
    R_1742_13d237f8 , 
    R_19b6_14b20778 , 
    R_c64_13c1fdf8 , 
    R_c18_12fc23b8 , 
    R_5f9_13b8f238 , 
    R_645_140b2118 , 
    R_1237_1162dad8 , 
    R_1283_14a18798 , 
    R_1856_117f4878 , 
    R_18a2_13d53998 , 
    R_f2d_100818f8 , 
    R_90e_11629898 , 
    R_94f_15888738 , 
    R_f6e_14a188d8 , 
    R_154c_14a147d8 , 
    R_158d_15ff0a08 , 
    R_9eb_117ef2d8 , 
    R_e91_1580e3d8 , 
    R_872_13c0c7f8 , 
    R_100a_117f81f8 , 
    R_14b0_124c2f58 , 
    R_1629_14a0b6d8 , 
    R_656_15886bb8 , 
    R_c75_156b0db8 , 
    R_c07_124c4cb8 , 
    R_5e8_1162f298 , 
    R_1226_13b8e018 , 
    R_1294_13b91ad8 , 
    R_1845_13cd83d8 , 
    R_18b3_13d1e118 , 
    R_ba0_156b4698 , 
    R_6bd_13c0ec38 , 
    R_581_13d1d8f8 , 
    R_cdc_13cd9378 , 
    R_11bf_123b6c98 , 
    R_12fb_150e3018 , 
    R_17de_14b20458 , 
    R_191a_123b2cd8 , 
    R_d5e_14a10278 , 
    R_b1e_13df7418 , 
    R_73f_1587b998 , 
    R_113d_13d58498 , 
    R_137d_14a11b78 , 
    R_175c_1587b218 , 
    R_199c_17017408 , 
    R_b09_15884f98 , 
    R_d73_1580b4f8 , 
    R_754_15811d58 , 
    R_1128_10084d78 , 
    R_1392_14a15db8 , 
    R_1747_17018588 , 
    R_19b1_13dd9f98 , 
    R_d35_14a11858 , 
    R_716_156b9c38 , 
    R_b47_140af4b8 , 
    R_1166_13ccdcf8 , 
    R_1354_13d41738 , 
    R_1785_1162d218 , 
    R_1973_14a18338 , 
    R_a2b_13c1e6d8 , 
    R_832_13df5c58 , 
    R_e51_156ab278 , 
    R_104a_14a108b8 , 
    R_1470_15887bf8 , 
    R_1669_158828d8 , 
    R_e81_1007dc58 , 
    R_9fb_1486fb58 , 
    R_862_156ab138 , 
    R_101a_13d5a798 , 
    R_14a0_13d38818 , 
    R_1639_1162abf8 , 
    R_ba5_140b4af8 , 
    R_6b8_1580d898 , 
    R_586_15ff8488 , 
    R_cd7_156b7e38 , 
    R_11c4_117ecad8 , 
    R_12f6_17015ba8 , 
    R_17e3_13c1dd78 , 
    R_1915_14a17f78 , 
    R_aff_140aba98 , 
    R_d7d_148714f8 , 
    R_75e_10084418 , 
    R_111e_11635918 , 
    R_139c_1580e0b8 , 
    R_173d_13deffd8 , 
    R_19bb_13df9df8 , 
    R_7dd_13d28898 , 
    R_dfc_156b9ff8 , 
    R_a80_13ddc8d8 , 
    R_109f_13cd2cf8 , 
    R_141b_12fc10f8 , 
    R_16be_13bf0098 , 
    R_1a3a_156b79d8 , 
    R_9d5_15ff1908 , 
    R_ea7_14a124d8 , 
    R_888_13deebd8 , 
    R_ff4_13cd7b18 , 
    R_14c6_13cd5d18 , 
    R_1613_123bc198 , 
    R_677_13c0c758 , 
    R_c96_13c0d838 , 
    R_be6_1162cf98 , 
    R_5c7_1162f1f8 , 
    R_1205_156b94b8 , 
    R_12b5_158816b8 , 
    R_1824_13c04f58 , 
    R_18d4_13beb958 , 
    R_f1a_124c4f38 , 
    R_8fb_13c1e9f8 , 
    R_962_14a15ef8 , 
    R_f81_1580d438 , 
    R_1539_14b267b8 , 
    R_15a0_15ff32a8 , 
    R_d28_156b3fb8 , 
    R_709_117ea4b8 , 
    R_b54_13c04c38 , 
    R_1173_15810778 , 
    R_1347_13dd5f38 , 
    R_1792_13d39858 , 
    R_1966_12fc2098 , 
    R_a1b_123c17d8 , 
    R_842_13bf4738 , 
    R_e61_13cd0958 , 
    R_103a_13ccdbb8 , 
    R_1480_117f1e98 , 
    R_1659_13c1fcb8 , 
    R_820_17013088 , 
    R_a3d_11c6bc78 , 
    R_e3f_123c0e78 , 
    R_105c_13dd87d8 , 
    R_145e_13d5a3d8 , 
    R_167b_14a19878 , 
    R_ebb_13def998 , 
    R_89c_1486e898 , 
    R_9c1_13cd04f8 , 
    R_fe0_15fee7a8 , 
    R_14da_13b95818 , 
    R_15ff_117f1538 , 
    R_8d0_13ccd078 , 
    R_98d_13cceab8 , 
    R_eef_15ff2308 , 
    R_fac_13df65b8 , 
    R_150e_13bed398 , 
    R_15cb_1580a558 , 
    R_663_13c24218 , 
    R_c82_11633bb8 , 
    R_bfa_117f1d58 , 
    R_5db_13c0d798 , 
    R_1219_156b0f98 , 
    R_12a1_15811e98 , 
    R_1838_123c2098 , 
    R_18c0_13ddb258 , 
    R_bbb_13c08dd8 , 
    R_6a2_14870cd8 , 
    R_59c_1700ffc8 , 
    R_cc1_13d5b0f8 , 
    R_11da_14b1dcf8 , 
    R_12e0_14b29c38 , 
    R_17f9_13ddb438 , 
    R_18ff_1162d538 , 
    R_ecc_123bde58 , 
    R_9b0_1587f458 , 
    R_8ad_10082e38 , 
    R_fcf_14a0e798 , 
    R_14eb_140ad258 , 
    R_15ee_117f3158 , 
    R_d13_13c25e38 , 
    R_6f4_156b4918 , 
    R_b69_11c6e8d8 , 
    R_1188_13cd35b8 , 
    R_1332_11637d58 , 
    R_17a7_117f6a38 , 
    R_1951_156b6b78 , 
    R_acf_13d503d8 , 
    R_dad_13cd3838 , 
    R_78e_13b929d8 , 
    R_10ee_1587c438 , 
    R_13cc_1587b3f8 , 
    R_170d_12fbf9d8 , 
    R_19eb_15ff53c8 , 
    R_8c8_12fbe038 , 
    R_ee7_13c03dd8 , 
    R_995_13d50518 , 
    R_fb4_156b0e58 , 
    R_1506_156b9e18 , 
    R_15d3_123b5ed8 , 
    R_b9b_13dfa118 , 
    R_6c2_14b1d618 , 
    R_57c_13d464b8 , 
    R_ce1_13d27358 , 
    R_11ba_13cda458 , 
    R_1300_13dec478 , 
    R_17d9_156af918 , 
    R_191f_14a0d578 , 
    R_7e4_117f6c18 , 
    R_e03_13b8c718 , 
    R_a79_13d52db8 , 
    R_1098_13cd2438 , 
    R_1422_13cd7f78 , 
    R_16b7_14b28518 , 
    R_1a41_150e4d78 , 
    R_ae5_17012048 , 
    R_d97_1162ab58 , 
    R_778_13d52098 , 
    R_1104_13dd7a18 , 
    R_13b6_14a17118 , 
    R_1723_13d50018 , 
    R_19d5_117edc58 , 
    R_d53_13c0ae58 , 
    R_b29_13b95c78 , 
    R_734_14a0f558 , 
    R_1148_117f6218 , 
    R_1372_11c6cd58 , 
    R_1767_11c691f8 , 
    R_1991_13cd58b8 , 
    R_f2c_15814d78 , 
    R_90d_158848b8 , 
    R_950_140b3798 , 
    R_f6f_14a1a318 , 
    R_154b_11632218 , 
    R_158e_14a0b1d8 , 
    R_ec6_13d37b98 , 
    R_8a7_1580e6f8 , 
    R_9b6_14a0cc18 , 
    R_fd5_1580cc18 , 
    R_14e5_13b8fd78 , 
    R_15f4_170165a8 , 
    R_7c0_100854f8 , 
    R_ddf_13b92898 , 
    R_a9d_1162c318 , 
    R_10bc_140b7d98 , 
    R_13fe_13cd60d8 , 
    R_16db_156aaf58 , 
    R_1a1d_13cd9ff8 , 
    R_7f5_13b9a1d8 , 
    R_e14_123bf078 , 
    R_a68_150dbbd8 , 
    R_1087_1587ad18 , 
    R_1433_13dd7978 , 
    R_16a6_13df8458 , 
    R_1a52_11c70778 , 
    R_646_156ad618 , 
    R_c65_10086538 , 
    R_c17_13ccb3b8 , 
    R_5f8_1580f418 , 
    R_1236_1587e558 , 
    R_1284_14a1a458 , 
    R_1855_10084a58 , 
    R_18a3_1700b1a8 , 
    R_69c_156b9058 , 
    R_bc1_13bee298 , 
    R_cbb_13ccbbd8 , 
    R_5a2_15813658 , 
    R_11e0_1587e878 , 
    R_12da_14b29d78 , 
    R_17ff_14a10b38 , 
    R_18f9_14a16718 , 
    R_adc_156ae6f8 , 
    R_da0_13bf5db8 , 
    R_781_13d42f98 , 
    R_10fb_10085778 , 
    R_13bf_123bf6b8 , 
    R_171a_150deb58 , 
    R_19de_117ef918 , 
    R_9e7_13d54578 , 
    R_e95_13d26ef8 , 
    R_876_13d41698 , 
    R_1006_13c08f18 , 
    R_14b4_1700e268 , 
    R_1625_13b96d58 , 
    R_807_13cd8478 , 
    R_e26_1700df48 , 
    R_a56_124c4ad8 , 
    R_1075_15883b98 , 
    R_1445_15880218 , 
    R_1694_13d218b8 , 
    R_1a64_13ccac38 , 
    R_a28_13cd9918 , 
    R_835_140b35b8 , 
    R_e54_14a179d8 , 
    R_1047_14b26df8 , 
    R_1473_156b60d8 , 
    R_1666_14a165d8 , 
    R_b0e_14a15818 , 
    R_d6e_14a0c998 , 
    R_74f_13c24678 , 
    R_112d_1162be18 , 
    R_138d_13b92258 , 
    R_174c_116339d8 , 
    R_19ac_14b1b4f8 , 
    R_bb5_13cd29d8 , 
    R_6a8_1162e618 , 
    R_596_13dd6398 , 
    R_cc7_123b4b78 , 
    R_11d4_15ff30c8 , 
    R_12e6_14a0ff58 , 
    R_17f3_13ddb578 , 
    R_1905_1486dfd8 , 
    R_baa_14a15278 , 
    R_6b3_17011288 , 
    R_58b_140b1c18 , 
    R_cd2_13d24dd8 , 
    R_11c9_14b25278 , 
    R_12f1_1587da18 , 
    R_17e8_1587c078 , 
    R_1910_12fc0978 , 
    R_66e_17014348 , 
    R_c8d_123b7ff8 , 
    R_bef_14a167b8 , 
    R_5d0_13c1db98 , 
    R_120e_13c0d518 , 
    R_12ac_13ccaf58 , 
    R_182d_140b0098 , 
    R_18cb_123b9e98 , 
    R_8b3_13c0d298 , 
    R_ed2_1580c538 , 
    R_9aa_124c51b8 , 
    R_fc9_13b8d118 , 
    R_14f1_150e8978 , 
    R_15e8_15884db8 , 
    R_8e2_13bf6858 , 
    R_97b_150e7a78 , 
    R_f01_14a13e78 , 
    R_f9a_116364f8 , 
    R_1520_1162d678 , 
    R_15b9_13d21a98 , 
    R_7fa_123bbbf8 , 
    R_e19_13d59ed8 , 
    R_a63_14a16678 , 
    R_1082_13c09d78 , 
    R_1438_13bf2398 , 
    R_16a1_14a16cb8 , 
    R_1a57_13c28a98 , 
    R_81d_1580d078 , 
    R_a40_123bcd78 , 
    R_e3c_117f2c58 , 
    R_105f_13de2558 , 
    R_145b_11633e38 , 
    R_167e_1486d858 , 
    R_7f0_13b90458 , 
    R_e0f_140ab138 , 
    R_a6d_117ee838 , 
    R_108c_13bf90f8 , 
    R_142e_11632538 , 
    R_16ab_140b8d38 , 
    R_1a4d_11c70bd8 , 
    R_7d6_14b1e3d8 , 
    R_df5_1580eab8 , 
    R_a87_14a10138 , 
    R_10a6_117efa58 , 
    R_1414_1162b9b8 , 
    R_16c5_14a10db8 , 
    R_1a33_1486ebb8 , 
    R_f0c_140b21b8 , 
    R_8ed_11636d18 , 
    R_970_13c0f818 , 
    R_f8f_11632fd8 , 
    R_152b_13beb778 , 
    R_15ae_123b2eb8 , 
    R_e6b_13b8ded8 , 
    R_a11_158133d8 , 
    R_84c_13bef918 , 
    R_1030_140b72f8 , 
    R_148a_140b0598 , 
    R_164f_13d52778 , 
    R_afa_123c0c98 , 
    R_d82_13cd1858 , 
    R_763_1580e298 , 
    R_1119_1587c118 , 
    R_13a1_158898b8 , 
    R_1738_11c6f878 , 
    R_19c0_1007ded8 , 
    R_e7d_15811538 , 
    R_9ff_13d245b8 , 
    R_85e_13cd3018 , 
    R_101e_13d5d8f8 , 
    R_149c_13d5a978 , 
    R_163d_13ccd438 , 
    R_b8d_156aae18 , 
    R_6d0_1162bb98 , 
    R_56e_10086e98 , 
    R_cef_14870eb8 , 
    R_11ac_13c24498 , 
    R_130e_14a17758 , 
    R_17cb_14a0e478 , 
    R_192d_123becb8 , 
    R_d32_13d20558 , 
    R_713_15882978 , 
    R_b4a_13d22cb8 , 
    R_1169_123b7c38 , 
    R_1351_14a14558 , 
    R_1788_13ccae18 , 
    R_1970_124c43f8 , 
    R_7cd_13d58df8 , 
    R_dec_156ae518 , 
    R_a90_13dd8058 , 
    R_10af_117f0818 , 
    R_140b_1580d1b8 , 
    R_16ce_117ebe58 , 
    R_1a2a_15810e58 , 
    R_e72_13c1e8b8 , 
    R_a0a_13d54438 , 
    R_853_123bd778 , 
    R_1029_13cd2898 , 
    R_1491_117f33d8 , 
    R_1648_15ff12c8 , 
    R_80f_13d449d8 , 
    R_a4e_13b8e798 , 
    R_e2e_13dd57b8 , 
    R_106d_13b8b598 , 
    R_144d_13cd65d8 , 
    R_168c_15ff1c28;
wire n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
     n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
     n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
     n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
     n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
     n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
     n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
     n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
     n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
     n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
     n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
     n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
     n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
     n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
     n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
     n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
     n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
     n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
     n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
     n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
     n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
     n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
     n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
     n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
     n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
     n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
     n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
     n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
     n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
     n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
     n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
     n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
     n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
     n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
     n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
     n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
     n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
     n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
     n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
     n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
     n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
     n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
     n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
     n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
     n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
     n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
     n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
     n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
     n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
     n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
     n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
     n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
     n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
     n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
     n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
     n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
     n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
     n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
     n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
     n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
     n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
     n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
     n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
     n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
     n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
     n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
     n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
     n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
     n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
     n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
     n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
     n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
     n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
     n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
     n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
     n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
     n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
     n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
     n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
     n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
     n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
     n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
     n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
     n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
     n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
     n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
     n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
     n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
     n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
     n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
     n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
     n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
     n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
     n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
     n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
     n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
     n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
     n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
     n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
     n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
     n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
     n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
     n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
     n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
     n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
     n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
     n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
     n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
     n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
     n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
     n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
     n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
     n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
     n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
     n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
     n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
     n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
     n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
     n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , 
     n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , 
     n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , 
     n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , 
     n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , 
     n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , 
     n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
     n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , 
     n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , 
     n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , 
     n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , 
     n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , 
     n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , 
     n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , 
     n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , 
     n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , 
     n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , 
     n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , 
     n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , 
     n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , 
     n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
     n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
     n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
     n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , 
     n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , 
     n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , 
     n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , 
     n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , 
     n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , 
     n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , 
     n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , 
     n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , 
     n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , 
     n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
     n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , 
     n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , 
     n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , 
     n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , 
     n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , 
     n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , 
     n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , 
     n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , 
     n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , 
     n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , 
     n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , 
     n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , 
     n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , 
     n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , 
     n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , 
     n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , 
     n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , 
     n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , 
     n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , 
     n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , 
     n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , 
     n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , 
     n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , 
     n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , 
     n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , 
     n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , 
     n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , 
     n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , 
     n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , 
     n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , 
     n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , 
     n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , 
     n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , 
     n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , 
     n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , 
     n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , 
     n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , 
     n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , 
     n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , 
     n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , 
     n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , 
     n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , 
     n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , 
     n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , 
     n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , 
     n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , 
     n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , 
     n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , 
     n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , 
     n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , 
     n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , 
     n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , 
     n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , 
     n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , 
     n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , 
     n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , 
     n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , 
     n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , 
     n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , 
     n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , 
     n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , 
     n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , 
     n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , 
     n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , 
     n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , 
     n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , 
     n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , 
     n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , 
     n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , 
     n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , 
     n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , 
     n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , 
     n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , 
     n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , 
     n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , 
     n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , 
     n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , 
     n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , 
     n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , 
     n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , 
     n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , 
     n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , 
     n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , 
     n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , 
     n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , 
     n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , 
     n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , 
     n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , 
     n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , 
     n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , 
     n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , 
     n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , 
     n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , 
     n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , 
     n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , 
     n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , 
     n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , 
     n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , 
     n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , 
     n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , 
     n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , 
     n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , 
     n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , 
     n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , 
     n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , 
     n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , 
     n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , 
     n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , 
     n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , 
     n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , 
     n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , 
     n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , 
     n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , 
     n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , 
     n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , 
     n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , 
     n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , 
     n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , 
     n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , 
     n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , 
     n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , 
     n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , 
     n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , 
     n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , 
     n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , 
     n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , 
     n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , 
     n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , 
     n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , 
     n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , 
     n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , 
     n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , 
     n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , 
     n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , 
     n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , 
     n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , 
     n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , 
     n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , 
     n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , 
     n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , 
     n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , 
     n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , 
     n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , 
     n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , 
     n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , 
     n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , 
     n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , 
     n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , 
     n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , 
     n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , 
     n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , 
     n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , 
     n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , 
     n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , 
     n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , 
     n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , 
     n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , 
     n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , 
     n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , 
     n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , 
     n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , 
     n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , 
     n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , 
     n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , 
     n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , 
     n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , 
     n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , 
     n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , 
     n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , 
     n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , 
     n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , 
     n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , 
     n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , 
     n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , 
     n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , 
     n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , 
     n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , 
     n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , 
     n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , 
     n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , 
     n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , 
     n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , 
     n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , 
     n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , 
     n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , 
     n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , 
     n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , 
     n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , 
     n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , 
     n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , 
     n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , 
     n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , 
     n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , 
     n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , 
     n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , 
     n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , 
     n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , 
     n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , 
     n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , 
     n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , 
     n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , 
     n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , 
     n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , 
     n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , 
     n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , 
     n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , 
     n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , 
     n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , 
     n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , 
     n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , 
     n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , 
     n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , 
     n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , 
     n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , 
     n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , 
     n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , 
     n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , 
     n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , 
     n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , 
     n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , 
     n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , 
     n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , 
     n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , 
     n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , 
     n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , 
     n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , 
     n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , 
     n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , 
     n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , 
     n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , 
     n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , 
     n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , 
     n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , 
     n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , 
     n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , 
     n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , 
     n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , 
     n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , 
     n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , 
     n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , 
     n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , 
     n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , 
     n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , 
     n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , 
     n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , 
     n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , 
     n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , 
     n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , 
     n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , 
     n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , 
     n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , 
     n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , 
     n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , 
     n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , 
     n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , 
     n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , 
     n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , 
     n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , 
     n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , 
     n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , 
     n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , 
     n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , 
     n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , 
     n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , 
     n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , 
     n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , 
     n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , 
     n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , 
     n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , 
     n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , 
     n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , 
     n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , 
     n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , 
     n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , 
     n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , 
     n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , 
     n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , 
     n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , 
     n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , 
     n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , 
     n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , 
     n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , 
     n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , 
     n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , 
     n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , 
     n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , 
     n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , 
     n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , 
     n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , 
     n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , 
     n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , 
     n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , 
     n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , 
     n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , 
     n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , 
     n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , 
     n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , 
     n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , 
     n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , 
     n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , 
     n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , 
     n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , 
     n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , 
     n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , 
     n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , 
     n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
     n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , 
     n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , 
     n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , 
     n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , 
     n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , 
     n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , 
     n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , 
     n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
     n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
     n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , 
     n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , 
     n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , 
     n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , 
     n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , 
     n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , 
     n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , 
     n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , 
     n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , 
     n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , 
     n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , 
     n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , 
     n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , 
     n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , 
     n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , 
     n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , 
     n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , 
     n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , 
     n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , 
     n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , 
     n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , 
     n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , 
     n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , 
     n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , 
     n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , 
     n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , 
     n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , 
     n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , 
     n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , 
     n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , 
     n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , 
     n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , 
     n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , 
     n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , 
     n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , 
     n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , 
     n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , 
     n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , 
     n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , 
     n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , 
     n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , 
     n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , 
     n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , 
     n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , 
     n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , 
     n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , 
     n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , 
     n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , 
     n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , 
     n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , 
     n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , 
     n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , 
     n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , 
     n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , 
     n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , 
     n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , 
     n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , 
     n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , 
     n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , 
     n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , 
     n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , 
     n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , 
     n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , 
     n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , 
     n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , 
     n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , 
     n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , 
     n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , 
     n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , 
     n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , 
     n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , 
     n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , 
     n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , 
     n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , 
     n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , 
     n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , 
     n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , 
     n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , 
     n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , 
     n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , 
     n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , 
     n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , 
     n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , 
     n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , 
     n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , 
     n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , 
     n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , 
     n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , 
     n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , 
     n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , 
     n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , 
     n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , 
     n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , 
     n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , 
     n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , 
     n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , 
     n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , 
     n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , 
     n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , 
     n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , 
     n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , 
     n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , 
     n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , 
     n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , 
     n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , 
     n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , 
     n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , 
     n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , 
     n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , 
     n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , 
     n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , 
     n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , 
     n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , 
     n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , 
     n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , 
     n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , 
     n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , 
     n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , 
     n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , 
     n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , 
     n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , 
     n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , 
     n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , 
     n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , 
     n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , 
     n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , 
     n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , 
     n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , 
     n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , 
     n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , 
     n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , 
     n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , 
     n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , 
     n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , 
     n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , 
     n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , 
     n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , 
     n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , 
     n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , 
     n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , 
     n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , 
     n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , 
     n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , 
     n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , 
     n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , 
     n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , 
     n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , 
     n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , 
     n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , 
     n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , 
     n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , 
     n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , 
     n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , 
     n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , 
     n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , 
     n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , 
     n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , 
     n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , 
     n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , 
     n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , 
     n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , 
     n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , 
     n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , 
     n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , 
     n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , 
     n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , 
     n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , 
     n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , 
     n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , 
     n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , 
     n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , 
     n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , 
     n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , 
     n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , 
     n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , 
     n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , 
     n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , 
     n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , 
     n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , 
     n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , 
     n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , 
     n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , 
     n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , 
     n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , 
     n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , 
     n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , 
     n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , 
     n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , 
     n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , 
     n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , 
     n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , 
     n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , 
     n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , 
     n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , 
     n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , 
     n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , 
     n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , 
     n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , 
     n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , 
     n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , 
     n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , 
     n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , 
     n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , 
     n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , 
     n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , 
     n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , 
     n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , 
     n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , 
     n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , 
     n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , 
     n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , 
     n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , 
     n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , 
     n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , 
     n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , 
     n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , 
     n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , 
     n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , 
     n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , 
     n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , 
     n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , 
     n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , 
     n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , 
     n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , 
     n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , 
     n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , 
     n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , 
     n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , 
     n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , 
     n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , 
     n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , 
     n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , 
     n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , 
     n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , 
     n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , 
     n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , 
     n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , 
     n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , 
     n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , 
     n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , 
     n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , 
     n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , 
     n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , 
     n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , 
     n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , 
     n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , 
     n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , 
     n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , 
     n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , 
     n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
     n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , 
     n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , 
     n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , 
     n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , 
     n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , 
     n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , 
     n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , 
     n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , 
     n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , 
     n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , 
     n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , 
     n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , 
     n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , 
     n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , 
     n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , 
     n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , 
     n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , 
     n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , 
     n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , 
     n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , 
     n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , 
     n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , 
     n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , 
     n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , 
     n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , 
     n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , 
     n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , 
     n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , 
     n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , 
     n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , 
     n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , 
     n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , 
     n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , 
     n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , 
     n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , 
     n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , 
     n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , 
     n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , 
     n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , 
     n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , 
     n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , 
     n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , 
     n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , 
     n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , 
     n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , 
     n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , 
     n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , 
     n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , 
     n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , 
     n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , 
     n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , 
     n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , 
     n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , 
     n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , 
     n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , 
     n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , 
     n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , 
     n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , 
     n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , 
     n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , 
     n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , 
     n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , 
     n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , 
     n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , 
     n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , 
     n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , 
     n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , 
     n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , 
     n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , 
     n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , 
     n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , 
     n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , 
     n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , 
     n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , 
     n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , 
     n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , 
     n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , 
     n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , 
     n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , 
     n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , 
     n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , 
     n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , 
     n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , 
     n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , 
     n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , 
     n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , 
     n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , 
     n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , 
     n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , 
     n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , 
     n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , 
     n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , 
     n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , 
     n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , 
     n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , 
     n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , 
     n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , 
     n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , 
     n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , 
     n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , 
     n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , 
     n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , 
     n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , 
     n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , 
     n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , 
     n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , 
     n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , 
     n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , 
     n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , 
     n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , 
     n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , 
     n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , 
     n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , 
     n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , 
     n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , 
     n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , 
     n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , 
     n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , 
     n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , 
     n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , 
     n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , 
     n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , 
     n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , 
     n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , 
     n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , 
     n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , 
     n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , 
     n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , 
     n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , 
     n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , 
     n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , 
     n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , 
     n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , 
     n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , 
     n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , 
     n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , 
     n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , 
     n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , 
     n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , 
     n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , 
     n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , 
     n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , 
     n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , 
     n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , 
     n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , 
     n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , 
     n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , 
     n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , 
     n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , 
     n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , 
     n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , 
     n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , 
     n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , 
     n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , 
     n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , 
     n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , 
     n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , 
     n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , 
     n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , 
     n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , 
     n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , 
     n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , 
     n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , 
     n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , 
     n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , 
     n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , 
     n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , 
     n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , 
     n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , 
     n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , 
     n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , 
     n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , 
     n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , 
     n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , 
     n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , 
     n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , 
     n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , 
     n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , 
     n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , 
     n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , 
     n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , 
     n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , 
     n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , 
     n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , 
     n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , 
     n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , 
     n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , 
     n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , 
     n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , 
     n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , 
     n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , 
     n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , 
     n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , 
     n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , 
     n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , 
     n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , 
     n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , 
     n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , 
     n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , 
     n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , 
     n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , 
     n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , 
     n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , 
     n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , 
     n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , 
     n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , 
     n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , 
     n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , 
     n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , 
     n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , 
     n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , 
     n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , 
     n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , 
     n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , 
     n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , 
     n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , 
     n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , 
     n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , 
     n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , 
     n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , 
     n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , 
     n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , 
     n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , 
     n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , 
     n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , 
     n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , 
     n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , 
     n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , 
     n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , 
     n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , 
     n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , 
     n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , 
     n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , 
     n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , 
     n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , 
     n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , 
     n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , 
     n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , 
     n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , 
     n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , 
     n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , 
     n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , 
     n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , 
     n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , 
     n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , 
     n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , 
     n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , 
     n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , 
     n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , 
     n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , 
     n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , 
     n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , 
     n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , 
     n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , 
     n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , 
     n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , 
     n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , 
     n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , 
     n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , 
     n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , 
     n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , 
     n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , 
     n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , 
     n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , 
     n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , 
     n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , 
     n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , 
     n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , 
     n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , 
     n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , 
     n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , 
     n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , 
     n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , 
     n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , 
     n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , 
     n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , 
     n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , 
     n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , 
     n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , 
     n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , 
     n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , 
     n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , 
     n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , 
     n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , 
     n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , 
     n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , 
     n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , 
     n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , 
     n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , 
     n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , 
     n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , 
     n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , 
     n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , 
     n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , 
     n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , 
     n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , 
     n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , 
     n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , 
     n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , 
     n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , 
     n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , 
     n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , 
     n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , 
     n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , 
     n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , 
     n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , 
     n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , 
     n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , 
     n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , 
     n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , 
     n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , 
     n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , 
     n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , 
     n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , 
     n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , 
     n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , 
     n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , 
     n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , 
     n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , 
     n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , 
     n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , 
     n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , 
     n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , 
     n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , 
     n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , 
     n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , 
     n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , 
     n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , 
     n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , 
     n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , 
     n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , 
     n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , 
     n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , 
     n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , 
     n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , 
     n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , 
     n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , 
     n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , 
     n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , 
     n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , 
     n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , 
     n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , 
     n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , 
     n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , 
     n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , 
     n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , 
     n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , 
     n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , 
     n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , 
     n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , 
     n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , 
     n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , 
     n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , 
     n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , 
     n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , 
     n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , 
     n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , 
     n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , 
     n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , 
     n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , 
     n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , 
     n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , 
     n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , 
     n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , 
     n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , 
     n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , 
     n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , 
     n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , 
     n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , 
     n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , 
     n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , 
     n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , 
     n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , 
     n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , 
     n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , 
     n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , 
     n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , 
     n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , 
     n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , 
     n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , 
     n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , 
     n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , 
     n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , 
     n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , 
     n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , 
     n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , 
     n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , 
     n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , 
     n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , 
     n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , 
     n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , 
     n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , 
     n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , 
     n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , 
     n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , 
     n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , 
     n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , 
     n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , 
     n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , 
     n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , 
     n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , 
     n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , 
     n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , 
     n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , 
     n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , 
     n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , 
     n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , 
     n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , 
     n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , 
     n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , 
     n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , 
     n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , 
     n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , 
     n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , 
     n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , 
     n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , 
     n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , 
     n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , 
     n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , 
     n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , 
     n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , 
     n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , 
     n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , 
     n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , 
     n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , 
     n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , 
     n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , 
     n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , 
     n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , 
     n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , 
     n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , 
     n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , 
     n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , 
     n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , 
     n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , 
     n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , 
     n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , 
     n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , 
     n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , 
     n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , 
     n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , 
     n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , 
     n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , 
     n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , 
     n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , 
     n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , 
     n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , 
     n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , 
     n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , 
     n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , 
     n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , 
     n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , 
     n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , 
     n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , 
     n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , 
     n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , 
     n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , 
     n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , 
     n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , 
     n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , 
     n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , 
     n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , 
     n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , 
     n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , 
     n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , 
     n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , 
     n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , 
     n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , 
     n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , 
     n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , 
     n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , 
     n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , 
     n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , 
     n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , 
     n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , 
     n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , 
     n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , 
     n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , 
     n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , 
     n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , 
     n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , 
     n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , 
     n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , 
     n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , 
     n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , 
     n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , 
     n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , 
     n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , 
     n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , 
     n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , 
     n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , 
     n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , 
     n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , 
     n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , 
     n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , 
     n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , 
     n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , 
     n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , 
     n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , 
     n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , 
     n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , 
     n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , 
     n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , 
     n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , 
     n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , 
     n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , 
     n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , 
     n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , 
     n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , 
     n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , 
     n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , 
     n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , 
     n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , 
     n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , 
     n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , 
     n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , 
     n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , 
     n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , 
     n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , 
     n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , 
     n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , 
     n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , 
     n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , 
     n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , 
     n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , 
     n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , 
     n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , 
     n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , 
     n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , 
     n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , 
     n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , 
     n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , 
     n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , 
     n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , 
     n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , 
     n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , 
     n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , 
     n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , 
     n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , 
     n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , 
     n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , 
     n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , 
     n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , 
     n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , 
     n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , 
     n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , 
     n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , 
     n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , 
     n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , 
     n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , 
     n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , 
     n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , 
     n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , 
     n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , 
     n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , 
     n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , 
     n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , 
     n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , 
     n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , 
     n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , 
     n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , 
     n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , 
     n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , 
     n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , 
     n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , 
     n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , 
     n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , 
     n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , 
     n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , 
     n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , 
     n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , 
     n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , 
     n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , 
     n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , 
     n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , 
     n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , 
     n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , 
     n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , 
     n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , 
     n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , 
     n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , 
     n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , 
     n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , 
     n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , 
     n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , 
     n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , 
     n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , 
     n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , 
     n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , 
     n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , 
     n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , 
     n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , 
     n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , 
     n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , 
     n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , 
     n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , 
     n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , 
     n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , 
     n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , 
     n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , 
     n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , 
     n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , 
     n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , 
     n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , 
     n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , 
     n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , 
     n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , 
     n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , 
     n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , 
     n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , 
     n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , 
     n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , 
     n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , 
     n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , 
     n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , 
     n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , 
     n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , 
     n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , 
     n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , 
     n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , 
     n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , 
     n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , 
     n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , 
     n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , 
     n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , 
     n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , 
     n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , 
     n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , 
     n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , 
     n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , 
     n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , 
     n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , 
     n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , 
     n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , 
     n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , 
     n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , 
     n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , 
     n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , 
     n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , 
     n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , 
     n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , 
     n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , 
     n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , 
     n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , 
     n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , 
     n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , 
     n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , 
     n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , 
     n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , 
     n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , 
     n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , 
     n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , 
     n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , 
     n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , 
     n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , 
     n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , 
     n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , 
     n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , 
     n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , 
     n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , 
     n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , 
     n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , 
     n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , 
     n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , 
     n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , 
     n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , 
     n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , 
     n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , 
     n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , 
     n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , 
     n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , 
     n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , 
     n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , 
     n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , 
     n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , 
     n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , 
     n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , 
     n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , 
     n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , 
     n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , 
     n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , 
     n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , 
     n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , 
     n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , 
     n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , 
     n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , 
     n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , 
     n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , 
     n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , 
     n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , 
     n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , 
     n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , 
     n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , 
     n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , 
     n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , 
     n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , 
     n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , 
     n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , 
     n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , 
     n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , 
     n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , 
     n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , 
     n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , 
     n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , 
     n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , 
     n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , 
     n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , 
     n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , 
     n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , 
     n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , 
     n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , 
     n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , 
     n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , 
     n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , 
     n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , 
     n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , 
     n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , 
     n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , 
     n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , 
     n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , 
     n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , 
     n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , 
     n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , 
     n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , 
     n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , 
     n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , 
     n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , 
     n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , 
     n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , 
     n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , 
     n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , 
     n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , 
     n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , 
     n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , 
     n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , 
     n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , 
     n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , 
     n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , 
     n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , 
     n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , 
     n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , 
     n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , 
     n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , 
     n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , 
     n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , 
     n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , 
     n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , 
     n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , 
     n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , 
     n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , 
     n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , 
     n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , 
     n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , 
     n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , 
     n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , 
     n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , 
     n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , 
     n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , 
     n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , 
     n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , 
     n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , 
     n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , 
     n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , 
     n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , 
     n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , 
     n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , 
     n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , 
     n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , 
     n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , 
     n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , 
     n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , 
     n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , 
     n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , 
     n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , 
     n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , 
     n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , 
     n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , 
     n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , 
     n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , 
     n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , 
     n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , 
     n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , 
     n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , 
     n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , 
     n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , 
     n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , 
     n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , 
     n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , 
     n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , 
     n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , 
     n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , 
     n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , 
     n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , 
     n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , 
     n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , 
     n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , 
     n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , 
     n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , 
     n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , 
     n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , 
     n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , 
     n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , 
     n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , 
     n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , 
     n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , 
     n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , 
     n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , 
     n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , 
     n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , 
     n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , 
     n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , 
     n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , 
     n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , 
     n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , 
     n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , 
     n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , 
     n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , 
     n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , 
     n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , 
     n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , 
     n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , 
     n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , 
     n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , 
     n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , 
     n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , 
     n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , 
     n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , 
     n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , 
     n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , 
     n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , 
     n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , 
     n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , 
     n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , 
     n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , 
     n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , 
     n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , 
     n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , 
     n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , 
     n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , 
     n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , 
     n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , 
     n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , 
     n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , 
     n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , 
     n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , 
     n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , 
     n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , 
     n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , 
     n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , 
     n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , 
     n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , 
     n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , 
     n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , 
     n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , 
     n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , 
     n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , 
     n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , 
     n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , 
     n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , 
     n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , 
     n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , 
     n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , 
     n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , 
     n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , 
     n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , 
     n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , 
     n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , 
     n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , 
     n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , 
     n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , 
     n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , 
     n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , 
     n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , 
     n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , 
     n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , 
     n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , 
     n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , 
     n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , 
     n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , 
     n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , 
     n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , 
     n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , 
     n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , 
     n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , 
     n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , 
     n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , 
     n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , 
     n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , 
     n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , 
     n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , 
     n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , 
     n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , 
     n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , 
     n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , 
     n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , 
     n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , 
     n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , 
     n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , 
     n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , 
     n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , 
     n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , 
     n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , 
     n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , 
     n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , 
     n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , 
     n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , 
     n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , 
     n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , 
     n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , 
     n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , 
     n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , 
     n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , 
     n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , 
     n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , 
     n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , 
     n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , 
     n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , 
     n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , 
     n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , 
     n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , 
     n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , 
     n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , 
     n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , 
     n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , 
     n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , 
     n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , 
     n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , 
     n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , 
     n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , 
     n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , 
     n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , 
     n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , 
     n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , 
     n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , 
     n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , 
     n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , 
     n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , 
     n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , 
     n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , 
     n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , 
     n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , 
     n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , 
     n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , 
     n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , 
     n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , 
     n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , 
     n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , 
     n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , 
     n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , 
     n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , 
     n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , 
     n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , 
     n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , 
     n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , 
     n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , 
     n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , 
     n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , 
     n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , 
     n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , 
     n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , 
     n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , 
     n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , 
     n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , 
     n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , 
     n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , 
     n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , 
     n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , 
     n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , 
     n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , 
     n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , 
     n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , 
     n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , 
     n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , 
     n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , 
     n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , 
     n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , 
     n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , 
     n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , 
     n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , 
     n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , 
     n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , 
     n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , 
     n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , 
     n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , 
     n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , 
     n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , 
     n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , 
     n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , 
     n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , 
     n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , 
     n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , 
     n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , 
     n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , 
     n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , 
     n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , 
     n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , 
     n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , 
     n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , 
     n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , 
     n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , 
     n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , 
     n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , 
     n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , 
     n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , 
     n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , 
     n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , 
     n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , 
     n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , 
     n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , 
     n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , 
     n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , 
     n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , 
     n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , 
     n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , 
     n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , 
     n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , 
     n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , 
     n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , 
     n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , 
     n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , 
     n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , 
     n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , 
     n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , 
     n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , 
     n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , 
     n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , 
     n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , 
     n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , 
     n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , 
     n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , 
     n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , 
     n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , 
     n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , 
     n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , 
     n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , 
     n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , 
     n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , 
     n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , 
     n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , 
     n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , 
     n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , 
     n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , 
     n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , 
     n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , 
     n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , 
     n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , 
     n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , 
     n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , 
     n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , 
     n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , 
     n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , 
     n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , 
     n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , 
     n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , 
     n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , 
     n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , 
     n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , 
     n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , 
     n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , 
     n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , 
     n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , 
     n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , 
     n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , 
     n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , 
     n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , 
     n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , 
     n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , 
     n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , 
     n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , 
     n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , 
     n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , 
     n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , 
     n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , 
     n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , 
     n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , 
     n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , 
     n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , 
     n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , 
     n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , 
     n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , 
     n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , 
     n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , 
     n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , 
     n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , 
     n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , 
     n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , 
     n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , 
     n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , 
     n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , 
     n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , 
     n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , 
     n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , 
     n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , 
     n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , 
     n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , 
     n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , 
     n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , 
     n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , 
     n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , 
     n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , 
     n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , 
     n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , 
     n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , 
     n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , 
     n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , 
     n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , 
     n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , 
     n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , 
     n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , 
     n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , 
     n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , 
     n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , 
     n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , 
     n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , 
     n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , 
     n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , 
     n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , 
     n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , 
     n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , 
     n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , 
     n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , 
     n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , 
     n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , 
     n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , 
     n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , 
     n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , 
     n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , 
     n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , 
     n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , 
     n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , 
     n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , 
     n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , 
     n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , 
     n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , 
     n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , 
     n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , 
     n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , 
     n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , 
     n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , 
     n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , 
     n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , 
     n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , 
     n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , 
     n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , 
     n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , 
     n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , 
     n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , 
     n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , 
     n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , 
     n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , 
     n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , 
     n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , 
     n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , 
     n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , 
     n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , 
     n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , 
     n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , 
     n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , 
     n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , 
     n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , 
     n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , 
     n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , 
     n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , 
     n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , 
     n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , 
     n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , 
     n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , 
     n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , 
     n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , 
     n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , 
     n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , 
     n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , 
     n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , 
     n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , 
     n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , 
     n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , 
     n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , 
     n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , 
     n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , 
     n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , 
     n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , 
     n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , 
     n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , 
     n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , 
     n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , 
     n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , 
     n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , 
     n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , 
     n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , 
     n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , 
     n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , 
     n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , 
     n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , 
     n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , 
     n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , 
     n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , 
     n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , 
     n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , 
     n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , 
     n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , 
     n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , 
     n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , 
     n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , 
     n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , 
     n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , 
     n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , 
     n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , 
     n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , 
     n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , 
     n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , 
     n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , 
     n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , 
     n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , 
     n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , 
     n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , 
     n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , 
     n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , 
     n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , 
     n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , 
     n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , 
     n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , 
     n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , 
     n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , 
     n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , 
     n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , 
     n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , 
     n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , 
     n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , 
     n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , 
     n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , 
     n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , 
     n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , 
     n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , 
     n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , 
     n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , 
     n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , 
     n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , 
     n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , 
     n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , 
     n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , 
     n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , 
     n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , 
     n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , 
     n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , 
     n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , 
     n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , 
     n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , 
     n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , 
     n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , 
     n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , 
     n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , 
     n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , 
     n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , 
     n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , 
     n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , 
     n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , 
     n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , 
     n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , 
     n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , 
     n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , 
     n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , 
     n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , 
     n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , 
     n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , 
     n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , 
     n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , 
     n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , 
     n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , 
     n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , 
     n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , 
     n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , 
     n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , 
     n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , 
     n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , 
     n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , 
     n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , 
     n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , 
     n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , 
     n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , 
     n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , 
     n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , 
     n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , 
     n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , 
     n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , 
     n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , 
     n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , 
     n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , 
     n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , 
     n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , 
     n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , 
     n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , 
     n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , 
     n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , 
     n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , 
     n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , 
     n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , 
     n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , 
     n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , 
     n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , 
     n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , 
     n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , 
     n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , 
     n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , 
     n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , 
     n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , 
     n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , 
     n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , 
     n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , 
     n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , 
     n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , 
     n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , 
     n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , 
     n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , 
     n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , 
     n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , 
     n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , 
     n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , 
     n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , 
     n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , 
     n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , 
     n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , 
     n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , 
     n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , 
     n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , 
     n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , 
     n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , 
     n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , 
     n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , 
     n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , 
     n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , 
     n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , 
     n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , 
     n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , 
     n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , 
     n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , 
     n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , 
     n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , 
     n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , 
     n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , 
     n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , 
     n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , 
     n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , 
     n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , 
     n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , 
     n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , 
     n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , 
     n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , 
     n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , 
     n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , 
     n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , 
     n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , 
     n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , 
     n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , 
     n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , 
     n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , 
     n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , 
     n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , 
     n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , 
     n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , 
     n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , 
     n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , 
     n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , 
     n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , 
     n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , 
     n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , 
     n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , 
     n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , 
     n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , 
     n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , 
     n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , 
     n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , 
     n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , 
     n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , 
     n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , 
     n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , 
     n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , 
     n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , 
     n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , 
     n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , 
     n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , 
     n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , 
     n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , 
     n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , 
     n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , 
     n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , 
     n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , 
     n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , 
     n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , 
     n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , 
     n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , 
     n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , 
     n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , 
     n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , 
     n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , 
     n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , 
     n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , 
     n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , 
     n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , 
     n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , 
     n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , 
     n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , 
     n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , 
     n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , 
     n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , 
     n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , 
     n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , 
     n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , 
     n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , 
     n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , 
     n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , 
     n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , 
     n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , 
     n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , 
     n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , 
     n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , 
     n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , 
     n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , 
     n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , 
     n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , 
     n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , 
     n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , 
     n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , 
     n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , 
     n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , 
     n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , 
     n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , 
     n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , 
     n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , 
     n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , 
     n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , 
     n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , 
     n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , 
     n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , 
     n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , 
     n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , 
     n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , 
     n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , 
     n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , 
     n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , 
     n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , 
     n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , 
     n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , 
     n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , 
     n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , 
     n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , 
     n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , 
     n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , 
     n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , 
     n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , 
     n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , 
     n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , 
     n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , 
     n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , 
     n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , 
     n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , 
     n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , 
     n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , 
     n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , 
     n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , 
     n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , 
     n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , 
     n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , 
     n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , 
     n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , 
     n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , 
     n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , 
     n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , 
     n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , 
     n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , 
     n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , 
     n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , 
     n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , 
     n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , 
     n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , 
     n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , 
     n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , 
     n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , 
     n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , 
     n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , 
     n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , 
     n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , 
     n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , 
     n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , 
     n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , 
     n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , 
     n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , 
     n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , 
     n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , 
     n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , 
     n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , 
     n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , 
     n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , 
     n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , 
     n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , 
     n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , 
     n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , 
     n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , 
     n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , 
     n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , 
     n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , 
     n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , 
     n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , 
     n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , 
     n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , 
     n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , 
     n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , 
     n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , 
     n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , 
     n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , 
     n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , 
     n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , 
     n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , 
     n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , 
     n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , 
     n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , 
     n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , 
     n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , 
     n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , 
     n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , 
     n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , 
     n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , 
     n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , 
     n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , 
     n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , 
     n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , 
     n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , 
     n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , 
     n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , 
     n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , 
     n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , 
     n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , 
     n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , 
     n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , 
     n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , 
     n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , 
     n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , 
     n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , 
     n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , 
     n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , 
     n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , 
     n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , 
     n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , 
     n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , 
     n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , 
     n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , 
     n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , 
     n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , 
     n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , 
     n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , 
     n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , 
     n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , 
     n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , 
     n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , 
     n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , 
     n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , 
     n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , 
     n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , 
     n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , 
     n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , 
     n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , 
     n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , 
     n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , 
     n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , 
     n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , 
     n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , 
     n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , 
     n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , 
     n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , 
     n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , 
     n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , 
     n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , 
     n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , 
     n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , 
     n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , 
     n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , 
     n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , 
     n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , 
     n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , 
     n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , 
     n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , 
     n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , 
     n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , 
     n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , 
     n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , 
     n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , 
     n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , 
     n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , 
     n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , 
     n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , 
     n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , 
     n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , 
     n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , 
     n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , 
     n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , 
     n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , 
     n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , 
     n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , 
     n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , 
     n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , 
     n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , 
     n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , 
     n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , 
     n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , 
     n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , 
     n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , 
     n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , 
     n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , 
     n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , 
     n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , 
     n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , 
     n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , 
     n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , 
     n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , 
     n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , 
     n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , 
     n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , 
     n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , 
     n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , 
     n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , 
     n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , 
     n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , 
     n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , 
     n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , 
     n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , 
     n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , 
     n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , 
     n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , 
     n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , 
     n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , 
     n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , 
     n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , 
     n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , 
     n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , 
     n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , 
     n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , 
     n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , 
     n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , 
     n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , 
     n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , 
     n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , 
     n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , 
     n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , 
     n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , 
     n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , 
     n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , 
     n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , 
     n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , 
     n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , 
     n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , 
     n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , 
     n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , 
     n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , 
     n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , 
     n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , 
     n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , 
     n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , 
     n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , 
     n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , 
     n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , 
     n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , 
     n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , 
     n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , 
     n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , 
     n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , 
     n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , 
     n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , 
     n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , 
     n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , 
     n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , 
     n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , 
     n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , 
     n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , 
     n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , 
     n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , 
     n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , 
     n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , 
     n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , 
     n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , 
     n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , 
     n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , 
     n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , 
     n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , 
     n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , 
     n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , 
     n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , 
     n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , 
     n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , 
     n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , 
     n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , 
     n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , 
     n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , 
     n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , 
     n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , 
     n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , 
     n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , 
     n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , 
     n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , 
     n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , 
     n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , 
     n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , 
     n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , 
     n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , 
     n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , 
     n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , 
     n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , 
     n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , 
     n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , 
     n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , 
     n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , 
     n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , 
     n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , 
     n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , 
     n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , 
     n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , 
     n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , 
     n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , 
     n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , 
     n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , 
     n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , 
     n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , 
     n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , 
     n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , 
     n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , 
     n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , 
     n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , 
     n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , 
     n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , 
     n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , 
     n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , 
     n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , 
     n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , 
     n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , 
     n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , 
     n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , 
     n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , 
     n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , 
     n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , 
     n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , 
     n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , 
     n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , 
     n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , 
     n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , 
     n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , 
     n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , 
     n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , 
     n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , 
     n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , 
     n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , 
     n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , 
     n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , 
     n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , 
     n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , 
     n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , 
     n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , 
     n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , 
     n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , 
     n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , 
     n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , 
     n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , 
     n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , 
     n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , 
     n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , 
     n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , 
     n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , 
     n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , 
     n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , 
     n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , 
     n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , 
     n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , 
     n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , 
     n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , 
     n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , 
     n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , 
     n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , 
     n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , 
     n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , 
     n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , 
     n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , 
     n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , 
     n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , 
     n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , 
     n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , 
     n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , 
     n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , 
     n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , 
     n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , 
     n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , 
     n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , 
     n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , 
     n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , 
     n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , 
     n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , 
     n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , 
     n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , 
     n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , 
     n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , 
     n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , 
     n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , 
     n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , 
     n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , 
     n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , 
     n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , 
     n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , 
     n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , 
     n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , 
     n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , 
     n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , 
     n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , 
     n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , 
     n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , 
     n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , 
     n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , 
     n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , 
     n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , 
     n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , 
     n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , 
     n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , 
     n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , 
     n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , 
     n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , 
     n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , 
     n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , 
     n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , 
     n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , 
     n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , 
     n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , 
     n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , 
     n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , 
     n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , 
     n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , 
     n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , 
     n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , 
     n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , 
     n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , 
     n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , 
     n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , 
     n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , 
     n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , 
     n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , 
     n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , 
     n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , 
     n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , 
     n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , 
     n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , 
     n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , 
     n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , 
     n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , 
     n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , 
     n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , 
     n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , 
     n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , 
     n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , 
     n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , 
     n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , 
     n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , 
     n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , 
     n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , 
     n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , 
     n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , 
     n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , 
     n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , 
     n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , 
     n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , 
     n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , 
     n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , 
     n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , 
     n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , 
     n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , 
     n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , 
     n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , 
     n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , 
     n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , 
     n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , 
     n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , 
     n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , 
     n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , 
     n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , 
     n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , 
     n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , 
     n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , 
     n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , 
     n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , 
     n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , 
     n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , 
     n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , 
     n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , 
     n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , 
     n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , 
     n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , 
     n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , 
     n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , 
     n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , 
     n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , 
     n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , 
     n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , 
     n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , 
     n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , 
     n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , 
     n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , 
     n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , 
     n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , 
     n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , 
     n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , 
     n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , 
     n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , 
     n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , 
     n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , 
     n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , 
     n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , 
     n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , 
     n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , 
     n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , 
     n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , 
     n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , 
     n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , 
     n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , 
     n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , 
     n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , 
     n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , 
     n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , 
     n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , 
     n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , 
     n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , 
     n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , 
     n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , 
     n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , 
     n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , 
     n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , 
     n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , 
     n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , 
     n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , 
     n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , 
     n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , 
     n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , 
     n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , 
     n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , 
     n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , 
     n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , 
     n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , 
     n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , 
     n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , 
     n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , 
     n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , 
     n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , 
     n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , 
     n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , 
     n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , 
     n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , 
     n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , 
     n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , 
     n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , 
     n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , 
     n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , 
     n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , 
     n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , 
     n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , 
     n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , 
     n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , 
     n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , 
     n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , 
     n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , 
     n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , 
     n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , 
     n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , 
     n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , 
     n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , 
     n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , 
     n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , 
     n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , 
     n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , 
     n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , 
     n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , 
     n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , 
     n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , 
     n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , 
     n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , 
     n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , 
     n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , 
     n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , 
     n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , 
     n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , 
     n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , 
     n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , 
     n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , 
     n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , 
     n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , 
     n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , 
     n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , 
     n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , 
     n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , 
     n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , 
     n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , 
     n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , 
     n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , 
     n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , 
     n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , 
     n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , 
     n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , 
     n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , 
     n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , 
     n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , 
     n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , 
     n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , 
     n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , 
     n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , 
     n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , 
     n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , 
     n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , 
     n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , 
     n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , 
     n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , 
     n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , 
     n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , 
     n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , 
     n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , 
     n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , 
     n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , 
     n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , 
     n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , 
     n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , 
     n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , 
     n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , 
     n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , 
     n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , 
     n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , 
     n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , 
     n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , 
     n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , 
     n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , 
     n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , 
     n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , 
     n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , 
     n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , 
     n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , 
     n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , 
     n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , 
     n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , 
     n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , 
     n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , 
     n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , 
     n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , 
     n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , 
     n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , 
     n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , 
     n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , 
     n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , 
     n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , 
     n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , 
     n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , 
     n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , 
     n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , 
     n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , 
     n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , 
     n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , 
     n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , 
     n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , 
     n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , 
     n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , 
     n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , 
     n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , 
     n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , 
     n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , 
     n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , 
     n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , 
     n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , 
     n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , 
     n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , 
     n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , 
     n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , 
     n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , 
     n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , 
     n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , 
     n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , 
     n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , 
     n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , 
     n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , 
     n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , 
     n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , 
     n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , 
     n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , 
     n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , 
     n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , 
     n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , 
     n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , 
     n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , 
     n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , 
     n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , 
     n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , 
     n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , 
     n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , 
     n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , 
     n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , 
     n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , 
     n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , 
     n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , 
     n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , 
     n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , 
     n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , 
     n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , 
     n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , 
     n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , 
     n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , 
     n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , 
     n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , 
     n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , 
     n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , 
     n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , 
     n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , 
     n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , 
     n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , 
     n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , 
     n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , 
     n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , 
     n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , 
     n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , 
     n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , 
     n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , 
     n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , 
     n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , 
     n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , 
     n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , 
     n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , 
     n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , 
     n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , 
     n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , 
     n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , 
     n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , 
     n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , 
     n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , 
     n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , 
     n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , 
     n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , 
     n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , 
     n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , 
     n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , 
     n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , 
     n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , 
     n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , 
     n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , 
     n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , 
     n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , 
     n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , 
     n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , 
     n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , 
     n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , 
     n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , 
     n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , 
     n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , 
     n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , 
     n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , 
     n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , 
     n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , 
     n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , 
     n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , 
     n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , 
     n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , 
     n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , 
     n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , 
     n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , 
     n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , 
     n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , 
     n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , 
     n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , 
     n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , 
     n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , 
     n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , 
     n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , 
     n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , 
     n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , 
     n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , 
     n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , 
     n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , 
     n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , 
     n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , 
     n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , 
     n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , 
     n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , 
     n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , 
     n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , 
     n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , 
     n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , 
     n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , 
     n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , 
     n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , 
     n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , 
     n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , 
     n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , 
     n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , 
     n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , 
     n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , 
     n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , 
     n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , 
     n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , 
     n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , 
     n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , 
     n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , 
     n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , 
     n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , 
     n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , 
     n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , 
     n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , 
     n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , 
     n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , 
     n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , 
     n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , 
     n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , 
     n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , 
     n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , 
     n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , 
     n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , 
     n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , 
     n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , 
     n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , 
     n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , 
     n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , 
     n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , 
     n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , 
     n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , 
     n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , 
     n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , 
     n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , 
     n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , 
     n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , 
     n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , 
     n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , 
     n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , 
     n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , 
     n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , 
     n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , 
     n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , 
     n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , 
     n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , 
     n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , 
     n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , 
     n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , 
     n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , 
     n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , 
     n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , 
     n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , 
     n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , 
     n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , 
     n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , 
     n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , 
     n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , 
     n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , 
     n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , 
     n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , 
     n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , 
     n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , 
     n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , 
     n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , 
     n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , 
     n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , 
     n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , 
     n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , 
     n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , 
     n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , 
     n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , 
     n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , 
     n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , 
     n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , 
     n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , 
     n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , 
     n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , 
     n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , 
     n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , 
     n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , 
     n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , 
     n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , 
     n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , 
     n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , 
     n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , 
     n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , 
     n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , 
     n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , 
     n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , 
     n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , 
     n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , 
     n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , 
     n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , 
     n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , 
     n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , 
     n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , 
     n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , 
     n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , 
     n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , 
     n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , 
     n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , 
     n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , 
     n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , 
     n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , 
     n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , 
     n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , 
     n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , 
     n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , 
     n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , 
     n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , 
     n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , 
     n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , 
     n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , 
     n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , 
     n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , 
     n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , 
     n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , 
     n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , 
     n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , 
     n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , 
     n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , 
     n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , 
     n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , 
     n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , 
     n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , 
     n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , 
     n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , 
     n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , 
     n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , 
     n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , 
     n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , 
     n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , 
     n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , 
     n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , 
     n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , 
     n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , 
     n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , 
     n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , 
     n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , 
     n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , 
     n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , 
     n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , 
     n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , 
     n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , 
     n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , 
     n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , 
     n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , 
     n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , 
     n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , 
     n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , 
     n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , 
     n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , 
     n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , 
     n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , 
     n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , 
     n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , 
     n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , 
     n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , 
     n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , 
     n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , 
     n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , 
     n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , 
     n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , 
     n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , 
     n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , 
     n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , 
     n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , 
     n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , 
     n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , 
     n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , 
     n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , 
     n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , 
     n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , 
     n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , 
     n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , 
     n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , 
     n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , 
     n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , 
     n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , 
     n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , 
     n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , 
     n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , 
     n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , 
     n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , 
     n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , 
     n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , 
     n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , 
     n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , 
     n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , 
     n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , 
     n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , 
     n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , 
     n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , 
     n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , 
     n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , 
     n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , 
     n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , 
     n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , 
     n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , 
     n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , 
     n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , 
     n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , 
     n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , 
     n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , 
     n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , 
     n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , 
     n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , 
     n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , 
     n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , 
     n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , 
     n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , 
     n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , 
     n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , 
     n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , 
     n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , 
     n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , 
     n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , 
     n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , 
     n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , 
     n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , 
     n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , 
     n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , 
     n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , 
     n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , 
     n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , 
     n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , 
     n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , 
     n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , 
     n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , 
     n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , 
     n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , 
     n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , 
     n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , 
     n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , 
     n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , 
     n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , 
     n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , 
     n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , 
     n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , 
     n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , 
     n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , 
     n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , 
     n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , 
     n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , 
     n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , 
     n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , 
     n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , 
     n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , 
     n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , 
     n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , 
     n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , 
     n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , 
     n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , 
     n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , 
     n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , 
     n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , 
     n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , 
     n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , 
     n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , 
     n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , 
     n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , 
     n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , 
     n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , 
     n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , 
     n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , 
     n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , 
     n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , 
     n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , 
     n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , 
     n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , 
     n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , 
     n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , 
     n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , 
     n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , 
     n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , 
     n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , 
     n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , 
     n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , 
     n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , 
     n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , 
     n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , 
     n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , 
     n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , 
     n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , 
     n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , 
     n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , 
     n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , 
     n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , 
     n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , 
     n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , 
     n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , 
     n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , 
     n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , 
     n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , 
     n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , 
     n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , 
     n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , 
     n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , 
     n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , 
     n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , 
     n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , 
     n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , 
     n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , 
     n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , 
     n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , 
     n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , 
     n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , 
     n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , 
     n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , 
     n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , 
     n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , 
     n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , 
     n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , 
     n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , 
     n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , 
     n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , 
     n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , 
     n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , 
     n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , 
     n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , 
     n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , 
     n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , 
     n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , 
     n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , 
     n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , 
     n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , 
     n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , 
     n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , 
     n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , 
     n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , 
     n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , 
     n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , 
     n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , 
     n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , 
     n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , 
     n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , 
     n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , 
     n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , 
     n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , 
     n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , 
     n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , 
     n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , 
     n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , 
     n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , 
     n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , 
     n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , 
     n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , 
     n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , 
     n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , 
     n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , 
     n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , 
     n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , 
     n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , 
     n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , 
     n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , 
     n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , 
     n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , 
     n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , 
     n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , 
     n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , 
     n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , 
     n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , 
     n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , 
     n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , 
     n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , 
     n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , 
     n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , 
     n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , 
     n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , 
     n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , 
     n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , 
     n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , 
     n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , 
     n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , 
     n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , 
     n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , 
     n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , 
     n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , 
     n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , 
     n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , 
     n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , 
     n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , 
     n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , 
     n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , 
     n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , 
     n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , 
     n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , 
     n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , 
     n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , 
     n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , 
     n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , 
     n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , 
     n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , 
     n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , 
     n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , 
     n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , 
     n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , 
     n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , 
     n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , 
     n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , 
     n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , 
     n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , 
     n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , 
     n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , 
     n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , 
     n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , 
     n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , 
     n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , 
     n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , 
     n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , 
     n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , 
     n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , 
     n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , 
     n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , 
     n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , 
     n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , 
     n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , 
     n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , 
     n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , 
     n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , 
     n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , 
     n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , 
     n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , 
     n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , 
     n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , 
     n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , 
     n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , 
     n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , 
     n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , 
     n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , 
     n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , 
     n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , 
     n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , 
     n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , 
     n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , 
     n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , 
     n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , 
     n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , 
     n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , 
     n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , 
     n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , 
     n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , 
     n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , 
     n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , 
     n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , 
     n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , 
     n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , 
     n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , 
     n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , 
     n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , 
     n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , 
     n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , 
     n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , 
     n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , 
     n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , 
     n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , 
     n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , 
     n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , 
     n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , 
     n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , 
     n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , 
     n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , 
     n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , 
     n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , 
     n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , 
     n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , 
     n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , 
     n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , 
     n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , 
     n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , 
     n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , 
     n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , 
     n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , 
     n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , 
     n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , 
     n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , 
     n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , 
     n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , 
     n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , 
     n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , 
     n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , 
     n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , 
     n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , 
     n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , 
     n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , 
     n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , 
     n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , 
     n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , 
     n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , 
     n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , 
     n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , 
     n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , 
     n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , 
     n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , 
     n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , 
     n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , 
     n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , 
     n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , 
     n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , 
     n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , 
     n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , 
     n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , 
     n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , 
     n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , 
     n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , 
     n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , 
     n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , 
     n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , 
     n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , 
     n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , 
     n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , 
     n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , 
     n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , 
     n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , 
     n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , 
     n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , 
     n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , 
     n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , 
     n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , 
     n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , 
     n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , 
     n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , 
     n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , 
     n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , 
     n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , 
     n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , 
     n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , 
     n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , 
     n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , 
     n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , 
     n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , 
     n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , 
     n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , 
     n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , 
     n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , 
     n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , 
     n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , 
     n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , 
     n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , 
     n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , 
     n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , 
     n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , 
     n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , 
     n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , 
     n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , 
     n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , 
     n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , 
     n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , 
     n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , 
     n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , 
     n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , 
     n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , 
     n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , 
     n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , 
     n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , 
     n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , 
     n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , 
     n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , 
     n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , 
     n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , 
     n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , 
     n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , 
     n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , 
     n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , 
     n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , 
     n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , 
     n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , 
     n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , 
     n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , 
     n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , 
     n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , 
     n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , 
     n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , 
     n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , 
     n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , 
     n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , 
     n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , 
     n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , 
     n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , 
     n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , 
     n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , 
     n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , 
     n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , 
     n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , 
     n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , 
     n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , 
     n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , 
     n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , 
     n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , 
     n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , 
     n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , 
     n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , 
     n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , 
     n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , 
     n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , 
     n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , 
     n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , 
     n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , 
     n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , 
     n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , 
     n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , 
     n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , 
     n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , 
     n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , 
     n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , 
     n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , 
     n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , 
     n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , 
     n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , 
     n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , 
     n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , 
     n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , 
     n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , 
     n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , 
     n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , 
     n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , 
     n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , 
     n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , 
     n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , 
     n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , 
     n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , 
     n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , 
     n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , 
     n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , 
     n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , 
     n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , 
     n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , 
     n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , 
     n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , 
     n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , 
     n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , 
     n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , 
     n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , 
     n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , 
     n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , 
     n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , 
     n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , 
     n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , 
     n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , 
     n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , 
     n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , 
     n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , 
     n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , 
     n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , 
     n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , 
     n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , 
     n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , 
     n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , 
     n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , 
     n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , 
     n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , 
     n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , 
     n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , 
     n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , 
     n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , 
     n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , 
     n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , 
     n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , 
     n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , 
     n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , 
     n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , 
     n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , 
     n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , 
     n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , 
     n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , 
     n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , 
     n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , 
     n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , 
     n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , 
     n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , 
     n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , 
     n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , 
     n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , 
     n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , 
     n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , 
     n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , 
     n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , 
     n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , 
     n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , 
     n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , 
     n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , 
     n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , 
     n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , 
     n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , 
     n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , 
     n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , 
     n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , 
     n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , 
     n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , 
     n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , 
     n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , 
     n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , 
     n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , 
     n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , 
     n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , 
     n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , 
     n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , 
     n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , 
     n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , 
     n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , 
     n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , 
     n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , 
     n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , 
     n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , 
     n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , 
     n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , 
     n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , 
     n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , 
     n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , 
     n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , 
     n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , 
     n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , 
     n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , 
     n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , 
     n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , 
     n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , 
     n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , 
     n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , 
     n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , 
     n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , 
     n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , 
     n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , 
     n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , 
     n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , 
     n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , 
     n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , 
     n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , 
     n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , 
     n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , 
     n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , 
     n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , 
     n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , 
     n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , 
     n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , 
     n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , 
     n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , 
     n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , 
     n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , 
     n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , 
     n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , 
     n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , 
     n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , 
     n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , 
     n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , 
     n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , 
     n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , 
     n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , 
     n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , 
     n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , 
     n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , 
     n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , 
     n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , 
     n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , 
     n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , 
     n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , 
     n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , 
     n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , 
     n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , 
     n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , 
     n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , 
     n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , 
     n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , 
     n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , 
     n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , 
     n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , 
     n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , 
     n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , 
     n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , 
     n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , 
     n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , 
     n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , 
     n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , 
     n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , 
     n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , 
     n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , 
     n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , 
     n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , 
     n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , 
     n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , 
     n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , 
     n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , 
     n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , 
     n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , 
     n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , 
     n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , 
     n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , 
     n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , 
     n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , 
     n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , 
     n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , 
     n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , 
     n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , 
     n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , 
     n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , 
     n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , 
     n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , 
     n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , 
     n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , 
     n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , 
     n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , 
     n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , 
     n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , 
     n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , 
     n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , 
     n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , 
     n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , 
     n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , 
     n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , 
     n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , 
     n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , 
     n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , 
     n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , 
     n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , 
     n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , 
     n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , 
     n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , 
     n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , 
     n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , 
     n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , 
     n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , 
     n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , 
     n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , 
     n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , 
     n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , 
     n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , 
     n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , 
     n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , 
     n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , 
     n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , 
     n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , 
     n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , 
     n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , 
     n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , 
     n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , 
     n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , 
     n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , 
     n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , 
     n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , 
     n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , 
     n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , 
     n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , 
     n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , 
     n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , 
     n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , 
     n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , 
     n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , 
     n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , 
     n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , 
     n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , 
     n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , 
     n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , 
     n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , 
     n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , 
     n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , 
     n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , 
     n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , 
     n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , 
     n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , 
     n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , 
     n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , 
     n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , 
     n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , 
     n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , 
     n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , 
     n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , 
     n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , 
     n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , 
     n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , 
     n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , 
     n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , 
     n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , 
     n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , 
     n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , 
     n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , 
     n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , 
     n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , 
     n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , 
     n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , 
     n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , 
     n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , 
     n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , 
     n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , 
     n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , 
     n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , 
     n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , 
     n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , 
     n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , 
     n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , 
     n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , 
     n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , 
     n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , 
     n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , 
     n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , 
     n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , 
     n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , 
     n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , 
     n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , 
     n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , 
     n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , 
     n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , 
     n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , 
     n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , 
     n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , 
     n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , 
     n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , 
     n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , 
     n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , 
     n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , 
     n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , 
     n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , 
     n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , 
     n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , 
     n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , 
     n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , 
     n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , 
     n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , 
     n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , 
     n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , 
     n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , 
     n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , 
     n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , 
     n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , 
     n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , 
     n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , 
     n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , 
     n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , 
     n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , 
     n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , 
     n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , 
     n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , 
     n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , 
     n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , 
     n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , 
     n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , 
     n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , 
     n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , 
     n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , 
     n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , 
     n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , 
     n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , 
     n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , 
     n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , 
     n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , 
     n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , 
     n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , 
     n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , 
     n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , 
     n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , 
     n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , 
     n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , 
     n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , 
     n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , 
     n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , 
     n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , 
     n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , 
     n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , 
     n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , 
     n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , 
     n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , 
     n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , 
     n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , 
     n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , 
     n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , 
     n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , 
     n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , 
     n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , 
     n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , 
     n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , 
     n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , 
     n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , 
     n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , 
     n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , 
     n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , 
     n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , 
     n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , 
     n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , 
     n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , 
     n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , 
     n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , 
     n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , 
     n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , 
     n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , 
     n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , 
     n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , 
     n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , 
     n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , 
     n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , 
     n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , 
     n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , 
     n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , 
     n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , 
     n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , 
     n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , 
     n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , 
     n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , 
     n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , 
     n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , 
     n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , 
     n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , 
     n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , 
     n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , 
     n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , 
     n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , 
     n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , 
     n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , 
     n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , 
     n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , 
     n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , 
     n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , 
     n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , 
     n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , 
     n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , 
     n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , 
     n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , 
     n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , 
     n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , 
     n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , 
     n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , 
     n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , 
     n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , 
     n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , 
     n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , 
     n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , 
     n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , 
     n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , 
     n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , 
     n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , 
     n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , 
     n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , 
     n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , 
     n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , 
     n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , 
     n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , 
     n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , 
     n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , 
     n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , 
     n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , 
     n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , 
     n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , 
     n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , 
     n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , 
     n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , 
     n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , 
     n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , 
     n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , 
     n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , 
     n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , 
     n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , 
     n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , 
     n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , 
     n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , 
     n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , 
     n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , 
     n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , 
     n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , 
     n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , 
     n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , 
     n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , 
     n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , 
     n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , 
     n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , 
     n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , 
     n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , 
     n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , 
     n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , 
     n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , 
     n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , 
     n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , 
     n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , 
     n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , 
     n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , 
     n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , 
     n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , 
     n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , 
     n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , 
     n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , 
     n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , 
     n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , 
     n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , 
     n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , 
     n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , 
     n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , 
     n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , 
     n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , 
     n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , 
     n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , 
     n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , 
     n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , 
     n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , 
     n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , 
     n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , 
     n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , 
     n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , 
     n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , 
     n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , 
     n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , 
     n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , 
     n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , 
     n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , 
     n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , 
     n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , 
     n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , 
     n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , 
     n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , 
     n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , 
     n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , 
     n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , 
     n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , 
     n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , 
     n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , 
     n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , 
     n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , 
     n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , 
     n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , 
     n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , 
     n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , 
     n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , 
     n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , 
     n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , 
     n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , 
     n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , 
     n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , 
     n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , 
     n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , 
     n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , 
     n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , 
     n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , 
     n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , 
     n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , 
     n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , 
     n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , 
     n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , 
     n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , 
     n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , 
     n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , 
     n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , 
     n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , 
     n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , 
     n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , 
     n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , 
     n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , 
     n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , 
     n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , 
     n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , 
     n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , 
     n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , 
     n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , 
     n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , 
     n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , 
     n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , 
     n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , 
     n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , 
     n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , 
     n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , 
     n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , 
     n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , 
     n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , 
     n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , 
     n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , 
     n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , 
     n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , 
     n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , 
     n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , 
     n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , 
     n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , 
     n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , 
     n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , 
     n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , 
     n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , 
     n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , 
     n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , 
     n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , 
     n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , 
     n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , 
     n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , 
     n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , 
     n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , 
     n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , 
     n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , 
     n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , 
     n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , 
     n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , 
     n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , 
     n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , 
     n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , 
     n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , 
     n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , 
     n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , 
     n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , 
     n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , 
     n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , 
     n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , 
     n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , 
     n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , 
     n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , 
     n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , 
     n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , 
     n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , 
     n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , 
     n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , 
     n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , 
     n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , 
     n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , 
     n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , 
     n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , 
     n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , 
     n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , 
     n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , 
     n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , 
     n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , 
     n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , 
     n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , 
     n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , 
     n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , 
     n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , 
     n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , 
     n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , 
     n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , 
     n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , 
     n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , 
     n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , 
     n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , 
     n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , 
     n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , 
     n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , 
     n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , 
     n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , 
     n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , 
     n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , 
     n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , 
     n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , 
     n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , 
     n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , 
     n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , 
     n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , 
     n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , 
     n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , 
     n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , 
     n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , 
     n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , 
     n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , 
     n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , 
     n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , 
     n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , 
     n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , 
     n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , 
     n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , 
     n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , 
     n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , 
     n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , 
     n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , 
     n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , 
     n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , 
     n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , 
     n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , 
     n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , 
     n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , 
     n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , 
     n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , 
     n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , 
     n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , 
     n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , 
     n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , 
     n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , 
     n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , 
     n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , 
     n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , 
     n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , 
     n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , 
     n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , 
     n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , 
     n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , 
     n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , 
     n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , 
     n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , 
     n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , 
     n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , 
     n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , 
     n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , 
     n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , 
     n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , 
     n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , 
     n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , 
     n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , 
     n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , 
     n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , 
     n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , 
     n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , 
     n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , 
     n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , 
     n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , 
     n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , 
     n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , 
     n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , 
     n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , 
     n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , 
     n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , 
     n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , 
     n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , 
     n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , 
     n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , 
     n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , 
     n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , 
     n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , 
     n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , 
     n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , 
     n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , 
     n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , 
     n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , 
     n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , 
     n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , 
     n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , 
     n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , 
     n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , 
     n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , 
     n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , 
     n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , 
     n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , 
     n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , 
     n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , 
     n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , 
     n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , 
     n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , 
     n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , 
     n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , 
     n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , 
     n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , 
     n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , 
     n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , 
     n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , 
     n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , 
     n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , 
     n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , 
     n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , 
     n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , 
     n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , 
     n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , 
     n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , 
     n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , 
     n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , 
     n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , 
     n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , 
     n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , 
     n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , 
     n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , 
     n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , 
     n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , 
     n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , 
     n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , 
     n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , 
     n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , 
     n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , 
     n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , 
     n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , 
     n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , 
     n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , 
     n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , 
     n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , 
     n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , 
     n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , 
     n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , 
     n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , 
     n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , 
     n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , 
     n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , 
     n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , 
     n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , 
     n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , 
     n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , 
     n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , 
     n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , 
     n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , 
     n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , 
     n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , 
     n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , 
     n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , 
     n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , 
     n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , 
     n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , 
     n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , 
     n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , 
     n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , 
     n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , 
     n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , 
     n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , 
     n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , 
     n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , 
     n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , 
     n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , 
     n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , 
     n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , 
     n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , 
     n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , 
     n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , 
     n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , 
     n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , 
     n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , 
     n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , 
     n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , 
     n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , 
     n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , 
     n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , 
     n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , 
     n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , 
     n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , 
     n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , 
     n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , 
     n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , 
     n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , 
     n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , 
     n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , 
     n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , 
     n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , 
     n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , 
     n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , 
     n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , 
     n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , 
     n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , 
     n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , 
     n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , 
     n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , 
     n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , 
     n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , 
     n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , 
     n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , 
     n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , 
     n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , 
     n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , 
     n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , 
     n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , 
     n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , 
     n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , 
     n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , 
     n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , 
     n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , 
     n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , 
     n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , 
     n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , 
     n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , 
     n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , 
     n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , 
     n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , 
     n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , 
     n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , 
     n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , 
     n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , 
     n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , 
     n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , 
     n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , 
     n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , 
     n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , 
     n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , 
     n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , 
     n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , 
     n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , 
     n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , 
     n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , 
     n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , 
     n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , 
     n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , 
     n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , 
     n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , 
     n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , 
     n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , 
     n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , 
     n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , 
     n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , 
     n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , 
     n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , 
     n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , 
     n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , 
     n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , 
     n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , 
     n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , 
     n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , 
     n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , 
     n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , 
     n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , 
     n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , 
     n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , 
     n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , 
     n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , 
     n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , 
     n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , 
     n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , 
     n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , 
     n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , 
     n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , 
     n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , 
     n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , 
     n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , 
     n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , 
     n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , 
     n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , 
     n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , 
     n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , 
     n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , 
     n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , 
     n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , 
     n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , 
     n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , 
     n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , 
     n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , 
     n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , 
     n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , 
     n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , 
     n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , 
     n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , 
     n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , 
     n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , 
     n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , 
     n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , 
     n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , 
     n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , 
     n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , 
     n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , 
     n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , 
     n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , 
     n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , 
     n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , 
     n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , 
     n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , 
     n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , 
     n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , 
     n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , 
     n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , 
     n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , 
     n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , 
     n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , 
     n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , 
     n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , 
     n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , 
     n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , 
     n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , 
     n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , 
     n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , 
     n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , 
     n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , 
     n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , 
     n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , 
     n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , 
     n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , 
     n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , 
     n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , 
     n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , 
     n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , 
     n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , 
     n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , 
     n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , 
     n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , 
     n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , 
     n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , 
     n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , 
     n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , 
     n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , 
     n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , 
     n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , 
     n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , 
     n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , 
     n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , 
     n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , 
     n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , 
     n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , 
     n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , 
     n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , 
     n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , 
     n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , 
     n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , 
     n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , 
     n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , 
     n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , 
     n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , 
     n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , 
     n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , 
     n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , 
     n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , 
     n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , 
     n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , 
     n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , 
     n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , 
     n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , 
     n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , 
     n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , 
     n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , 
     n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , 
     n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , 
     n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , 
     n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , 
     n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , 
     n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , 
     n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , 
     n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , 
     n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , 
     n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , 
     n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , 
     n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , 
     n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , 
     n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , 
     n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , 
     n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , 
     n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , 
     n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , 
     n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , 
     n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , 
     n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , 
     n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , 
     n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , 
     n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , 
     n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , 
     n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , 
     n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , 
     n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , 
     n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , 
     n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , 
     n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , 
     n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , 
     n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , 
     n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , 
     n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , 
     n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , 
     n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , 
     n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , 
     n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , 
     n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , 
     n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , 
     n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , 
     n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , 
     n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , 
     n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , 
     n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , 
     n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , 
     n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , 
     n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , 
     n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , 
     n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , 
     n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , 
     n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , 
     n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , 
     n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , 
     n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , 
     n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , 
     n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , 
     n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , 
     n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , 
     n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , 
     n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , 
     n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , 
     n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , 
     n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , 
     n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , 
     n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , 
     n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , 
     n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , 
     n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , 
     n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , 
     n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , 
     n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , 
     n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , 
     n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , 
     n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , 
     n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , 
     n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , 
     n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , 
     n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , 
     n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , 
     n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , 
     n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , 
     n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , 
     n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , 
     n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , 
     n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , 
     n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , 
     n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , 
     n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , 
     n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , 
     n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , 
     n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , 
     n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , 
     n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , 
     n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , 
     n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , 
     n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , 
     n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , 
     n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , 
     n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , 
     n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , 
     n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , 
     n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , 
     n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , 
     n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , 
     n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , 
     n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , 
     n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , 
     n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , 
     n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , 
     n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , 
     n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , 
     n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , 
     n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , 
     n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , 
     n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , 
     n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , 
     n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , 
     n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , 
     n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , 
     n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , 
     n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , 
     n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , 
     n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , 
     n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , 
     n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , 
     n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , 
     n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , 
     n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , 
     n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , 
     n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , 
     n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , 
     n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , 
     n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , 
     n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , 
     n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , 
     n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , 
     n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , 
     n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , 
     n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , 
     n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , 
     n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , 
     n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , 
     n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , 
     n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , 
     n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , 
     n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , 
     n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , 
     n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , 
     n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , 
     n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , 
     n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , 
     n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , 
     n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , 
     n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , 
     n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , 
     n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , 
     n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , 
     n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , 
     n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , 
     n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , 
     n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , 
     n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , 
     n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , 
     n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , 
     n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , 
     n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , 
     n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , 
     n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , 
     n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , 
     n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , 
     n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , 
     n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , 
     n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , 
     n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , 
     n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , 
     n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , 
     n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , 
     n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , 
     n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , 
     n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , 
     n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , 
     n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , 
     n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , 
     n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , 
     n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , 
     n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , 
     n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , 
     n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , 
     n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , 
     n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , 
     n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , 
     n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , 
     n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , 
     n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , 
     n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , 
     n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , 
     n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , 
     n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , 
     n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , 
     n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , 
     n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , 
     n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , 
     n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , 
     n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , 
     n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , 
     n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , 
     n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , 
     n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , 
     n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , 
     n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , 
     n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , 
     n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , 
     n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , 
     n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , 
     n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , 
     n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , 
     n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , 
     n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , 
     n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , 
     n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , 
     n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , 
     n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , 
     n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , 
     n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , 
     n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , 
     n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , 
     n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , 
     n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , 
     n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , 
     n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , 
     n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , 
     n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , 
     n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , 
     n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , 
     n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , 
     n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , 
     n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , 
     n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , 
     n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , 
     n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , 
     n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , 
     n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , 
     n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , 
     n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , 
     n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , 
     n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , 
     n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , 
     n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , 
     n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , 
     n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , 
     n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , 
     n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , 
     n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , 
     n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , 
     n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , 
     n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , 
     n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , 
     n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , 
     n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , 
     n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , 
     n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , 
     n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , 
     n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , 
     n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , 
     n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , 
     n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , 
     n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , 
     n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , 
     n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , 
     n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , 
     n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , 
     n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , 
     n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , 
     n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , 
     n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , 
     n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , 
     n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , 
     n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , 
     n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , 
     n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , 
     n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , 
     n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , 
     n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , 
     n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , 
     n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , 
     n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , 
     n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , 
     n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , 
     n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , 
     n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , 
     n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , 
     n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , 
     n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , 
     n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , 
     n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , 
     n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , 
     n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , 
     n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , 
     n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , 
     n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , 
     n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , 
     n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , 
     n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , 
     n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , 
     n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , 
     n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , 
     n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , 
     n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , 
     n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , 
     n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , 
     n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , 
     n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , 
     n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , 
     n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , 
     n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , 
     n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , 
     n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , 
     n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , 
     n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , 
     n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , 
     n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , 
     n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , 
     n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , 
     n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , 
     n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , 
     n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , 
     n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , 
     n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , 
     n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , 
     n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , 
     n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , 
     n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , 
     n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , 
     n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , 
     n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , 
     n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , 
     n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , 
     n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , 
     n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , 
     n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , 
     n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , 
     n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , 
     n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , 
     n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , 
     n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , 
     n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , 
     n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , 
     n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , 
     n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , 
     n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , 
     n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , 
     n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , 
     n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , 
     n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , 
     n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , 
     n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , 
     n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , 
     n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , 
     n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , 
     n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , 
     n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , 
     n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , 
     n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , 
     n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , 
     n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , 
     n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , 
     n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , 
     n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , 
     n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , 
     n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , 
     n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , 
     n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , 
     n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , 
     n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , 
     n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , 
     n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , 
     n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , 
     n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , 
     n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , 
     n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , 
     n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , 
     n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , 
     n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , 
     n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , 
     n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , 
     n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , 
     n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , 
     n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , 
     n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , 
     n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , 
     n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , 
     n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , 
     n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , 
     n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , 
     n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , 
     n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , 
     n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , 
     n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , 
     n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , 
     n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , 
     n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , 
     n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , 
     n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , 
     n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , 
     n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , 
     n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , 
     n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , 
     n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , 
     n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , 
     n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , 
     n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , 
     n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , 
     n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , 
     n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , 
     n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , 
     n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , 
     n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , 
     n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , 
     n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , 
     n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , 
     n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , 
     n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , 
     n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , 
     n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , 
     n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , 
     n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , 
     n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , 
     n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , 
     n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , 
     n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , 
     n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , 
     n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , 
     n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , 
     n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , 
     n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , 
     n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , 
     n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , 
     n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , 
     n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , 
     n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , 
     n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , 
     n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , 
     n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , 
     n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , 
     n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , 
     n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , 
     n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , 
     n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , 
     n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , 
     n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , 
     n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , 
     n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , 
     n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , 
     n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , 
     n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , 
     n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , 
     n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , 
     n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , 
     n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , 
     n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , 
     n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , 
     n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , 
     n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , 
     n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , 
     n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , 
     n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , 
     n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , 
     n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , 
     n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , 
     n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , 
     n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , 
     n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , 
     n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , 
     n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , 
     n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , 
     n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , 
     n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , 
     n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , 
     n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , 
     n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , 
     n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , 
     n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , 
     n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , 
     n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , 
     n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , 
     n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , 
     n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , 
     n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , 
     n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , 
     n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , 
     n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , 
     n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , 
     n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , 
     n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , 
     n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , 
     n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , 
     n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , 
     n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , 
     n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , 
     n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , 
     n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , 
     n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , 
     n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , 
     n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , 
     n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , 
     n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , 
     n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , 
     n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , 
     n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , 
     n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , 
     n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , 
     n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , 
     n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , 
     n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , 
     n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , 
     n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , 
     n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , 
     n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , 
     n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , 
     n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , 
     n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , 
     n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , 
     n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , 
     n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , 
     n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , 
     n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , 
     n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , 
     n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , 
     n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , 
     n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , 
     n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , 
     n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , 
     n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , 
     n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , 
     n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , 
     n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , 
     n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , 
     n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , 
     n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , 
     n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , 
     n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , 
     n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , 
     n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , 
     n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , 
     n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , 
     n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , 
     n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , 
     n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , 
     n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , 
     n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , 
     n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , 
     n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , 
     n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , 
     n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , 
     n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , 
     n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , 
     n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , 
     n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , 
     n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , 
     n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , 
     n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , 
     n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , 
     n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , 
     n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , 
     n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , 
     n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , 
     n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , 
     n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , 
     n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , 
     n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , 
     n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , 
     n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , 
     n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , 
     n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , 
     n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , 
     n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , 
     n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , 
     n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , 
     n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , 
     n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , 
     n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , 
     n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , 
     n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , 
     n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , 
     n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , 
     n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , 
     n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , 
     n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , 
     n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , 
     n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , 
     n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , 
     n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , 
     n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , 
     n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , 
     n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , 
     n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , 
     n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , 
     n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , 
     n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , 
     n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , 
     n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , 
     n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , 
     n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , 
     n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , 
     n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , 
     n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , 
     n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , 
     n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , 
     n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , 
     n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , 
     n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , 
     n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , 
     n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , 
     n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , 
     n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , 
     n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , 
     n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , 
     n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , 
     n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , 
     n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , 
     n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , 
     n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , 
     n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , 
     n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , 
     n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , 
     n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , 
     n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , 
     n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , 
     n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , 
     n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , 
     n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , 
     n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , 
     n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , 
     n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , 
     n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , 
     n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , 
     n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , 
     n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , 
     n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , 
     n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , 
     n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , 
     n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , 
     n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , 
     n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , 
     n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , 
     n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , 
     n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , 
     n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , 
     n64901 , n64902 , n64903 , n64904 , n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , 
     n64911 , n64912 , n64913 , n64914 , n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , 
     n64921 , n64922 , n64923 , n64924 , n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , 
     n64931 , n64932 , n64933 , n64934 , n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , 
     n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , 
     n64951 , n64952 , n64953 , n64954 , n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , 
     n64961 , n64962 , n64963 , n64964 , n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , 
     n64971 , n64972 , n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , 
     n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , 
     n64991 , n64992 , n64993 , n64994 , n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , 
     n65001 , n65002 , n65003 , n65004 , n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , 
     n65011 , n65012 , n65013 , n65014 , n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , 
     n65021 , n65022 , n65023 , n65024 , n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , 
     n65031 , n65032 , n65033 , n65034 , n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , 
     n65041 , n65042 , n65043 , n65044 , n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , 
     n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , 
     n65061 , n65062 , n65063 , n65064 , n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , 
     n65071 , n65072 , n65073 , n65074 , n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , 
     n65081 , n65082 , n65083 , n65084 , n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , 
     n65091 , n65092 , n65093 , n65094 , n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , 
     n65101 , n65102 , n65103 , n65104 , n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , 
     n65111 , n65112 , n65113 , n65114 , n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , 
     n65121 , n65122 , n65123 , n65124 , n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , 
     n65131 , n65132 , n65133 , n65134 , n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , 
     n65141 , n65142 , n65143 , n65144 , n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , 
     n65151 , n65152 , n65153 , n65154 , n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , 
     n65161 , n65162 , n65163 , n65164 , n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , 
     n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , 
     n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , 
     n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , 
     n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , 
     n65211 , n65212 , n65213 , n65214 , n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , 
     n65221 , n65222 , n65223 , n65224 , n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , 
     n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , 
     n65241 , n65242 , n65243 , n65244 , n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , 
     n65251 , n65252 , n65253 , n65254 , n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , 
     n65261 , n65262 , n65263 , n65264 , n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , 
     n65271 , n65272 , n65273 , n65274 , n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , 
     n65281 , n65282 , n65283 , n65284 , n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , 
     n65291 , n65292 , n65293 , n65294 , n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , 
     n65301 , n65302 , n65303 , n65304 , n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , 
     n65311 , n65312 , n65313 , n65314 , n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , 
     n65321 , n65322 , n65323 , n65324 , n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , 
     n65331 , n65332 , n65333 , n65334 , n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , 
     n65341 , n65342 , n65343 , n65344 , n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , 
     n65351 , n65352 , n65353 , n65354 , n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , 
     n65361 , n65362 , n65363 , n65364 , n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , 
     n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , 
     n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , 
     n65391 , n65392 , n65393 , n65394 , n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , 
     n65401 , n65402 , n65403 , n65404 , n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , 
     n65411 , n65412 , n65413 , n65414 , n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , 
     n65421 , n65422 , n65423 , n65424 , n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , 
     n65431 , n65432 , n65433 , n65434 , n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , 
     n65441 , n65442 , n65443 , n65444 , n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , 
     n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , 
     n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , 
     n65471 , n65472 , n65473 , n65474 , n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , 
     n65481 , n65482 , n65483 , n65484 , n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , 
     n65491 , n65492 , n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , 
     n65501 , n65502 , n65503 , n65504 , n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , 
     n65511 , n65512 , n65513 , n65514 , n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , 
     n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , 
     n65531 , n65532 , n65533 , n65534 , n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , 
     n65541 , n65542 , n65543 , n65544 , n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , 
     n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , 
     n65561 , n65562 , n65563 , n65564 , n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , 
     n65571 , n65572 , n65573 , n65574 , n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , 
     n65581 , n65582 , n65583 , n65584 , n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , 
     n65591 , n65592 , n65593 , n65594 , n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , 
     n65601 , n65602 , n65603 , n65604 , n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , 
     n65611 , n65612 , n65613 , n65614 , n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , 
     n65621 , n65622 , n65623 , n65624 , n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , 
     n65631 , n65632 , n65633 , n65634 , n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , 
     n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , 
     n65651 , n65652 , n65653 , n65654 , n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , 
     n65661 , n65662 , n65663 , n65664 , n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , 
     n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , 
     n65681 , n65682 , n65683 , n65684 , n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , 
     n65691 , n65692 , n65693 , n65694 , n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , 
     n65701 , n65702 , n65703 , n65704 , n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , 
     n65711 , n65712 , n65713 , n65714 , n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , 
     n65721 , n65722 , n65723 , n65724 , n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , 
     n65731 , n65732 , n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , 
     n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , 
     n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , 
     n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , 
     n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , 
     n65781 , n65782 , n65783 , n65784 , n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , 
     n65791 , n65792 , n65793 , n65794 , n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , 
     n65801 , n65802 , n65803 , n65804 , n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , 
     n65811 , n65812 , n65813 , n65814 , n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , 
     n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , 
     n65831 , n65832 , n65833 , n65834 , n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , 
     n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , 
     n65851 , n65852 , n65853 , n65854 , n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , 
     n65861 , n65862 , n65863 , n65864 , n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , 
     n65871 , n65872 , n65873 , n65874 , n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , 
     n65881 , n65882 , n65883 , n65884 , n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , 
     n65891 , n65892 , n65893 , n65894 , n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , 
     n65901 , n65902 , n65903 , n65904 , n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , 
     n65911 , n65912 , n65913 , n65914 , n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , 
     n65921 , n65922 , n65923 , n65924 , n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , 
     n65931 , n65932 , n65933 , n65934 , n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , 
     n65941 , n65942 , n65943 , n65944 , n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , 
     n65951 , n65952 , n65953 , n65954 , n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , 
     n65961 , n65962 , n65963 , n65964 , n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , 
     n65971 , n65972 , n65973 , n65974 , n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , 
     n65981 , n65982 , n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , 
     n65991 , n65992 , n65993 , n65994 , n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , 
     n66001 , n66002 , n66003 , n66004 , n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , 
     n66011 , n66012 , n66013 , n66014 , n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , 
     n66021 , n66022 , n66023 , n66024 , n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , 
     n66031 , n66032 , n66033 , n66034 , n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , 
     n66041 , n66042 , n66043 , n66044 , n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , 
     n66051 , n66052 , n66053 , n66054 , n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , 
     n66061 , n66062 , n66063 , n66064 , n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , 
     n66071 , n66072 , n66073 , n66074 , n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , 
     n66081 , n66082 , n66083 , n66084 , n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , 
     n66091 , n66092 , n66093 , n66094 , n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , 
     n66101 , n66102 , n66103 , n66104 , n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , 
     n66111 , n66112 , n66113 , n66114 , n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , 
     n66121 , n66122 , n66123 , n66124 , n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , 
     n66131 , n66132 , n66133 , n66134 , n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , 
     n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , 
     n66151 , n66152 , n66153 , n66154 , n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , 
     n66161 , n66162 , n66163 , n66164 , n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , 
     n66171 , n66172 , n66173 , n66174 , n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , 
     n66181 , n66182 , n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , 
     n66191 , n66192 , n66193 , n66194 , n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , 
     n66201 , n66202 , n66203 , n66204 , n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , 
     n66211 , n66212 , n66213 , n66214 , n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , 
     n66221 , n66222 , n66223 , n66224 , n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , 
     n66231 , n66232 , n66233 , n66234 , n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , 
     n66241 , n66242 , n66243 , n66244 , n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , 
     n66251 , n66252 , n66253 , n66254 , n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , 
     n66261 , n66262 , n66263 , n66264 , n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , 
     n66271 , n66272 , n66273 , n66274 , n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , 
     n66281 , n66282 , n66283 , n66284 , n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , 
     n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , 
     n66301 , n66302 , n66303 , n66304 , n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , 
     n66311 , n66312 , n66313 , n66314 , n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , 
     n66321 , n66322 , n66323 , n66324 , n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , 
     n66331 , n66332 , n66333 , n66334 , n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , 
     n66341 , n66342 , n66343 , n66344 , n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , 
     n66351 , n66352 , n66353 , n66354 , n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , 
     n66361 , n66362 , n66363 , n66364 , n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , 
     n66371 , n66372 , n66373 , n66374 , n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , 
     n66381 , n66382 , n66383 , n66384 , n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , 
     n66391 , n66392 , n66393 , n66394 , n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , 
     n66401 , n66402 , n66403 , n66404 , n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , 
     n66411 , n66412 , n66413 , n66414 , n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , 
     n66421 , n66422 , n66423 , n66424 , n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , 
     n66431 , n66432 , n66433 , n66434 , n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , 
     n66441 , n66442 , n66443 , n66444 , n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , 
     n66451 , n66452 , n66453 , n66454 , n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , 
     n66461 , n66462 , n66463 , n66464 , n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , 
     n66471 , n66472 , n66473 , n66474 , n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , 
     n66481 , n66482 , n66483 , n66484 , n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , 
     n66491 , n66492 , n66493 , n66494 , n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , 
     n66501 , n66502 , n66503 , n66504 , n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , 
     n66511 , n66512 , n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , 
     n66521 , n66522 , n66523 , n66524 , n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , 
     n66531 , n66532 , n66533 , n66534 , n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , 
     n66541 , n66542 , n66543 , n66544 , n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , 
     n66551 , n66552 , n66553 , n66554 , n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , 
     n66561 , n66562 , n66563 , n66564 , n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , 
     n66571 , n66572 , n66573 , n66574 , n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , 
     n66581 , n66582 , n66583 , n66584 , n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , 
     n66591 , n66592 , n66593 , n66594 , n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , 
     n66601 , n66602 , n66603 , n66604 , n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , 
     n66611 , n66612 , n66613 , n66614 , n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , 
     n66621 , n66622 , n66623 , n66624 , n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , 
     n66631 , n66632 , n66633 , n66634 , n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , 
     n66641 , n66642 , n66643 , n66644 , n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , 
     n66651 , n66652 , n66653 , n66654 , n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , 
     n66661 , n66662 , n66663 , n66664 , n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , 
     n66671 , n66672 , n66673 , n66674 , n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , 
     n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , 
     n66691 , n66692 , n66693 , n66694 , n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , 
     n66701 , n66702 , n66703 , n66704 , n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , 
     n66711 , n66712 , n66713 , n66714 , n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , 
     n66721 , n66722 , n66723 , n66724 , n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , 
     n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , 
     n66741 , n66742 , n66743 , n66744 , n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , 
     n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , 
     n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , 
     n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , 
     n66781 , n66782 , n66783 , n66784 , n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , 
     n66791 , n66792 , n66793 , n66794 , n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , 
     n66801 , n66802 , n66803 , n66804 , n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , 
     n66811 , n66812 , n66813 , n66814 , n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , 
     n66821 , n66822 , n66823 , n66824 , n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , 
     n66831 , n66832 , n66833 , n66834 , n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , 
     n66841 , n66842 , n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , 
     n66851 , n66852 , n66853 , n66854 , n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , 
     n66861 , n66862 , n66863 , n66864 , n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , 
     n66871 , n66872 , n66873 , n66874 , n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , 
     n66881 , n66882 , n66883 , n66884 , n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , 
     n66891 , n66892 , n66893 , n66894 , n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , 
     n66901 , n66902 , n66903 , n66904 , n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , 
     n66911 , n66912 , n66913 , n66914 , n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , 
     n66921 , n66922 , n66923 , n66924 , n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , 
     n66931 , n66932 , n66933 , n66934 , n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , 
     n66941 , n66942 , n66943 , n66944 , n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , 
     n66951 , n66952 , n66953 , n66954 , n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , 
     n66961 , n66962 , n66963 , n66964 , n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , 
     n66971 , n66972 , n66973 , n66974 , n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , 
     n66981 , n66982 , n66983 , n66984 , n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , 
     n66991 , n66992 , n66993 , n66994 , n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , 
     n67001 , n67002 , n67003 , n67004 , n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , 
     n67011 , n67012 , n67013 , n67014 , n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , 
     n67021 , n67022 , n67023 , n67024 , n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , 
     n67031 , n67032 , n67033 , n67034 , n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , 
     n67041 , n67042 , n67043 , n67044 , n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , 
     n67051 , n67052 , n67053 , n67054 , n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , 
     n67061 , n67062 , n67063 , n67064 , n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , 
     n67071 , n67072 , n67073 , n67074 , n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , 
     n67081 , n67082 , n67083 , n67084 , n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , 
     n67091 , n67092 , n67093 , n67094 , n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , 
     n67101 , n67102 , n67103 , n67104 , n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , 
     n67111 , n67112 , n67113 , n67114 , n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , 
     n67121 , n67122 , n67123 , n67124 , n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , 
     n67131 , n67132 , n67133 , n67134 , n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , 
     n67141 , n67142 , n67143 , n67144 , n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , 
     n67151 , n67152 , n67153 , n67154 , n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , 
     n67161 , n67162 , n67163 , n67164 , n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , 
     n67171 , n67172 , n67173 , n67174 , n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , 
     n67181 , n67182 , n67183 , n67184 , n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , 
     n67191 , n67192 , n67193 , n67194 , n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , 
     n67201 , n67202 , n67203 , n67204 , n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , 
     n67211 , n67212 , n67213 , n67214 , n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , 
     n67221 , n67222 , n67223 , n67224 , n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , 
     n67231 , n67232 , n67233 , n67234 , n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , 
     n67241 , n67242 , n67243 , n67244 , n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , 
     n67251 , n67252 , n67253 , n67254 , n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , 
     n67261 , n67262 , n67263 , n67264 , n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , 
     n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , 
     n67281 , n67282 , n67283 , n67284 , n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , 
     n67291 , n67292 , n67293 , n67294 , n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , 
     n67301 , n67302 , n67303 , n67304 , n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , 
     n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , 
     n67321 , n67322 , n67323 , n67324 , n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , 
     n67331 , n67332 , n67333 , n67334 , n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , 
     n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , 
     n67351 , n67352 , n67353 , n67354 , n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , 
     n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , 
     n67371 , n67372 , n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , 
     n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , 
     n67391 , n67392 , n67393 , n67394 , n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , 
     n67401 , n67402 , n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , 
     n67411 , n67412 , n67413 , n67414 , n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , 
     n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , 
     n67431 , n67432 , n67433 , n67434 , n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , 
     n67441 , n67442 , n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , 
     n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , 
     n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , 
     n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , 
     n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , 
     n67491 , n67492 , n67493 , n67494 , n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , 
     n67501 , n67502 , n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , 
     n67511 , n67512 , n67513 , n67514 , n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , 
     n67521 , n67522 , n67523 , n67524 , n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , 
     n67531 , n67532 , n67533 , n67534 , n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , 
     n67541 , n67542 , n67543 , n67544 , n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , 
     n67551 , n67552 , n67553 , n67554 , n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , 
     n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , 
     n67571 , n67572 , n67573 , n67574 , n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , 
     n67581 , n67582 , n67583 , n67584 , n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , 
     n67591 , n67592 , n67593 , n67594 , n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , 
     n67601 , n67602 , n67603 , n67604 , n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , 
     n67611 , n67612 , n67613 , n67614 , n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , 
     n67621 , n67622 , n67623 , n67624 , n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , 
     n67631 , n67632 , n67633 , n67634 , n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , 
     n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , 
     n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , 
     n67661 , n67662 , n67663 , n67664 , n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , 
     n67671 , n67672 , n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , 
     n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , 
     n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , 
     n67701 , n67702 , n67703 , n67704 , n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , 
     n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , 
     n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , 
     n67731 , n67732 , n67733 , n67734 , n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , 
     n67741 , n67742 , n67743 , n67744 , n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , 
     n67751 , n67752 , n67753 , n67754 , n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , 
     n67761 , n67762 , n67763 , n67764 , n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , 
     n67771 , n67772 , n67773 , n67774 , n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , 
     n67781 , n67782 , n67783 , n67784 , n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , 
     n67791 , n67792 , n67793 , n67794 , n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , 
     n67801 , n67802 , n67803 , n67804 , n67805 , n67806 , n67807 , n67808 , n67809 , n67810 , 
     n67811 , n67812 , n67813 , n67814 , n67815 , n67816 , n67817 , n67818 , n67819 , n67820 , 
     n67821 , n67822 , n67823 , n67824 , n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , 
     n67831 , n67832 , n67833 , n67834 , n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , 
     n67841 , n67842 , n67843 , n67844 , n67845 , n67846 , n67847 , n67848 , n67849 , n67850 , 
     n67851 , n67852 , n67853 , n67854 , n67855 , n67856 , n67857 , n67858 , n67859 , n67860 , 
     n67861 , n67862 , n67863 , n67864 , n67865 , n67866 , n67867 , n67868 , n67869 , n67870 , 
     n67871 , n67872 , n67873 , n67874 , n67875 , n67876 , n67877 , n67878 , n67879 , n67880 , 
     n67881 , n67882 , n67883 , n67884 , n67885 , n67886 , n67887 , n67888 , n67889 , n67890 , 
     n67891 , n67892 , n67893 , n67894 , n67895 , n67896 , n67897 , n67898 , n67899 , n67900 , 
     n67901 , n67902 , n67903 , n67904 , n67905 , n67906 , n67907 , n67908 , n67909 , n67910 , 
     n67911 , n67912 , n67913 , n67914 , n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , 
     n67921 , n67922 , n67923 , n67924 , n67925 , n67926 , n67927 , n67928 , n67929 , n67930 , 
     n67931 , n67932 , n67933 , n67934 , n67935 , n67936 , n67937 , n67938 , n67939 , n67940 , 
     n67941 , n67942 , n67943 , n67944 , n67945 , n67946 , n67947 , n67948 , n67949 , n67950 , 
     n67951 , n67952 , n67953 , n67954 , n67955 , n67956 , n67957 , n67958 , n67959 , n67960 , 
     n67961 , n67962 , n67963 , n67964 , n67965 , n67966 , n67967 , n67968 , n67969 , n67970 , 
     n67971 , n67972 , n67973 , n67974 , n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , 
     n67981 , n67982 , n67983 , n67984 , n67985 , n67986 , n67987 , n67988 , n67989 , n67990 , 
     n67991 , n67992 , n67993 , n67994 , n67995 , n67996 , n67997 , n67998 , n67999 , n68000 , 
     n68001 , n68002 , n68003 , n68004 , n68005 , n68006 , n68007 , n68008 , n68009 , n68010 , 
     n68011 , n68012 , n68013 , n68014 , n68015 , n68016 , n68017 , n68018 , n68019 , n68020 , 
     n68021 , n68022 , n68023 , n68024 , n68025 , n68026 , n68027 , n68028 , n68029 , n68030 , 
     n68031 , n68032 , n68033 , n68034 , n68035 , n68036 , n68037 , n68038 , n68039 , n68040 , 
     n68041 , n68042 , n68043 , n68044 , n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , 
     n68051 , n68052 , n68053 , n68054 , n68055 , n68056 , n68057 , n68058 , n68059 , n68060 , 
     n68061 , n68062 , n68063 , n68064 , n68065 , n68066 , n68067 , n68068 , n68069 , n68070 , 
     n68071 , n68072 , n68073 , n68074 , n68075 , n68076 , n68077 , n68078 , n68079 , n68080 , 
     n68081 , n68082 , n68083 , n68084 , n68085 , n68086 , n68087 , n68088 , n68089 , n68090 , 
     n68091 , n68092 , n68093 , n68094 , n68095 , n68096 , n68097 , n68098 , n68099 , n68100 , 
     n68101 , n68102 , n68103 , n68104 , n68105 , n68106 , n68107 , n68108 , n68109 , n68110 , 
     n68111 , n68112 , n68113 , n68114 , n68115 , n68116 , n68117 , n68118 , n68119 , n68120 , 
     n68121 , n68122 , n68123 , n68124 , n68125 , n68126 , n68127 , n68128 , n68129 , n68130 , 
     n68131 , n68132 , n68133 , n68134 , n68135 , n68136 , n68137 , n68138 , n68139 , n68140 , 
     n68141 , n68142 , n68143 , n68144 , n68145 , n68146 , n68147 , n68148 , n68149 , n68150 , 
     n68151 , n68152 , n68153 , n68154 , n68155 , n68156 , n68157 , n68158 , n68159 , n68160 , 
     n68161 , n68162 , n68163 , n68164 , n68165 , n68166 , n68167 , n68168 , n68169 , n68170 , 
     n68171 , n68172 , n68173 , n68174 , n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , 
     n68181 , n68182 , n68183 , n68184 , n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , 
     n68191 , n68192 , n68193 , n68194 , n68195 , n68196 , n68197 , n68198 , n68199 , n68200 , 
     n68201 , n68202 , n68203 , n68204 , n68205 , n68206 , n68207 , n68208 , n68209 , n68210 , 
     n68211 , n68212 , n68213 , n68214 , n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , 
     n68221 , n68222 , n68223 , n68224 , n68225 , n68226 , n68227 , n68228 , n68229 , n68230 , 
     n68231 , n68232 , n68233 , n68234 , n68235 , n68236 , n68237 , n68238 , n68239 , n68240 , 
     n68241 , n68242 , n68243 , n68244 , n68245 , n68246 , n68247 , n68248 , n68249 , n68250 , 
     n68251 , n68252 , n68253 , n68254 , n68255 , n68256 , n68257 , n68258 , n68259 , n68260 , 
     n68261 , n68262 , n68263 , n68264 , n68265 , n68266 , n68267 , n68268 , n68269 , n68270 , 
     n68271 , n68272 , n68273 , n68274 , n68275 , n68276 , n68277 , n68278 , n68279 , n68280 , 
     n68281 , n68282 , n68283 , n68284 , n68285 , n68286 , n68287 , n68288 , n68289 , n68290 , 
     n68291 , n68292 , n68293 , n68294 , n68295 , n68296 , n68297 , n68298 , n68299 , n68300 , 
     n68301 , n68302 , n68303 , n68304 , n68305 , n68306 , n68307 , n68308 , n68309 , n68310 , 
     n68311 , n68312 , n68313 , n68314 , n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , 
     n68321 , n68322 , n68323 , n68324 , n68325 , n68326 , n68327 , n68328 , n68329 , n68330 , 
     n68331 , n68332 , n68333 , n68334 , n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , 
     n68341 , n68342 , n68343 , n68344 , n68345 , n68346 , n68347 , n68348 , n68349 , n68350 , 
     n68351 , n68352 , n68353 , n68354 , n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , 
     n68361 , n68362 , n68363 , n68364 , n68365 , n68366 , n68367 , n68368 , n68369 , n68370 , 
     n68371 , n68372 , n68373 , n68374 , n68375 , n68376 , n68377 , n68378 , n68379 , n68380 , 
     n68381 , n68382 , n68383 , n68384 , n68385 , n68386 , n68387 , n68388 , n68389 , n68390 , 
     n68391 , n68392 , n68393 , n68394 , n68395 , n68396 , n68397 , n68398 , n68399 , n68400 , 
     n68401 , n68402 , n68403 , n68404 , n68405 , n68406 , n68407 , n68408 , n68409 , n68410 , 
     n68411 , n68412 , n68413 , n68414 , n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , 
     n68421 , n68422 , n68423 , n68424 , n68425 , n68426 , n68427 , n68428 , n68429 , n68430 , 
     n68431 , n68432 , n68433 , n68434 , n68435 , n68436 , n68437 , n68438 , n68439 , n68440 , 
     n68441 , n68442 , n68443 , n68444 , n68445 , n68446 , n68447 , n68448 , n68449 , n68450 , 
     n68451 , n68452 , n68453 , n68454 , n68455 , n68456 , n68457 , n68458 , n68459 , n68460 , 
     n68461 , n68462 , n68463 , n68464 , n68465 , n68466 , n68467 , n68468 , n68469 , n68470 , 
     n68471 , n68472 , n68473 , n68474 , n68475 , n68476 , n68477 , n68478 , n68479 , n68480 , 
     n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , n68487 , n68488 , n68489 , n68490 , 
     n68491 , n68492 , n68493 , n68494 , n68495 , n68496 , n68497 , n68498 , n68499 , n68500 , 
     n68501 , n68502 , n68503 , n68504 , n68505 , n68506 , n68507 , n68508 , n68509 , n68510 , 
     n68511 , n68512 , n68513 , n68514 , n68515 , n68516 , n68517 , n68518 , n68519 , n68520 , 
     n68521 , n68522 , n68523 , n68524 , n68525 , n68526 , n68527 , n68528 , n68529 , n68530 , 
     n68531 , n68532 , n68533 , n68534 , n68535 , n68536 , n68537 , n68538 , n68539 , n68540 , 
     n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , n68547 , n68548 , n68549 , n68550 , 
     n68551 , n68552 , n68553 , n68554 , n68555 , n68556 , n68557 , n68558 , n68559 , n68560 , 
     n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , n68567 , n68568 , n68569 , n68570 , 
     n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , n68579 , n68580 , 
     n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , n68587 , n68588 , n68589 , n68590 , 
     n68591 , n68592 , n68593 , n68594 , n68595 , n68596 , n68597 , n68598 , n68599 , n68600 , 
     n68601 , n68602 , n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , n68609 , n68610 , 
     n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , n68619 , n68620 , 
     n68621 , n68622 , n68623 , n68624 , n68625 , n68626 , n68627 , n68628 , n68629 , n68630 , 
     n68631 , n68632 , n68633 , n68634 , n68635 , n68636 , n68637 , n68638 , n68639 , n68640 , 
     n68641 , n68642 , n68643 , n68644 , n68645 , n68646 , n68647 , n68648 , n68649 , n68650 , 
     n68651 , n68652 , n68653 , n68654 , n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , 
     n68661 , n68662 , n68663 , n68664 , n68665 , n68666 , n68667 , n68668 , n68669 , n68670 , 
     n68671 , n68672 , n68673 , n68674 , n68675 , n68676 , n68677 , n68678 , n68679 , n68680 , 
     n68681 , n68682 , n68683 , n68684 , n68685 , n68686 , n68687 , n68688 , n68689 , n68690 , 
     n68691 , n68692 , n68693 , n68694 , n68695 , n68696 , n68697 , n68698 , n68699 , n68700 , 
     n68701 , n68702 , n68703 , n68704 , n68705 , n68706 , n68707 , n68708 , n68709 , n68710 , 
     n68711 , n68712 , n68713 , n68714 , n68715 , n68716 , n68717 , n68718 , n68719 , n68720 , 
     n68721 , n68722 , n68723 , n68724 , n68725 , n68726 , n68727 , n68728 , n68729 , n68730 , 
     n68731 , n68732 , n68733 , n68734 , n68735 , n68736 , n68737 , n68738 , n68739 , n68740 , 
     n68741 , n68742 , n68743 , n68744 , n68745 , n68746 , n68747 , n68748 , n68749 , n68750 , 
     n68751 , n68752 , n68753 , n68754 , n68755 , n68756 , n68757 , n68758 , n68759 , n68760 , 
     n68761 , n68762 , n68763 , n68764 , n68765 , n68766 , n68767 , n68768 , n68769 , n68770 , 
     n68771 , n68772 , n68773 , n68774 , n68775 , n68776 , n68777 , n68778 , n68779 , n68780 , 
     n68781 , n68782 , n68783 , n68784 , n68785 , n68786 , n68787 , n68788 , n68789 , n68790 , 
     n68791 , n68792 , n68793 , n68794 , n68795 , n68796 , n68797 , n68798 , n68799 , n68800 , 
     n68801 , n68802 , n68803 , n68804 , n68805 , n68806 , n68807 , n68808 , n68809 , n68810 , 
     n68811 , n68812 , n68813 , n68814 , n68815 , n68816 , n68817 , n68818 , n68819 , n68820 , 
     n68821 , n68822 , n68823 , n68824 , n68825 , n68826 , n68827 , n68828 , n68829 , n68830 , 
     n68831 , n68832 , n68833 , n68834 , n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , 
     n68841 , n68842 , n68843 , n68844 , n68845 , n68846 , n68847 , n68848 , n68849 , n68850 , 
     n68851 , n68852 , n68853 , n68854 , n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , 
     n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , n68867 , n68868 , n68869 , n68870 , 
     n68871 , n68872 , n68873 , n68874 , n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , 
     n68881 , n68882 , n68883 , n68884 , n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , 
     n68891 , n68892 , n68893 , n68894 , n68895 , n68896 , n68897 , n68898 , n68899 , n68900 , 
     n68901 , n68902 , n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , 
     n68911 , n68912 , n68913 , n68914 , n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , 
     n68921 , n68922 , n68923 , n68924 , n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , 
     n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , 
     n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , 
     n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , 
     n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , 
     n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , 
     n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , 
     n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , 
     n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , 
     n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , 
     n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , 
     n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , 
     n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , 
     n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , 
     n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , 
     n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , 
     n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , 
     n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , 
     n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , 
     n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , 
     n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , 
     n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , n69139 , n69140 , 
     n69141 , n69142 , n69143 , n69144 , n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , 
     n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , 
     n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , 
     n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , 
     n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , 
     n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , n69197 , n69198 , n69199 , n69200 , 
     n69201 , n69202 , n69203 , n69204 , n69205 , n69206 , n69207 , n69208 , n69209 , n69210 , 
     n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , 
     n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , 
     n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , 
     n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , 
     n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , 
     n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , 
     n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , 
     n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , 
     n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , 
     n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , 
     n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , 
     n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , 
     n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , 
     n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , 
     n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , 
     n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , 
     n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , 
     n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , 
     n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , 
     n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , 
     n69411 , n69412 , n69413 , n69414 , n69415 , n69416 , n69417 , n69418 , n69419 , n69420 , 
     n69421 , n69422 , n69423 , n69424 , n69425 , n69426 , n69427 , n69428 , n69429 , n69430 , 
     n69431 , n69432 , n69433 , n69434 , n69435 , n69436 , n69437 , n69438 , n69439 , n69440 , 
     n69441 , n69442 , n69443 , n69444 , n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , 
     n69451 , n69452 , n69453 , n69454 , n69455 , n69456 , n69457 , n69458 , n69459 , n69460 , 
     n69461 , n69462 , n69463 , n69464 , n69465 , n69466 , n69467 , n69468 , n69469 , n69470 , 
     n69471 , n69472 , n69473 , n69474 , n69475 , n69476 , n69477 , n69478 , n69479 , n69480 , 
     n69481 , n69482 , n69483 , n69484 , n69485 , n69486 , n69487 , n69488 , n69489 , n69490 , 
     n69491 , n69492 , n69493 , n69494 , n69495 , n69496 , n69497 , n69498 , n69499 , n69500 , 
     n69501 , n69502 , n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , 
     n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , 
     n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , 
     n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , 
     n69541 , n69542 , n69543 , n69544 , n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , 
     n69551 , n69552 , n69553 , n69554 , n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , 
     n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , 
     n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , 
     n69581 , n69582 , n69583 , n69584 , n69585 , n69586 , n69587 , n69588 , n69589 , n69590 , 
     n69591 , n69592 , n69593 , n69594 , n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , 
     n69601 , n69602 , n69603 , n69604 , n69605 , n69606 , n69607 , n69608 , n69609 , n69610 , 
     n69611 , n69612 , n69613 , n69614 , n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , 
     n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , 
     n69631 , n69632 , n69633 , n69634 , n69635 , n69636 , n69637 , n69638 , n69639 , n69640 , 
     n69641 , n69642 , n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , n69649 , n69650 , 
     n69651 , n69652 , n69653 , n69654 , n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , 
     n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , n69667 , n69668 , n69669 , n69670 , 
     n69671 , n69672 , n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , 
     n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , 
     n69691 , n69692 , n69693 , n69694 , n69695 , n69696 , n69697 , n69698 , n69699 , n69700 , 
     n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , 
     n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n69719 , n69720 , 
     n69721 , n69722 , n69723 , n69724 , n69725 , n69726 , n69727 , n69728 , n69729 , n69730 , 
     n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , 
     n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , 
     n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , n69759 , n69760 , 
     n69761 , n69762 , n69763 , n69764 , n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , 
     n69771 , n69772 , n69773 , n69774 , n69775 , n69776 , n69777 , n69778 , n69779 , n69780 , 
     n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , 
     n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , 
     n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , 
     n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , 
     n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , 
     n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , 
     n69841 , n69842 , n69843 , n69844 , n69845 , n69846 , n69847 , n69848 , n69849 , n69850 , 
     n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , n69859 , n69860 , 
     n69861 , n69862 , n69863 , n69864 , n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , 
     n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , 
     n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , 
     n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , 
     n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , n69909 , n69910 , 
     n69911 , n69912 , n69913 , n69914 , n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , 
     n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , 
     n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , n69937 , n69938 , n69939 , n69940 , 
     n69941 , n69942 , n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , 
     n69951 , n69952 , n69953 , n69954 , n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , 
     n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , 
     n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , 
     n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , 
     n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , 
     n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , 
     n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , 
     n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , 
     n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , 
     n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , 
     n70051 , n70052 , n70053 , n70054 , n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , 
     n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , 
     n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , 
     n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , 
     n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , 
     n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , 
     n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , 
     n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , 
     n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , 
     n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , 
     n70151 , n70152 , n70153 , n70154 , n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , 
     n70161 , n70162 , n70163 , n70164 , n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , 
     n70171 , n70172 , n70173 , n70174 , n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , 
     n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , 
     n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , 
     n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , 
     n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , 
     n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , 
     n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , 
     n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , 
     n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , 
     n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , 
     n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , 
     n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , 
     n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , 
     n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , 
     n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , 
     n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , 
     n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , 
     n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , 
     n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , 
     n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , 
     n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , 
     n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , 
     n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , 
     n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , 
     n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , 
     n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , 
     n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , 
     n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , 
     n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , 
     n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , 
     n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , 
     n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , 
     n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , 
     n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , 
     n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , 
     n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , 
     n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , 
     n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , 
     n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , 
     n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , 
     n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , 
     n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , 
     n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , 
     n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , 
     n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , 
     n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , 
     n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , 
     n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , 
     n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , 
     n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , 
     n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , 
     n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , 
     n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , 
     n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , 
     n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , 
     n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , 
     n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , 
     n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , 
     n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , 
     n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , 
     n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , 
     n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , 
     n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , 
     n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , 
     n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , 
     n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , 
     n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , 
     n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , 
     n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , 
     n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , 
     n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , 
     n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , 
     n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , 
     n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , n70909 , n70910 , 
     n70911 , n70912 , n70913 , n70914 , n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , 
     n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , 
     n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , 
     n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , 
     n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , 
     n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , 
     n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , 
     n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , 
     n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , 
     n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , 
     n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , n71019 , n71020 , 
     n71021 , n71022 , n71023 , n71024 , n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , 
     n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , 
     n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , 
     n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , 
     n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , 
     n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , 
     n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , 
     n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , 
     n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , 
     n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , 
     n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , 
     n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , 
     n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , 
     n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , 
     n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , 
     n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , 
     n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , 
     n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , 
     n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , n71209 , n71210 , 
     n71211 , n71212 , n71213 , n71214 , n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , 
     n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , 
     n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , 
     n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , 
     n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , 
     n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , n71267 , n71268 , n71269 , n71270 , 
     n71271 , n71272 , n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , 
     n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , 
     n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , 
     n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , 
     n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , 
     n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , 
     n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , 
     n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , 
     n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , 
     n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , 
     n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , 
     n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , 
     n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , 
     n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , 
     n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , 
     n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , 
     n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , n71439 , n71440 , 
     n71441 , n71442 , n71443 , n71444 , n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , 
     n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , 
     n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , 
     n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , 
     n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , 
     n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , 
     n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , 
     n71511 , n71512 , n71513 , n71514 , n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , 
     n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , 
     n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , 
     n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , 
     n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , 
     n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , 
     n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , 
     n71581 , n71582 , n71583 , n71584 , n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , 
     n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , 
     n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , 
     n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , 
     n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , 
     n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , 
     n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , 
     n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , 
     n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , 
     n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , 
     n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , 
     n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , 
     n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , 
     n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , 
     n71721 , n71722 , n71723 , n71724 , n71725 , n71726 , n71727 , n71728 , n71729 , n71730 , 
     n71731 , n71732 , n71733 , n71734 , n71735 , n71736 , n71737 , n71738 , n71739 , n71740 , 
     n71741 , n71742 , n71743 , n71744 , n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , 
     n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , 
     n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , n71769 , n71770 , 
     n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , 
     n71781 , n71782 , n71783 , n71784 , n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , 
     n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , 
     n71801 , n71802 , n71803 , n71804 , n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , 
     n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , n71819 , n71820 , 
     n71821 , n71822 , n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , 
     n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , n71839 , n71840 , 
     n71841 , n71842 , n71843 , n71844 , n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , 
     n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , 
     n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , 
     n71871 , n71872 , n71873 , n71874 , n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , 
     n71881 , n71882 , n71883 , n71884 , n71885 , n71886 , n71887 , n71888 , n71889 , n71890 , 
     n71891 , n71892 , n71893 , n71894 , n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , 
     n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , 
     n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , 
     n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , 
     n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , 
     n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , 
     n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , 
     n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , 
     n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , 
     n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , 
     n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , 
     n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , 
     n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , 
     n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , n72028 , n72029 , n72030 , 
     n72031 , n72032 , n72033 , n72034 , n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , 
     n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , 
     n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , 
     n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , 
     n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , 
     n72081 , n72082 , n72083 , n72084 , n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , 
     n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , 
     n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , 
     n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , 
     n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , 
     n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , 
     n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , 
     n72151 , n72152 , n72153 , n72154 , n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , 
     n72161 , n72162 , n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , 
     n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , 
     n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , 
     n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , 
     n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , 
     n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , n72217 , n72218 , n72219 , n72220 , 
     n72221 , n72222 , n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , 
     n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , 
     n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , 
     n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , 
     n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , 
     n72271 , n72272 , n72273 , n72274 , n72275 , n72276 , n72277 , n72278 , n72279 , n72280 , 
     n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , 
     n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , 
     n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , 
     n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , 
     n72321 , n72322 , n72323 , n72324 , n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , 
     n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , 
     n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , 
     n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , 
     n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , 
     n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , 
     n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , 
     n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , 
     n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , 
     n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , 
     n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , 
     n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , 
     n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , 
     n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , 
     n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , 
     n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , 
     n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , 
     n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , 
     n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , 
     n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , 
     n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , 
     n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , 
     n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , 
     n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , 
     n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , 
     n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , 
     n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , 
     n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , 
     n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , 
     n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , 
     n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , 
     n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , 
     n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , 
     n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , 
     n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , 
     n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , 
     n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , 
     n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , 
     n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , 
     n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , 
     n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , 
     n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , 
     n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , 
     n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , 
     n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , 
     n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , 
     n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , 
     n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , 
     n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , 
     n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , 
     n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , 
     n72831 , n72832 , n72833 , n72834 , n72835 , n72836 , n72837 , n72838 , n72839 , n72840 , 
     n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , 
     n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , 
     n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , 
     n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , 
     n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , 
     n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , 
     n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , 
     n72911 , n72912 , n72913 , n72914 , n72915 , n72916 , n72917 , n72918 , n72919 , n72920 , 
     n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , 
     n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , 
     n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , 
     n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , 
     n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , 
     n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , 
     n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , 
     n72991 , n72992 , n72993 , n72994 , n72995 , n72996 , n72997 , n72998 , n72999 , n73000 , 
     n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , 
     n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , 
     n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , 
     n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , 
     n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , 
     n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , 
     n73061 , n73062 , n73063 , n73064 , n73065 , n73066 , n73067 , n73068 , n73069 , n73070 , 
     n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , 
     n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , 
     n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , 
     n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , 
     n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , 
     n73121 , n73122 , n73123 , n73124 , n73125 , n73126 , n73127 , n73128 , n73129 , n73130 , 
     n73131 , n73132 , n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , 
     n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , 
     n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , 
     n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , 
     n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , 
     n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , 
     n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , 
     n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , 
     n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , 
     n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , 
     n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , 
     n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , 
     n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , 
     n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , 
     n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , n73277 , n73278 , n73279 , n73280 , 
     n73281 , n73282 , n73283 , n73284 , n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , 
     n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , 
     n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , 
     n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , 
     n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , 
     n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , 
     n73341 , n73342 , n73343 , n73344 , n73345 , n73346 , n73347 , n73348 , n73349 , n73350 , 
     n73351 , n73352 , n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , 
     n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , 
     n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , 
     n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , 
     n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , 
     n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , 
     n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , 
     n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , 
     n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , 
     n73441 , n73442 , n73443 , n73444 , n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , 
     n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , 
     n73461 , n73462 , n73463 , n73464 , n73465 , n73466 , n73467 , n73468 , n73469 , n73470 , 
     n73471 , n73472 , n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , 
     n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , n73489 , n73490 , 
     n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , 
     n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , 
     n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , 
     n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , n73527 , n73528 , n73529 , n73530 , 
     n73531 , n73532 , n73533 , n73534 , n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , 
     n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , 
     n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , 
     n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , 
     n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , 
     n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , 
     n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , 
     n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , 
     n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , 
     n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , 
     n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , 
     n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , 
     n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , 
     n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , 
     n73671 , n73672 , n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , 
     n73681 , n73682 , n73683 , n73684 , n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , 
     n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , 
     n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , 
     n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , 
     n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , 
     n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , 
     n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , 
     n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , n73757 , n73758 , n73759 , n73760 , 
     n73761 , n73762 , n73763 , n73764 , n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , 
     n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , n73779 , n73780 , 
     n73781 , n73782 , n73783 , n73784 , n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , 
     n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , 
     n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , 
     n73811 , n73812 , n73813 , n73814 , n73815 , n73816 , n73817 , n73818 , n73819 , n73820 , 
     n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , 
     n73831 , n73832 , n73833 , n73834 , n73835 , n73836 , n73837 , n73838 , n73839 , n73840 , 
     n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , 
     n73851 , n73852 , n73853 , n73854 , n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , 
     n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , 
     n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , 
     n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , n73887 , n73888 , n73889 , n73890 , 
     n73891 , n73892 , n73893 , n73894 , n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , 
     n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , 
     n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , 
     n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , 
     n73931 , n73932 , n73933 , n73934 , n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , 
     n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , 
     n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , 
     n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , n73967 , n73968 , n73969 , n73970 , 
     n73971 , n73972 , n73973 , n73974 , n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , 
     n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , 
     n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , 
     n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , 
     n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , 
     n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , 
     n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , 
     n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , 
     n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , n74059 , n74060 , 
     n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , 
     n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , n74079 , n74080 , 
     n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , 
     n74091 , n74092 , n74093 , n74094 , n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , 
     n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , n74109 , n74110 , 
     n74111 , n74112 , n74113 , n74114 , n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , 
     n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , n74127 , n74128 , n74129 , n74130 , 
     n74131 , n74132 , n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , 
     n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , n74149 , n74150 , 
     n74151 , n74152 , n74153 , n74154 , n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , 
     n74161 , n74162 , n74163 , n74164 , n74165 , n74166 , n74167 , n74168 , n74169 , n74170 , 
     n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , 
     n74181 , n74182 , n74183 , n74184 , n74185 , n74186 , n74187 , n74188 , n74189 , n74190 , 
     n74191 , n74192 , n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , 
     n74201 , n74202 , n74203 , n74204 , n74205 , n74206 , n74207 , n74208 , n74209 , n74210 , 
     n74211 , n74212 , n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , 
     n74221 , n74222 , n74223 , n74224 , n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , 
     n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , 
     n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , 
     n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , 
     n74261 , n74262 , n74263 , n74264 , n74265 , n74266 , n74267 , n74268 , n74269 , n74270 , 
     n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , 
     n74281 , n74282 , n74283 , n74284 , n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , 
     n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , 
     n74301 , n74302 , n74303 , n74304 , n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , 
     n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , 
     n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , 
     n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , n74337 , n74338 , n74339 , n74340 , 
     n74341 , n74342 , n74343 , n74344 , n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , 
     n74351 , n74352 , n74353 , n74354 , n74355 , n74356 , n74357 , n74358 , n74359 , n74360 , 
     n74361 , n74362 , n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , 
     n74371 , n74372 , n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , n74379 , n74380 , 
     n74381 , n74382 , n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , 
     n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , 
     n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , 
     n74411 , n74412 , n74413 , n74414 , n74415 , n74416 , n74417 , n74418 , n74419 , n74420 , 
     n74421 , n74422 , n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , 
     n74431 , n74432 , n74433 , n74434 , n74435 , n74436 , n74437 , n74438 , n74439 , n74440 , 
     n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , n74449 , n74450 , 
     n74451 , n74452 , n74453 , n74454 , n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , 
     n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , 
     n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , 
     n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , 
     n74491 , n74492 , n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , 
     n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , 
     n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , 
     n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , 
     n74531 , n74532 , n74533 , n74534 , n74535 , n74536 , n74537 , n74538 , n74539 , n74540 , 
     n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , 
     n74551 , n74552 , n74553 , n74554 , n74555 , n74556 , n74557 , n74558 , n74559 , n74560 , 
     n74561 , n74562 , n74563 , n74564 , n74565 , n74566 , n74567 , n74568 , n74569 , n74570 , 
     n74571 , n74572 , n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , n74579 , n74580 , 
     n74581 , n74582 , n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , 
     n74591 , n74592 , n74593 , n74594 , n74595 , n74596 , n74597 , n74598 , n74599 , n74600 , 
     n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , 
     n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , 
     n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , 
     n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , n74637 , n74638 , n74639 , n74640 , 
     n74641 , n74642 , n74643 , n74644 , n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , 
     n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , n74657 , n74658 , n74659 , n74660 , 
     n74661 , n74662 , n74663 , n74664 , n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , 
     n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , n74677 , n74678 , n74679 , n74680 , 
     n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , 
     n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , 
     n74701 , n74702 , n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , 
     n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n74719 , n74720 , 
     n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , 
     n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , 
     n74741 , n74742 , n74743 , n74744 , n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , 
     n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , n74759 , n74760 , 
     n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , 
     n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , n74777 , n74778 , n74779 , n74780 , 
     n74781 , n74782 , n74783 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , 
     n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , n74799 , n74800 , 
     n74801 , n74802 , n74803 , n74804 , n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , 
     n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , n74819 , n74820 , 
     n74821 , n74822 , n74823 , n74824 , n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , 
     n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , 
     n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , 
     n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , n74859 , n74860 , 
     n74861 , n74862 , n74863 , n74864 , n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , 
     n74871 , n74872 , n74873 , n74874 , n74875 , n74876 , n74877 , n74878 , n74879 , n74880 , 
     n74881 , n74882 , n74883 , n74884 , n74885 , n74886 , n74887 , n74888 , n74889 , n74890 , 
     n74891 , n74892 , n74893 , n74894 , n74895 , n74896 , n74897 , n74898 , n74899 , n74900 , 
     n74901 , n74902 , n74903 , n74904 , n74905 , n74906 , n74907 , n74908 , n74909 , n74910 , 
     n74911 , n74912 , n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , 
     n74921 , n74922 , n74923 , n74924 , n74925 , n74926 , n74927 , n74928 , n74929 , n74930 , 
     n74931 , n74932 , n74933 , n74934 , n74935 , n74936 , n74937 , n74938 , n74939 , n74940 , 
     n74941 , n74942 , n74943 , n74944 , n74945 , n74946 , n74947 , n74948 , n74949 , n74950 , 
     n74951 , n74952 , n74953 , n74954 , n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , 
     n74961 , n74962 , n74963 , n74964 , n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , 
     n74971 , n74972 , n74973 , n74974 , n74975 , n74976 , n74977 , n74978 , n74979 , n74980 , 
     n74981 , n74982 , n74983 , n74984 , n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , 
     n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , n74997 , n74998 , n74999 , n75000 , 
     n75001 , n75002 , n75003 , n75004 , n75005 , n75006 , n75007 , n75008 , n75009 , n75010 , 
     n75011 , n75012 , n75013 , n75014 , n75015 , n75016 , n75017 , n75018 , n75019 , n75020 , 
     n75021 , n75022 , n75023 , n75024 , n75025 , n75026 , n75027 , n75028 , n75029 , n75030 , 
     n75031 , n75032 , n75033 , n75034 , n75035 , n75036 , n75037 , n75038 , n75039 , n75040 , 
     n75041 , n75042 , n75043 , n75044 , n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , 
     n75051 , n75052 , n75053 , n75054 , n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , 
     n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , 
     n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n75077 , n75078 , n75079 , n75080 , 
     n75081 , n75082 , n75083 , n75084 , n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , 
     n75091 , n75092 , n75093 , n75094 , n75095 , n75096 , n75097 , n75098 , n75099 , n75100 , 
     n75101 , n75102 , n75103 , n75104 , n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , 
     n75111 , n75112 , n75113 , n75114 , n75115 , n75116 , n75117 , n75118 , n75119 , n75120 , 
     n75121 , n75122 , n75123 , n75124 , n75125 , n75126 , n75127 , n75128 , n75129 , n75130 , 
     n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , 
     n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , 
     n75151 , n75152 , n75153 , n75154 , n75155 , n75156 , n75157 , n75158 , n75159 , n75160 , 
     n75161 , n75162 , n75163 , n75164 , n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , 
     n75171 , n75172 , n75173 , n75174 , n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , 
     n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , 
     n75191 , n75192 , n75193 , n75194 , n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , 
     n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , 
     n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , 
     n75221 , n75222 , n75223 , n75224 , n75225 , n75226 , n75227 , n75228 , n75229 , n75230 , 
     n75231 , n75232 , n75233 , n75234 , n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , 
     n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , 
     n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , 
     n75261 , n75262 , n75263 , n75264 , n75265 , n75266 , n75267 , n75268 , n75269 , n75270 , 
     n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , 
     n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , 
     n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , 
     n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , 
     n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , 
     n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , 
     n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , 
     n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , 
     n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , 
     n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , 
     n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , 
     n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , 
     n75391 , n75392 , n75393 , n75394 , n75395 , n75396 , n75397 , n75398 , n75399 , n75400 , 
     n75401 , n75402 , n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , 
     n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , 
     n75421 , n75422 , n75423 , n75424 , n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , 
     n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , 
     n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , 
     n75451 , n75452 , n75453 , n75454 , n75455 , n75456 , n75457 , n75458 , n75459 , n75460 , 
     n75461 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , 
     n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , 
     n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , 
     n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , 
     n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , 
     n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , 
     n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , 
     n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , 
     n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , 
     n75551 , n75552 , n75553 , n75554 , n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , 
     n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , 
     n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , 
     n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , 
     n75591 , n75592 , n75593 , n75594 , n75595 , n75596 , n75597 , n75598 , n75599 , n75600 , 
     n75601 , n75602 , n75603 , n75604 , n75605 , n75606 , n75607 , n75608 , n75609 , n75610 , 
     n75611 , n75612 , n75613 , n75614 , n75615 , n75616 , n75617 , n75618 , n75619 , n75620 , 
     n75621 , n75622 , n75623 , n75624 , n75625 , n75626 , n75627 , n75628 , n75629 , n75630 , 
     n75631 , n75632 , n75633 , n75634 , n75635 , n75636 , n75637 , n75638 , n75639 , n75640 , 
     n75641 , n75642 , n75643 , n75644 , n75645 , n75646 , n75647 , n75648 , n75649 , n75650 , 
     n75651 , n75652 , n75653 , n75654 , n75655 , n75656 , n75657 , n75658 , n75659 , n75660 , 
     n75661 , n75662 , n75663 , n75664 , n75665 , n75666 , n75667 , n75668 , n75669 , n75670 , 
     n75671 , n75672 , n75673 , n75674 , n75675 , n75676 , n75677 , n75678 , n75679 , n75680 , 
     n75681 , n75682 , n75683 , n75684 , n75685 , n75686 , n75687 , n75688 , n75689 , n75690 , 
     n75691 , n75692 , n75693 , n75694 , n75695 , n75696 , n75697 , n75698 , n75699 , n75700 , 
     n75701 , n75702 , n75703 , n75704 , n75705 , n75706 , n75707 , n75708 , n75709 , n75710 , 
     n75711 , n75712 , n75713 , n75714 , n75715 , n75716 , n75717 , n75718 , n75719 , n75720 , 
     n75721 , n75722 , n75723 , n75724 , n75725 , n75726 , n75727 , n75728 , n75729 , n75730 , 
     n75731 , n75732 , n75733 , n75734 , n75735 , n75736 , n75737 , n75738 , n75739 , n75740 , 
     n75741 , n75742 , n75743 , n75744 , n75745 , n75746 , n75747 , n75748 , n75749 , n75750 , 
     n75751 , n75752 , n75753 , n75754 , n75755 , n75756 , n75757 , n75758 , n75759 , n75760 , 
     n75761 , n75762 , n75763 , n75764 , n75765 , n75766 , n75767 , n75768 , n75769 , n75770 , 
     n75771 , n75772 , n75773 , n75774 , n75775 , n75776 , n75777 , n75778 , n75779 , n75780 , 
     n75781 , n75782 , n75783 , n75784 , n75785 , n75786 , n75787 , n75788 , n75789 , n75790 , 
     n75791 , n75792 , n75793 , n75794 , n75795 , n75796 , n75797 , n75798 , n75799 , n75800 , 
     n75801 , n75802 , n75803 , n75804 , n75805 , n75806 , n75807 , n75808 , n75809 , n75810 , 
     n75811 , n75812 , n75813 , n75814 , n75815 , n75816 , n75817 , n75818 , n75819 , n75820 , 
     n75821 , n75822 , n75823 , n75824 , n75825 , n75826 , n75827 , n75828 , n75829 , n75830 , 
     n75831 , n75832 , n75833 , n75834 , n75835 , n75836 , n75837 , n75838 , n75839 , n75840 , 
     n75841 , n75842 , n75843 , n75844 , n75845 , n75846 , n75847 , n75848 , n75849 , n75850 , 
     n75851 , n75852 , n75853 , n75854 , n75855 , n75856 , n75857 , n75858 , n75859 , n75860 , 
     n75861 , n75862 , n75863 , n75864 , n75865 , n75866 , n75867 , n75868 , n75869 , n75870 , 
     n75871 , n75872 , n75873 , n75874 , n75875 , n75876 , n75877 , n75878 , n75879 , n75880 , 
     n75881 , n75882 , n75883 , n75884 , n75885 , n75886 , n75887 , n75888 , n75889 , n75890 , 
     n75891 , n75892 , n75893 , n75894 , n75895 , n75896 , n75897 , n75898 , n75899 , n75900 , 
     n75901 , n75902 , n75903 , n75904 , n75905 , n75906 , n75907 , n75908 , n75909 , n75910 , 
     n75911 , n75912 , n75913 , n75914 , n75915 , n75916 , n75917 , n75918 , n75919 , n75920 , 
     n75921 , n75922 , n75923 , n75924 , n75925 , n75926 , n75927 , n75928 , n75929 , n75930 , 
     n75931 , n75932 , n75933 , n75934 , n75935 , n75936 , n75937 , n75938 , n75939 , n75940 , 
     n75941 , n75942 , n75943 , n75944 , n75945 , n75946 , n75947 , n75948 , n75949 , n75950 , 
     n75951 , n75952 , n75953 , n75954 , n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , 
     n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , n75969 , n75970 , 
     n75971 , n75972 , n75973 , n75974 , n75975 , n75976 , n75977 , n75978 , n75979 , n75980 , 
     n75981 , n75982 , n75983 , n75984 , n75985 , n75986 , n75987 , n75988 , n75989 , n75990 , 
     n75991 , n75992 , n75993 , n75994 , n75995 , n75996 , n75997 , n75998 , n75999 , n76000 , 
     n76001 , n76002 , n76003 , n76004 , n76005 , n76006 , n76007 , n76008 , n76009 , n76010 , 
     n76011 , n76012 , n76013 , n76014 , n76015 , n76016 , n76017 , n76018 , n76019 , n76020 , 
     n76021 , n76022 , n76023 , n76024 , n76025 , n76026 , n76027 , n76028 , n76029 , n76030 , 
     n76031 , n76032 , n76033 , n76034 , n76035 , n76036 , n76037 , n76038 , n76039 , n76040 , 
     n76041 , n76042 , n76043 , n76044 , n76045 , n76046 , n76047 , n76048 , n76049 , n76050 , 
     n76051 , n76052 , n76053 , n76054 , n76055 , n76056 , n76057 , n76058 , n76059 , n76060 , 
     n76061 , n76062 , n76063 , n76064 , n76065 , n76066 , n76067 , n76068 , n76069 , n76070 , 
     n76071 , n76072 , n76073 , n76074 , n76075 , n76076 , n76077 , n76078 , n76079 , n76080 , 
     n76081 , n76082 , n76083 , n76084 , n76085 , n76086 , n76087 , n76088 , n76089 , n76090 , 
     n76091 , n76092 , n76093 , n76094 , n76095 , n76096 , n76097 , n76098 , n76099 , n76100 , 
     n76101 , n76102 , n76103 , n76104 , n76105 , n76106 , n76107 , n76108 , n76109 , n76110 , 
     n76111 , n76112 , n76113 , n76114 , n76115 , n76116 , n76117 , n76118 , n76119 , n76120 , 
     n76121 , n76122 , n76123 , n76124 , n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , 
     n76131 , n76132 , n76133 , n76134 , n76135 , n76136 , n76137 , n76138 , n76139 , n76140 , 
     n76141 , n76142 , n76143 , n76144 , n76145 , n76146 , n76147 , n76148 , n76149 , n76150 , 
     n76151 , n76152 , n76153 , n76154 , n76155 , n76156 , n76157 , n76158 , n76159 , n76160 , 
     n76161 , n76162 , n76163 , n76164 , n76165 , n76166 , n76167 , n76168 , n76169 , n76170 , 
     n76171 , n76172 , n76173 , n76174 , n76175 , n76176 , n76177 , n76178 , n76179 , n76180 , 
     n76181 , n76182 , n76183 , n76184 , n76185 , n76186 , n76187 , n76188 , n76189 , n76190 , 
     n76191 , n76192 , n76193 , n76194 , n76195 , n76196 , n76197 , n76198 , n76199 , n76200 , 
     n76201 , n76202 , n76203 , n76204 , n76205 , n76206 , n76207 , n76208 , n76209 , n76210 , 
     n76211 , n76212 , n76213 , n76214 , n76215 , n76216 , n76217 , n76218 , n76219 , n76220 , 
     n76221 , n76222 , n76223 , n76224 , n76225 , n76226 , n76227 , n76228 , n76229 , n76230 , 
     n76231 , n76232 , n76233 , n76234 , n76235 , n76236 , n76237 , n76238 , n76239 , n76240 , 
     n76241 , n76242 , n76243 , n76244 , n76245 , n76246 , n76247 , n76248 , n76249 , n76250 , 
     n76251 , n76252 , n76253 , n76254 , n76255 , n76256 , n76257 , n76258 , n76259 , n76260 , 
     n76261 , n76262 , n76263 , n76264 , n76265 , n76266 , n76267 , n76268 , n76269 , n76270 , 
     n76271 , n76272 , n76273 , n76274 , n76275 , n76276 , n76277 , n76278 , n76279 , n76280 , 
     n76281 , n76282 , n76283 , n76284 , n76285 , n76286 , n76287 , n76288 , n76289 , n76290 , 
     n76291 , n76292 , n76293 , n76294 , n76295 , n76296 , n76297 , n76298 , n76299 , n76300 , 
     n76301 , n76302 , n76303 , n76304 , n76305 , n76306 , n76307 , n76308 , n76309 , n76310 , 
     n76311 , n76312 , n76313 , n76314 , n76315 , n76316 , n76317 , n76318 , n76319 , n76320 , 
     n76321 , n76322 , n76323 , n76324 , n76325 , n76326 , n76327 , n76328 , n76329 , n76330 , 
     n76331 , n76332 , n76333 , n76334 , n76335 , n76336 , n76337 , n76338 , n76339 , n76340 , 
     n76341 , n76342 , n76343 , n76344 , n76345 , n76346 , n76347 , n76348 , n76349 , n76350 , 
     n76351 , n76352 , n76353 , n76354 , n76355 , n76356 , n76357 , n76358 , n76359 , n76360 , 
     n76361 , n76362 , n76363 , n76364 , n76365 , n76366 , n76367 , n76368 , n76369 , n76370 , 
     n76371 , n76372 , n76373 , n76374 , n76375 , n76376 , n76377 , n76378 , n76379 , n76380 , 
     n76381 , n76382 , n76383 , n76384 , n76385 , n76386 , n76387 , n76388 , n76389 , n76390 , 
     n76391 , n76392 , n76393 , n76394 , n76395 , n76396 , n76397 , n76398 , n76399 , n76400 , 
     n76401 , n76402 , n76403 , n76404 , n76405 , n76406 , n76407 , n76408 , n76409 , n76410 , 
     n76411 , n76412 , n76413 , n76414 , n76415 , n76416 , n76417 , n76418 , n76419 , n76420 , 
     n76421 , n76422 , n76423 , n76424 , n76425 , n76426 , n76427 , n76428 , n76429 , n76430 , 
     n76431 , n76432 , n76433 , n76434 , n76435 , n76436 , n76437 , n76438 , n76439 , n76440 , 
     n76441 , n76442 , n76443 , n76444 , n76445 , n76446 , n76447 , n76448 , n76449 , n76450 , 
     n76451 , n76452 , n76453 , n76454 , n76455 , n76456 , n76457 , n76458 , n76459 , n76460 , 
     n76461 , n76462 , n76463 , n76464 , n76465 , n76466 , n76467 , n76468 , n76469 , n76470 , 
     n76471 , n76472 , n76473 , n76474 , n76475 , n76476 , n76477 , n76478 , n76479 , n76480 , 
     n76481 , n76482 , n76483 , n76484 , n76485 , n76486 , n76487 , n76488 , n76489 , n76490 , 
     n76491 , n76492 , n76493 , n76494 , n76495 , n76496 , n76497 , n76498 , n76499 , n76500 , 
     n76501 , n76502 , n76503 , n76504 , n76505 , n76506 , n76507 , n76508 , n76509 , n76510 , 
     n76511 , n76512 , n76513 , n76514 , n76515 , n76516 , n76517 , n76518 , n76519 , n76520 , 
     n76521 , n76522 , n76523 , n76524 , n76525 , n76526 , n76527 , n76528 , n76529 , n76530 , 
     n76531 , n76532 , n76533 , n76534 , n76535 , n76536 , n76537 , n76538 , n76539 , n76540 , 
     n76541 , n76542 , n76543 , n76544 , n76545 , n76546 , n76547 , n76548 , n76549 , n76550 , 
     n76551 , n76552 , n76553 , n76554 , n76555 , n76556 , n76557 , n76558 , n76559 , n76560 , 
     n76561 , n76562 , n76563 , n76564 , n76565 , n76566 , n76567 , n76568 , n76569 , n76570 , 
     n76571 , n76572 , n76573 , n76574 , n76575 , n76576 , n76577 , n76578 , n76579 , n76580 , 
     n76581 , n76582 , n76583 , n76584 , n76585 , n76586 , n76587 , n76588 , n76589 , n76590 , 
     n76591 , n76592 , n76593 , n76594 , n76595 , n76596 , n76597 , n76598 , n76599 , n76600 , 
     n76601 , n76602 , n76603 , n76604 , n76605 , n76606 , n76607 , n76608 , n76609 , n76610 , 
     n76611 , n76612 , n76613 , n76614 , n76615 , n76616 , n76617 , n76618 , n76619 , n76620 , 
     n76621 , n76622 , n76623 , n76624 , n76625 , n76626 , n76627 , n76628 , n76629 , n76630 , 
     n76631 , n76632 , n76633 , n76634 , n76635 , n76636 , n76637 , n76638 , n76639 , n76640 , 
     n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , n76649 , n76650 , 
     n76651 , n76652 , n76653 , n76654 , n76655 , n76656 , n76657 , n76658 , n76659 , n76660 , 
     n76661 , n76662 , n76663 , n76664 , n76665 , n76666 , n76667 , n76668 , n76669 , n76670 , 
     n76671 , n76672 , n76673 , n76674 , n76675 , n76676 , n76677 , n76678 , n76679 , n76680 , 
     n76681 , n76682 , n76683 , n76684 , n76685 , n76686 , n76687 , n76688 , n76689 , n76690 , 
     n76691 , n76692 , n76693 , n76694 , n76695 , n76696 , n76697 , n76698 , n76699 , n76700 , 
     n76701 , n76702 , n76703 , n76704 , n76705 , n76706 , n76707 , n76708 , n76709 , n76710 , 
     n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , 
     n76721 , n76722 , n76723 , n76724 , n76725 , n76726 , n76727 , n76728 , n76729 , n76730 , 
     n76731 , n76732 , n76733 , n76734 , n76735 , n76736 , n76737 , n76738 , n76739 , n76740 , 
     n76741 , n76742 , n76743 , n76744 , n76745 , n76746 , n76747 , n76748 , n76749 , n76750 , 
     n76751 , n76752 , n76753 , n76754 , n76755 , n76756 , n76757 , n76758 , n76759 , n76760 , 
     n76761 , n76762 , n76763 , n76764 , n76765 , n76766 , n76767 , n76768 , n76769 , n76770 , 
     n76771 , n76772 , n76773 , n76774 , n76775 , n76776 , n76777 , n76778 , n76779 , n76780 , 
     n76781 , n76782 , n76783 , n76784 , n76785 , n76786 , n76787 , n76788 , n76789 , n76790 , 
     n76791 , n76792 , n76793 , n76794 , n76795 , n76796 , n76797 , n76798 , n76799 , n76800 , 
     n76801 , n76802 , n76803 , n76804 , n76805 , n76806 , n76807 , n76808 , n76809 , n76810 , 
     n76811 , n76812 , n76813 , n76814 , n76815 , n76816 , n76817 , n76818 , n76819 , n76820 , 
     n76821 , n76822 , n76823 , n76824 , n76825 , n76826 , n76827 , n76828 , n76829 , n76830 , 
     n76831 , n76832 , n76833 , n76834 , n76835 , n76836 , n76837 , n76838 , n76839 , n76840 , 
     n76841 , n76842 , n76843 , n76844 , n76845 , n76846 , n76847 , n76848 , n76849 , n76850 , 
     n76851 , n76852 , n76853 , n76854 , n76855 , n76856 , n76857 , n76858 , n76859 , n76860 , 
     n76861 , n76862 , n76863 , n76864 , n76865 , n76866 , n76867 , n76868 , n76869 , n76870 , 
     n76871 , n76872 , n76873 , n76874 , n76875 , n76876 , n76877 , n76878 , n76879 , n76880 , 
     n76881 , n76882 , n76883 , n76884 , n76885 , n76886 , n76887 , n76888 , n76889 , n76890 , 
     n76891 , n76892 , n76893 , n76894 , n76895 , n76896 , n76897 , n76898 , n76899 , n76900 , 
     n76901 , n76902 , n76903 , n76904 , n76905 , n76906 , n76907 , n76908 , n76909 , n76910 , 
     n76911 , n76912 , n76913 , n76914 , n76915 , n76916 , n76917 , n76918 , n76919 , n76920 , 
     n76921 , n76922 , n76923 , n76924 , n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , 
     n76931 , n76932 , n76933 , n76934 , n76935 , n76936 , n76937 , n76938 , n76939 , n76940 , 
     n76941 , n76942 , n76943 , n76944 , n76945 , n76946 , n76947 , n76948 , n76949 , n76950 , 
     n76951 , n76952 , n76953 , n76954 , n76955 , n76956 , n76957 , n76958 , n76959 , n76960 , 
     n76961 , n76962 , n76963 , n76964 , n76965 , n76966 , n76967 , n76968 , n76969 , n76970 , 
     n76971 , n76972 , n76973 , n76974 , n76975 , n76976 , n76977 , n76978 , n76979 , n76980 , 
     n76981 , n76982 , n76983 , n76984 , n76985 , n76986 , n76987 , n76988 , n76989 , n76990 , 
     n76991 , n76992 , n76993 , n76994 , n76995 , n76996 , n76997 , n76998 , n76999 , n77000 , 
     n77001 , n77002 , n77003 , n77004 , n77005 , n77006 , n77007 , n77008 , n77009 , n77010 , 
     n77011 , n77012 , n77013 , n77014 , n77015 , n77016 , n77017 , n77018 , n77019 , n77020 , 
     n77021 , n77022 , n77023 , n77024 , n77025 , n77026 , n77027 , n77028 , n77029 , n77030 , 
     n77031 , n77032 , n77033 , n77034 , n77035 , n77036 , n77037 , n77038 , n77039 , n77040 , 
     n77041 , n77042 , n77043 , n77044 , n77045 , n77046 , n77047 , n77048 , n77049 , n77050 , 
     n77051 , n77052 , n77053 , n77054 , n77055 , n77056 , n77057 , n77058 , n77059 , n77060 , 
     n77061 , n77062 , n77063 , n77064 , n77065 , n77066 , n77067 , n77068 , n77069 , n77070 , 
     n77071 , n77072 , n77073 , n77074 , n77075 , n77076 , n77077 , n77078 , n77079 , n77080 , 
     n77081 , n77082 , n77083 , n77084 , n77085 , n77086 , n77087 , n77088 , n77089 , n77090 , 
     n77091 , n77092 , n77093 , n77094 , n77095 , n77096 , n77097 , n77098 , n77099 , n77100 , 
     n77101 , n77102 , n77103 , n77104 , n77105 , n77106 , n77107 , n77108 , n77109 , n77110 , 
     n77111 , n77112 , n77113 , n77114 , n77115 , n77116 , n77117 , n77118 , n77119 , n77120 , 
     n77121 , n77122 , n77123 , n77124 , n77125 , n77126 , n77127 , n77128 , n77129 , n77130 , 
     n77131 , n77132 , n77133 , n77134 , n77135 , n77136 , n77137 , n77138 , n77139 , n77140 , 
     n77141 , n77142 , n77143 , n77144 , n77145 , n77146 , n77147 , n77148 , n77149 , n77150 , 
     n77151 , n77152 , n77153 , n77154 , n77155 , n77156 , n77157 , n77158 , n77159 , n77160 , 
     n77161 , n77162 , n77163 , n77164 , n77165 , n77166 , n77167 , n77168 , n77169 , n77170 , 
     n77171 , n77172 , n77173 , n77174 , n77175 , n77176 , n77177 , n77178 , n77179 , n77180 , 
     n77181 , n77182 , n77183 , n77184 , n77185 , n77186 , n77187 , n77188 , n77189 , n77190 , 
     n77191 , n77192 , n77193 , n77194 , n77195 , n77196 , n77197 , n77198 , n77199 , n77200 , 
     n77201 , n77202 , n77203 , n77204 , n77205 , n77206 , n77207 , n77208 , n77209 , n77210 , 
     n77211 , n77212 , n77213 , n77214 , n77215 , n77216 , n77217 , n77218 , n77219 , n77220 , 
     n77221 , n77222 , n77223 , n77224 , n77225 , n77226 , n77227 , n77228 , n77229 , n77230 , 
     n77231 , n77232 , n77233 , n77234 , n77235 , n77236 , n77237 , n77238 , n77239 , n77240 , 
     n77241 , n77242 , n77243 , n77244 , n77245 , n77246 , n77247 , n77248 , n77249 , n77250 , 
     n77251 , n77252 , n77253 , n77254 , n77255 , n77256 , n77257 , n77258 , n77259 , n77260 , 
     n77261 , n77262 , n77263 , n77264 , n77265 , n77266 , n77267 , n77268 , n77269 , n77270 , 
     n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , 
     n77281 , n77282 , n77283 , n77284 , n77285 , n77286 , n77287 , n77288 , n77289 , n77290 , 
     n77291 , n77292 , n77293 , n77294 , n77295 , n77296 , n77297 , n77298 , n77299 , n77300 , 
     n77301 , n77302 , n77303 , n77304 , n77305 , n77306 , n77307 , n77308 , n77309 , n77310 , 
     n77311 , n77312 , n77313 , n77314 , n77315 , n77316 , n77317 , n77318 , n77319 , n77320 , 
     n77321 , n77322 , n77323 , n77324 , n77325 , n77326 , n77327 , n77328 , n77329 , n77330 , 
     n77331 , n77332 , n77333 , n77334 , n77335 , n77336 , n77337 , n77338 , n77339 , n77340 , 
     n77341 , n77342 , n77343 , n77344 , n77345 , n77346 , n77347 , n77348 , n77349 , n77350 , 
     n77351 , n77352 , n77353 , n77354 , n77355 , n77356 , n77357 , n77358 , n77359 , n77360 , 
     n77361 , n77362 , n77363 , n77364 , n77365 , n77366 , n77367 , n77368 , n77369 , n77370 , 
     n77371 , n77372 , n77373 , n77374 , n77375 , n77376 , n77377 , n77378 , n77379 , n77380 , 
     n77381 , n77382 , n77383 , n77384 , n77385 , n77386 , n77387 , n77388 , n77389 , n77390 , 
     n77391 , n77392 , n77393 , n77394 , n77395 , n77396 , n77397 , n77398 , n77399 , n77400 , 
     n77401 , n77402 , n77403 , n77404 , n77405 , n77406 , n77407 , n77408 , n77409 , n77410 , 
     n77411 , n77412 , n77413 , n77414 , n77415 , n77416 , n77417 , n77418 , n77419 , n77420 , 
     n77421 , n77422 , n77423 , n77424 , n77425 , n77426 , n77427 , n77428 , n77429 , n77430 , 
     n77431 , n77432 , n77433 , n77434 , n77435 , n77436 , n77437 , n77438 , n77439 , n77440 , 
     n77441 , n77442 , n77443 , n77444 , n77445 , n77446 , n77447 , n77448 , n77449 , n77450 , 
     n77451 , n77452 , n77453 , n77454 , n77455 , n77456 , n77457 , n77458 , n77459 , n77460 , 
     n77461 , n77462 , n77463 , n77464 , n77465 , n77466 , n77467 , n77468 , n77469 , n77470 , 
     n77471 , n77472 , n77473 , n77474 , n77475 , n77476 , n77477 , n77478 , n77479 , n77480 , 
     n77481 , n77482 , n77483 , n77484 , n77485 , n77486 , n77487 , n77488 , n77489 , n77490 , 
     n77491 , n77492 , n77493 , n77494 , n77495 , n77496 , n77497 , n77498 , n77499 , n77500 , 
     n77501 , n77502 , n77503 , n77504 , n77505 , n77506 , n77507 , n77508 , n77509 , n77510 , 
     n77511 , n77512 , n77513 , n77514 , n77515 , n77516 , n77517 , n77518 , n77519 , n77520 , 
     n77521 , n77522 , n77523 , n77524 , n77525 , n77526 , n77527 , n77528 , n77529 , n77530 , 
     n77531 , n77532 , n77533 , n77534 , n77535 , n77536 , n77537 , n77538 , n77539 , n77540 , 
     n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , 
     n77551 , n77552 , n77553 , n77554 , n77555 , n77556 , n77557 , n77558 , n77559 , n77560 , 
     n77561 , n77562 , n77563 , n77564 , n77565 , n77566 , n77567 , n77568 , n77569 , n77570 , 
     n77571 , n77572 , n77573 , n77574 , n77575 , n77576 , n77577 , n77578 , n77579 , n77580 , 
     n77581 , n77582 , n77583 , n77584 , n77585 , n77586 , n77587 , n77588 , n77589 , n77590 , 
     n77591 , n77592 , n77593 , n77594 , n77595 , n77596 , n77597 , n77598 , n77599 , n77600 , 
     n77601 , n77602 , n77603 , n77604 , n77605 , n77606 , n77607 , n77608 , n77609 , n77610 , 
     n77611 , n77612 , n77613 , n77614 , n77615 , n77616 , n77617 , n77618 , n77619 , n77620 , 
     n77621 , n77622 , n77623 , n77624 , n77625 , n77626 , n77627 , n77628 , n77629 , n77630 , 
     n77631 , n77632 , n77633 , n77634 , n77635 , n77636 , n77637 , n77638 , n77639 , n77640 , 
     n77641 , n77642 , n77643 , n77644 , n77645 , n77646 , n77647 , n77648 , n77649 , n77650 , 
     n77651 , n77652 , n77653 , n77654 , n77655 , n77656 , n77657 , n77658 , n77659 , n77660 , 
     n77661 , n77662 , n77663 , n77664 , n77665 , n77666 , n77667 , n77668 , n77669 , n77670 , 
     n77671 , n77672 , n77673 , n77674 , n77675 , n77676 , n77677 , n77678 , n77679 , n77680 , 
     n77681 , n77682 , n77683 , n77684 , n77685 , n77686 , n77687 , n77688 , n77689 , n77690 , 
     n77691 , n77692 , n77693 , n77694 , n77695 , n77696 , n77697 , n77698 , n77699 , n77700 , 
     n77701 , n77702 , n77703 , n77704 , n77705 , n77706 , n77707 , n77708 , n77709 , n77710 , 
     n77711 , n77712 , n77713 , n77714 , n77715 , n77716 , n77717 , n77718 , n77719 , n77720 , 
     n77721 , n77722 , n77723 , n77724 , n77725 , n77726 , n77727 , n77728 , n77729 , n77730 , 
     n77731 , n77732 , n77733 , n77734 , n77735 , n77736 , n77737 , n77738 , n77739 , n77740 , 
     n77741 , n77742 , n77743 , n77744 , n77745 , n77746 , n77747 , n77748 , n77749 , n77750 , 
     n77751 , n77752 , n77753 , n77754 , n77755 , n77756 , n77757 , n77758 , n77759 , n77760 , 
     n77761 , n77762 , n77763 , n77764 , n77765 , n77766 , n77767 , n77768 , n77769 , n77770 , 
     n77771 , n77772 , n77773 , n77774 , n77775 , n77776 , n77777 , n77778 , n77779 , n77780 , 
     n77781 , n77782 , n77783 , n77784 , n77785 , n77786 , n77787 , n77788 , n77789 , n77790 , 
     n77791 , n77792 , n77793 , n77794 , n77795 , n77796 , n77797 , n77798 , n77799 , n77800 , 
     n77801 , n77802 , n77803 , n77804 , n77805 , n77806 , n77807 , n77808 , n77809 , n77810 , 
     n77811 , n77812 , n77813 , n77814 , n77815 , n77816 , n77817 , n77818 , n77819 , n77820 , 
     n77821 , n77822 , n77823 , n77824 , n77825 , n77826 , n77827 , n77828 , n77829 , n77830 , 
     n77831 , n77832 , n77833 , n77834 , n77835 , n77836 , n77837 , n77838 , n77839 , n77840 , 
     n77841 , n77842 , n77843 , n77844 , n77845 , n77846 , n77847 , n77848 , n77849 , n77850 , 
     n77851 , n77852 , n77853 , n77854 , n77855 , n77856 , n77857 , n77858 , n77859 , n77860 , 
     n77861 , n77862 , n77863 , n77864 , n77865 , n77866 , n77867 , n77868 , n77869 , n77870 , 
     n77871 , n77872 , n77873 , n77874 , n77875 , n77876 , n77877 , n77878 , n77879 , n77880 , 
     n77881 , n77882 , n77883 , n77884 , n77885 , n77886 , n77887 , n77888 , n77889 , n77890 , 
     n77891 , n77892 , n77893 , n77894 , n77895 , n77896 , n77897 , n77898 , n77899 , n77900 , 
     n77901 , n77902 , n77903 , n77904 , n77905 , n77906 , n77907 , n77908 , n77909 , n77910 , 
     n77911 , n77912 , n77913 , n77914 , n77915 , n77916 , n77917 , n77918 , n77919 , n77920 , 
     n77921 , n77922 , n77923 , n77924 , n77925 , n77926 , n77927 , n77928 , n77929 , n77930 , 
     n77931 , n77932 , n77933 , n77934 , n77935 , n77936 , n77937 , n77938 , n77939 , n77940 , 
     n77941 , n77942 , n77943 , n77944 , n77945 , n77946 , n77947 , n77948 , n77949 , n77950 , 
     n77951 , n77952 , n77953 , n77954 , n77955 , n77956 , n77957 , n77958 , n77959 , n77960 , 
     n77961 , n77962 , n77963 , n77964 , n77965 , n77966 , n77967 , n77968 , n77969 , n77970 , 
     n77971 , n77972 , n77973 , n77974 , n77975 , n77976 , n77977 , n77978 , n77979 , n77980 , 
     n77981 , n77982 , n77983 , n77984 , n77985 , n77986 , n77987 , n77988 , n77989 , n77990 , 
     n77991 , n77992 , n77993 , n77994 , n77995 , n77996 , n77997 , n77998 , n77999 , n78000 , 
     n78001 , n78002 , n78003 , n78004 , n78005 , n78006 , n78007 , n78008 , n78009 , n78010 , 
     n78011 , n78012 , n78013 , n78014 , n78015 , n78016 , n78017 , n78018 , n78019 , n78020 , 
     n78021 , n78022 , n78023 , n78024 , n78025 , n78026 , n78027 , n78028 , n78029 , n78030 , 
     n78031 , n78032 , n78033 , n78034 , n78035 , n78036 , n78037 , n78038 , n78039 , n78040 , 
     n78041 , n78042 , n78043 , n78044 , n78045 , n78046 , n78047 , n78048 , n78049 , n78050 , 
     n78051 , n78052 , n78053 , n78054 , n78055 , n78056 , n78057 , n78058 , n78059 , n78060 , 
     n78061 , n78062 , n78063 , n78064 , n78065 , n78066 , n78067 , n78068 , n78069 , n78070 , 
     n78071 , n78072 , n78073 , n78074 , n78075 , n78076 , n78077 , n78078 , n78079 , n78080 , 
     n78081 , n78082 , n78083 , n78084 , n78085 , n78086 , n78087 , n78088 , n78089 , n78090 , 
     n78091 , n78092 , n78093 , n78094 , n78095 , n78096 , n78097 , n78098 , n78099 , n78100 , 
     n78101 , n78102 , n78103 , n78104 , n78105 , n78106 , n78107 , n78108 , n78109 , n78110 , 
     n78111 , n78112 , n78113 , n78114 , n78115 , n78116 , n78117 , n78118 , n78119 , n78120 , 
     n78121 , n78122 , n78123 , n78124 , n78125 , n78126 , n78127 , n78128 , n78129 , n78130 , 
     n78131 , n78132 , n78133 , n78134 , n78135 , n78136 , n78137 , n78138 , n78139 , n78140 , 
     n78141 , n78142 , n78143 , n78144 , n78145 , n78146 , n78147 , n78148 , n78149 , n78150 , 
     n78151 , n78152 , n78153 , n78154 , n78155 , n78156 , n78157 , n78158 , n78159 , n78160 , 
     n78161 , n78162 , n78163 , n78164 , n78165 , n78166 , n78167 , n78168 , n78169 , n78170 , 
     n78171 , n78172 , n78173 , n78174 , n78175 , n78176 , n78177 , n78178 , n78179 , n78180 , 
     n78181 , n78182 , n78183 , n78184 , n78185 , n78186 , n78187 , n78188 , n78189 , n78190 , 
     n78191 , n78192 , n78193 , n78194 , n78195 , n78196 , n78197 , n78198 , n78199 , n78200 , 
     n78201 , n78202 , n78203 , n78204 , n78205 , n78206 , n78207 , n78208 , n78209 , n78210 , 
     n78211 , n78212 , n78213 , n78214 , n78215 , n78216 , n78217 , n78218 , n78219 , n78220 , 
     n78221 , n78222 , n78223 , n78224 , n78225 , n78226 , n78227 , n78228 , n78229 , n78230 , 
     n78231 , n78232 , n78233 , n78234 , n78235 , n78236 , n78237 , n78238 , n78239 , n78240 , 
     n78241 , n78242 , n78243 , n78244 , n78245 , n78246 , n78247 , n78248 , n78249 , n78250 , 
     n78251 , n78252 , n78253 , n78254 , n78255 , n78256 , n78257 , n78258 , n78259 , n78260 , 
     n78261 , n78262 , n78263 , n78264 , n78265 , n78266 , n78267 , n78268 , n78269 , n78270 , 
     n78271 , n78272 , n78273 , n78274 , n78275 , n78276 , n78277 , n78278 , n78279 , n78280 , 
     n78281 , n78282 , n78283 , n78284 , n78285 , n78286 , n78287 , n78288 , n78289 , n78290 , 
     n78291 , n78292 , n78293 , n78294 , n78295 , n78296 , n78297 , n78298 , n78299 , n78300 , 
     n78301 , n78302 , n78303 , n78304 , n78305 , n78306 , n78307 , n78308 , n78309 , n78310 , 
     n78311 , n78312 , n78313 , n78314 , n78315 , n78316 , n78317 , n78318 , n78319 , n78320 , 
     n78321 , n78322 , n78323 , n78324 , n78325 , n78326 , n78327 , n78328 , n78329 , n78330 , 
     n78331 , n78332 , n78333 , n78334 , n78335 , n78336 , n78337 , n78338 , n78339 , n78340 , 
     n78341 , n78342 , n78343 , n78344 , n78345 , n78346 , n78347 , n78348 , n78349 , n78350 , 
     n78351 , n78352 , n78353 , n78354 , n78355 , n78356 , n78357 , n78358 , n78359 , n78360 , 
     n78361 , n78362 , n78363 , n78364 , n78365 , n78366 , n78367 , n78368 , n78369 , n78370 , 
     n78371 , n78372 , n78373 , n78374 , n78375 , n78376 , n78377 , n78378 , n78379 , n78380 , 
     n78381 , n78382 , n78383 , n78384 , n78385 , n78386 , n78387 , n78388 , n78389 , n78390 , 
     n78391 , n78392 , n78393 , n78394 , n78395 , n78396 , n78397 , n78398 , n78399 , n78400 , 
     n78401 , n78402 , n78403 , n78404 , n78405 , n78406 , n78407 , n78408 , n78409 , n78410 , 
     n78411 , n78412 , n78413 , n78414 , n78415 , n78416 , n78417 , n78418 , n78419 , n78420 , 
     n78421 , n78422 , n78423 , n78424 , n78425 , n78426 , n78427 , n78428 , n78429 , n78430 , 
     n78431 , n78432 , n78433 , n78434 , n78435 , n78436 , n78437 , n78438 , n78439 , n78440 , 
     n78441 , n78442 , n78443 , n78444 , n78445 , n78446 , n78447 , n78448 , n78449 , n78450 , 
     n78451 , n78452 , n78453 , n78454 , n78455 , n78456 , n78457 , n78458 , n78459 , n78460 , 
     n78461 , n78462 , n78463 , n78464 , n78465 , n78466 , n78467 , n78468 , n78469 , n78470 , 
     n78471 , n78472 , n78473 , n78474 , n78475 , n78476 , n78477 , n78478 , n78479 , n78480 , 
     n78481 , n78482 , n78483 , n78484 , n78485 , n78486 , n78487 , n78488 , n78489 , n78490 , 
     n78491 , n78492 , n78493 , n78494 , n78495 , n78496 , n78497 , n78498 , n78499 , n78500 , 
     n78501 , n78502 , n78503 , n78504 , n78505 , n78506 , n78507 , n78508 , n78509 , n78510 , 
     n78511 , n78512 , n78513 , n78514 , n78515 , n78516 , n78517 , n78518 , n78519 , n78520 , 
     n78521 , n78522 , n78523 , n78524 , n78525 , n78526 , n78527 , n78528 , n78529 , n78530 , 
     n78531 , n78532 , n78533 , n78534 , n78535 , n78536 , n78537 , n78538 , n78539 , n78540 , 
     n78541 , n78542 , n78543 , n78544 , n78545 , n78546 , n78547 , n78548 , n78549 , n78550 , 
     n78551 , n78552 , n78553 , n78554 , n78555 , n78556 , n78557 , n78558 , n78559 , n78560 , 
     n78561 , n78562 , n78563 , n78564 , n78565 , n78566 , n78567 , n78568 , n78569 , n78570 , 
     n78571 , n78572 , n78573 , n78574 , n78575 , n78576 , n78577 , n78578 , n78579 , n78580 , 
     n78581 , n78582 , n78583 , n78584 , n78585 , n78586 , n78587 , n78588 , n78589 , n78590 , 
     n78591 , n78592 , n78593 , n78594 , n78595 , n78596 , n78597 , n78598 , n78599 , n78600 , 
     n78601 , n78602 , n78603 , n78604 , n78605 , n78606 , n78607 , n78608 , n78609 , n78610 , 
     n78611 , n78612 , n78613 , n78614 , n78615 , n78616 , n78617 , n78618 , n78619 , n78620 , 
     n78621 , n78622 , n78623 , n78624 , n78625 , n78626 , n78627 , n78628 , n78629 , n78630 , 
     n78631 , n78632 , n78633 , n78634 , n78635 , n78636 , n78637 , n78638 , n78639 , n78640 , 
     n78641 , n78642 , n78643 , n78644 , n78645 , n78646 , n78647 , n78648 , n78649 , n78650 , 
     n78651 , n78652 , n78653 , n78654 , n78655 , n78656 , n78657 , n78658 , n78659 , n78660 , 
     n78661 , n78662 , n78663 , n78664 , n78665 , n78666 , n78667 , n78668 , n78669 , n78670 , 
     n78671 , n78672 , n78673 , n78674 , n78675 , n78676 , n78677 , n78678 , n78679 , n78680 , 
     n78681 , n78682 , n78683 , n78684 , n78685 , n78686 , n78687 , n78688 , n78689 , n78690 , 
     n78691 , n78692 , n78693 , n78694 , n78695 , n78696 , n78697 , n78698 , n78699 , n78700 , 
     n78701 , n78702 , n78703 , n78704 , n78705 , n78706 , n78707 , n78708 , n78709 , n78710 , 
     n78711 , n78712 , n78713 , n78714 , n78715 , n78716 , n78717 , n78718 , n78719 , n78720 , 
     n78721 , n78722 , n78723 , n78724 , n78725 , n78726 , n78727 , n78728 , n78729 , n78730 , 
     n78731 , n78732 , n78733 , n78734 , n78735 , n78736 , n78737 , n78738 , n78739 , n78740 , 
     n78741 , n78742 , n78743 , n78744 , n78745 , n78746 , n78747 , n78748 , n78749 , n78750 , 
     n78751 , n78752 , n78753 , n78754 , n78755 , n78756 , n78757 , n78758 , n78759 , n78760 , 
     n78761 , n78762 , n78763 , n78764 , n78765 , n78766 , n78767 , n78768 , n78769 , n78770 , 
     n78771 , n78772 , n78773 , n78774 , n78775 , n78776 , n78777 , n78778 , n78779 , n78780 , 
     n78781 , n78782 , n78783 , n78784 , n78785 , n78786 , n78787 , n78788 , n78789 , n78790 , 
     n78791 , n78792 , n78793 , n78794 , n78795 , n78796 , n78797 , n78798 , n78799 , n78800 , 
     n78801 , n78802 , n78803 , n78804 , n78805 , n78806 , n78807 , n78808 , n78809 , n78810 , 
     n78811 , n78812 , n78813 , n78814 , n78815 , n78816 , n78817 , n78818 , n78819 , n78820 , 
     n78821 , n78822 , n78823 , n78824 , n78825 , n78826 , n78827 , n78828 , n78829 , n78830 , 
     n78831 , n78832 , n78833 , n78834 , n78835 , n78836 , n78837 , n78838 , n78839 , n78840 , 
     n78841 , n78842 , n78843 , n78844 , n78845 , n78846 , n78847 , n78848 , n78849 , n78850 , 
     n78851 , n78852 , n78853 , n78854 , n78855 , n78856 , n78857 , n78858 , n78859 , n78860 , 
     n78861 , n78862 , n78863 , n78864 , n78865 , n78866 , n78867 , n78868 , n78869 , n78870 , 
     n78871 , n78872 , n78873 , n78874 , n78875 , n78876 , n78877 , n78878 , n78879 , n78880 , 
     n78881 , n78882 , n78883 , n78884 , n78885 , n78886 , n78887 , n78888 , n78889 , n78890 , 
     n78891 , n78892 , n78893 , n78894 , n78895 , n78896 , n78897 , n78898 , n78899 , n78900 , 
     n78901 , n78902 , n78903 , n78904 , n78905 , n78906 , n78907 , n78908 , n78909 , n78910 , 
     n78911 , n78912 , n78913 , n78914 , n78915 , n78916 , n78917 , n78918 , n78919 , n78920 , 
     n78921 , n78922 , n78923 , n78924 , n78925 , n78926 , n78927 , n78928 , n78929 , n78930 , 
     n78931 , n78932 , n78933 , n78934 , n78935 , n78936 , n78937 , n78938 , n78939 , n78940 , 
     n78941 , n78942 , n78943 , n78944 , n78945 , n78946 , n78947 , n78948 , n78949 , n78950 , 
     n78951 , n78952 , n78953 , n78954 , n78955 , n78956 , n78957 , n78958 , n78959 , n78960 , 
     n78961 , n78962 , n78963 , n78964 , n78965 , n78966 , n78967 , n78968 , n78969 , n78970 , 
     n78971 , n78972 , n78973 , n78974 , n78975 , n78976 , n78977 , n78978 , n78979 , n78980 , 
     n78981 , n78982 , n78983 , n78984 , n78985 , n78986 , n78987 , n78988 , n78989 , n78990 , 
     n78991 , n78992 , n78993 , n78994 , n78995 , n78996 , n78997 , n78998 , n78999 , n79000 , 
     n79001 , n79002 , n79003 , n79004 , n79005 , n79006 , n79007 , n79008 , n79009 , n79010 , 
     n79011 , n79012 , n79013 , n79014 , n79015 , n79016 , n79017 , n79018 , n79019 , n79020 , 
     n79021 , n79022 , n79023 , n79024 , n79025 , n79026 , n79027 , n79028 , n79029 , n79030 , 
     n79031 , n79032 , n79033 , n79034 , n79035 , n79036 , n79037 , n79038 , n79039 , n79040 , 
     n79041 , n79042 , n79043 , n79044 , n79045 , n79046 , n79047 , n79048 , n79049 , n79050 , 
     n79051 , n79052 , n79053 , n79054 , n79055 , n79056 , n79057 , n79058 , n79059 , n79060 , 
     n79061 , n79062 , n79063 , n79064 , n79065 , n79066 , n79067 , n79068 , n79069 , n79070 , 
     n79071 , n79072 , n79073 , n79074 , n79075 , n79076 , n79077 , n79078 , n79079 , n79080 , 
     n79081 , n79082 , n79083 , n79084 , n79085 , n79086 , n79087 , n79088 , n79089 , n79090 , 
     n79091 , n79092 , n79093 , n79094 , n79095 , n79096 , n79097 , n79098 , n79099 , n79100 , 
     n79101 , n79102 , n79103 , n79104 , n79105 , n79106 , n79107 , n79108 , n79109 , n79110 , 
     n79111 , n79112 , n79113 , n79114 , n79115 , n79116 , n79117 , n79118 , n79119 , n79120 , 
     n79121 , n79122 , n79123 , n79124 , n79125 , n79126 , n79127 , n79128 , n79129 , n79130 , 
     n79131 , n79132 , n79133 , n79134 , n79135 , n79136 , n79137 , n79138 , n79139 , n79140 , 
     n79141 , n79142 , n79143 , n79144 , n79145 , n79146 , n79147 , n79148 , n79149 , n79150 , 
     n79151 , n79152 , n79153 , n79154 , n79155 , n79156 , n79157 , n79158 , n79159 , n79160 , 
     n79161 , n79162 , n79163 , n79164 , n79165 , n79166 , n79167 , n79168 , n79169 , n79170 , 
     n79171 , n79172 , n79173 , n79174 , n79175 , n79176 , n79177 , n79178 , n79179 , n79180 , 
     n79181 , n79182 , n79183 , n79184 , n79185 , n79186 , n79187 , n79188 , n79189 , n79190 , 
     n79191 , n79192 , n79193 , n79194 , n79195 , n79196 , n79197 , n79198 , n79199 , n79200 , 
     n79201 , n79202 , n79203 , n79204 , n79205 , n79206 , n79207 , n79208 , n79209 , n79210 , 
     n79211 , n79212 , n79213 , n79214 , n79215 , n79216 , n79217 , n79218 , n79219 , n79220 , 
     n79221 , n79222 , n79223 , n79224 , n79225 , n79226 , n79227 , n79228 , n79229 , n79230 , 
     n79231 , n79232 , n79233 , n79234 , n79235 , n79236 , n79237 , n79238 , n79239 , n79240 , 
     n79241 , n79242 , n79243 , n79244 , n79245 , n79246 , n79247 , n79248 , n79249 , n79250 , 
     n79251 , n79252 , n79253 , n79254 , n79255 , n79256 , n79257 , n79258 , n79259 , n79260 , 
     n79261 , n79262 , n79263 , n79264 , n79265 , n79266 , n79267 , n79268 , n79269 , n79270 , 
     n79271 , n79272 , n79273 , n79274 , n79275 , n79276 , n79277 , n79278 , n79279 , n79280 , 
     n79281 , n79282 , n79283 , n79284 , n79285 , n79286 , n79287 , n79288 , n79289 , n79290 , 
     n79291 , n79292 , n79293 , n79294 , n79295 , n79296 , n79297 , n79298 , n79299 , n79300 , 
     n79301 , n79302 , n79303 , n79304 , n79305 , n79306 , n79307 , n79308 , n79309 , n79310 , 
     n79311 , n79312 , n79313 , n79314 , n79315 , n79316 , n79317 , n79318 , n79319 , n79320 , 
     n79321 , n79322 , n79323 , n79324 , n79325 , n79326 , n79327 , n79328 , n79329 , n79330 , 
     n79331 , n79332 , n79333 , n79334 , n79335 , n79336 , n79337 , n79338 , n79339 , n79340 , 
     n79341 , n79342 , n79343 , n79344 , n79345 , n79346 , n79347 , n79348 , n79349 , n79350 , 
     n79351 , n79352 , n79353 , n79354 , n79355 , n79356 , n79357 , n79358 , n79359 , n79360 , 
     n79361 , n79362 , n79363 , n79364 , n79365 , n79366 , n79367 , n79368 , n79369 , n79370 , 
     n79371 , n79372 , n79373 , n79374 , n79375 , n79376 , n79377 , n79378 , n79379 , n79380 , 
     n79381 , n79382 , n79383 , n79384 , n79385 , n79386 , n79387 , n79388 , n79389 , n79390 , 
     n79391 , n79392 , n79393 , n79394 , n79395 , n79396 , n79397 , n79398 , n79399 , n79400 , 
     n79401 , n79402 , n79403 , n79404 , n79405 , n79406 , n79407 , n79408 , n79409 , n79410 , 
     n79411 , n79412 , n79413 , n79414 , n79415 , n79416 , n79417 , n79418 , n79419 , n79420 , 
     n79421 , n79422 , n79423 , n79424 , n79425 , n79426 , n79427 , n79428 , n79429 , n79430 , 
     n79431 , n79432 , n79433 , n79434 , n79435 , n79436 , n79437 , n79438 , n79439 , n79440 , 
     n79441 , n79442 , n79443 , n79444 , n79445 , n79446 , n79447 , n79448 , n79449 , n79450 , 
     n79451 , n79452 , n79453 , n79454 , n79455 , n79456 , n79457 , n79458 , n79459 , n79460 , 
     n79461 , n79462 , n79463 , n79464 , n79465 , n79466 , n79467 , n79468 , n79469 , n79470 , 
     n79471 , n79472 , n79473 , n79474 , n79475 , n79476 , n79477 , n79478 , n79479 , n79480 , 
     n79481 , n79482 , n79483 , n79484 , n79485 , n79486 , n79487 , n79488 , n79489 , n79490 , 
     n79491 , n79492 , n79493 , n79494 , n79495 , n79496 , n79497 , n79498 , n79499 , n79500 , 
     n79501 , n79502 , n79503 , n79504 , n79505 , n79506 , n79507 , n79508 , n79509 , n79510 , 
     n79511 , n79512 , n79513 , n79514 , n79515 , n79516 , n79517 , n79518 , n79519 , n79520 , 
     n79521 , n79522 , n79523 , n79524 , n79525 , n79526 , n79527 , n79528 , n79529 , n79530 , 
     n79531 , n79532 , n79533 , n79534 , n79535 , n79536 , n79537 , n79538 , n79539 , n79540 , 
     n79541 , n79542 , n79543 , n79544 , n79545 , n79546 , n79547 , n79548 , n79549 , n79550 , 
     n79551 , n79552 , n79553 , n79554 , n79555 , n79556 , n79557 , n79558 , n79559 , n79560 , 
     n79561 , n79562 , n79563 , n79564 , n79565 , n79566 , n79567 , n79568 , n79569 , n79570 , 
     n79571 , n79572 , n79573 , n79574 , n79575 , n79576 , n79577 , n79578 , n79579 , n79580 , 
     n79581 , n79582 , n79583 , n79584 , n79585 , n79586 , n79587 , n79588 , n79589 , n79590 , 
     n79591 , n79592 , n79593 , n79594 , n79595 , n79596 , n79597 , n79598 , n79599 , n79600 , 
     n79601 , n79602 , n79603 , n79604 , n79605 , n79606 , n79607 , n79608 , n79609 , n79610 , 
     n79611 , n79612 , n79613 , n79614 , n79615 , n79616 , n79617 , n79618 , n79619 , n79620 , 
     n79621 , n79622 , n79623 , n79624 , n79625 , n79626 , n79627 , n79628 , n79629 , n79630 , 
     n79631 , n79632 , n79633 , n79634 , n79635 , n79636 , n79637 , n79638 , n79639 , n79640 , 
     n79641 , n79642 , n79643 , n79644 , n79645 , n79646 , n79647 , n79648 , n79649 , n79650 , 
     n79651 , n79652 , n79653 , n79654 , n79655 , n79656 , n79657 , n79658 , n79659 , n79660 , 
     n79661 , n79662 , n79663 , n79664 , n79665 , n79666 , n79667 , n79668 , n79669 , n79670 , 
     n79671 , n79672 , n79673 , n79674 , n79675 , n79676 , n79677 , n79678 , n79679 , n79680 , 
     n79681 , n79682 , n79683 , n79684 , n79685 , n79686 , n79687 , n79688 , n79689 , n79690 , 
     n79691 , n79692 , n79693 , n79694 , n79695 , n79696 , n79697 , n79698 , n79699 , n79700 , 
     n79701 , n79702 , n79703 , n79704 , n79705 , n79706 , n79707 , n79708 , n79709 , n79710 , 
     n79711 , n79712 , n79713 , n79714 , n79715 , n79716 , n79717 , n79718 , n79719 , n79720 , 
     n79721 , n79722 , n79723 , n79724 , n79725 , n79726 , n79727 , n79728 , n79729 , n79730 , 
     n79731 , n79732 , n79733 , n79734 , n79735 , n79736 , n79737 , n79738 , n79739 , n79740 , 
     n79741 , n79742 , n79743 , n79744 , n79745 , n79746 , n79747 , n79748 , n79749 , n79750 , 
     n79751 , n79752 , n79753 , n79754 , n79755 , n79756 , n79757 , n79758 , n79759 , n79760 , 
     n79761 , n79762 , n79763 , n79764 , n79765 , n79766 , n79767 , n79768 , n79769 , n79770 , 
     n79771 , n79772 , n79773 , n79774 , n79775 , n79776 , n79777 , n79778 , n79779 , n79780 , 
     n79781 , n79782 , n79783 , n79784 , n79785 , n79786 , n79787 , n79788 , n79789 , n79790 , 
     n79791 , n79792 , n79793 , n79794 , n79795 , n79796 , n79797 , n79798 , n79799 , n79800 , 
     n79801 , n79802 , n79803 , n79804 , n79805 , n79806 , n79807 , n79808 , n79809 , n79810 , 
     n79811 , n79812 , n79813 , n79814 , n79815 , n79816 , n79817 , n79818 , n79819 , n79820 , 
     n79821 , n79822 , n79823 , n79824 , n79825 , n79826 , n79827 , n79828 , n79829 , n79830 , 
     n79831 , n79832 , n79833 , n79834 , n79835 , n79836 , n79837 , n79838 , n79839 , n79840 , 
     n79841 , n79842 , n79843 , n79844 , n79845 , n79846 , n79847 , n79848 , n79849 , n79850 , 
     n79851 , n79852 , n79853 , n79854 , n79855 , n79856 , n79857 , n79858 , n79859 , n79860 , 
     n79861 , n79862 , n79863 , n79864 , n79865 , n79866 , n79867 , n79868 , n79869 , n79870 , 
     n79871 , n79872 , n79873 , n79874 , n79875 , n79876 , n79877 , n79878 , n79879 , n79880 , 
     n79881 , n79882 , n79883 , n79884 , n79885 , n79886 , n79887 , n79888 , n79889 , n79890 , 
     n79891 , n79892 , n79893 , n79894 , n79895 , n79896 , n79897 , n79898 , n79899 , n79900 , 
     n79901 , n79902 , n79903 , n79904 , n79905 , n79906 , n79907 , n79908 , n79909 , n79910 , 
     n79911 , n79912 , n79913 , n79914 , n79915 , n79916 , n79917 , n79918 , n79919 , n79920 , 
     n79921 , n79922 , n79923 , n79924 , n79925 , n79926 , n79927 , n79928 , n79929 , n79930 , 
     n79931 , n79932 , n79933 , n79934 , n79935 , n79936 , n79937 , n79938 , n79939 , n79940 , 
     n79941 , n79942 , n79943 , n79944 , n79945 , n79946 , n79947 , n79948 , n79949 , n79950 , 
     n79951 , n79952 , n79953 , n79954 , n79955 , n79956 , n79957 , n79958 , n79959 , n79960 , 
     n79961 , n79962 , n79963 , n79964 , n79965 , n79966 , n79967 , n79968 , n79969 , n79970 , 
     n79971 , n79972 , n79973 , n79974 , n79975 , n79976 , n79977 , n79978 , n79979 , n79980 , 
     n79981 , n79982 , n79983 , n79984 , n79985 , n79986 , n79987 , n79988 , n79989 , n79990 , 
     n79991 , n79992 , n79993 , n79994 , n79995 , n79996 , n79997 , n79998 , n79999 , n80000 , 
     n80001 , n80002 , n80003 , n80004 , n80005 , n80006 , n80007 , n80008 , n80009 , n80010 , 
     n80011 , n80012 , n80013 , n80014 , n80015 , n80016 , n80017 , n80018 , n80019 , n80020 , 
     n80021 , n80022 , n80023 , n80024 , n80025 , n80026 , n80027 , n80028 , n80029 , n80030 , 
     n80031 , n80032 , n80033 , n80034 , n80035 , n80036 , n80037 , n80038 , n80039 , n80040 , 
     n80041 , n80042 , n80043 , n80044 , n80045 , n80046 , n80047 , n80048 , n80049 , n80050 , 
     n80051 , n80052 , n80053 , n80054 , n80055 , n80056 , n80057 , n80058 , n80059 , n80060 , 
     n80061 , n80062 , n80063 , n80064 , n80065 , n80066 , n80067 , n80068 , n80069 , n80070 , 
     n80071 , n80072 , n80073 , n80074 , n80075 , n80076 , n80077 , n80078 , n80079 , n80080 , 
     n80081 , n80082 , n80083 , n80084 , n80085 , n80086 , n80087 , n80088 , n80089 , n80090 , 
     n80091 , n80092 , n80093 , n80094 , n80095 , n80096 , n80097 , n80098 , n80099 , n80100 , 
     n80101 , n80102 , n80103 , n80104 , n80105 , n80106 , n80107 , n80108 , n80109 , n80110 , 
     n80111 , n80112 , n80113 , n80114 , n80115 , n80116 , n80117 , n80118 , n80119 , n80120 , 
     n80121 , n80122 , n80123 , n80124 , n80125 , n80126 , n80127 , n80128 , n80129 , n80130 , 
     n80131 , n80132 , n80133 , n80134 , n80135 , n80136 , n80137 , n80138 , n80139 , n80140 , 
     n80141 , n80142 , n80143 , n80144 , n80145 , n80146 , n80147 , n80148 , n80149 , n80150 , 
     n80151 , n80152 , n80153 , n80154 , n80155 , n80156 , n80157 , n80158 , n80159 , n80160 , 
     n80161 , n80162 , n80163 , n80164 , n80165 , n80166 , n80167 , n80168 , n80169 , n80170 , 
     n80171 , n80172 , n80173 , n80174 , n80175 , n80176 , n80177 , n80178 , n80179 , n80180 , 
     n80181 , n80182 , n80183 , n80184 , n80185 , n80186 , n80187 , n80188 , n80189 , n80190 , 
     n80191 , n80192 , n80193 , n80194 , n80195 , n80196 , n80197 , n80198 , n80199 , n80200 , 
     n80201 , n80202 , n80203 , n80204 , n80205 , n80206 , n80207 , n80208 , n80209 , n80210 , 
     n80211 , n80212 , n80213 , n80214 , n80215 , n80216 , n80217 , n80218 , n80219 , n80220 , 
     n80221 , n80222 , n80223 , n80224 , n80225 , n80226 , n80227 , n80228 , n80229 , n80230 , 
     n80231 , n80232 , n80233 , n80234 , n80235 , n80236 , n80237 , n80238 , n80239 , n80240 , 
     n80241 , n80242 , n80243 , n80244 , n80245 , n80246 , n80247 , n80248 , n80249 , n80250 , 
     n80251 , n80252 , n80253 , n80254 , n80255 , n80256 , n80257 , n80258 , n80259 , n80260 , 
     n80261 , n80262 , n80263 , n80264 , n80265 , n80266 , n80267 , n80268 , n80269 , n80270 , 
     n80271 , n80272 , n80273 , n80274 , n80275 , n80276 , n80277 , n80278 , n80279 , n80280 , 
     n80281 , n80282 , n80283 , n80284 , n80285 , n80286 , n80287 , n80288 , n80289 , n80290 , 
     n80291 , n80292 , n80293 , n80294 , n80295 , n80296 , n80297 , n80298 , n80299 , n80300 , 
     n80301 , n80302 , n80303 , n80304 , n80305 , n80306 , n80307 , n80308 , n80309 , n80310 , 
     n80311 , n80312 , n80313 , n80314 , n80315 , n80316 , n80317 , n80318 , n80319 , n80320 , 
     n80321 , n80322 , n80323 , n80324 , n80325 , n80326 , n80327 , n80328 , n80329 , n80330 , 
     n80331 , n80332 , n80333 , n80334 , n80335 , n80336 , n80337 , n80338 , n80339 , n80340 , 
     n80341 , n80342 , n80343 , n80344 , n80345 , n80346 , n80347 , n80348 , n80349 , n80350 , 
     n80351 , n80352 , n80353 , n80354 , n80355 , n80356 , n80357 , n80358 , n80359 , n80360 , 
     n80361 , n80362 , n80363 , n80364 , n80365 , n80366 , n80367 , n80368 , n80369 , n80370 , 
     n80371 , n80372 , n80373 , n80374 , n80375 , n80376 , n80377 , n80378 , n80379 , n80380 , 
     n80381 , n80382 , n80383 , n80384 , n80385 , n80386 , n80387 , n80388 , n80389 , n80390 , 
     n80391 , n80392 , n80393 , n80394 , n80395 , n80396 , n80397 , n80398 , n80399 , n80400 , 
     n80401 , n80402 , n80403 , n80404 , n80405 , n80406 , n80407 , n80408 , n80409 , n80410 , 
     n80411 , n80412 , n80413 , n80414 , n80415 , n80416 , n80417 , n80418 , n80419 , n80420 , 
     n80421 , n80422 , n80423 , n80424 , n80425 , n80426 , n80427 , n80428 , n80429 , n80430 , 
     n80431 , n80432 , n80433 , n80434 , n80435 , n80436 , n80437 , n80438 , n80439 , n80440 , 
     n80441 , n80442 , n80443 , n80444 , n80445 , n80446 , n80447 , n80448 , n80449 , n80450 , 
     n80451 , n80452 , n80453 , n80454 , n80455 , n80456 , n80457 , n80458 , n80459 , n80460 , 
     n80461 , n80462 , n80463 , n80464 , n80465 , n80466 , n80467 , n80468 , n80469 , n80470 , 
     n80471 , n80472 , n80473 , n80474 , n80475 , n80476 , n80477 , n80478 , n80479 , n80480 , 
     n80481 , n80482 , n80483 , n80484 , n80485 , n80486 , n80487 , n80488 , n80489 , n80490 , 
     n80491 , n80492 , n80493 , n80494 , n80495 , n80496 , n80497 , n80498 , n80499 , n80500 , 
     n80501 , n80502 , n80503 , n80504 , n80505 , n80506 , n80507 , n80508 , n80509 , n80510 , 
     n80511 , n80512 , n80513 , n80514 , n80515 , n80516 , n80517 , n80518 , n80519 , n80520 , 
     n80521 , n80522 , n80523 , n80524 , n80525 , n80526 , n80527 , n80528 , n80529 , n80530 , 
     n80531 , n80532 , n80533 , n80534 , n80535 , n80536 , n80537 , n80538 , n80539 , n80540 , 
     n80541 , n80542 , n80543 , n80544 , n80545 , n80546 , n80547 , n80548 , n80549 , n80550 , 
     n80551 , n80552 , n80553 , n80554 , n80555 , n80556 , n80557 , n80558 , n80559 , n80560 , 
     n80561 , n80562 , n80563 , n80564 , n80565 , n80566 , n80567 , n80568 , n80569 , n80570 , 
     n80571 , n80572 , n80573 , n80574 , n80575 , n80576 , n80577 , n80578 , n80579 , n80580 , 
     n80581 , n80582 , n80583 , n80584 , n80585 , n80586 , n80587 , n80588 , n80589 , n80590 , 
     n80591 , n80592 , n80593 , n80594 , n80595 , n80596 , n80597 , n80598 , n80599 , n80600 , 
     n80601 , n80602 , n80603 , n80604 , n80605 , n80606 , n80607 , n80608 , n80609 , n80610 , 
     n80611 , n80612 , n80613 , n80614 , n80615 , n80616 , n80617 , n80618 , n80619 , n80620 , 
     n80621 , n80622 , n80623 , n80624 , n80625 , n80626 , n80627 , n80628 , n80629 , n80630 , 
     n80631 , n80632 , n80633 , n80634 , n80635 , n80636 , n80637 , n80638 , n80639 , n80640 , 
     n80641 , n80642 , n80643 , n80644 , n80645 , n80646 , n80647 , n80648 , n80649 , n80650 , 
     n80651 , n80652 , n80653 , n80654 , n80655 , n80656 , n80657 , n80658 , n80659 , n80660 , 
     n80661 , n80662 , n80663 , n80664 , n80665 , n80666 , n80667 , n80668 , n80669 , n80670 , 
     n80671 , n80672 , n80673 , n80674 , n80675 , n80676 , n80677 , n80678 , n80679 , n80680 , 
     n80681 , n80682 , n80683 , n80684 , n80685 , n80686 , n80687 , n80688 , n80689 , n80690 , 
     n80691 , n80692 , n80693 , n80694 , n80695 , n80696 , n80697 , n80698 , n80699 , n80700 , 
     n80701 , n80702 , n80703 , n80704 , n80705 , n80706 , n80707 , n80708 , n80709 , n80710 , 
     n80711 , n80712 , n80713 , n80714 , n80715 , n80716 , n80717 , n80718 , n80719 , n80720 , 
     n80721 , n80722 , n80723 , n80724 , n80725 , n80726 , n80727 , n80728 , n80729 , n80730 , 
     n80731 , n80732 , n80733 , n80734 , n80735 , n80736 , n80737 , n80738 , n80739 , n80740 , 
     n80741 , n80742 , n80743 , n80744 , n80745 , n80746 , n80747 , n80748 , n80749 , n80750 , 
     n80751 , n80752 , n80753 , n80754 , n80755 , n80756 , n80757 , n80758 , n80759 , n80760 , 
     n80761 , n80762 , n80763 , n80764 , n80765 , n80766 , n80767 , n80768 , n80769 , n80770 , 
     n80771 , n80772 , n80773 , n80774 , n80775 , n80776 , n80777 , n80778 , n80779 , n80780 , 
     n80781 , n80782 , n80783 , n80784 , n80785 , n80786 , n80787 , n80788 , n80789 , n80790 , 
     n80791 , n80792 , n80793 , n80794 , n80795 , n80796 , n80797 , n80798 , n80799 , n80800 , 
     n80801 , n80802 , n80803 , n80804 , n80805 , n80806 , n80807 , n80808 , n80809 , n80810 , 
     n80811 , n80812 , n80813 , n80814 , n80815 , n80816 , n80817 , n80818 , n80819 , n80820 , 
     n80821 , n80822 , n80823 , n80824 , n80825 , n80826 , n80827 , n80828 , n80829 , n80830 , 
     n80831 , n80832 , n80833 , n80834 , n80835 , n80836 , n80837 , n80838 , n80839 , n80840 , 
     n80841 , n80842 , n80843 , n80844 , n80845 , n80846 , n80847 , n80848 , n80849 , n80850 , 
     n80851 , n80852 , n80853 , n80854 , n80855 , n80856 , n80857 , n80858 , n80859 , n80860 , 
     n80861 , n80862 , n80863 , n80864 , n80865 , n80866 , n80867 , n80868 , n80869 , n80870 , 
     n80871 , n80872 , n80873 , n80874 , n80875 , n80876 , n80877 , n80878 , n80879 , n80880 , 
     n80881 , n80882 , n80883 , n80884 , n80885 , n80886 , n80887 , n80888 , n80889 , n80890 , 
     n80891 , n80892 , n80893 , n80894 , n80895 , n80896 , n80897 , n80898 , n80899 , n80900 , 
     n80901 , n80902 , n80903 , n80904 , n80905 , n80906 , n80907 , n80908 , n80909 , n80910 , 
     n80911 , n80912 , n80913 , n80914 , n80915 , n80916 , n80917 , n80918 , n80919 , n80920 , 
     n80921 , n80922 , n80923 , n80924 , n80925 , n80926 , n80927 , n80928 , n80929 , n80930 , 
     n80931 , n80932 , n80933 , n80934 , n80935 , n80936 , n80937 , n80938 , n80939 , n80940 , 
     n80941 , n80942 , n80943 , n80944 , n80945 , n80946 , n80947 , n80948 , n80949 , n80950 , 
     n80951 , n80952 , n80953 , n80954 , n80955 , n80956 , n80957 , n80958 , n80959 , n80960 , 
     n80961 , n80962 , n80963 , n80964 , n80965 , n80966 , n80967 , n80968 , n80969 , n80970 , 
     n80971 , n80972 , n80973 , n80974 , n80975 , n80976 , n80977 , n80978 , n80979 , n80980 , 
     n80981 , n80982 , n80983 , n80984 , n80985 , n80986 , n80987 , n80988 , n80989 , n80990 , 
     n80991 , n80992 , n80993 , n80994 , n80995 , n80996 , n80997 , n80998 , n80999 , n81000 , 
     n81001 , n81002 , n81003 , n81004 , n81005 , n81006 , n81007 , n81008 , n81009 , n81010 , 
     n81011 , n81012 , n81013 , n81014 , n81015 , n81016 , n81017 , n81018 , n81019 , n81020 , 
     n81021 , n81022 , n81023 , n81024 , n81025 , n81026 , n81027 , n81028 , n81029 , n81030 , 
     n81031 , n81032 , n81033 , n81034 , n81035 , n81036 , n81037 , n81038 , n81039 , n81040 , 
     n81041 , n81042 , n81043 , n81044 , n81045 , n81046 , n81047 , n81048 , n81049 , n81050 , 
     n81051 , n81052 , n81053 , n81054 , n81055 , n81056 , n81057 , n81058 , n81059 , n81060 , 
     n81061 , n81062 , n81063 , n81064 , n81065 , n81066 , n81067 , n81068 , n81069 , n81070 , 
     n81071 , n81072 , n81073 , n81074 , n81075 , n81076 , n81077 , n81078 , n81079 , n81080 , 
     n81081 , n81082 , n81083 , n81084 , n81085 , n81086 , n81087 , n81088 , n81089 , n81090 , 
     n81091 , n81092 , n81093 , n81094 , n81095 , n81096 , n81097 , n81098 , n81099 , n81100 , 
     n81101 , n81102 , n81103 , n81104 , n81105 , n81106 , n81107 , n81108 , n81109 , n81110 , 
     n81111 , n81112 , n81113 , n81114 , n81115 , n81116 , n81117 , n81118 , n81119 , n81120 , 
     n81121 , n81122 , n81123 , n81124 , n81125 , n81126 , n81127 , n81128 , n81129 , n81130 , 
     n81131 , n81132 , n81133 , n81134 , n81135 , n81136 , n81137 , n81138 , n81139 , n81140 , 
     n81141 , n81142 , n81143 , n81144 , n81145 , n81146 , n81147 , n81148 , n81149 , n81150 , 
     n81151 , n81152 , n81153 , n81154 , n81155 , n81156 , n81157 , n81158 , n81159 , n81160 , 
     n81161 , n81162 , n81163 , n81164 , n81165 , n81166 , n81167 , n81168 , n81169 , n81170 , 
     n81171 , n81172 , n81173 , n81174 , n81175 , n81176 , n81177 , n81178 , n81179 , n81180 , 
     n81181 , n81182 , n81183 , n81184 , n81185 , n81186 , n81187 , n81188 , n81189 , n81190 , 
     n81191 , n81192 , n81193 , n81194 , n81195 , n81196 , n81197 , n81198 , n81199 , n81200 , 
     n81201 , n81202 , n81203 , n81204 , n81205 , n81206 , n81207 , n81208 , n81209 , n81210 , 
     n81211 , n81212 , n81213 , n81214 , n81215 , n81216 , n81217 , n81218 , n81219 , n81220 , 
     n81221 , n81222 , n81223 , n81224 , n81225 , n81226 , n81227 , n81228 , n81229 , n81230 , 
     n81231 , n81232 , n81233 , n81234 , n81235 , n81236 , n81237 , n81238 , n81239 , n81240 , 
     n81241 , n81242 , n81243 , n81244 , n81245 , n81246 , n81247 , n81248 , n81249 , n81250 , 
     n81251 , n81252 , n81253 , n81254 , n81255 , n81256 , n81257 , n81258 , n81259 , n81260 , 
     n81261 , n81262 , n81263 , n81264 , n81265 , n81266 , n81267 , n81268 , n81269 , n81270 , 
     n81271 , n81272 , n81273 , n81274 , n81275 , n81276 , n81277 , n81278 , n81279 , n81280 , 
     n81281 , n81282 , n81283 , n81284 , n81285 , n81286 , n81287 , n81288 , n81289 , n81290 , 
     n81291 , n81292 , n81293 , n81294 , n81295 , n81296 , n81297 , n81298 , n81299 , n81300 , 
     n81301 , n81302 , n81303 , n81304 , n81305 , n81306 , n81307 , n81308 , n81309 , n81310 , 
     n81311 , n81312 , n81313 , n81314 , n81315 , n81316 , n81317 , n81318 , n81319 , n81320 , 
     n81321 , n81322 , n81323 , n81324 , n81325 , n81326 , n81327 , n81328 , n81329 , n81330 , 
     n81331 , n81332 , n81333 , n81334 , n81335 , n81336 , n81337 , n81338 , n81339 , n81340 , 
     n81341 , n81342 , n81343 , n81344 , n81345 , n81346 , n81347 , n81348 , n81349 , n81350 , 
     n81351 , n81352 , n81353 , n81354 , n81355 , n81356 , n81357 , n81358 , n81359 , n81360 , 
     n81361 , n81362 , n81363 , n81364 , n81365 , n81366 , n81367 , n81368 , n81369 , n81370 , 
     n81371 , n81372 , n81373 , n81374 , n81375 , n81376 , n81377 , n81378 , n81379 , n81380 , 
     n81381 , n81382 , n81383 , n81384 , n81385 , n81386 , n81387 , n81388 , n81389 , n81390 , 
     n81391 , n81392 , n81393 , n81394 , n81395 , n81396 , n81397 , n81398 , n81399 , n81400 , 
     n81401 , n81402 , n81403 , n81404 , n81405 , n81406 , n81407 , n81408 , n81409 , n81410 , 
     n81411 , n81412 , n81413 , n81414 , n81415 , n81416 , n81417 , n81418 , n81419 , n81420 , 
     n81421 , n81422 , n81423 , n81424 , n81425 , n81426 , n81427 , n81428 , n81429 , n81430 , 
     n81431 , n81432 , n81433 , n81434 , n81435 , n81436 , n81437 , n81438 , n81439 , n81440 , 
     n81441 , n81442 , n81443 , n81444 , n81445 , n81446 , n81447 , n81448 , n81449 , n81450 , 
     n81451 , n81452 , n81453 , n81454 , n81455 , n81456 , n81457 , n81458 , n81459 , n81460 , 
     n81461 , n81462 , n81463 , n81464 , n81465 , n81466 , n81467 , n81468 , n81469 , n81470 , 
     n81471 , n81472 , n81473 , n81474 , n81475 , n81476 , n81477 , n81478 , n81479 , n81480 , 
     n81481 , n81482 , n81483 , n81484 , n81485 , n81486 , n81487 , n81488 , n81489 , n81490 , 
     n81491 , n81492 , n81493 , n81494 , n81495 , n81496 , n81497 , n81498 , n81499 , n81500 , 
     n81501 , n81502 , n81503 , n81504 , n81505 , n81506 , n81507 , n81508 , n81509 , n81510 , 
     n81511 , n81512 , n81513 , n81514 , n81515 , n81516 , n81517 , n81518 , n81519 , n81520 , 
     n81521 , n81522 , n81523 , n81524 , n81525 , n81526 , n81527 , n81528 , n81529 , n81530 , 
     n81531 , n81532 , n81533 , n81534 , n81535 , n81536 , n81537 , n81538 , n81539 , n81540 , 
     n81541 , n81542 , n81543 , n81544 , n81545 , n81546 , n81547 , n81548 , n81549 , n81550 , 
     n81551 , n81552 , n81553 , n81554 , n81555 , n81556 , n81557 , n81558 , n81559 , n81560 , 
     n81561 , n81562 , n81563 , n81564 , n81565 , n81566 , n81567 , n81568 , n81569 , n81570 , 
     n81571 , n81572 , n81573 , n81574 , n81575 , n81576 , n81577 , n81578 , n81579 , n81580 , 
     n81581 , n81582 , n81583 , n81584 , n81585 , n81586 , n81587 , n81588 , n81589 , n81590 , 
     n81591 , n81592 , n81593 , n81594 , n81595 , n81596 , n81597 , n81598 , n81599 , n81600 , 
     n81601 , n81602 , n81603 , n81604 , n81605 , n81606 , n81607 , n81608 , n81609 , n81610 , 
     n81611 , n81612 , n81613 , n81614 , n81615 , n81616 , n81617 , n81618 , n81619 , n81620 , 
     n81621 , n81622 , n81623 , n81624 , n81625 , n81626 , n81627 , n81628 , n81629 , n81630 , 
     n81631 , n81632 , n81633 , n81634 , n81635 , n81636 , n81637 , n81638 , n81639 , n81640 , 
     n81641 , n81642 , n81643 , n81644 , n81645 , n81646 , n81647 , n81648 , n81649 , n81650 , 
     n81651 , n81652 , n81653 , n81654 , n81655 , n81656 , n81657 , n81658 , n81659 , n81660 , 
     n81661 , n81662 , n81663 , n81664 , n81665 , n81666 , n81667 , n81668 , n81669 , n81670 , 
     n81671 , n81672 , n81673 , n81674 , n81675 , n81676 , n81677 , n81678 , n81679 , n81680 , 
     n81681 , n81682 , n81683 , n81684 , n81685 , n81686 , n81687 , n81688 , n81689 , n81690 , 
     n81691 , n81692 , n81693 , n81694 , n81695 , n81696 , n81697 , n81698 , n81699 , n81700 , 
     n81701 , n81702 , n81703 , n81704 , n81705 , n81706 , n81707 , n81708 , n81709 , n81710 , 
     n81711 , n81712 , n81713 , n81714 , n81715 , n81716 , n81717 , n81718 , n81719 , n81720 , 
     n81721 , n81722 , n81723 , n81724 , n81725 , n81726 , n81727 , n81728 , n81729 , n81730 , 
     n81731 , n81732 , n81733 , n81734 , n81735 , n81736 , n81737 , n81738 , n81739 , n81740 , 
     n81741 , n81742 , n81743 , n81744 , n81745 , n81746 , n81747 , n81748 , n81749 , n81750 , 
     n81751 , n81752 , n81753 , n81754 , n81755 , n81756 , n81757 , n81758 , n81759 , n81760 , 
     n81761 , n81762 , n81763 , n81764 , n81765 , n81766 , n81767 , n81768 , n81769 , n81770 , 
     n81771 , n81772 , n81773 , n81774 , n81775 , n81776 , n81777 , n81778 , n81779 , n81780 , 
     n81781 , n81782 , n81783 , n81784 , n81785 , n81786 , n81787 , n81788 , n81789 , n81790 , 
     n81791 , n81792 , n81793 , n81794 , n81795 , n81796 , n81797 , n81798 , n81799 , n81800 , 
     n81801 , n81802 , n81803 , n81804 , n81805 , n81806 , n81807 , n81808 , n81809 , n81810 , 
     n81811 , n81812 , n81813 , n81814 , n81815 , n81816 , n81817 , n81818 , n81819 , n81820 , 
     n81821 , n81822 , n81823 , n81824 , n81825 , n81826 , n81827 , n81828 , n81829 , n81830 , 
     n81831 , n81832 , n81833 , n81834 , n81835 , n81836 , n81837 , n81838 , n81839 , n81840 , 
     n81841 , n81842 , n81843 , n81844 , n81845 , n81846 , n81847 , n81848 , n81849 , n81850 , 
     n81851 , n81852 , n81853 , n81854 , n81855 , n81856 , n81857 , n81858 , n81859 , n81860 , 
     n81861 , n81862 , n81863 , n81864 , n81865 , n81866 , n81867 , n81868 , n81869 , n81870 , 
     n81871 , n81872 , n81873 , n81874 , n81875 , n81876 , n81877 , n81878 , n81879 , n81880 , 
     n81881 , n81882 , n81883 , n81884 , n81885 , n81886 , n81887 , n81888 , n81889 , n81890 , 
     n81891 , n81892 , n81893 , n81894 , n81895 , n81896 , n81897 , n81898 , n81899 , n81900 , 
     n81901 , n81902 , n81903 , n81904 , n81905 , n81906 , n81907 , n81908 , n81909 , n81910 , 
     n81911 , n81912 , n81913 , n81914 , n81915 , n81916 , n81917 , n81918 , n81919 , n81920 , 
     n81921 , n81922 , n81923 , n81924 , n81925 , n81926 , n81927 , n81928 , n81929 , n81930 , 
     n81931 , n81932 , n81933 , n81934 , n81935 , n81936 , n81937 , n81938 , n81939 , n81940 , 
     n81941 , n81942 , n81943 , n81944 , n81945 , n81946 , n81947 , n81948 , n81949 , n81950 , 
     n81951 , n81952 , n81953 , n81954 , n81955 , n81956 , n81957 , n81958 , n81959 , n81960 , 
     n81961 , n81962 , n81963 , n81964 , n81965 , n81966 , n81967 , n81968 , n81969 , n81970 , 
     n81971 , n81972 , n81973 , n81974 , n81975 , n81976 , n81977 , n81978 , n81979 , n81980 , 
     n81981 , n81982 , n81983 , n81984 , n81985 , n81986 , n81987 , n81988 , n81989 , n81990 , 
     n81991 , n81992 , n81993 , n81994 , n81995 , n81996 , n81997 , n81998 , n81999 , n82000 , 
     n82001 , n82002 , n82003 , n82004 , n82005 , n82006 , n82007 , n82008 , n82009 , n82010 , 
     n82011 , n82012 , n82013 , n82014 , n82015 , n82016 , n82017 , n82018 , n82019 , n82020 , 
     n82021 , n82022 , n82023 , n82024 , n82025 , n82026 , n82027 , n82028 , n82029 , n82030 , 
     n82031 , n82032 , n82033 , n82034 , n82035 , n82036 , n82037 , n82038 , n82039 , n82040 , 
     n82041 , n82042 , n82043 , n82044 , n82045 , n82046 , n82047 , n82048 , n82049 , n82050 , 
     n82051 , n82052 , n82053 , n82054 , n82055 , n82056 , n82057 , n82058 , n82059 , n82060 , 
     n82061 , n82062 , n82063 , n82064 , n82065 , n82066 , n82067 , n82068 , n82069 , n82070 , 
     n82071 , n82072 , n82073 , n82074 , n82075 , n82076 , n82077 , n82078 , n82079 , n82080 , 
     n82081 , n82082 , n82083 , n82084 , n82085 , n82086 , n82087 , n82088 , n82089 , n82090 , 
     n82091 , n82092 , n82093 , n82094 , n82095 , n82096 , n82097 , n82098 , n82099 , n82100 , 
     n82101 , n82102 , n82103 , n82104 , n82105 , n82106 , n82107 , n82108 , n82109 , n82110 , 
     n82111 , n82112 , n82113 , n82114 , n82115 , n82116 , n82117 , n82118 , n82119 , n82120 , 
     n82121 , n82122 , n82123 , n82124 , n82125 , n82126 , n82127 , n82128 , n82129 , n82130 , 
     n82131 , n82132 , n82133 , n82134 , n82135 , n82136 , n82137 , n82138 , n82139 , n82140 , 
     n82141 , n82142 , n82143 , n82144 , n82145 , n82146 , n82147 , n82148 , n82149 , n82150 , 
     n82151 , n82152 , n82153 , n82154 , n82155 , n82156 , n82157 , n82158 , n82159 , n82160 , 
     n82161 , n82162 , n82163 , n82164 , n82165 , n82166 , n82167 , n82168 , n82169 , n82170 , 
     n82171 , n82172 , n82173 , n82174 , n82175 , n82176 , n82177 , n82178 , n82179 , n82180 , 
     n82181 , n82182 , n82183 , n82184 , n82185 , n82186 , n82187 , n82188 , n82189 , n82190 , 
     n82191 , n82192 , n82193 , n82194 , n82195 , n82196 , n82197 , n82198 , n82199 , n82200 , 
     n82201 , n82202 , n82203 , n82204 , n82205 , n82206 , n82207 , n82208 , n82209 , n82210 , 
     n82211 , n82212 , n82213 , n82214 , n82215 , n82216 , n82217 , n82218 , n82219 , n82220 , 
     n82221 , n82222 , n82223 , n82224 , n82225 , n82226 , n82227 , n82228 , n82229 , n82230 , 
     n82231 , n82232 , n82233 , n82234 , n82235 , n82236 , n82237 , n82238 , n82239 , n82240 , 
     n82241 , n82242 , n82243 , n82244 , n82245 , n82246 , n82247 , n82248 , n82249 , n82250 , 
     n82251 , n82252 , n82253 , n82254 , n82255 , n82256 , n82257 , n82258 , n82259 , n82260 , 
     n82261 , n82262 , n82263 , n82264 , n82265 , n82266 , n82267 , n82268 , n82269 , n82270 , 
     n82271 , n82272 , n82273 , n82274 , n82275 , n82276 , n82277 , n82278 , n82279 , n82280 , 
     n82281 , n82282 , n82283 , n82284 , n82285 , n82286 , n82287 , n82288 , n82289 , n82290 , 
     n82291 , n82292 , n82293 , n82294 , n82295 , n82296 , n82297 , n82298 , n82299 , n82300 , 
     n82301 , n82302 , n82303 , n82304 , n82305 , n82306 , n82307 , n82308 , n82309 , n82310 , 
     n82311 , n82312 , n82313 , n82314 , n82315 , n82316 , n82317 , n82318 , n82319 , n82320 , 
     n82321 , n82322 , n82323 , n82324 , n82325 , n82326 , n82327 , n82328 , n82329 , n82330 , 
     n82331 , n82332 , n82333 , n82334 , n82335 , n82336 , n82337 , n82338 , n82339 , n82340 , 
     n82341 , n82342 , n82343 , n82344 , n82345 , n82346 , n82347 , n82348 , n82349 , n82350 , 
     n82351 , n82352 , n82353 , n82354 , n82355 , n82356 , n82357 , n82358 , n82359 , n82360 , 
     n82361 , n82362 , n82363 , n82364 , n82365 , n82366 , n82367 , n82368 , n82369 , n82370 , 
     n82371 , n82372 , n82373 , n82374 , n82375 , n82376 , n82377 , n82378 , n82379 , n82380 , 
     n82381 , n82382 , n82383 , n82384 , n82385 , n82386 , n82387 , n82388 , n82389 , n82390 , 
     n82391 , n82392 , n82393 , n82394 , n82395 , n82396 , n82397 , n82398 , n82399 , n82400 , 
     n82401 , n82402 , n82403 , n82404 , n82405 , n82406 , n82407 , n82408 , n82409 , n82410 , 
     n82411 , n82412 , n82413 , n82414 , n82415 , n82416 , n82417 , n82418 , n82419 , n82420 , 
     n82421 , n82422 , n82423 , n82424 , n82425 , n82426 , n82427 , n82428 , n82429 , n82430 , 
     n82431 , n82432 , n82433 , n82434 , n82435 , n82436 , n82437 , n82438 , n82439 , n82440 , 
     n82441 , n82442 , n82443 , n82444 , n82445 , n82446 , n82447 , n82448 , n82449 , n82450 , 
     n82451 , n82452 , n82453 , n82454 , n82455 , n82456 , n82457 , n82458 , n82459 , n82460 , 
     n82461 , n82462 , n82463 , n82464 , n82465 , n82466 , n82467 , n82468 , n82469 , n82470 , 
     n82471 , n82472 , n82473 , n82474 , n82475 , n82476 , n82477 , n82478 , n82479 , n82480 , 
     n82481 , n82482 , n82483 , n82484 , n82485 , n82486 , n82487 , n82488 , n82489 , n82490 , 
     n82491 , n82492 , n82493 , n82494 , n82495 , n82496 , n82497 , n82498 , n82499 , n82500 , 
     n82501 , n82502 , n82503 , n82504 , n82505 , n82506 , n82507 , n82508 , n82509 , n82510 , 
     n82511 , n82512 , n82513 , n82514 , n82515 , n82516 , n82517 , n82518 , n82519 , n82520 , 
     n82521 , n82522 , n82523 , n82524 , n82525 , n82526 , n82527 , n82528 , n82529 , n82530 , 
     n82531 , n82532 , n82533 , n82534 , n82535 , n82536 , n82537 , n82538 , n82539 , n82540 , 
     n82541 , n82542 , n82543 , n82544 , n82545 , n82546 , n82547 , n82548 , n82549 , n82550 , 
     n82551 , n82552 , n82553 , n82554 , n82555 , n82556 , n82557 , n82558 , n82559 , n82560 , 
     n82561 , n82562 , n82563 , n82564 , n82565 , n82566 , n82567 , n82568 , n82569 , n82570 , 
     n82571 , n82572 , n82573 , n82574 , n82575 , n82576 , n82577 , n82578 , n82579 , n82580 , 
     n82581 , n82582 , n82583 , n82584 , n82585 , n82586 , n82587 , n82588 , n82589 , n82590 , 
     n82591 , n82592 , n82593 , n82594 , n82595 , n82596 , n82597 , n82598 , n82599 , n82600 , 
     n82601 , n82602 , n82603 , n82604 , n82605 , n82606 , n82607 , n82608 , n82609 , n82610 , 
     n82611 , n82612 , n82613 , n82614 , n82615 , n82616 , n82617 , n82618 , n82619 , n82620 , 
     n82621 , n82622 , n82623 , n82624 , n82625 , n82626 , n82627 , n82628 , n82629 , n82630 , 
     n82631 , n82632 , n82633 , n82634 , n82635 , n82636 , n82637 , n82638 , n82639 , n82640 , 
     n82641 , n82642 , n82643 , n82644 , n82645 , n82646 , n82647 , n82648 , n82649 , n82650 , 
     n82651 , n82652 , n82653 , n82654 , n82655 , n82656 , n82657 , n82658 , n82659 , n82660 , 
     n82661 , n82662 , n82663 , n82664 , n82665 , n82666 , n82667 , n82668 , n82669 , n82670 , 
     n82671 , n82672 , n82673 , n82674 , n82675 , n82676 , n82677 , n82678 , n82679 , n82680 , 
     n82681 , n82682 , n82683 , n82684 , n82685 , n82686 , n82687 , n82688 , n82689 , n82690 , 
     n82691 , n82692 , n82693 , n82694 , n82695 , n82696 , n82697 , n82698 , n82699 , n82700 , 
     n82701 , n82702 , n82703 , n82704 , n82705 , n82706 , n82707 , n82708 , n82709 , n82710 , 
     n82711 , n82712 , n82713 , n82714 , n82715 , n82716 , n82717 , n82718 , n82719 , n82720 , 
     n82721 , n82722 , n82723 , n82724 , n82725 , n82726 , n82727 , n82728 , n82729 , n82730 , 
     n82731 , n82732 , n82733 , n82734 , n82735 , n82736 , n82737 , n82738 , n82739 , n82740 , 
     n82741 , n82742 , n82743 , n82744 , n82745 , n82746 , n82747 , n82748 , n82749 , n82750 , 
     n82751 , n82752 , n82753 , n82754 , n82755 , n82756 , n82757 , n82758 , n82759 , n82760 , 
     n82761 , n82762 , n82763 , n82764 , n82765 , n82766 , n82767 , n82768 , n82769 , n82770 , 
     n82771 , n82772 , n82773 , n82774 , n82775 , n82776 , n82777 , n82778 , n82779 , n82780 , 
     n82781 , n82782 , n82783 , n82784 , n82785 , n82786 , n82787 , n82788 , n82789 , n82790 , 
     n82791 , n82792 , n82793 , n82794 , n82795 , n82796 , n82797 , n82798 , n82799 , n82800 , 
     n82801 , n82802 , n82803 , n82804 , n82805 , n82806 , n82807 , n82808 , n82809 , n82810 , 
     n82811 , n82812 , n82813 , n82814 , n82815 , n82816 , n82817 , n82818 , n82819 , n82820 , 
     n82821 , n82822 , n82823 , n82824 , n82825 , n82826 , n82827 , n82828 , n82829 , n82830 , 
     n82831 , n82832 , n82833 , n82834 , n82835 , n82836 , n82837 , n82838 , n82839 , n82840 , 
     n82841 , n82842 , n82843 , n82844 , n82845 , n82846 , n82847 , n82848 , n82849 , n82850 , 
     n82851 , n82852 , n82853 , n82854 , n82855 , n82856 , n82857 , n82858 , n82859 , n82860 , 
     n82861 , n82862 , n82863 , n82864 , n82865 , n82866 , n82867 , n82868 , n82869 , n82870 , 
     n82871 , n82872 , n82873 , n82874 , n82875 , n82876 , n82877 , n82878 , n82879 , n82880 , 
     n82881 , n82882 , n82883 , n82884 , n82885 , n82886 , n82887 , n82888 , n82889 , n82890 , 
     n82891 , n82892 , n82893 , n82894 , n82895 , n82896 , n82897 , n82898 , n82899 , n82900 , 
     n82901 , n82902 , n82903 , n82904 , n82905 , n82906 , n82907 , n82908 , n82909 , n82910 , 
     n82911 , n82912 , n82913 , n82914 , n82915 , n82916 , n82917 , n82918 , n82919 , n82920 , 
     n82921 , n82922 , n82923 , n82924 , n82925 , n82926 , n82927 , n82928 , n82929 , n82930 , 
     n82931 , n82932 , n82933 , n82934 , n82935 , n82936 , n82937 , n82938 , n82939 , n82940 , 
     n82941 , n82942 , n82943 , n82944 , n82945 , n82946 , n82947 , n82948 , n82949 , n82950 , 
     n82951 , n82952 , n82953 , n82954 , n82955 , n82956 , n82957 , n82958 , n82959 , n82960 , 
     n82961 , n82962 , n82963 , n82964 , n82965 , n82966 , n82967 , n82968 , n82969 , n82970 , 
     n82971 , n82972 , n82973 , n82974 , n82975 , n82976 , n82977 , n82978 , n82979 , n82980 , 
     n82981 , n82982 , n82983 , n82984 , n82985 , n82986 , n82987 , n82988 , n82989 , n82990 , 
     n82991 , n82992 , n82993 , n82994 , n82995 , n82996 , n82997 , n82998 , n82999 , n83000 , 
     n83001 , n83002 , n83003 , n83004 , n83005 , n83006 , n83007 , n83008 , n83009 , n83010 , 
     n83011 , n83012 , n83013 , n83014 , n83015 , n83016 , n83017 , n83018 , n83019 , n83020 , 
     n83021 , n83022 , n83023 , n83024 , n83025 , n83026 , n83027 , n83028 , n83029 , n83030 , 
     n83031 , n83032 , n83033 , n83034 , n83035 , n83036 , n83037 , n83038 , n83039 , n83040 , 
     n83041 , n83042 , n83043 , n83044 , n83045 , n83046 , n83047 , n83048 , n83049 , n83050 , 
     n83051 , n83052 , n83053 , n83054 , n83055 , n83056 , n83057 , n83058 , n83059 , n83060 , 
     n83061 , n83062 , n83063 , n83064 , n83065 , n83066 , n83067 , n83068 , n83069 , n83070 , 
     n83071 , n83072 , n83073 , n83074 , n83075 , n83076 , n83077 , n83078 , n83079 , n83080 , 
     n83081 , n83082 , n83083 , n83084 , n83085 , n83086 , n83087 , n83088 , n83089 , n83090 , 
     n83091 , n83092 , n83093 , n83094 , n83095 , n83096 , n83097 , n83098 , n83099 , n83100 , 
     n83101 , n83102 , n83103 , n83104 , n83105 , n83106 , n83107 , n83108 , n83109 , n83110 , 
     n83111 , n83112 , n83113 , n83114 , n83115 , n83116 , n83117 , n83118 , n83119 , n83120 , 
     n83121 , n83122 , n83123 , n83124 , n83125 , n83126 , n83127 , n83128 , n83129 , n83130 , 
     n83131 , n83132 , n83133 , n83134 , n83135 , n83136 , n83137 , n83138 , n83139 , n83140 , 
     n83141 , n83142 , n83143 , n83144 , n83145 , n83146 , n83147 , n83148 , n83149 , n83150 , 
     n83151 , n83152 , n83153 , n83154 , n83155 , n83156 , n83157 , n83158 , n83159 , n83160 , 
     n83161 , n83162 , n83163 , n83164 , n83165 , n83166 , n83167 , n83168 , n83169 , n83170 , 
     n83171 , n83172 , n83173 , n83174 , n83175 , n83176 , n83177 , n83178 , n83179 , n83180 , 
     n83181 , n83182 , n83183 , n83184 , n83185 , n83186 , n83187 , n83188 , n83189 , n83190 , 
     n83191 , n83192 , n83193 , n83194 , n83195 , n83196 , n83197 , n83198 , n83199 , n83200 , 
     n83201 , n83202 , n83203 , n83204 , n83205 , n83206 , n83207 , n83208 , n83209 , n83210 , 
     n83211 , n83212 , n83213 , n83214 , n83215 , n83216 , n83217 , n83218 , n83219 , n83220 , 
     n83221 , n83222 , n83223 , n83224 , n83225 , n83226 , n83227 , n83228 , n83229 , n83230 , 
     n83231 , n83232 , n83233 , n83234 , n83235 , n83236 , n83237 , n83238 , n83239 , n83240 , 
     n83241 , n83242 , n83243 , n83244 , n83245 , n83246 , n83247 , n83248 , n83249 , n83250 , 
     n83251 , n83252 , n83253 , n83254 , n83255 , n83256 , n83257 , n83258 , n83259 , n83260 , 
     n83261 , n83262 , n83263 , n83264 , n83265 , n83266 , n83267 , n83268 , n83269 , n83270 , 
     n83271 , n83272 , n83273 , n83274 , n83275 , n83276 , n83277 , n83278 , n83279 , n83280 , 
     n83281 , n83282 , n83283 , n83284 , n83285 , n83286 , n83287 , n83288 , n83289 , n83290 , 
     n83291 , n83292 , n83293 , n83294 , n83295 , n83296 , n83297 , n83298 , n83299 , n83300 , 
     n83301 , n83302 , n83303 , n83304 , n83305 , n83306 , n83307 , n83308 , n83309 , n83310 , 
     n83311 , n83312 , n83313 , n83314 , n83315 , n83316 , n83317 , n83318 , n83319 , n83320 , 
     n83321 , n83322 , n83323 , n83324 , n83325 , n83326 , n83327 , n83328 , n83329 , n83330 , 
     n83331 , n83332 , n83333 , n83334 , n83335 , n83336 , n83337 , n83338 , n83339 , n83340 , 
     n83341 , n83342 , n83343 , n83344 , n83345 , n83346 , n83347 , n83348 , n83349 , n83350 , 
     n83351 , n83352 , n83353 , n83354 , n83355 , n83356 , n83357 , n83358 , n83359 , n83360 , 
     n83361 , n83362 , n83363 , n83364 , n83365 , n83366 , n83367 , n83368 , n83369 , n83370 , 
     n83371 , n83372 , n83373 , n83374 , n83375 , n83376 , n83377 , n83378 , n83379 , n83380 , 
     n83381 , n83382 , n83383 , n83384 , n83385 , n83386 , n83387 , n83388 , n83389 , n83390 , 
     n83391 , n83392 , n83393 , n83394 , n83395 , n83396 , n83397 , n83398 , n83399 , n83400 , 
     n83401 , n83402 , n83403 , n83404 , n83405 , n83406 , n83407 , n83408 , n83409 , n83410 , 
     n83411 , n83412 , n83413 , n83414 , n83415 , n83416 , n83417 , n83418 , n83419 , n83420 , 
     n83421 , n83422 , n83423 , n83424 , n83425 , n83426 , n83427 , n83428 , n83429 , n83430 , 
     n83431 , n83432 , n83433 , n83434 , n83435 , n83436 , n83437 , n83438 , n83439 , n83440 , 
     n83441 , n83442 , n83443 , n83444 , n83445 , n83446 , n83447 , n83448 , n83449 , n83450 , 
     n83451 , n83452 , n83453 , n83454 , n83455 , n83456 , n83457 , n83458 , n83459 , n83460 , 
     n83461 , n83462 , n83463 , n83464 , n83465 , n83466 , n83467 , n83468 , n83469 , n83470 , 
     n83471 , n83472 , n83473 , n83474 , n83475 , n83476 , n83477 , n83478 , n83479 , n83480 , 
     n83481 , n83482 , n83483 , n83484 , n83485 , n83486 , n83487 , n83488 , n83489 , n83490 , 
     n83491 , n83492 , n83493 , n83494 , n83495 , n83496 , n83497 , n83498 , n83499 , n83500 , 
     n83501 , n83502 , n83503 , n83504 , n83505 , n83506 , n83507 , n83508 , n83509 , n83510 , 
     n83511 , n83512 , n83513 , n83514 , n83515 , n83516 , n83517 , n83518 , n83519 , n83520 , 
     n83521 , n83522 , n83523 , n83524 , n83525 , n83526 , n83527 , n83528 , n83529 , n83530 , 
     n83531 , n83532 , n83533 , n83534 , n83535 , n83536 , n83537 , n83538 , n83539 , n83540 , 
     n83541 , n83542 , n83543 , n83544 , n83545 , n83546 , n83547 , n83548 , n83549 , n83550 , 
     n83551 , n83552 , n83553 , n83554 , n83555 , n83556 , n83557 , n83558 , n83559 , n83560 , 
     n83561 , n83562 , n83563 , n83564 , n83565 , n83566 , n83567 , n83568 , n83569 , n83570 , 
     n83571 , n83572 , n83573 , n83574 , n83575 , n83576 , n83577 , n83578 , n83579 , n83580 , 
     n83581 , n83582 , n83583 , n83584 , n83585 , n83586 , n83587 , n83588 , n83589 , n83590 , 
     n83591 , n83592 , n83593 , n83594 , n83595 , n83596 , n83597 , n83598 , n83599 , n83600 , 
     n83601 , n83602 , n83603 , n83604 , n83605 , n83606 , n83607 , n83608 , n83609 , n83610 , 
     n83611 , n83612 , n83613 , n83614 , n83615 , n83616 , n83617 , n83618 , n83619 , n83620 , 
     n83621 , n83622 , n83623 , n83624 , n83625 , n83626 , n83627 , n83628 , n83629 , n83630 , 
     n83631 , n83632 , n83633 , n83634 , n83635 , n83636 , n83637 , n83638 , n83639 , n83640 , 
     n83641 , n83642 , n83643 , n83644 , n83645 , n83646 , n83647 , n83648 , n83649 , n83650 , 
     n83651 , n83652 , n83653 , n83654 , n83655 , n83656 , n83657 , n83658 , n83659 , n83660 , 
     n83661 , n83662 , n83663 , n83664 , n83665 , n83666 , n83667 , n83668 , n83669 , n83670 , 
     n83671 , n83672 , n83673 , n83674 , n83675 , n83676 , n83677 , n83678 , n83679 , n83680 , 
     n83681 , n83682 , n83683 , n83684 , n83685 , n83686 , n83687 , n83688 , n83689 , n83690 , 
     n83691 , n83692 , n83693 , n83694 , n83695 , n83696 , n83697 , n83698 , n83699 , n83700 , 
     n83701 , n83702 , n83703 , n83704 , n83705 , n83706 , n83707 , n83708 , n83709 , n83710 , 
     n83711 , n83712 , n83713 , n83714 , n83715 , n83716 , n83717 , n83718 , n83719 , n83720 , 
     n83721 , n83722 , n83723 , n83724 , n83725 , n83726 , n83727 , n83728 , n83729 , n83730 , 
     n83731 , n83732 , n83733 , n83734 , n83735 , n83736 , n83737 , n83738 , n83739 , n83740 , 
     n83741 , n83742 , n83743 , n83744 , n83745 , n83746 , n83747 , n83748 , n83749 , n83750 , 
     n83751 , n83752 , n83753 , n83754 , n83755 , n83756 , n83757 , n83758 , n83759 , n83760 , 
     n83761 , n83762 , n83763 , n83764 , n83765 , n83766 , n83767 , n83768 , n83769 , n83770 , 
     n83771 , n83772 , n83773 , n83774 , n83775 , n83776 , n83777 , n83778 , n83779 , n83780 , 
     n83781 , n83782 , n83783 , n83784 , n83785 , n83786 , n83787 , n83788 , n83789 , n83790 , 
     n83791 , n83792 , n83793 , n83794 , n83795 , n83796 , n83797 , n83798 , n83799 , n83800 , 
     n83801 , n83802 , n83803 , n83804 , n83805 , n83806 , n83807 , n83808 , n83809 , n83810 , 
     n83811 , n83812 , n83813 , n83814 , n83815 , n83816 , n83817 , n83818 , n83819 , n83820 , 
     n83821 , n83822 , n83823 , n83824 , n83825 , n83826 , n83827 , n83828 , n83829 , n83830 , 
     n83831 , n83832 , n83833 , n83834 , n83835 , n83836 , n83837 , n83838 , n83839 , n83840 , 
     n83841 , n83842 , n83843 , n83844 , n83845 , n83846 , n83847 , n83848 , n83849 , n83850 , 
     n83851 , n83852 , n83853 , n83854 , n83855 , n83856 , n83857 , n83858 , n83859 , n83860 , 
     n83861 , n83862 , n83863 , n83864 , n83865 , n83866 , n83867 , n83868 , n83869 , n83870 , 
     n83871 , n83872 , n83873 , n83874 , n83875 , n83876 , n83877 , n83878 , n83879 , n83880 , 
     n83881 , n83882 , n83883 , n83884 , n83885 , n83886 , n83887 , n83888 , n83889 , n83890 , 
     n83891 , n83892 , n83893 , n83894 , n83895 , n83896 , n83897 , n83898 , n83899 , n83900 , 
     n83901 , n83902 , n83903 , n83904 , n83905 , n83906 , n83907 , n83908 , n83909 , n83910 , 
     n83911 , n83912 , n83913 , n83914 , n83915 , n83916 , n83917 , n83918 , n83919 , n83920 , 
     n83921 , n83922 , n83923 , n83924 , n83925 , n83926 , n83927 , n83928 , n83929 , n83930 , 
     n83931 , n83932 , n83933 , n83934 , n83935 , n83936 , n83937 , n83938 , n83939 , n83940 , 
     n83941 , n83942 , n83943 , n83944 , n83945 , n83946 , n83947 , n83948 , n83949 , n83950 , 
     n83951 , n83952 , n83953 , n83954 , n83955 , n83956 , n83957 , n83958 , n83959 , n83960 , 
     n83961 , n83962 , n83963 , n83964 , n83965 , n83966 , n83967 , n83968 , n83969 , n83970 , 
     n83971 , n83972 , n83973 , n83974 , n83975 , n83976 , n83977 , n83978 , n83979 , n83980 , 
     n83981 , n83982 , n83983 , n83984 , n83985 , n83986 , n83987 , n83988 , n83989 , n83990 , 
     n83991 , n83992 , n83993 , n83994 , n83995 , n83996 , n83997 , n83998 , n83999 , n84000 , 
     n84001 , n84002 , n84003 , n84004 , n84005 , n84006 , n84007 , n84008 , n84009 , n84010 , 
     n84011 , n84012 , n84013 , n84014 , n84015 , n84016 , n84017 , n84018 , n84019 , n84020 , 
     n84021 , n84022 , n84023 , n84024 , n84025 , n84026 , n84027 , n84028 , n84029 , n84030 , 
     n84031 , n84032 , n84033 , n84034 , n84035 , n84036 , n84037 , n84038 , n84039 , n84040 , 
     n84041 , n84042 , n84043 , n84044 , n84045 , n84046 , n84047 , n84048 , n84049 , n84050 , 
     n84051 , n84052 , n84053 , n84054 , n84055 , n84056 , n84057 , n84058 , n84059 , n84060 , 
     n84061 , n84062 , n84063 , n84064 , n84065 , n84066 , n84067 , n84068 , n84069 , n84070 , 
     n84071 , n84072 , n84073 , n84074 , n84075 , n84076 , n84077 , n84078 , n84079 , n84080 , 
     n84081 , n84082 , n84083 , n84084 , n84085 , n84086 , n84087 , n84088 , n84089 , n84090 , 
     n84091 , n84092 , n84093 , n84094 , n84095 , n84096 , n84097 , n84098 , n84099 , n84100 , 
     n84101 , n84102 , n84103 , n84104 , n84105 , n84106 , n84107 , n84108 , n84109 , n84110 , 
     n84111 , n84112 , n84113 , n84114 , n84115 , n84116 , n84117 , n84118 , n84119 , n84120 , 
     n84121 , n84122 , n84123 , n84124 , n84125 , n84126 , n84127 , n84128 , n84129 , n84130 , 
     n84131 , n84132 , n84133 , n84134 , n84135 , n84136 , n84137 , n84138 , n84139 , n84140 , 
     n84141 , n84142 , n84143 , n84144 , n84145 , n84146 , n84147 , n84148 , n84149 , n84150 , 
     n84151 , n84152 , n84153 , n84154 , n84155 , n84156 , n84157 , n84158 , n84159 , n84160 , 
     n84161 , n84162 , n84163 , n84164 , n84165 , n84166 , n84167 , n84168 , n84169 , n84170 , 
     n84171 , n84172 , n84173 , n84174 , n84175 , n84176 , n84177 , n84178 , n84179 , n84180 , 
     n84181 , n84182 , n84183 , n84184 , n84185 , n84186 , n84187 , n84188 , n84189 , n84190 , 
     n84191 , n84192 , n84193 , n84194 , n84195 , n84196 , n84197 , n84198 , n84199 , n84200 , 
     n84201 , n84202 , n84203 , n84204 , n84205 , n84206 , n84207 , n84208 , n84209 , n84210 , 
     n84211 , n84212 , n84213 , n84214 , n84215 , n84216 , n84217 , n84218 , n84219 , n84220 , 
     n84221 , n84222 , n84223 , n84224 , n84225 , n84226 , n84227 , n84228 , n84229 , n84230 , 
     n84231 , n84232 , n84233 , n84234 , n84235 , n84236 , n84237 , n84238 , n84239 , n84240 , 
     n84241 , n84242 , n84243 , n84244 , n84245 , n84246 , n84247 , n84248 , n84249 , n84250 , 
     n84251 , n84252 , n84253 , n84254 , n84255 , n84256 , n84257 , n84258 , n84259 , n84260 , 
     n84261 , n84262 , n84263 , n84264 , n84265 , n84266 , n84267 , n84268 , n84269 , n84270 , 
     n84271 , n84272 , n84273 , n84274 , n84275 , n84276 , n84277 , n84278 , n84279 , n84280 , 
     n84281 , n84282 , n84283 , n84284 , n84285 , n84286 , n84287 , n84288 , n84289 , n84290 , 
     n84291 , n84292 , n84293 , n84294 , n84295 , n84296 , n84297 , n84298 , n84299 , n84300 , 
     n84301 , n84302 , n84303 , n84304 , n84305 , n84306 , n84307 , n84308 , n84309 , n84310 , 
     n84311 , n84312 , n84313 , n84314 , n84315 , n84316 , n84317 , n84318 , n84319 , n84320 , 
     n84321 , n84322 , n84323 , n84324 , n84325 , n84326 , n84327 , n84328 , n84329 , n84330 , 
     n84331 , n84332 , n84333 , n84334 , n84335 , n84336 , n84337 , n84338 , n84339 , n84340 , 
     n84341 , n84342 , n84343 , n84344 , n84345 , n84346 , n84347 , n84348 , n84349 , n84350 , 
     n84351 , n84352 , n84353 , n84354 , n84355 , n84356 , n84357 , n84358 , n84359 , n84360 , 
     n84361 , n84362 , n84363 , n84364 , n84365 , n84366 , n84367 , n84368 , n84369 , n84370 , 
     n84371 , n84372 , n84373 , n84374 , n84375 , n84376 , n84377 , n84378 , n84379 , n84380 , 
     n84381 , n84382 , n84383 , n84384 , n84385 , n84386 , n84387 , n84388 , n84389 , n84390 , 
     n84391 , n84392 , n84393 , n84394 , n84395 , n84396 , n84397 , n84398 , n84399 , n84400 , 
     n84401 , n84402 , n84403 , n84404 , n84405 , n84406 , n84407 , n84408 , n84409 , n84410 , 
     n84411 , n84412 , n84413 , n84414 , n84415 , n84416 , n84417 , n84418 , n84419 , n84420 , 
     n84421 , n84422 , n84423 , n84424 , n84425 , n84426 , n84427 , n84428 , n84429 , n84430 , 
     n84431 , n84432 , n84433 , n84434 , n84435 , n84436 , n84437 , n84438 , n84439 , n84440 , 
     n84441 , n84442 , n84443 , n84444 , n84445 , n84446 , n84447 , n84448 , n84449 , n84450 , 
     n84451 , n84452 , n84453 , n84454 , n84455 , n84456 , n84457 , n84458 , n84459 , n84460 , 
     n84461 , n84462 , n84463 , n84464 , n84465 , n84466 , n84467 , n84468 , n84469 , n84470 , 
     n84471 , n84472 , n84473 , n84474 , n84475 , n84476 , n84477 , n84478 , n84479 , n84480 , 
     n84481 , n84482 , n84483 , n84484 , n84485 , n84486 , n84487 , n84488 , n84489 , n84490 , 
     n84491 , n84492 , n84493 , n84494 , n84495 , n84496 , n84497 , n84498 , n84499 , n84500 , 
     n84501 , n84502 , n84503 , n84504 , n84505 , n84506 , n84507 , n84508 , n84509 , n84510 , 
     n84511 , n84512 , n84513 , n84514 , n84515 , n84516 , n84517 , n84518 , n84519 , n84520 , 
     n84521 , n84522 , n84523 , n84524 , n84525 , n84526 , n84527 , n84528 , n84529 , n84530 , 
     n84531 , n84532 , n84533 , n84534 , n84535 , n84536 , n84537 , n84538 , n84539 , n84540 , 
     n84541 , n84542 , n84543 , n84544 , n84545 , n84546 , n84547 , n84548 , n84549 , n84550 , 
     n84551 , n84552 , n84553 , n84554 , n84555 , n84556 , n84557 , n84558 , n84559 , n84560 , 
     n84561 , n84562 , n84563 , n84564 , n84565 , n84566 , n84567 , n84568 , n84569 , n84570 , 
     n84571 , n84572 , n84573 , n84574 , n84575 , n84576 , n84577 , n84578 , n84579 , n84580 , 
     n84581 , n84582 , n84583 , n84584 , n84585 , n84586 , n84587 , n84588 , n84589 , n84590 , 
     n84591 , n84592 , n84593 , n84594 , n84595 , n84596 , n84597 , n84598 , n84599 , n84600 , 
     n84601 , n84602 , n84603 , n84604 , n84605 , n84606 , n84607 , n84608 , n84609 , n84610 , 
     n84611 , n84612 , n84613 , n84614 , n84615 , n84616 , n84617 , n84618 , n84619 , n84620 , 
     n84621 , n84622 , n84623 , n84624 , n84625 , n84626 , n84627 , n84628 , n84629 , n84630 , 
     n84631 , n84632 , n84633 , n84634 , n84635 , n84636 , n84637 , n84638 , n84639 , n84640 , 
     n84641 , n84642 , n84643 , n84644 , n84645 , n84646 , n84647 , n84648 , n84649 , n84650 , 
     n84651 , n84652 , n84653 , n84654 , n84655 , n84656 , n84657 , n84658 , n84659 , n84660 , 
     n84661 , n84662 , n84663 , n84664 , n84665 , n84666 , n84667 , n84668 , n84669 , n84670 , 
     n84671 , n84672 , n84673 , n84674 , n84675 , n84676 , n84677 , n84678 , n84679 , n84680 , 
     n84681 , n84682 , n84683 , n84684 , n84685 , n84686 , n84687 , n84688 , n84689 , n84690 , 
     n84691 , n84692 , n84693 , n84694 , n84695 , n84696 , n84697 , n84698 , n84699 , n84700 , 
     n84701 , n84702 , n84703 , n84704 , n84705 , n84706 , n84707 , n84708 , n84709 , n84710 , 
     n84711 , n84712 , n84713 , n84714 , n84715 , n84716 , n84717 , n84718 , n84719 , n84720 , 
     n84721 , n84722 , n84723 , n84724 , n84725 , n84726 , n84727 , n84728 , n84729 , n84730 , 
     n84731 , n84732 , n84733 , n84734 , n84735 , n84736 , n84737 , n84738 , n84739 , n84740 , 
     n84741 , n84742 , n84743 , n84744 , n84745 , n84746 , n84747 , n84748 , n84749 , n84750 , 
     n84751 , n84752 , n84753 , n84754 , n84755 , n84756 , n84757 , n84758 , n84759 , n84760 , 
     n84761 , n84762 , n84763 , n84764 , n84765 , n84766 , n84767 , n84768 , n84769 , n84770 , 
     n84771 , n84772 , n84773 , n84774 , n84775 , n84776 , n84777 , n84778 , n84779 , n84780 , 
     n84781 , n84782 , n84783 , n84784 , n84785 , n84786 , n84787 , n84788 , n84789 , n84790 , 
     n84791 , n84792 , n84793 , n84794 , n84795 , n84796 , n84797 , n84798 , n84799 , n84800 , 
     n84801 , n84802 , n84803 , n84804 , n84805 , n84806 , n84807 , n84808 , n84809 , n84810 , 
     n84811 , n84812 , n84813 , n84814 , n84815 , n84816 , n84817 , n84818 , n84819 , n84820 , 
     n84821 , n84822 , n84823 , n84824 , n84825 , n84826 , n84827 , n84828 , n84829 , n84830 , 
     n84831 , n84832 , n84833 , n84834 , n84835 , n84836 , n84837 , n84838 , n84839 , n84840 , 
     n84841 , n84842 , n84843 , n84844 , n84845 , n84846 , n84847 , n84848 , n84849 , n84850 , 
     n84851 , n84852 , n84853 , n84854 , n84855 , n84856 , n84857 , n84858 , n84859 , n84860 , 
     n84861 , n84862 , n84863 , n84864 , n84865 , n84866 , n84867 , n84868 , n84869 , n84870 , 
     n84871 , n84872 , n84873 , n84874 , n84875 , n84876 , n84877 , n84878 , n84879 , n84880 , 
     n84881 , n84882 , n84883 , n84884 , n84885 , n84886 , n84887 , n84888 , n84889 , n84890 , 
     n84891 , n84892 , n84893 , n84894 , n84895 , n84896 , n84897 , n84898 , n84899 , n84900 , 
     n84901 , n84902 , n84903 , n84904 , n84905 , n84906 , n84907 , n84908 , n84909 , n84910 , 
     n84911 , n84912 , n84913 , n84914 , n84915 , n84916 , n84917 , n84918 , n84919 , n84920 , 
     n84921 , n84922 , n84923 , n84924 , n84925 , n84926 , n84927 , n84928 , n84929 , n84930 , 
     n84931 , n84932 , n84933 , n84934 , n84935 , n84936 , n84937 , n84938 , n84939 , n84940 , 
     n84941 , n84942 , n84943 , n84944 , n84945 , n84946 , n84947 , n84948 , n84949 , n84950 , 
     n84951 , n84952 , n84953 , n84954 , n84955 , n84956 , n84957 , n84958 , n84959 , n84960 , 
     n84961 , n84962 , n84963 , n84964 , n84965 , n84966 , n84967 , n84968 , n84969 , n84970 , 
     n84971 , n84972 , n84973 , n84974 , n84975 , n84976 , n84977 , n84978 , n84979 , n84980 , 
     n84981 , n84982 , n84983 , n84984 , n84985 , n84986 , n84987 , n84988 , n84989 , n84990 , 
     n84991 , n84992 , n84993 , n84994 , n84995 , n84996 , n84997 , n84998 , n84999 , n85000 , 
     n85001 , n85002 , n85003 , n85004 , n85005 , n85006 , n85007 , n85008 , n85009 , n85010 , 
     n85011 , n85012 , n85013 , n85014 , n85015 , n85016 , n85017 , n85018 , n85019 , n85020 , 
     n85021 , n85022 , n85023 , n85024 , n85025 , n85026 , n85027 , n85028 , n85029 , n85030 , 
     n85031 , n85032 , n85033 , n85034 , n85035 , n85036 , n85037 , n85038 , n85039 , n85040 , 
     n85041 , n85042 , n85043 , n85044 , n85045 , n85046 , n85047 , n85048 , n85049 , n85050 , 
     n85051 , n85052 , n85053 , n85054 , n85055 , n85056 , n85057 , n85058 , n85059 , n85060 , 
     n85061 , n85062 , n85063 , n85064 , n85065 , n85066 , n85067 , n85068 , n85069 , n85070 , 
     n85071 , n85072 , n85073 , n85074 , n85075 , n85076 , n85077 , n85078 , n85079 , n85080 , 
     n85081 , n85082 , n85083 , n85084 , n85085 , n85086 , n85087 , n85088 , n85089 , n85090 , 
     n85091 , n85092 , n85093 , n85094 , n85095 , n85096 , n85097 , n85098 , n85099 , n85100 , 
     n85101 , n85102 , n85103 , n85104 , n85105 , n85106 , n85107 , n85108 , n85109 , n85110 , 
     n85111 , n85112 , n85113 , n85114 , n85115 , n85116 , n85117 , n85118 , n85119 , n85120 , 
     n85121 , n85122 , n85123 , n85124 , n85125 , n85126 , n85127 , n85128 , n85129 , n85130 , 
     n85131 , n85132 , n85133 , n85134 , n85135 , n85136 , n85137 , n85138 , n85139 , n85140 , 
     n85141 , n85142 , n85143 , n85144 , n85145 , n85146 , n85147 , n85148 , n85149 , n85150 , 
     n85151 , n85152 , n85153 , n85154 , n85155 , n85156 , n85157 , n85158 , n85159 , n85160 , 
     n85161 , n85162 , n85163 , n85164 , n85165 , n85166 , n85167 , n85168 , n85169 , n85170 , 
     n85171 , n85172 , n85173 , n85174 , n85175 , n85176 , n85177 , n85178 , n85179 , n85180 , 
     n85181 , n85182 , n85183 , n85184 , n85185 , n85186 , n85187 , n85188 , n85189 , n85190 , 
     n85191 , n85192 , n85193 , n85194 , n85195 , n85196 , n85197 , n85198 , n85199 , n85200 , 
     n85201 , n85202 , n85203 , n85204 , n85205 , n85206 , n85207 , n85208 , n85209 , n85210 , 
     n85211 , n85212 , n85213 , n85214 , n85215 , n85216 , n85217 , n85218 , n85219 , n85220 , 
     n85221 , n85222 , n85223 , n85224 , n85225 , n85226 , n85227 , n85228 , n85229 , n85230 , 
     n85231 , n85232 , n85233 , n85234 , n85235 , n85236 , n85237 , n85238 , n85239 , n85240 , 
     n85241 , n85242 , n85243 , n85244 , n85245 , n85246 , n85247 , n85248 , n85249 , n85250 , 
     n85251 , n85252 , n85253 , n85254 , n85255 , n85256 , n85257 , n85258 , n85259 , n85260 , 
     n85261 , n85262 , n85263 , n85264 , n85265 , n85266 , n85267 , n85268 , n85269 , n85270 , 
     n85271 , n85272 , n85273 , n85274 , n85275 , n85276 , n85277 , n85278 , n85279 , n85280 , 
     n85281 , n85282 , n85283 , n85284 , n85285 , n85286 , n85287 , n85288 , n85289 , n85290 , 
     n85291 , n85292 , n85293 , n85294 , n85295 , n85296 , n85297 , n85298 , n85299 , n85300 , 
     n85301 , n85302 , n85303 , n85304 , n85305 , n85306 , n85307 , n85308 , n85309 , n85310 , 
     n85311 , n85312 , n85313 , n85314 , n85315 , n85316 , n85317 , n85318 , n85319 , n85320 , 
     n85321 , n85322 , n85323 , n85324 , n85325 , n85326 , n85327 , n85328 , n85329 , n85330 , 
     n85331 , n85332 , n85333 , n85334 , n85335 , n85336 , n85337 , n85338 , n85339 , n85340 , 
     n85341 , n85342 , n85343 , n85344 , n85345 , n85346 , n85347 , n85348 , n85349 , n85350 , 
     n85351 , n85352 , n85353 , n85354 , n85355 , n85356 , n85357 , n85358 , n85359 , n85360 , 
     n85361 , n85362 , n85363 , n85364 , n85365 , n85366 , n85367 , n85368 , n85369 , n85370 , 
     n85371 , n85372 , n85373 , n85374 , n85375 , n85376 , n85377 , n85378 , n85379 , n85380 , 
     n85381 , n85382 , n85383 , n85384 , n85385 , n85386 , n85387 , n85388 , n85389 , n85390 , 
     n85391 , n85392 , n85393 , n85394 , n85395 , n85396 , n85397 , n85398 , n85399 , n85400 , 
     n85401 , n85402 , n85403 , n85404 , n85405 , n85406 , n85407 , n85408 , n85409 , n85410 , 
     n85411 , n85412 , n85413 , n85414 , n85415 , n85416 , n85417 , n85418 , n85419 , n85420 , 
     n85421 , n85422 , n85423 , n85424 , n85425 , n85426 , n85427 , n85428 , n85429 , n85430 , 
     n85431 , n85432 , n85433 , n85434 , n85435 , n85436 , n85437 , n85438 , n85439 , n85440 , 
     n85441 , n85442 , n85443 , n85444 , n85445 , n85446 , n85447 , n85448 , n85449 , n85450 , 
     n85451 , n85452 , n85453 , n85454 , n85455 , n85456 , n85457 , n85458 , n85459 , n85460 , 
     n85461 , n85462 , n85463 , n85464 , n85465 , n85466 , n85467 , n85468 , n85469 , n85470 , 
     n85471 , n85472 , n85473 , n85474 , n85475 , n85476 , n85477 , n85478 , n85479 , n85480 , 
     n85481 , n85482 , n85483 , n85484 , n85485 , n85486 , n85487 , n85488 , n85489 , n85490 , 
     n85491 , n85492 , n85493 , n85494 , n85495 , n85496 , n85497 , n85498 , n85499 , n85500 , 
     n85501 , n85502 , n85503 , n85504 , n85505 , n85506 , n85507 , n85508 , n85509 , n85510 , 
     n85511 , n85512 , n85513 , n85514 , n85515 , n85516 , n85517 , n85518 , n85519 , n85520 , 
     n85521 , n85522 , n85523 , n85524 , n85525 , n85526 , n85527 , n85528 , n85529 , n85530 , 
     n85531 , n85532 , n85533 , n85534 , n85535 , n85536 , n85537 , n85538 , n85539 , n85540 , 
     n85541 , n85542 , n85543 , n85544 , n85545 , n85546 , n85547 , n85548 , n85549 , n85550 , 
     n85551 , n85552 , n85553 , n85554 , n85555 , n85556 , n85557 , n85558 , n85559 , n85560 , 
     n85561 , n85562 , n85563 , n85564 , n85565 , n85566 , n85567 , n85568 , n85569 , n85570 , 
     n85571 , n85572 , n85573 , n85574 , n85575 , n85576 , n85577 , n85578 , n85579 , n85580 , 
     n85581 , n85582 , n85583 , n85584 , n85585 , n85586 , n85587 , n85588 , n85589 , n85590 , 
     n85591 , n85592 , n85593 , n85594 , n85595 , n85596 , n85597 , n85598 , n85599 , n85600 , 
     n85601 , n85602 , n85603 , n85604 , n85605 , n85606 , n85607 , n85608 , n85609 , n85610 , 
     n85611 , n85612 , n85613 , n85614 , n85615 , n85616 , n85617 , n85618 , n85619 , n85620 , 
     n85621 , n85622 , n85623 , n85624 , n85625 , n85626 , n85627 , n85628 , n85629 , n85630 , 
     n85631 , n85632 , n85633 , n85634 , n85635 , n85636 , n85637 , n85638 , n85639 , n85640 , 
     n85641 , n85642 , n85643 , n85644 , n85645 , n85646 , n85647 , n85648 , n85649 , n85650 , 
     n85651 , n85652 , n85653 , n85654 , n85655 , n85656 , n85657 , n85658 , n85659 , n85660 , 
     n85661 , n85662 , n85663 , n85664 , n85665 , n85666 , n85667 , n85668 , n85669 , n85670 , 
     n85671 , n85672 , n85673 , n85674 , n85675 , n85676 , n85677 , n85678 , n85679 , n85680 , 
     n85681 , n85682 , n85683 , n85684 , n85685 , n85686 , n85687 , n85688 , n85689 , n85690 , 
     n85691 , n85692 , n85693 , n85694 , n85695 , n85696 , n85697 , n85698 , n85699 , n85700 , 
     n85701 , n85702 , n85703 , n85704 , n85705 , n85706 , n85707 , n85708 , n85709 , n85710 , 
     n85711 , n85712 , n85713 , n85714 , n85715 , n85716 , n85717 , n85718 , n85719 , n85720 , 
     n85721 , n85722 , n85723 , n85724 , n85725 , n85726 , n85727 , n85728 , n85729 , n85730 , 
     n85731 , n85732 , n85733 , n85734 , n85735 , n85736 , n85737 , n85738 , n85739 , n85740 , 
     n85741 , n85742 , n85743 , n85744 , n85745 , n85746 , n85747 , n85748 , n85749 , n85750 , 
     n85751 , n85752 , n85753 , n85754 , n85755 , n85756 , n85757 , n85758 , n85759 , n85760 , 
     n85761 , n85762 , n85763 , n85764 , n85765 , n85766 , n85767 , n85768 , n85769 , n85770 , 
     n85771 , n85772 , n85773 , n85774 , n85775 , n85776 , n85777 , n85778 , n85779 , n85780 , 
     n85781 , n85782 , n85783 , n85784 , n85785 , n85786 , n85787 , n85788 , n85789 , n85790 , 
     n85791 , n85792 , n85793 , n85794 , n85795 , n85796 , n85797 , n85798 , n85799 , n85800 , 
     n85801 , n85802 , n85803 , n85804 , n85805 , n85806 , n85807 , n85808 , n85809 , n85810 , 
     n85811 , n85812 , n85813 , n85814 , n85815 , n85816 , n85817 , n85818 , n85819 , n85820 , 
     n85821 , n85822 , n85823 , n85824 , n85825 , n85826 , n85827 , n85828 , n85829 , n85830 , 
     n85831 , n85832 , n85833 , n85834 , n85835 , n85836 , n85837 , n85838 , n85839 , n85840 , 
     n85841 , n85842 , n85843 , n85844 , n85845 , n85846 , n85847 , n85848 , n85849 , n85850 , 
     n85851 , n85852 , n85853 , n85854 , n85855 , n85856 , n85857 , n85858 , n85859 , n85860 , 
     n85861 , n85862 , n85863 , n85864 , n85865 , n85866 , n85867 , n85868 , n85869 , n85870 , 
     n85871 , n85872 , n85873 , n85874 , n85875 , n85876 , n85877 , n85878 , n85879 , n85880 , 
     n85881 , n85882 , n85883 , n85884 , n85885 , n85886 , n85887 , n85888 , n85889 , n85890 , 
     n85891 , n85892 , n85893 , n85894 , n85895 , n85896 , n85897 , n85898 , n85899 , n85900 , 
     n85901 , n85902 , n85903 , n85904 , n85905 , n85906 , n85907 , n85908 , n85909 , n85910 , 
     n85911 , n85912 , n85913 , n85914 , n85915 , n85916 , n85917 , n85918 , n85919 , n85920 , 
     n85921 , n85922 , n85923 , n85924 , n85925 , n85926 , n85927 , n85928 , n85929 , n85930 , 
     n85931 , n85932 , n85933 , n85934 , n85935 , n85936 , n85937 , n85938 , n85939 , n85940 , 
     n85941 , n85942 , n85943 , n85944 , n85945 , n85946 , n85947 , n85948 , n85949 , n85950 , 
     n85951 , n85952 , n85953 , n85954 , n85955 , n85956 , n85957 , n85958 , n85959 , n85960 , 
     n85961 , n85962 , n85963 , n85964 , n85965 , n85966 , n85967 , n85968 , n85969 , n85970 , 
     n85971 , n85972 , n85973 , n85974 , n85975 , n85976 , n85977 , n85978 , n85979 , n85980 , 
     n85981 , n85982 , n85983 , n85984 , n85985 , n85986 , n85987 , n85988 , n85989 , n85990 , 
     n85991 , n85992 , n85993 , n85994 , n85995 , n85996 , n85997 , n85998 , n85999 , n86000 , 
     n86001 , n86002 , n86003 , n86004 , n86005 , n86006 , n86007 , n86008 , n86009 , n86010 , 
     n86011 , n86012 , n86013 , n86014 , n86015 , n86016 , n86017 , n86018 , n86019 , n86020 , 
     n86021 , n86022 , n86023 , n86024 , n86025 , n86026 , n86027 , n86028 , n86029 , n86030 , 
     n86031 , n86032 , n86033 , n86034 , n86035 , n86036 , n86037 , n86038 , n86039 , n86040 , 
     n86041 , n86042 , n86043 , n86044 , n86045 , n86046 , n86047 , n86048 , n86049 , n86050 , 
     n86051 , n86052 , n86053 , n86054 , n86055 , n86056 , n86057 , n86058 , n86059 , n86060 , 
     n86061 , n86062 , n86063 , n86064 , n86065 , n86066 , n86067 , n86068 , n86069 , n86070 , 
     n86071 , n86072 , n86073 , n86074 , n86075 , n86076 , n86077 , n86078 , n86079 , n86080 , 
     n86081 , n86082 , n86083 , n86084 , n86085 , n86086 , n86087 , n86088 , n86089 , n86090 , 
     n86091 , n86092 , n86093 , n86094 , n86095 , n86096 , n86097 , n86098 , n86099 , n86100 , 
     n86101 , n86102 , n86103 , n86104 , n86105 , n86106 , n86107 , n86108 , n86109 , n86110 , 
     n86111 , n86112 , n86113 , n86114 , n86115 , n86116 , n86117 , n86118 , n86119 , n86120 , 
     n86121 , n86122 , n86123 , n86124 , n86125 , n86126 , n86127 , n86128 , n86129 , n86130 , 
     n86131 , n86132 , n86133 , n86134 , n86135 , n86136 , n86137 , n86138 , n86139 , n86140 , 
     n86141 , n86142 , n86143 , n86144 , n86145 , n86146 , n86147 , n86148 , n86149 , n86150 , 
     n86151 , n86152 , n86153 , n86154 , n86155 , n86156 , n86157 , n86158 , n86159 , n86160 , 
     n86161 , n86162 , n86163 , n86164 , n86165 , n86166 , n86167 , n86168 , n86169 , n86170 , 
     n86171 , n86172 , n86173 , n86174 , n86175 , n86176 , n86177 , n86178 , n86179 , n86180 , 
     n86181 , n86182 , n86183 , n86184 , n86185 , n86186 , n86187 , n86188 , n86189 , n86190 , 
     n86191 , n86192 , n86193 , n86194 , n86195 , n86196 , n86197 , n86198 , n86199 , n86200 , 
     n86201 , n86202 , n86203 , n86204 , n86205 , n86206 , n86207 , n86208 , n86209 , n86210 , 
     n86211 , n86212 , n86213 , n86214 , n86215 , n86216 , n86217 , n86218 , n86219 , n86220 , 
     n86221 , n86222 , n86223 , n86224 , n86225 , n86226 , n86227 , n86228 , n86229 , n86230 , 
     n86231 , n86232 , n86233 , n86234 , n86235 , n86236 , n86237 , n86238 , n86239 , n86240 , 
     n86241 , n86242 , n86243 , n86244 , n86245 , n86246 , n86247 , n86248 , n86249 , n86250 , 
     n86251 , n86252 , n86253 , n86254 , n86255 , n86256 , n86257 , n86258 , n86259 , n86260 , 
     n86261 , n86262 , n86263 , n86264 , n86265 , n86266 , n86267 , n86268 , n86269 , n86270 , 
     n86271 , n86272 , n86273 , n86274 , n86275 , n86276 , n86277 , n86278 , n86279 , n86280 , 
     n86281 , n86282 , n86283 , n86284 , n86285 , n86286 , n86287 , n86288 , n86289 , n86290 , 
     n86291 , n86292 , n86293 , n86294 , n86295 , n86296 , n86297 , n86298 , n86299 , n86300 , 
     n86301 , n86302 , n86303 , n86304 , n86305 , n86306 , n86307 , n86308 , n86309 , n86310 , 
     n86311 , n86312 , n86313 , n86314 , n86315 , n86316 , n86317 , n86318 , n86319 , n86320 , 
     n86321 , n86322 , n86323 , n86324 , n86325 , n86326 , n86327 , n86328 , n86329 , n86330 , 
     n86331 , n86332 , n86333 , n86334 , n86335 , n86336 , n86337 , n86338 , n86339 , n86340 , 
     n86341 , n86342 , n86343 , n86344 , n86345 , n86346 , n86347 , n86348 , n86349 , n86350 , 
     n86351 , n86352 , n86353 , n86354 , n86355 , n86356 , n86357 , n86358 , n86359 , n86360 , 
     n86361 , n86362 , n86363 , n86364 , n86365 , n86366 , n86367 , n86368 , n86369 , n86370 , 
     n86371 , n86372 , n86373 , n86374 , n86375 , n86376 , n86377 , n86378 , n86379 , n86380 , 
     n86381 , n86382 , n86383 , n86384 , n86385 , n86386 , n86387 , n86388 , n86389 , n86390 , 
     n86391 , n86392 , n86393 , n86394 , n86395 , n86396 , n86397 , n86398 , n86399 , n86400 , 
     n86401 , n86402 , n86403 , n86404 , n86405 , n86406 , n86407 , n86408 , n86409 , n86410 , 
     n86411 , n86412 , n86413 , n86414 , n86415 , n86416 , n86417 , n86418 , n86419 , n86420 , 
     n86421 , n86422 , n86423 , n86424 , n86425 , n86426 , n86427 , n86428 , n86429 , n86430 , 
     n86431 , n86432 , n86433 , n86434 , n86435 , n86436 , n86437 , n86438 , n86439 , n86440 , 
     n86441 , n86442 , n86443 , n86444 , n86445 , n86446 , n86447 , n86448 , n86449 , n86450 , 
     n86451 , n86452 , n86453 , n86454 , n86455 , n86456 , n86457 , n86458 , n86459 , n86460 , 
     n86461 , n86462 , n86463 , n86464 , n86465 , n86466 , n86467 , n86468 , n86469 , n86470 , 
     n86471 , n86472 , n86473 , n86474 , n86475 , n86476 , n86477 , n86478 , n86479 , n86480 , 
     n86481 , n86482 , n86483 , n86484 , n86485 , n86486 , n86487 , n86488 , n86489 , n86490 , 
     n86491 , n86492 , n86493 , n86494 , n86495 , n86496 , n86497 , n86498 , n86499 , n86500 , 
     n86501 , n86502 , n86503 , n86504 , n86505 , n86506 , n86507 , n86508 , n86509 , n86510 , 
     n86511 , n86512 , n86513 , n86514 , n86515 , n86516 , n86517 , n86518 , n86519 , n86520 , 
     n86521 , n86522 , n86523 , n86524 , n86525 , n86526 , n86527 , n86528 , n86529 , n86530 , 
     n86531 , n86532 , n86533 , n86534 , n86535 , n86536 , n86537 , n86538 , n86539 , n86540 , 
     n86541 , n86542 , n86543 , n86544 , n86545 , n86546 , n86547 , n86548 , n86549 , n86550 , 
     n86551 , n86552 , n86553 , n86554 , n86555 , n86556 , n86557 , n86558 , n86559 , n86560 , 
     n86561 , n86562 , n86563 , n86564 , n86565 , n86566 , n86567 , n86568 , n86569 , n86570 , 
     n86571 , n86572 , n86573 , n86574 , n86575 , n86576 , n86577 , n86578 , n86579 , n86580 , 
     n86581 , n86582 , n86583 , n86584 , n86585 , n86586 , n86587 , n86588 , n86589 , n86590 , 
     n86591 , n86592 , n86593 , n86594 , n86595 , n86596 , n86597 , n86598 , n86599 , n86600 , 
     n86601 , n86602 , n86603 , n86604 , n86605 , n86606 , n86607 , n86608 , n86609 , n86610 , 
     n86611 , n86612 , n86613 , n86614 , n86615 , n86616 , n86617 , n86618 , n86619 , n86620 , 
     n86621 , n86622 , n86623 , n86624 , n86625 , n86626 , n86627 , n86628 , n86629 , n86630 , 
     n86631 , n86632 , n86633 , n86634 , n86635 , n86636 , n86637 , n86638 , n86639 , n86640 , 
     n86641 , n86642 , n86643 , n86644 , n86645 , n86646 , n86647 , n86648 , n86649 , n86650 , 
     n86651 , n86652 , n86653 , n86654 , n86655 , n86656 , n86657 , n86658 , n86659 , n86660 , 
     n86661 , n86662 , n86663 , n86664 , n86665 , n86666 , n86667 , n86668 , n86669 , n86670 , 
     n86671 , n86672 , n86673 , n86674 , n86675 , n86676 , n86677 , n86678 , n86679 , n86680 , 
     n86681 , n86682 , n86683 , n86684 , n86685 , n86686 , n86687 , n86688 , n86689 , n86690 , 
     n86691 , n86692 , n86693 , n86694 , n86695 , n86696 , n86697 , n86698 , n86699 , n86700 , 
     n86701 , n86702 , n86703 , n86704 , n86705 , n86706 , n86707 , n86708 , n86709 , n86710 , 
     n86711 , n86712 , n86713 , n86714 , n86715 , n86716 , n86717 , n86718 , n86719 , n86720 , 
     n86721 , n86722 , n86723 , n86724 , n86725 , n86726 , n86727 , n86728 , n86729 , n86730 , 
     n86731 , n86732 , n86733 , n86734 , n86735 , n86736 , n86737 , n86738 , n86739 , n86740 , 
     n86741 , n86742 , n86743 , n86744 , n86745 , n86746 , n86747 , n86748 , n86749 , n86750 , 
     n86751 , n86752 , n86753 , n86754 , n86755 , n86756 , n86757 , n86758 , n86759 , n86760 , 
     n86761 , n86762 , n86763 , n86764 , n86765 , n86766 , n86767 , n86768 , n86769 , n86770 , 
     n86771 , n86772 , n86773 , n86774 , n86775 , n86776 , n86777 , n86778 , n86779 , n86780 , 
     n86781 , n86782 , n86783 , n86784 , n86785 , n86786 , n86787 , n86788 , n86789 , n86790 , 
     n86791 , n86792 , n86793 , n86794 , n86795 , n86796 , n86797 , n86798 , n86799 , n86800 , 
     n86801 , n86802 , n86803 , n86804 , n86805 , n86806 , n86807 , n86808 , n86809 , n86810 , 
     n86811 , n86812 , n86813 , n86814 , n86815 , n86816 , n86817 , n86818 , n86819 , n86820 , 
     n86821 , n86822 , n86823 , n86824 , n86825 , n86826 , n86827 , n86828 , n86829 , n86830 , 
     n86831 , n86832 , n86833 , n86834 , n86835 , n86836 , n86837 , n86838 , n86839 , n86840 , 
     n86841 , n86842 , n86843 , n86844 , n86845 , n86846 , n86847 , n86848 , n86849 , n86850 , 
     n86851 , n86852 , n86853 , n86854 , n86855 , n86856 , n86857 , n86858 , n86859 , n86860 , 
     n86861 , n86862 , n86863 , n86864 , n86865 , n86866 , n86867 , n86868 , n86869 , n86870 , 
     n86871 , n86872 , n86873 , n86874 , n86875 , n86876 , n86877 , n86878 , n86879 , n86880 , 
     n86881 , n86882 , n86883 , n86884 , n86885 , n86886 , n86887 , n86888 , n86889 , n86890 , 
     n86891 , n86892 , n86893 , n86894 , n86895 , n86896 , n86897 , n86898 , n86899 , n86900 , 
     n86901 , n86902 , n86903 , n86904 , n86905 , n86906 , n86907 , n86908 , n86909 , n86910 , 
     n86911 , n86912 , n86913 , n86914 , n86915 , n86916 , n86917 , n86918 , n86919 , n86920 , 
     n86921 , n86922 , n86923 , n86924 , n86925 , n86926 , n86927 , n86928 , n86929 , n86930 , 
     n86931 , n86932 , n86933 , n86934 , n86935 , n86936 , n86937 , n86938 , n86939 , n86940 , 
     n86941 , n86942 , n86943 , n86944 , n86945 , n86946 , n86947 , n86948 , n86949 , n86950 , 
     n86951 , n86952 , n86953 , n86954 , n86955 , n86956 , n86957 , n86958 , n86959 , n86960 , 
     n86961 , n86962 , n86963 , n86964 , n86965 , n86966 , n86967 , n86968 , n86969 , n86970 , 
     n86971 , n86972 , n86973 , n86974 , n86975 , n86976 , n86977 , n86978 , n86979 , n86980 , 
     n86981 , n86982 , n86983 , n86984 , n86985 , n86986 , n86987 , n86988 , n86989 , n86990 , 
     n86991 , n86992 , n86993 , n86994 , n86995 , n86996 , n86997 , n86998 , n86999 , n87000 , 
     n87001 , n87002 , n87003 , n87004 , n87005 , n87006 , n87007 , n87008 , n87009 , n87010 , 
     n87011 , n87012 , n87013 , n87014 , n87015 , n87016 , n87017 , n87018 , n87019 , n87020 , 
     n87021 , n87022 , n87023 , n87024 , n87025 , n87026 , n87027 , n87028 , n87029 , n87030 , 
     n87031 , n87032 , n87033 , n87034 , n87035 , n87036 , n87037 , n87038 , n87039 , n87040 , 
     n87041 , n87042 , n87043 , n87044 , n87045 , n87046 , n87047 , n87048 , n87049 , n87050 , 
     n87051 , n87052 , n87053 , n87054 , n87055 , n87056 , n87057 , n87058 , n87059 , n87060 , 
     n87061 , n87062 , n87063 , n87064 , n87065 , n87066 , n87067 , n87068 , n87069 , n87070 , 
     n87071 , n87072 , n87073 , n87074 , n87075 , n87076 , n87077 , n87078 , n87079 , n87080 , 
     n87081 , n87082 , n87083 , n87084 , n87085 , n87086 , n87087 , n87088 , n87089 , n87090 , 
     n87091 , n87092 , n87093 , n87094 , n87095 , n87096 , n87097 , n87098 , n87099 , n87100 , 
     n87101 , n87102 , n87103 , n87104 , n87105 , n87106 , n87107 , n87108 , n87109 , n87110 , 
     n87111 , n87112 , n87113 , n87114 , n87115 , n87116 , n87117 , n87118 , n87119 , n87120 , 
     n87121 , n87122 , n87123 , n87124 , n87125 , n87126 , n87127 , n87128 , n87129 , n87130 , 
     n87131 , n87132 , n87133 , n87134 , n87135 , n87136 , n87137 , n87138 , n87139 , n87140 , 
     n87141 , n87142 , n87143 , n87144 , n87145 , n87146 , n87147 , n87148 , n87149 , n87150 , 
     n87151 , n87152 , n87153 , n87154 , n87155 , n87156 , n87157 , n87158 , n87159 , n87160 , 
     n87161 , n87162 , n87163 , n87164 , n87165 , n87166 , n87167 , n87168 , n87169 , n87170 , 
     n87171 , n87172 , n87173 , n87174 , n87175 , n87176 , n87177 , n87178 , n87179 , n87180 , 
     n87181 , n87182 , n87183 , n87184 , n87185 , n87186 , n87187 , n87188 , n87189 , n87190 , 
     n87191 , n87192 , n87193 , n87194 , n87195 , n87196 , n87197 , n87198 , n87199 , n87200 , 
     n87201 , n87202 , n87203 , n87204 , n87205 , n87206 , n87207 , n87208 , n87209 , n87210 , 
     n87211 , n87212 , n87213 , n87214 , n87215 , n87216 , n87217 , n87218 , n87219 , n87220 , 
     n87221 , n87222 , n87223 , n87224 , n87225 , n87226 , n87227 , n87228 , n87229 , n87230 , 
     n87231 , n87232 , n87233 , n87234 , n87235 , n87236 , n87237 , n87238 , n87239 , n87240 , 
     n87241 , n87242 , n87243 , n87244 , n87245 , n87246 , n87247 , n87248 , n87249 , n87250 , 
     n87251 , n87252 , n87253 , n87254 , n87255 , n87256 , n87257 , n87258 , n87259 , n87260 , 
     n87261 , n87262 , n87263 , n87264 , n87265 , n87266 , n87267 , n87268 , n87269 , n87270 , 
     n87271 , n87272 , n87273 , n87274 , n87275 , n87276 , n87277 , n87278 , n87279 , n87280 , 
     n87281 , n87282 , n87283 , n87284 , n87285 , n87286 , n87287 , n87288 , n87289 , n87290 , 
     n87291 , n87292 , n87293 , n87294 , n87295 , n87296 , n87297 , n87298 , n87299 , n87300 , 
     n87301 , n87302 , n87303 , n87304 , n87305 , n87306 , n87307 , n87308 , n87309 , n87310 , 
     n87311 , n87312 , n87313 , n87314 , n87315 , n87316 , n87317 , n87318 , n87319 , n87320 , 
     n87321 , n87322 , n87323 , n87324 , n87325 , n87326 , n87327 , n87328 , n87329 , n87330 , 
     n87331 , n87332 , n87333 , n87334 , n87335 , n87336 , n87337 , n87338 , n87339 , n87340 , 
     n87341 , n87342 , n87343 , n87344 , n87345 , n87346 , n87347 , n87348 , n87349 , n87350 , 
     n87351 , n87352 , n87353 , n87354 , n87355 , n87356 , n87357 , n87358 , n87359 , n87360 , 
     n87361 , n87362 , n87363 , n87364 , n87365 , n87366 , n87367 , n87368 , n87369 , n87370 , 
     n87371 , n87372 , n87373 , n87374 , n87375 , n87376 , n87377 , n87378 , n87379 , n87380 , 
     n87381 , n87382 , n87383 , n87384 , n87385 , n87386 , n87387 , n87388 , n87389 , n87390 , 
     n87391 , n87392 , n87393 , n87394 , n87395 , n87396 , n87397 , n87398 , n87399 , n87400 , 
     n87401 , n87402 , n87403 , n87404 , n87405 , n87406 , n87407 , n87408 , n87409 , n87410 , 
     n87411 , n87412 , n87413 , n87414 , n87415 , n87416 , n87417 , n87418 , n87419 , n87420 , 
     n87421 , n87422 , n87423 , n87424 , n87425 , n87426 , n87427 , n87428 , n87429 , n87430 , 
     n87431 , n87432 , n87433 , n87434 , n87435 , n87436 , n87437 , n87438 , n87439 , n87440 , 
     n87441 , n87442 , n87443 , n87444 , n87445 , n87446 , n87447 , n87448 , n87449 , n87450 , 
     n87451 , n87452 , n87453 , n87454 , n87455 , n87456 , n87457 , n87458 , n87459 , n87460 , 
     n87461 , n87462 , n87463 , n87464 , n87465 , n87466 , n87467 , n87468 , n87469 , n87470 , 
     n87471 , n87472 , n87473 , n87474 , n87475 , n87476 , n87477 , n87478 , n87479 , n87480 , 
     n87481 , n87482 , n87483 , n87484 , n87485 , n87486 , n87487 , n87488 , n87489 , n87490 , 
     n87491 , n87492 , n87493 , n87494 , n87495 , n87496 , n87497 , n87498 , n87499 , n87500 , 
     n87501 , n87502 , n87503 , n87504 , n87505 , n87506 , n87507 , n87508 , n87509 , n87510 , 
     n87511 , n87512 , n87513 , n87514 , n87515 , n87516 , n87517 , n87518 , n87519 , n87520 , 
     n87521 , n87522 , n87523 , n87524 , n87525 , n87526 , n87527 , n87528 , n87529 , n87530 , 
     n87531 , n87532 , n87533 , n87534 , n87535 , n87536 , n87537 , n87538 , n87539 , n87540 , 
     n87541 , n87542 , n87543 , n87544 , n87545 , n87546 , n87547 , n87548 , n87549 , n87550 , 
     n87551 , n87552 , n87553 , n87554 , n87555 , n87556 , n87557 , n87558 , n87559 , n87560 , 
     n87561 , n87562 , n87563 , n87564 , n87565 , n87566 , n87567 , n87568 , n87569 , n87570 , 
     n87571 , n87572 , n87573 , n87574 , n87575 , n87576 , n87577 , n87578 , n87579 , n87580 , 
     n87581 , n87582 , n87583 , n87584 , n87585 , n87586 , n87587 , n87588 , n87589 , n87590 , 
     n87591 , n87592 , n87593 , n87594 , n87595 , n87596 , n87597 , n87598 , n87599 , n87600 , 
     n87601 , n87602 , n87603 , n87604 , n87605 , n87606 , n87607 , n87608 , n87609 , n87610 , 
     n87611 , n87612 , n87613 , n87614 , n87615 , n87616 , n87617 , n87618 , n87619 , n87620 , 
     n87621 , n87622 , n87623 , n87624 , n87625 , n87626 , n87627 , n87628 , n87629 , n87630 , 
     n87631 , n87632 , n87633 , n87634 , n87635 , n87636 , n87637 , n87638 , n87639 , n87640 , 
     n87641 , n87642 , n87643 , n87644 , n87645 , n87646 , n87647 , n87648 , n87649 , n87650 , 
     n87651 , n87652 , n87653 , n87654 , n87655 , n87656 , n87657 , n87658 , n87659 , n87660 , 
     n87661 , n87662 , n87663 , n87664 , n87665 , n87666 , n87667 , n87668 , n87669 , n87670 , 
     n87671 , n87672 , n87673 , n87674 , n87675 , n87676 , n87677 , n87678 , n87679 , n87680 , 
     n87681 , n87682 , n87683 , n87684 , n87685 , n87686 , n87687 , n87688 , n87689 , n87690 , 
     n87691 , n87692 , n87693 , n87694 , n87695 , n87696 , n87697 , n87698 , n87699 , n87700 , 
     n87701 , n87702 , n87703 , n87704 , n87705 , n87706 , n87707 , n87708 , n87709 , n87710 , 
     n87711 , n87712 , n87713 , n87714 , n87715 , n87716 , n87717 , n87718 , n87719 , n87720 , 
     n87721 , n87722 , n87723 , n87724 , n87725 , n87726 , n87727 , n87728 , n87729 , n87730 , 
     n87731 , n87732 , n87733 , n87734 , n87735 , n87736 , n87737 , n87738 , n87739 , n87740 , 
     n87741 , n87742 , n87743 , n87744 , n87745 , n87746 , n87747 , n87748 , n87749 , n87750 , 
     n87751 , n87752 , n87753 , n87754 , n87755 , n87756 , n87757 , n87758 , n87759 , n87760 , 
     n87761 , n87762 , n87763 , n87764 , n87765 , n87766 , n87767 , n87768 , n87769 , n87770 , 
     n87771 , n87772 , n87773 , n87774 , n87775 , n87776 , n87777 , n87778 , n87779 , n87780 , 
     n87781 , n87782 , n87783 , n87784 , n87785 , n87786 , n87787 , n87788 , n87789 , n87790 , 
     n87791 , n87792 , n87793 , n87794 , n87795 , n87796 , n87797 , n87798 , n87799 , n87800 , 
     n87801 , n87802 , n87803 , n87804 , n87805 , n87806 , n87807 , n87808 , n87809 , n87810 , 
     n87811 , n87812 , n87813 , n87814 , n87815 , n87816 , n87817 , n87818 , n87819 , n87820 , 
     n87821 , n87822 , n87823 , n87824 , n87825 , n87826 , n87827 , n87828 , n87829 , n87830 , 
     n87831 , n87832 , n87833 , n87834 , n87835 , n87836 , n87837 , n87838 , n87839 , n87840 , 
     n87841 , n87842 , n87843 , n87844 , n87845 , n87846 , n87847 , n87848 , n87849 , n87850 , 
     n87851 , n87852 , n87853 , n87854 , n87855 , n87856 , n87857 , n87858 , n87859 , n87860 , 
     n87861 , n87862 , n87863 , n87864 , n87865 , n87866 , n87867 , n87868 , n87869 , n87870 , 
     n87871 , n87872 , n87873 , n87874 , n87875 , n87876 , n87877 , n87878 , n87879 , n87880 , 
     n87881 , n87882 , n87883 , n87884 , n87885 , n87886 , n87887 , n87888 , n87889 , n87890 , 
     n87891 , n87892 , n87893 , n87894 , n87895 , n87896 , n87897 , n87898 , n87899 , n87900 , 
     n87901 , n87902 , n87903 , n87904 , n87905 , n87906 , n87907 , n87908 , n87909 , n87910 , 
     n87911 , n87912 , n87913 , n87914 , n87915 , n87916 , n87917 , n87918 , n87919 , n87920 , 
     n87921 , n87922 , n87923 , n87924 , n87925 , n87926 , n87927 , n87928 , n87929 , n87930 , 
     n87931 , n87932 , n87933 , n87934 , n87935 , n87936 , n87937 , n87938 , n87939 , n87940 , 
     n87941 , n87942 , n87943 , n87944 , n87945 , n87946 , n87947 , n87948 , n87949 , n87950 , 
     n87951 , n87952 , n87953 , n87954 , n87955 , n87956 , n87957 , n87958 , n87959 , n87960 , 
     n87961 , n87962 , n87963 , n87964 , n87965 , n87966 , n87967 , n87968 , n87969 , n87970 , 
     n87971 , n87972 , n87973 , n87974 , n87975 , n87976 , n87977 , n87978 , n87979 , n87980 , 
     n87981 , n87982 , n87983 , n87984 , n87985 , n87986 , n87987 , n87988 , n87989 , n87990 , 
     n87991 , n87992 , n87993 , n87994 , n87995 , n87996 , n87997 , n87998 , n87999 , n88000 , 
     n88001 , n88002 , n88003 , n88004 , n88005 , n88006 , n88007 , n88008 , n88009 , n88010 , 
     n88011 , n88012 , n88013 , n88014 , n88015 , n88016 , n88017 , n88018 , n88019 , n88020 , 
     n88021 , n88022 , n88023 , n88024 , n88025 , n88026 , n88027 , n88028 , n88029 , n88030 , 
     n88031 , n88032 , n88033 , n88034 , n88035 , n88036 , n88037 , n88038 , n88039 , n88040 , 
     n88041 , n88042 , n88043 , n88044 , n88045 , n88046 , n88047 , n88048 , n88049 , n88050 , 
     n88051 , n88052 , n88053 , n88054 , n88055 , n88056 , n88057 , n88058 , n88059 , n88060 , 
     n88061 , n88062 , n88063 , n88064 , n88065 , n88066 , n88067 , n88068 , n88069 , n88070 , 
     n88071 , n88072 , n88073 , n88074 , n88075 , n88076 , n88077 , n88078 , n88079 , n88080 , 
     n88081 , n88082 , n88083 , n88084 , n88085 , n88086 , n88087 , n88088 , n88089 , n88090 , 
     n88091 , n88092 , n88093 , n88094 , n88095 , n88096 , n88097 , n88098 , n88099 , n88100 , 
     n88101 , n88102 , n88103 , n88104 , n88105 , n88106 , n88107 , n88108 , n88109 , n88110 , 
     n88111 , n88112 , n88113 , n88114 , n88115 , n88116 , n88117 , n88118 , n88119 , n88120 , 
     n88121 , n88122 , n88123 , n88124 , n88125 , n88126 , n88127 , n88128 , n88129 , n88130 , 
     n88131 , n88132 , n88133 , n88134 , n88135 , n88136 , n88137 , n88138 , n88139 , n88140 , 
     n88141 , n88142 , n88143 , n88144 , n88145 , n88146 , n88147 , n88148 , n88149 , n88150 , 
     n88151 , n88152 , n88153 , n88154 , n88155 , n88156 , n88157 , n88158 , n88159 , n88160 , 
     n88161 , n88162 , n88163 , n88164 , n88165 , n88166 , n88167 , n88168 , n88169 , n88170 , 
     n88171 , n88172 , n88173 , n88174 , n88175 , n88176 , n88177 , n88178 , n88179 , n88180 , 
     n88181 , n88182 , n88183 , n88184 , n88185 , n88186 , n88187 , n88188 , n88189 , n88190 , 
     n88191 , n88192 , n88193 , n88194 , n88195 , n88196 , n88197 , n88198 , n88199 , n88200 , 
     n88201 , n88202 , n88203 , n88204 , n88205 , n88206 , n88207 , n88208 , n88209 , n88210 , 
     n88211 , n88212 , n88213 , n88214 , n88215 , n88216 , n88217 , n88218 , n88219 , n88220 , 
     n88221 , n88222 , n88223 , n88224 , n88225 , n88226 , n88227 , n88228 , n88229 , n88230 , 
     n88231 , n88232 , n88233 , n88234 , n88235 , n88236 , n88237 , n88238 , n88239 , n88240 , 
     n88241 , n88242 , n88243 , n88244 , n88245 , n88246 , n88247 , n88248 , n88249 , n88250 , 
     n88251 , n88252 , n88253 , n88254 , n88255 , n88256 , n88257 , n88258 , n88259 , n88260 , 
     n88261 , n88262 , n88263 , n88264 , n88265 , n88266 , n88267 , n88268 , n88269 , n88270 , 
     n88271 , n88272 , n88273 , n88274 , n88275 , n88276 , n88277 , n88278 , n88279 , n88280 , 
     n88281 , n88282 , n88283 , n88284 , n88285 , n88286 , n88287 , n88288 , n88289 , n88290 , 
     n88291 , n88292 , n88293 , n88294 , n88295 , n88296 , n88297 , n88298 , n88299 , n88300 , 
     n88301 , n88302 , n88303 , n88304 , n88305 , n88306 , n88307 , n88308 , n88309 , n88310 , 
     n88311 , n88312 , n88313 , n88314 , n88315 , n88316 , n88317 , n88318 , n88319 , n88320 , 
     n88321 , n88322 , n88323 , n88324 , n88325 , n88326 , n88327 , n88328 , n88329 , n88330 , 
     n88331 , n88332 , n88333 , n88334 , n88335 , n88336 , n88337 , n88338 , n88339 , n88340 , 
     n88341 , n88342 , n88343 , n88344 , n88345 , n88346 , n88347 , n88348 , n88349 , n88350 , 
     n88351 , n88352 , n88353 , n88354 , n88355 , n88356 , n88357 , n88358 , n88359 , n88360 , 
     n88361 , n88362 , n88363 , n88364 , n88365 , n88366 , n88367 , n88368 , n88369 , n88370 , 
     n88371 , n88372 , n88373 , n88374 , n88375 , n88376 , n88377 , n88378 , n88379 , n88380 , 
     n88381 , n88382 , n88383 , n88384 , n88385 , n88386 , n88387 , n88388 , n88389 , n88390 , 
     n88391 , n88392 , n88393 , n88394 , n88395 , n88396 , n88397 , n88398 , n88399 , n88400 , 
     n88401 , n88402 , n88403 , n88404 , n88405 , n88406 , n88407 , n88408 , n88409 , n88410 , 
     n88411 , n88412 , n88413 , n88414 , n88415 , n88416 , n88417 , n88418 , n88419 , n88420 , 
     n88421 , n88422 , n88423 , n88424 , n88425 , n88426 , n88427 , n88428 , n88429 , n88430 , 
     n88431 , n88432 , n88433 , n88434 , n88435 , n88436 , n88437 , n88438 , n88439 , n88440 , 
     n88441 , n88442 , n88443 , n88444 , n88445 , n88446 , n88447 , n88448 , n88449 , n88450 , 
     n88451 , n88452 , n88453 , n88454 , n88455 , n88456 , n88457 , n88458 , n88459 , n88460 , 
     n88461 , n88462 , n88463 , n88464 , n88465 , n88466 , n88467 , n88468 , n88469 , n88470 , 
     n88471 , n88472 , n88473 , n88474 , n88475 , n88476 , n88477 , n88478 , n88479 , n88480 , 
     n88481 , n88482 , n88483 , n88484 , n88485 , n88486 , n88487 , n88488 , n88489 , n88490 , 
     n88491 , n88492 , n88493 , n88494 , n88495 , n88496 , n88497 , n88498 , n88499 , n88500 , 
     n88501 , n88502 , n88503 , n88504 , n88505 , n88506 , n88507 , n88508 , n88509 , n88510 , 
     n88511 , n88512 , n88513 , n88514 , n88515 , n88516 , n88517 , n88518 , n88519 , n88520 , 
     n88521 , n88522 , n88523 , n88524 , n88525 , n88526 , n88527 , n88528 , n88529 , n88530 , 
     n88531 , n88532 , n88533 , n88534 , n88535 , n88536 , n88537 , n88538 , n88539 , n88540 , 
     n88541 , n88542 , n88543 , n88544 , n88545 , n88546 , n88547 , n88548 , n88549 , n88550 , 
     n88551 , n88552 , n88553 , n88554 , n88555 , n88556 , n88557 , n88558 , n88559 , n88560 , 
     n88561 , n88562 , n88563 , n88564 , n88565 , n88566 , n88567 , n88568 , n88569 , n88570 , 
     n88571 , n88572 , n88573 , n88574 , n88575 , n88576 , n88577 , n88578 , n88579 , n88580 , 
     n88581 , n88582 , n88583 , n88584 , n88585 , n88586 , n88587 , n88588 , n88589 , n88590 , 
     n88591 , n88592 , n88593 , n88594 , n88595 , n88596 , n88597 , n88598 , n88599 , n88600 , 
     n88601 , n88602 , n88603 , n88604 , n88605 , n88606 , n88607 , n88608 , n88609 , n88610 , 
     n88611 , n88612 , n88613 , n88614 , n88615 , n88616 , n88617 , n88618 , n88619 , n88620 , 
     n88621 , n88622 , n88623 , n88624 , n88625 , n88626 , n88627 , n88628 , n88629 , n88630 , 
     n88631 , n88632 , n88633 , n88634 , n88635 , n88636 , n88637 , n88638 , n88639 , n88640 , 
     n88641 , n88642 , n88643 , n88644 , n88645 , n88646 , n88647 , n88648 , n88649 , n88650 , 
     n88651 , n88652 , n88653 , n88654 , n88655 , n88656 , n88657 , n88658 , n88659 , n88660 , 
     n88661 , n88662 , n88663 , n88664 , n88665 , n88666 , n88667 , n88668 , n88669 , n88670 , 
     n88671 , n88672 , n88673 , n88674 , n88675 , n88676 , n88677 , n88678 , n88679 , n88680 , 
     n88681 , n88682 , n88683 , n88684 , n88685 , n88686 , n88687 , n88688 , n88689 , n88690 , 
     n88691 , n88692 , n88693 , n88694 , n88695 , n88696 , n88697 , n88698 , n88699 , n88700 , 
     n88701 , n88702 , n88703 , n88704 , n88705 , n88706 , n88707 , n88708 , n88709 , n88710 , 
     n88711 , n88712 , n88713 , n88714 , n88715 , n88716 , n88717 , n88718 , n88719 , n88720 , 
     n88721 , n88722 , n88723 , n88724 , n88725 , n88726 , n88727 , n88728 , n88729 , n88730 , 
     n88731 , n88732 , n88733 , n88734 , n88735 , n88736 , n88737 , n88738 , n88739 , n88740 , 
     n88741 , n88742 , n88743 , n88744 , n88745 , n88746 , n88747 , n88748 , n88749 , n88750 , 
     n88751 , n88752 , n88753 , n88754 , n88755 , n88756 , n88757 , n88758 , n88759 , n88760 , 
     n88761 , n88762 , n88763 , n88764 , n88765 , n88766 , n88767 , n88768 , n88769 , n88770 , 
     n88771 , n88772 , n88773 , n88774 , n88775 , n88776 , n88777 , n88778 , n88779 , n88780 , 
     n88781 , n88782 , n88783 , n88784 , n88785 , n88786 , n88787 , n88788 , n88789 , n88790 , 
     n88791 , n88792 , n88793 , n88794 , n88795 , n88796 , n88797 , n88798 , n88799 , n88800 , 
     n88801 , n88802 , n88803 , n88804 , n88805 , n88806 , n88807 , n88808 , n88809 , n88810 , 
     n88811 , n88812 , n88813 , n88814 , n88815 , n88816 , n88817 , n88818 , n88819 , n88820 , 
     n88821 , n88822 , n88823 , n88824 , n88825 , n88826 , n88827 , n88828 , n88829 , n88830 , 
     n88831 , n88832 , n88833 , n88834 , n88835 , n88836 , n88837 , n88838 , n88839 , n88840 , 
     n88841 , n88842 , n88843 , n88844 , n88845 , n88846 , n88847 , n88848 , n88849 , n88850 , 
     n88851 , n88852 , n88853 , n88854 , n88855 , n88856 , n88857 , n88858 , n88859 , n88860 , 
     n88861 , n88862 , n88863 , n88864 , n88865 , n88866 , n88867 , n88868 , n88869 , n88870 , 
     n88871 , n88872 , n88873 , n88874 , n88875 , n88876 , n88877 , n88878 , n88879 , n88880 , 
     n88881 , n88882 , n88883 , n88884 , n88885 , n88886 , n88887 , n88888 , n88889 , n88890 , 
     n88891 , n88892 , n88893 , n88894 , n88895 , n88896 , n88897 , n88898 , n88899 , n88900 , 
     n88901 , n88902 , n88903 , n88904 , n88905 , n88906 , n88907 , n88908 , n88909 , n88910 , 
     n88911 , n88912 , n88913 , n88914 , n88915 , n88916 , n88917 , n88918 , n88919 , n88920 , 
     n88921 , n88922 , n88923 , n88924 , n88925 , n88926 , n88927 , n88928 , n88929 , n88930 , 
     n88931 , n88932 , n88933 , n88934 , n88935 , n88936 , n88937 , n88938 , n88939 , n88940 , 
     n88941 , n88942 , n88943 , n88944 , n88945 , n88946 , n88947 , n88948 , n88949 , n88950 , 
     n88951 , n88952 , n88953 , n88954 , n88955 , n88956 , n88957 , n88958 , n88959 , n88960 , 
     n88961 , n88962 , n88963 , n88964 , n88965 , n88966 , n88967 , n88968 , n88969 , n88970 , 
     n88971 , n88972 , n88973 , n88974 , n88975 , n88976 , n88977 , n88978 , n88979 , n88980 , 
     n88981 , n88982 , n88983 , n88984 , n88985 , n88986 , n88987 , n88988 , n88989 , n88990 , 
     n88991 , n88992 , n88993 , n88994 , n88995 , n88996 , n88997 , n88998 , n88999 , n89000 , 
     n89001 , n89002 , n89003 , n89004 , n89005 , n89006 , n89007 , n89008 , n89009 , n89010 , 
     n89011 , n89012 , n89013 , n89014 , n89015 , n89016 , n89017 , n89018 , n89019 , n89020 , 
     n89021 , n89022 , n89023 , n89024 , n89025 , n89026 , n89027 , n89028 , n89029 , n89030 , 
     n89031 , n89032 , n89033 , n89034 , n89035 , n89036 , n89037 , n89038 , n89039 , n89040 , 
     n89041 , n89042 , n89043 , n89044 , n89045 , n89046 , n89047 , n89048 , n89049 , n89050 , 
     n89051 , n89052 , n89053 , n89054 , n89055 , n89056 , n89057 , n89058 , n89059 , n89060 , 
     n89061 , n89062 , n89063 , n89064 , n89065 , n89066 , n89067 , n89068 , n89069 , n89070 , 
     n89071 , n89072 , n89073 , n89074 , n89075 , n89076 , n89077 , n89078 , n89079 , n89080 , 
     n89081 , n89082 , n89083 , n89084 , n89085 , n89086 , n89087 , n89088 , n89089 , n89090 , 
     n89091 , n89092 , n89093 , n89094 , n89095 , n89096 , n89097 , n89098 , n89099 , n89100 , 
     n89101 , n89102 , n89103 , n89104 , n89105 , n89106 , n89107 , n89108 , n89109 , n89110 , 
     n89111 , n89112 , n89113 , n89114 , n89115 , n89116 , n89117 , n89118 , n89119 , n89120 , 
     n89121 , n89122 , n89123 , n89124 , n89125 , n89126 , n89127 , n89128 , n89129 , n89130 , 
     n89131 , n89132 , n89133 , n89134 , n89135 , n89136 , n89137 , n89138 , n89139 , n89140 , 
     n89141 , n89142 , n89143 , n89144 , n89145 , n89146 , n89147 , n89148 , n89149 , n89150 , 
     n89151 , n89152 , n89153 , n89154 , n89155 , n89156 , n89157 , n89158 , n89159 , n89160 , 
     n89161 , n89162 , n89163 , n89164 , n89165 , n89166 , n89167 , n89168 , n89169 , n89170 , 
     n89171 , n89172 , n89173 , n89174 , n89175 , n89176 , n89177 , n89178 , n89179 , n89180 , 
     n89181 , n89182 , n89183 , n89184 , n89185 , n89186 , n89187 , n89188 , n89189 , n89190 , 
     n89191 , n89192 , n89193 , n89194 , n89195 , n89196 , n89197 , n89198 , n89199 , n89200 , 
     n89201 , n89202 , n89203 , n89204 , n89205 , n89206 , n89207 , n89208 , n89209 , n89210 , 
     n89211 , n89212 , n89213 , n89214 , n89215 , n89216 , n89217 , n89218 , n89219 , n89220 , 
     n89221 , n89222 , n89223 , n89224 , n89225 , n89226 , n89227 , n89228 , n89229 , n89230 , 
     n89231 , n89232 , n89233 , n89234 , n89235 , n89236 , n89237 , n89238 , n89239 , n89240 , 
     n89241 , n89242 , n89243 , n89244 , n89245 , n89246 , n89247 , n89248 , n89249 , n89250 , 
     n89251 , n89252 , n89253 , n89254 , n89255 , n89256 , n89257 , n89258 , n89259 , n89260 , 
     n89261 , n89262 , n89263 , n89264 , n89265 , n89266 , n89267 , n89268 , n89269 , n89270 , 
     n89271 , n89272 , n89273 , n89274 , n89275 , n89276 , n89277 , n89278 , n89279 , n89280 , 
     n89281 , n89282 , n89283 , n89284 , n89285 , n89286 , n89287 , n89288 , n89289 , n89290 , 
     n89291 , n89292 , n89293 , n89294 , n89295 , n89296 , n89297 , n89298 , n89299 , n89300 , 
     n89301 , n89302 , n89303 , n89304 , n89305 , n89306 , n89307 , n89308 , n89309 , n89310 , 
     n89311 , n89312 , n89313 , n89314 , n89315 , n89316 , n89317 , n89318 , n89319 , n89320 , 
     n89321 , n89322 , n89323 , n89324 , n89325 , n89326 , n89327 , n89328 , n89329 , n89330 , 
     n89331 , n89332 , n89333 , n89334 , n89335 , n89336 , n89337 , n89338 , n89339 , n89340 , 
     n89341 , n89342 , n89343 , n89344 , n89345 , n89346 , n89347 , n89348 , n89349 , n89350 , 
     n89351 , n89352 , n89353 , n89354 , n89355 , n89356 , n89357 , n89358 , n89359 , n89360 , 
     n89361 , n89362 , n89363 , n89364 , n89365 , n89366 , n89367 , n89368 , n89369 , n89370 , 
     n89371 , n89372 , n89373 , n89374 , n89375 , n89376 , n89377 , n89378 , n89379 , n89380 , 
     n89381 , n89382 , n89383 , n89384 , n89385 , n89386 , n89387 , n89388 , n89389 , n89390 , 
     n89391 , n89392 , n89393 , n89394 , n89395 , n89396 , n89397 , n89398 , n89399 , n89400 , 
     n89401 , n89402 , n89403 , n89404 , n89405 , n89406 , n89407 , n89408 , n89409 , n89410 , 
     n89411 , n89412 , n89413 , n89414 , n89415 , n89416 , n89417 , n89418 , n89419 , n89420 , 
     n89421 , n89422 , n89423 , n89424 , n89425 , n89426 , n89427 , n89428 , n89429 , n89430 , 
     n89431 , n89432 , n89433 , n89434 , n89435 , n89436 , n89437 , n89438 , n89439 , n89440 , 
     n89441 , n89442 , n89443 , n89444 , n89445 , n89446 , n89447 , n89448 , n89449 , n89450 , 
     n89451 , n89452 , n89453 , n89454 , n89455 , n89456 , n89457 , n89458 , n89459 , n89460 , 
     n89461 , n89462 , n89463 , n89464 , n89465 , n89466 , n89467 , n89468 , n89469 , n89470 , 
     n89471 , n89472 , n89473 , n89474 , n89475 , n89476 , n89477 , n89478 , n89479 , n89480 , 
     n89481 , n89482 , n89483 , n89484 , n89485 , n89486 , n89487 , n89488 , n89489 , n89490 , 
     n89491 , n89492 , n89493 , n89494 , n89495 , n89496 , n89497 , n89498 , n89499 , n89500 , 
     n89501 , n89502 , n89503 , n89504 , n89505 , n89506 , n89507 , n89508 , n89509 , n89510 , 
     n89511 , n89512 , n89513 , n89514 , n89515 , n89516 , n89517 , n89518 , n89519 , n89520 , 
     n89521 , n89522 , n89523 , n89524 , n89525 , n89526 , n89527 , n89528 , n89529 , n89530 , 
     n89531 , n89532 , n89533 , n89534 , n89535 , n89536 , n89537 , n89538 , n89539 , n89540 , 
     n89541 , n89542 , n89543 , n89544 , n89545 , n89546 , n89547 , n89548 , n89549 , n89550 , 
     n89551 , n89552 , n89553 , n89554 , n89555 , n89556 , n89557 , n89558 , n89559 , n89560 , 
     n89561 , n89562 , n89563 , n89564 , n89565 , n89566 , n89567 , n89568 , n89569 , n89570 , 
     n89571 , n89572 , n89573 , n89574 , n89575 , n89576 , n89577 , n89578 , n89579 , n89580 , 
     n89581 , n89582 , n89583 , n89584 , n89585 , n89586 , n89587 , n89588 , n89589 , n89590 , 
     n89591 , n89592 , n89593 , n89594 , n89595 , n89596 , n89597 , n89598 , n89599 , n89600 , 
     n89601 , n89602 , n89603 , n89604 , n89605 , n89606 , n89607 , n89608 , n89609 , n89610 , 
     n89611 , n89612 , n89613 , n89614 , n89615 , n89616 , n89617 , n89618 , n89619 , n89620 , 
     n89621 , n89622 , n89623 , n89624 , n89625 , n89626 , n89627 , n89628 , n89629 , n89630 , 
     n89631 , n89632 , n89633 , n89634 , n89635 , n89636 , n89637 , n89638 , n89639 , n89640 , 
     n89641 , n89642 , n89643 , n89644 , n89645 , n89646 , n89647 , n89648 , n89649 , n89650 , 
     n89651 , n89652 , n89653 , n89654 , n89655 , n89656 , n89657 , n89658 , n89659 , n89660 , 
     n89661 , n89662 , n89663 , n89664 , n89665 , n89666 , n89667 , n89668 , n89669 , n89670 , 
     n89671 , n89672 , n89673 , n89674 , n89675 , n89676 , n89677 , n89678 , n89679 , n89680 , 
     n89681 , n89682 , n89683 , n89684 , n89685 , n89686 , n89687 , n89688 , n89689 , n89690 , 
     n89691 , n89692 , n89693 , n89694 , n89695 , n89696 , n89697 , n89698 , n89699 , n89700 , 
     n89701 , n89702 , n89703 , n89704 , n89705 , n89706 , n89707 , n89708 , n89709 , n89710 , 
     n89711 , n89712 , n89713 , n89714 , n89715 , n89716 , n89717 , n89718 , n89719 , n89720 , 
     n89721 , n89722 , n89723 , n89724 , n89725 , n89726 , n89727 , n89728 , n89729 , n89730 , 
     n89731 , n89732 , n89733 , n89734 , n89735 , n89736 , n89737 , n89738 , n89739 , n89740 , 
     n89741 , n89742 , n89743 , n89744 , n89745 , n89746 , n89747 , n89748 , n89749 , n89750 , 
     n89751 , n89752 , n89753 , n89754 , n89755 , n89756 , n89757 , n89758 , n89759 , n89760 , 
     n89761 , n89762 , n89763 , n89764 , n89765 , n89766 , n89767 , n89768 , n89769 , n89770 , 
     n89771 , n89772 , n89773 , n89774 , n89775 , n89776 , n89777 , n89778 , n89779 , n89780 , 
     n89781 , n89782 , n89783 , n89784 , n89785 , n89786 , n89787 , n89788 , n89789 , n89790 , 
     n89791 , n89792 , n89793 , n89794 , n89795 , n89796 , n89797 , n89798 , n89799 , n89800 , 
     n89801 , n89802 , n89803 , n89804 , n89805 , n89806 , n89807 , n89808 , n89809 , n89810 , 
     n89811 , n89812 , n89813 , n89814 , n89815 , n89816 , n89817 , n89818 , n89819 , n89820 , 
     n89821 , n89822 , n89823 , n89824 , n89825 , n89826 , n89827 , n89828 , n89829 , n89830 , 
     n89831 , n89832 , n89833 , n89834 , n89835 , n89836 , n89837 , n89838 , n89839 , n89840 , 
     n89841 , n89842 , n89843 , n89844 , n89845 , n89846 , n89847 , n89848 , n89849 , n89850 , 
     n89851 , n89852 , n89853 , n89854 , n89855 , n89856 , n89857 , n89858 , n89859 , n89860 , 
     n89861 , n89862 , n89863 , n89864 , n89865 , n89866 , n89867 , n89868 , n89869 , n89870 , 
     n89871 , n89872 , n89873 , n89874 , n89875 , n89876 , n89877 , n89878 , n89879 , n89880 , 
     n89881 , n89882 , n89883 , n89884 , n89885 , n89886 , n89887 , n89888 , n89889 , n89890 , 
     n89891 , n89892 , n89893 , n89894 , n89895 , n89896 , n89897 , n89898 , n89899 , n89900 , 
     n89901 , n89902 , n89903 , n89904 , n89905 , n89906 , n89907 , n89908 , n89909 , n89910 , 
     n89911 , n89912 , n89913 , n89914 , n89915 , n89916 , n89917 , n89918 , n89919 , n89920 , 
     n89921 , n89922 , n89923 , n89924 , n89925 , n89926 , n89927 , n89928 , n89929 , n89930 , 
     n89931 , n89932 , n89933 , n89934 , n89935 , n89936 , n89937 , n89938 , n89939 , n89940 , 
     n89941 , n89942 , n89943 , n89944 , n89945 , n89946 , n89947 , n89948 , n89949 , n89950 , 
     n89951 , n89952 , n89953 , n89954 , n89955 , n89956 , n89957 , n89958 , n89959 , n89960 , 
     n89961 , n89962 , n89963 , n89964 , n89965 , n89966 , n89967 , n89968 , n89969 , n89970 , 
     n89971 , n89972 , n89973 , n89974 , n89975 , n89976 , n89977 , n89978 , n89979 , n89980 , 
     n89981 , n89982 , n89983 , n89984 , n89985 , n89986 , n89987 , n89988 , n89989 , n89990 , 
     n89991 , n89992 , n89993 , n89994 , n89995 , n89996 , n89997 , n89998 , n89999 , n90000 , 
     n90001 , n90002 , n90003 , n90004 , n90005 , n90006 , n90007 , n90008 , n90009 , n90010 , 
     n90011 , n90012 , n90013 , n90014 , n90015 , n90016 , n90017 , n90018 , n90019 , n90020 , 
     n90021 , n90022 , n90023 , n90024 , n90025 , n90026 , n90027 , n90028 , n90029 , n90030 , 
     n90031 , n90032 , n90033 , n90034 , n90035 , n90036 , n90037 , n90038 , n90039 , n90040 , 
     n90041 , n90042 , n90043 , n90044 , n90045 , n90046 , n90047 , n90048 , n90049 , n90050 , 
     n90051 , n90052 , n90053 , n90054 , n90055 , n90056 , n90057 , n90058 , n90059 , n90060 , 
     n90061 , n90062 , n90063 , n90064 , n90065 , n90066 , n90067 , n90068 , n90069 , n90070 , 
     n90071 , n90072 , n90073 , n90074 , n90075 , n90076 , n90077 , n90078 , n90079 , n90080 , 
     n90081 , n90082 , n90083 , n90084 , n90085 , n90086 , n90087 , n90088 , n90089 , n90090 , 
     n90091 , n90092 , n90093 , n90094 , n90095 , n90096 , n90097 , n90098 , n90099 , n90100 , 
     n90101 , n90102 , n90103 , n90104 , n90105 , n90106 , n90107 , n90108 , n90109 , n90110 , 
     n90111 , n90112 , n90113 , n90114 , n90115 , n90116 , n90117 , n90118 , n90119 , n90120 , 
     n90121 , n90122 , n90123 , n90124 , n90125 , n90126 , n90127 , n90128 , n90129 , n90130 , 
     n90131 , n90132 , n90133 , n90134 , n90135 , n90136 , n90137 , n90138 , n90139 , n90140 , 
     n90141 , n90142 , n90143 , n90144 , n90145 , n90146 , n90147 , n90148 , n90149 , n90150 , 
     n90151 , n90152 , n90153 , n90154 , n90155 , n90156 , n90157 , n90158 , n90159 , n90160 , 
     n90161 , n90162 , n90163 , n90164 , n90165 , n90166 , n90167 , n90168 , n90169 , n90170 , 
     n90171 , n90172 , n90173 , n90174 , n90175 , n90176 , n90177 , n90178 , n90179 , n90180 , 
     n90181 , n90182 , n90183 , n90184 , n90185 , n90186 , n90187 , n90188 , n90189 , n90190 , 
     n90191 , n90192 , n90193 , n90194 , n90195 , n90196 , n90197 , n90198 , n90199 , n90200 , 
     n90201 , n90202 , n90203 , n90204 , n90205 , n90206 , n90207 , n90208 , n90209 , n90210 , 
     n90211 , n90212 , n90213 , n90214 , n90215 , n90216 , n90217 , n90218 , n90219 , n90220 , 
     n90221 , n90222 , n90223 , n90224 , n90225 , n90226 , n90227 , n90228 , n90229 , n90230 , 
     n90231 , n90232 , n90233 , n90234 , n90235 , n90236 , n90237 , n90238 , n90239 , n90240 , 
     n90241 , n90242 , n90243 , n90244 , n90245 , n90246 , n90247 , n90248 , n90249 , n90250 , 
     n90251 , n90252 , n90253 , n90254 , n90255 , n90256 , n90257 , n90258 , n90259 , n90260 , 
     n90261 , n90262 , n90263 , n90264 , n90265 , n90266 , n90267 , n90268 , n90269 , n90270 , 
     n90271 , n90272 , n90273 , n90274 , n90275 , n90276 , n90277 , n90278 , n90279 , n90280 , 
     n90281 , n90282 , n90283 , n90284 , n90285 , n90286 , n90287 , n90288 , n90289 , n90290 , 
     n90291 , n90292 , n90293 , n90294 , n90295 , n90296 , n90297 , n90298 , n90299 , n90300 , 
     n90301 , n90302 , n90303 , n90304 , n90305 , n90306 , n90307 , n90308 , n90309 , n90310 , 
     n90311 , n90312 , n90313 , n90314 , n90315 , n90316 , n90317 , n90318 , n90319 , n90320 , 
     n90321 , n90322 , n90323 , n90324 , n90325 , n90326 , n90327 , n90328 , n90329 , n90330 , 
     n90331 , n90332 , n90333 , n90334 , n90335 , n90336 , n90337 , n90338 , n90339 , n90340 , 
     n90341 , n90342 , n90343 , n90344 , n90345 , n90346 , n90347 , n90348 , n90349 , n90350 , 
     n90351 , n90352 , n90353 , n90354 , n90355 , n90356 , n90357 , n90358 , n90359 , n90360 , 
     n90361 , n90362 , n90363 , n90364 , n90365 , n90366 , n90367 , n90368 , n90369 , n90370 , 
     n90371 , n90372 , n90373 , n90374 , n90375 , n90376 , n90377 , n90378 , n90379 , n90380 , 
     n90381 , n90382 , n90383 , n90384 , n90385 , n90386 , n90387 , n90388 , n90389 , n90390 , 
     n90391 , n90392 , n90393 , n90394 , n90395 , n90396 , n90397 , n90398 , n90399 , n90400 , 
     n90401 , n90402 , n90403 , n90404 , n90405 , n90406 , n90407 , n90408 , n90409 , n90410 , 
     n90411 , n90412 , n90413 , n90414 , n90415 , n90416 , n90417 , n90418 , n90419 , n90420 , 
     n90421 , n90422 , n90423 , n90424 , n90425 , n90426 , n90427 , n90428 , n90429 , n90430 , 
     n90431 , n90432 , n90433 , n90434 , n90435 , n90436 , n90437 , n90438 , n90439 , n90440 , 
     n90441 , n90442 , n90443 , n90444 , n90445 , n90446 , n90447 , n90448 , n90449 , n90450 , 
     n90451 , n90452 , n90453 , n90454 , n90455 , n90456 , n90457 , n90458 , n90459 , n90460 , 
     n90461 , n90462 , n90463 , n90464 , n90465 , n90466 , n90467 , n90468 , n90469 , n90470 , 
     n90471 , n90472 , n90473 , n90474 , n90475 , n90476 , n90477 , n90478 , n90479 , n90480 , 
     n90481 , n90482 , n90483 , n90484 , n90485 , n90486 , n90487 , n90488 , n90489 , n90490 , 
     n90491 , n90492 , n90493 , n90494 , n90495 , n90496 , n90497 , n90498 , n90499 , n90500 , 
     n90501 , n90502 , n90503 , n90504 , n90505 , n90506 , n90507 , n90508 , n90509 , n90510 , 
     n90511 , n90512 , n90513 , n90514 , n90515 , n90516 , n90517 , n90518 , n90519 , n90520 , 
     n90521 , n90522 , n90523 , n90524 , n90525 , n90526 , n90527 , n90528 , n90529 , n90530 , 
     n90531 , n90532 , n90533 , n90534 , n90535 , n90536 , n90537 , n90538 , n90539 , n90540 , 
     n90541 , n90542 , n90543 , n90544 , n90545 , n90546 , n90547 , n90548 , n90549 , n90550 , 
     n90551 , n90552 , n90553 , n90554 , n90555 , n90556 , n90557 , n90558 , n90559 , n90560 , 
     n90561 , n90562 , n90563 , n90564 , n90565 , n90566 , n90567 , n90568 , n90569 , n90570 , 
     n90571 , n90572 , n90573 , n90574 , n90575 , n90576 , n90577 , n90578 , n90579 , n90580 , 
     n90581 , n90582 , n90583 , n90584 , n90585 , n90586 , n90587 , n90588 , n90589 , n90590 , 
     n90591 , n90592 , n90593 , n90594 , n90595 , n90596 , n90597 , n90598 , n90599 , n90600 , 
     n90601 , n90602 , n90603 , n90604 , n90605 , n90606 , n90607 , n90608 , n90609 , n90610 , 
     n90611 , n90612 , n90613 , n90614 , n90615 , n90616 , n90617 , n90618 , n90619 , n90620 , 
     n90621 , n90622 , n90623 , n90624 , n90625 , n90626 , n90627 , n90628 , n90629 , n90630 , 
     n90631 , n90632 , n90633 , n90634 , n90635 , n90636 , n90637 , n90638 , n90639 , n90640 , 
     n90641 , n90642 , n90643 , n90644 , n90645 , n90646 , n90647 , n90648 , n90649 , n90650 , 
     n90651 , n90652 , n90653 , n90654 , n90655 , n90656 , n90657 , n90658 , n90659 , n90660 , 
     n90661 , n90662 , n90663 , n90664 , n90665 , n90666 , n90667 , n90668 , n90669 , n90670 , 
     n90671 , n90672 , n90673 , n90674 , n90675 , n90676 , n90677 , n90678 , n90679 , n90680 , 
     n90681 , n90682 , n90683 , n90684 , n90685 , n90686 , n90687 , n90688 , n90689 , n90690 , 
     n90691 , n90692 , n90693 , n90694 , n90695 , n90696 , n90697 , n90698 , n90699 , n90700 , 
     n90701 , n90702 , n90703 , n90704 , n90705 , n90706 , n90707 , n90708 , n90709 , n90710 , 
     n90711 , n90712 , n90713 , n90714 , n90715 , n90716 , n90717 , n90718 , n90719 , n90720 , 
     n90721 , n90722 , n90723 , n90724 , n90725 , n90726 , n90727 , n90728 , n90729 , n90730 , 
     n90731 , n90732 , n90733 , n90734 , n90735 , n90736 , n90737 , n90738 , n90739 , n90740 , 
     n90741 , n90742 , n90743 , n90744 , n90745 , n90746 , n90747 , n90748 , n90749 , n90750 , 
     n90751 , n90752 , n90753 , n90754 , n90755 , n90756 , n90757 , n90758 , n90759 , n90760 , 
     n90761 , n90762 , n90763 , n90764 , n90765 , n90766 , n90767 , n90768 , n90769 , n90770 , 
     n90771 , n90772 , n90773 , n90774 , n90775 , n90776 , n90777 , n90778 , n90779 , n90780 , 
     n90781 , n90782 , n90783 , n90784 , n90785 , n90786 , n90787 , n90788 , n90789 , n90790 , 
     n90791 , n90792 , n90793 , n90794 , n90795 , n90796 , n90797 , n90798 , n90799 , n90800 , 
     n90801 , n90802 , n90803 , n90804 , n90805 , n90806 , n90807 , n90808 , n90809 , n90810 , 
     n90811 , n90812 , n90813 , n90814 , n90815 , n90816 , n90817 , n90818 , n90819 , n90820 , 
     n90821 , n90822 , n90823 , n90824 , n90825 , n90826 , n90827 , n90828 , n90829 , n90830 , 
     n90831 , n90832 , n90833 , n90834 , n90835 , n90836 , n90837 , n90838 , n90839 , n90840 , 
     n90841 , n90842 , n90843 , n90844 , n90845 , n90846 , n90847 , n90848 , n90849 , n90850 , 
     n90851 , n90852 , n90853 , n90854 , n90855 , n90856 , n90857 , n90858 , n90859 , n90860 , 
     n90861 , n90862 , n90863 , n90864 , n90865 , n90866 , n90867 , n90868 , n90869 , n90870 , 
     n90871 , n90872 , n90873 , n90874 , n90875 , n90876 , n90877 , n90878 , n90879 , n90880 , 
     n90881 , n90882 , n90883 , n90884 , n90885 , n90886 , n90887 , n90888 , n90889 , n90890 , 
     n90891 , n90892 , n90893 , n90894 , n90895 , n90896 , n90897 , n90898 , n90899 , n90900 , 
     n90901 , n90902 , n90903 , n90904 , n90905 , n90906 , n90907 , n90908 , n90909 , n90910 , 
     n90911 , n90912 , n90913 , n90914 , n90915 , n90916 , n90917 , n90918 , n90919 , n90920 , 
     n90921 , n90922 , n90923 , n90924 , n90925 , n90926 , n90927 , n90928 , n90929 , n90930 , 
     n90931 , n90932 , n90933 , n90934 , n90935 , n90936 , n90937 , n90938 , n90939 , n90940 , 
     n90941 , n90942 , n90943 , n90944 , n90945 , n90946 , n90947 , n90948 , n90949 , n90950 , 
     n90951 , n90952 , n90953 , n90954 , n90955 , n90956 , n90957 , n90958 , n90959 , n90960 , 
     n90961 , n90962 , n90963 , n90964 , n90965 , n90966 , n90967 , n90968 , n90969 , n90970 , 
     n90971 , n90972 , n90973 , n90974 , n90975 , n90976 , n90977 , n90978 , n90979 , n90980 , 
     n90981 , n90982 , n90983 , n90984 , n90985 , n90986 , n90987 , n90988 , n90989 , n90990 , 
     n90991 , n90992 , n90993 , n90994 , n90995 , n90996 , n90997 , n90998 , n90999 , n91000 , 
     n91001 , n91002 , n91003 , n91004 , n91005 , n91006 , n91007 , n91008 , n91009 , n91010 , 
     n91011 , n91012 , n91013 , n91014 , n91015 , n91016 , n91017 , n91018 , n91019 , n91020 , 
     n91021 , n91022 , n91023 , n91024 , n91025 , n91026 , n91027 , n91028 , n91029 , n91030 , 
     n91031 , n91032 , n91033 , n91034 , n91035 , n91036 , n91037 , n91038 , n91039 , n91040 , 
     n91041 , n91042 , n91043 , n91044 , n91045 , n91046 , n91047 , n91048 , n91049 , n91050 , 
     n91051 , n91052 , n91053 , n91054 , n91055 , n91056 , n91057 , n91058 , n91059 , n91060 , 
     n91061 , n91062 , n91063 , n91064 , n91065 , n91066 , n91067 , n91068 , n91069 , n91070 , 
     n91071 , n91072 , n91073 , n91074 , n91075 , n91076 , n91077 , n91078 , n91079 , n91080 , 
     n91081 , n91082 , n91083 , n91084 , n91085 , n91086 , n91087 , n91088 , n91089 , n91090 , 
     n91091 , n91092 , n91093 , n91094 , n91095 , n91096 , n91097 , n91098 , n91099 , n91100 , 
     n91101 , n91102 , n91103 , n91104 , n91105 , n91106 , n91107 , n91108 , n91109 , n91110 , 
     n91111 , n91112 , n91113 , n91114 , n91115 , n91116 , n91117 , n91118 , n91119 , n91120 , 
     n91121 , n91122 , n91123 , n91124 , n91125 , n91126 , n91127 , n91128 , n91129 , n91130 , 
     n91131 , n91132 , n91133 , n91134 , n91135 , n91136 , n91137 , n91138 , n91139 , n91140 , 
     n91141 , n91142 , n91143 , n91144 , n91145 , n91146 , n91147 , n91148 , n91149 , n91150 , 
     n91151 , n91152 , n91153 , n91154 , n91155 , n91156 , n91157 , n91158 , n91159 , n91160 , 
     n91161 , n91162 , n91163 , n91164 , n91165 , n91166 , n91167 , n91168 , n91169 , n91170 , 
     n91171 , n91172 , n91173 , n91174 , n91175 , n91176 , n91177 , n91178 , n91179 , n91180 , 
     n91181 , n91182 , n91183 , n91184 , n91185 , n91186 , n91187 , n91188 , n91189 , n91190 , 
     n91191 , n91192 , n91193 , n91194 , n91195 , n91196 , n91197 , n91198 , n91199 , n91200 , 
     n91201 , n91202 , n91203 , n91204 , n91205 , n91206 , n91207 , n91208 , n91209 , n91210 , 
     n91211 , n91212 , n91213 , n91214 , n91215 , n91216 , n91217 , n91218 , n91219 , n91220 , 
     n91221 , n91222 , n91223 , n91224 , n91225 , n91226 , n91227 , n91228 , n91229 , n91230 , 
     n91231 , n91232 , n91233 , n91234 , n91235 , n91236 , n91237 , n91238 , n91239 , n91240 , 
     n91241 , n91242 , n91243 , n91244 , n91245 , n91246 , n91247 , n91248 , n91249 , n91250 , 
     n91251 , n91252 , n91253 , n91254 , n91255 , n91256 , n91257 , n91258 , n91259 , n91260 , 
     n91261 , n91262 , n91263 , n91264 , n91265 , n91266 , n91267 , n91268 , n91269 , n91270 , 
     n91271 , n91272 , n91273 , n91274 , n91275 , n91276 , n91277 , n91278 , n91279 , n91280 , 
     n91281 , n91282 , n91283 , n91284 , n91285 , n91286 , n91287 , n91288 , n91289 , n91290 , 
     n91291 , n91292 , n91293 , n91294 , n91295 , n91296 , n91297 , n91298 , n91299 , n91300 , 
     n91301 , n91302 , n91303 , n91304 , n91305 , n91306 , n91307 , n91308 , n91309 , n91310 , 
     n91311 , n91312 , n91313 , n91314 , n91315 , n91316 , n91317 , n91318 , n91319 , n91320 , 
     n91321 , n91322 , n91323 , n91324 , n91325 , n91326 , n91327 , n91328 , n91329 , n91330 , 
     n91331 , n91332 , n91333 , n91334 , n91335 , n91336 , n91337 , n91338 , n91339 , n91340 , 
     n91341 , n91342 , n91343 , n91344 , n91345 , n91346 , n91347 , n91348 , n91349 , n91350 , 
     n91351 , n91352 , n91353 , n91354 , n91355 , n91356 , n91357 , n91358 , n91359 , n91360 , 
     n91361 , n91362 , n91363 , n91364 , n91365 , n91366 , n91367 , n91368 , n91369 , n91370 , 
     n91371 , n91372 , n91373 , n91374 , n91375 , n91376 , n91377 , n91378 , n91379 , n91380 , 
     n91381 , n91382 , n91383 , n91384 , n91385 , n91386 , n91387 , n91388 , n91389 , n91390 , 
     n91391 , n91392 , n91393 , n91394 , n91395 , n91396 , n91397 , n91398 , n91399 , n91400 , 
     n91401 , n91402 , n91403 , n91404 , n91405 , n91406 , n91407 , n91408 , n91409 , n91410 , 
     n91411 , n91412 , n91413 , n91414 , n91415 , n91416 , n91417 , n91418 , n91419 , n91420 , 
     n91421 , n91422 , n91423 , n91424 , n91425 , n91426 , n91427 , n91428 , n91429 , n91430 , 
     n91431 , n91432 , n91433 , n91434 , n91435 , n91436 , n91437 , n91438 , n91439 , n91440 , 
     n91441 , n91442 , n91443 , n91444 , n91445 , n91446 , n91447 , n91448 , n91449 , n91450 , 
     n91451 , n91452 , n91453 , n91454 , n91455 , n91456 , n91457 , n91458 , n91459 , n91460 , 
     n91461 , n91462 , n91463 , n91464 , n91465 , n91466 , n91467 , n91468 , n91469 , n91470 , 
     n91471 , n91472 , n91473 , n91474 , n91475 , n91476 , n91477 , n91478 , n91479 , n91480 , 
     n91481 , n91482 , n91483 , n91484 , n91485 , n91486 , n91487 , n91488 , n91489 , n91490 , 
     n91491 , n91492 , n91493 , n91494 , n91495 , n91496 , n91497 , n91498 , n91499 , n91500 , 
     n91501 , n91502 , n91503 , n91504 , n91505 , n91506 , n91507 , n91508 , n91509 , n91510 , 
     n91511 , n91512 , n91513 , n91514 , n91515 , n91516 , n91517 , n91518 , n91519 , n91520 , 
     n91521 , n91522 , n91523 , n91524 , n91525 , n91526 , n91527 , n91528 , n91529 , n91530 , 
     n91531 , n91532 , n91533 , n91534 , n91535 , n91536 , n91537 , n91538 , n91539 , n91540 , 
     n91541 , n91542 , n91543 , n91544 , n91545 , n91546 , n91547 , n91548 , n91549 , n91550 , 
     n91551 , n91552 , n91553 , n91554 , n91555 , n91556 , n91557 , n91558 , n91559 , n91560 , 
     n91561 , n91562 , n91563 , n91564 , n91565 , n91566 , n91567 , n91568 , n91569 , n91570 , 
     n91571 , n91572 , n91573 , n91574 , n91575 , n91576 , n91577 , n91578 , n91579 , n91580 , 
     n91581 , n91582 , n91583 , n91584 , n91585 , n91586 , n91587 , n91588 , n91589 , n91590 , 
     n91591 , n91592 , n91593 , n91594 , n91595 , n91596 , n91597 , n91598 , n91599 , n91600 , 
     n91601 , n91602 , n91603 , n91604 , n91605 , n91606 , n91607 , n91608 , n91609 , n91610 , 
     n91611 , n91612 , n91613 , n91614 , n91615 , n91616 , n91617 , n91618 , n91619 , n91620 , 
     n91621 , n91622 , n91623 , n91624 , n91625 , n91626 , n91627 , n91628 , n91629 , n91630 , 
     n91631 , n91632 , n91633 , n91634 , n91635 , n91636 , n91637 , n91638 , n91639 , n91640 , 
     n91641 , n91642 , n91643 , n91644 , n91645 , n91646 , n91647 , n91648 , n91649 , n91650 , 
     n91651 , n91652 , n91653 , n91654 , n91655 , n91656 , n91657 , n91658 , n91659 , n91660 , 
     n91661 , n91662 , n91663 , n91664 , n91665 , n91666 , n91667 , n91668 , n91669 , n91670 , 
     n91671 , n91672 , n91673 , n91674 , n91675 , n91676 , n91677 , n91678 , n91679 , n91680 , 
     n91681 , n91682 , n91683 , n91684 , n91685 , n91686 , n91687 , n91688 , n91689 , n91690 , 
     n91691 , n91692 , n91693 , n91694 , n91695 , n91696 , n91697 , n91698 , n91699 , n91700 , 
     n91701 , n91702 , n91703 , n91704 , n91705 , n91706 , n91707 , n91708 , n91709 , n91710 , 
     n91711 , n91712 , n91713 , n91714 , n91715 , n91716 , n91717 , n91718 , n91719 , n91720 , 
     n91721 , n91722 , n91723 , n91724 , n91725 , n91726 , n91727 , n91728 , n91729 , n91730 , 
     n91731 , n91732 , n91733 , n91734 , n91735 , n91736 , n91737 , n91738 , n91739 , n91740 , 
     n91741 , n91742 , n91743 , n91744 , n91745 , n91746 , n91747 , n91748 , n91749 , n91750 , 
     n91751 , n91752 , n91753 , n91754 , n91755 , n91756 , n91757 , n91758 , n91759 , n91760 , 
     n91761 , n91762 , n91763 , n91764 , n91765 , n91766 , n91767 , n91768 , n91769 , n91770 , 
     n91771 , n91772 , n91773 , n91774 , n91775 , n91776 , n91777 , n91778 , n91779 , n91780 , 
     n91781 , n91782 , n91783 , n91784 , n91785 , n91786 , n91787 , n91788 , n91789 , n91790 , 
     n91791 , n91792 , n91793 , n91794 , n91795 , n91796 , n91797 , n91798 , n91799 , n91800 , 
     n91801 , n91802 , n91803 , n91804 , n91805 , n91806 , n91807 , n91808 , n91809 , n91810 , 
     n91811 , n91812 , n91813 , n91814 , n91815 , n91816 , n91817 , n91818 , n91819 , n91820 , 
     n91821 , n91822 , n91823 , n91824 , n91825 , n91826 , n91827 , n91828 , n91829 , n91830 , 
     n91831 , n91832 , n91833 , n91834 , n91835 , n91836 , n91837 , n91838 , n91839 , n91840 , 
     n91841 , n91842 , n91843 , n91844 , n91845 , n91846 , n91847 , n91848 , n91849 , n91850 , 
     n91851 , n91852 , n91853 , n91854 , n91855 , n91856 , n91857 , n91858 , n91859 , n91860 , 
     n91861 , n91862 , n91863 , n91864 , n91865 , n91866 , n91867 , n91868 , n91869 , n91870 , 
     n91871 , n91872 , n91873 , n91874 , n91875 , n91876 , n91877 , n91878 , n91879 , n91880 , 
     n91881 , n91882 , n91883 , n91884 , n91885 , n91886 , n91887 , n91888 , n91889 , n91890 , 
     n91891 , n91892 , n91893 , n91894 , n91895 , n91896 , n91897 , n91898 , n91899 , n91900 , 
     n91901 , n91902 , n91903 , n91904 , n91905 , n91906 , n91907 , n91908 , n91909 , n91910 , 
     n91911 , n91912 , n91913 , n91914 , n91915 , n91916 , n91917 , n91918 , n91919 , n91920 , 
     n91921 , n91922 , n91923 , n91924 , n91925 , n91926 , n91927 , n91928 , n91929 , n91930 , 
     n91931 , n91932 , n91933 , n91934 , n91935 , n91936 , n91937 , n91938 , n91939 , n91940 , 
     n91941 , n91942 , n91943 , n91944 , n91945 , n91946 , n91947 , n91948 , n91949 , n91950 , 
     n91951 , n91952 , n91953 , n91954 , n91955 , n91956 , n91957 , n91958 , n91959 , n91960 , 
     n91961 , n91962 , n91963 , n91964 , n91965 , n91966 , n91967 , n91968 , n91969 , n91970 , 
     n91971 , n91972 , n91973 , n91974 , n91975 , n91976 , n91977 , n91978 , n91979 , n91980 , 
     n91981 , n91982 , n91983 , n91984 , n91985 , n91986 , n91987 , n91988 , n91989 , n91990 , 
     n91991 , n91992 , n91993 , n91994 , n91995 , n91996 , n91997 , n91998 , n91999 , n92000 , 
     n92001 , n92002 , n92003 , n92004 , n92005 , n92006 , n92007 , n92008 , n92009 , n92010 , 
     n92011 , n92012 , n92013 , n92014 , n92015 , n92016 , n92017 , n92018 , n92019 , n92020 , 
     n92021 , n92022 , n92023 , n92024 , n92025 , n92026 , n92027 , n92028 , n92029 , n92030 , 
     n92031 , n92032 , n92033 , n92034 , n92035 , n92036 , n92037 , n92038 , n92039 , n92040 , 
     n92041 , n92042 , n92043 , n92044 , n92045 , n92046 , n92047 , n92048 , n92049 , n92050 , 
     n92051 , n92052 , n92053 , n92054 , n92055 , n92056 , n92057 , n92058 , n92059 , n92060 , 
     n92061 , n92062 , n92063 , n92064 , n92065 , n92066 , n92067 , n92068 , n92069 , n92070 , 
     n92071 , n92072 , n92073 , n92074 , n92075 , n92076 , n92077 , n92078 , n92079 , n92080 , 
     n92081 , n92082 , n92083 , n92084 , n92085 , n92086 , n92087 , n92088 , n92089 , n92090 , 
     n92091 , n92092 , n92093 , n92094 , n92095 , n92096 , n92097 , n92098 , n92099 , n92100 , 
     n92101 , n92102 , n92103 , n92104 , n92105 , n92106 , n92107 , n92108 , n92109 , n92110 , 
     n92111 , n92112 , n92113 , n92114 , n92115 , n92116 , n92117 , n92118 , n92119 , n92120 , 
     n92121 , n92122 , n92123 , n92124 , n92125 , n92126 , n92127 , n92128 , n92129 , n92130 , 
     n92131 , n92132 , n92133 , n92134 , n92135 , n92136 , n92137 , n92138 , n92139 , n92140 , 
     n92141 , n92142 , n92143 , n92144 , n92145 , n92146 , n92147 , n92148 , n92149 , n92150 , 
     n92151 , n92152 , n92153 , n92154 , n92155 , n92156 , n92157 , n92158 , n92159 , n92160 , 
     n92161 , n92162 , n92163 , n92164 , n92165 , n92166 , n92167 , n92168 , n92169 , n92170 , 
     n92171 , n92172 , n92173 , n92174 , n92175 , n92176 , n92177 , n92178 , n92179 , n92180 , 
     n92181 , n92182 , n92183 , n92184 , n92185 , n92186 , n92187 , n92188 , n92189 , n92190 , 
     n92191 , n92192 , n92193 , n92194 , n92195 , n92196 , n92197 , n92198 , n92199 , n92200 , 
     n92201 , n92202 , n92203 , n92204 , n92205 , n92206 , n92207 , n92208 , n92209 , n92210 , 
     n92211 , n92212 , n92213 , n92214 , n92215 , n92216 , n92217 , n92218 , n92219 , n92220 , 
     n92221 , n92222 , n92223 , n92224 , n92225 , n92226 , n92227 , n92228 , n92229 , n92230 , 
     n92231 , n92232 , n92233 , n92234 , n92235 , n92236 , n92237 , n92238 , n92239 , n92240 , 
     n92241 , n92242 , n92243 , n92244 , n92245 , n92246 , n92247 , n92248 , n92249 , n92250 , 
     n92251 , n92252 , n92253 , n92254 , n92255 , n92256 , n92257 , n92258 , n92259 , n92260 , 
     n92261 , n92262 , n92263 , n92264 , n92265 , n92266 , n92267 , n92268 , n92269 , n92270 , 
     n92271 , n92272 , n92273 , n92274 , n92275 , n92276 , n92277 , n92278 , n92279 , n92280 , 
     n92281 , n92282 , n92283 , n92284 , n92285 , n92286 , n92287 , n92288 , n92289 , n92290 , 
     n92291 , n92292 , n92293 , n92294 , n92295 , n92296 , n92297 , n92298 , n92299 , n92300 , 
     n92301 , n92302 , n92303 , n92304 , n92305 , n92306 , n92307 , n92308 , n92309 , n92310 , 
     n92311 , n92312 , n92313 , n92314 , n92315 , n92316 , n92317 , n92318 , n92319 , n92320 , 
     n92321 , n92322 , n92323 , n92324 , n92325 , n92326 , n92327 , n92328 , n92329 , n92330 , 
     n92331 , n92332 , n92333 , n92334 , n92335 , n92336 , n92337 , n92338 , n92339 , n92340 , 
     n92341 , n92342 , n92343 , n92344 , n92345 , n92346 , n92347 , n92348 , n92349 , n92350 , 
     n92351 , n92352 , n92353 , n92354 , n92355 , n92356 , n92357 , n92358 , n92359 , n92360 , 
     n92361 , n92362 , n92363 , n92364 , n92365 , n92366 , n92367 , n92368 , n92369 , n92370 , 
     n92371 , n92372 , n92373 , n92374 , n92375 , n92376 , n92377 , n92378 , n92379 , n92380 , 
     n92381 , n92382 , n92383 , n92384 , n92385 , n92386 , n92387 , n92388 , n92389 , n92390 , 
     n92391 , n92392 , n92393 , n92394 , n92395 , n92396 , n92397 , n92398 , n92399 , n92400 , 
     n92401 , n92402 , n92403 , n92404 , n92405 , n92406 , n92407 , n92408 , n92409 , n92410 , 
     n92411 , n92412 , n92413 , n92414 , n92415 , n92416 , n92417 , n92418 , n92419 , n92420 , 
     n92421 , n92422 , n92423 , n92424 , n92425 , n92426 , n92427 , n92428 , n92429 , n92430 , 
     n92431 , n92432 , n92433 , n92434 , n92435 , n92436 , n92437 , n92438 , n92439 , n92440 , 
     n92441 , n92442 , n92443 , n92444 , n92445 , n92446 , n92447 , n92448 , n92449 , n92450 , 
     n92451 , n92452 , n92453 , n92454 , n92455 , n92456 , n92457 , n92458 , n92459 , n92460 , 
     n92461 , n92462 , n92463 , n92464 , n92465 , n92466 , n92467 , n92468 , n92469 , n92470 , 
     n92471 , n92472 , n92473 , n92474 , n92475 , n92476 , n92477 , n92478 , n92479 , n92480 , 
     n92481 , n92482 , n92483 , n92484 , n92485 , n92486 , n92487 , n92488 , n92489 , n92490 , 
     n92491 , n92492 , n92493 , n92494 , n92495 , n92496 , n92497 , n92498 , n92499 , n92500 , 
     n92501 , n92502 , n92503 , n92504 , n92505 , n92506 , n92507 , n92508 , n92509 , n92510 , 
     n92511 , n92512 , n92513 , n92514 , n92515 , n92516 , n92517 , n92518 , n92519 , n92520 , 
     n92521 , n92522 , n92523 , n92524 , n92525 , n92526 , n92527 , n92528 , n92529 , n92530 , 
     n92531 , n92532 , n92533 , n92534 , n92535 , n92536 , n92537 , n92538 , n92539 , n92540 , 
     n92541 , n92542 , n92543 , n92544 , n92545 , n92546 , n92547 , n92548 , n92549 , n92550 , 
     n92551 , n92552 , n92553 , n92554 , n92555 , n92556 , n92557 , n92558 , n92559 , n92560 , 
     n92561 , n92562 , n92563 , n92564 , n92565 , n92566 , n92567 , n92568 , n92569 , n92570 , 
     n92571 , n92572 , n92573 , n92574 , n92575 , n92576 , n92577 , n92578 , n92579 , n92580 , 
     n92581 , n92582 , n92583 , n92584 , n92585 , n92586 , n92587 , n92588 , n92589 , n92590 , 
     n92591 , n92592 , n92593 , n92594 , n92595 , n92596 , n92597 , n92598 , n92599 , n92600 , 
     n92601 , n92602 , n92603 , n92604 , n92605 , n92606 , n92607 , n92608 , n92609 , n92610 , 
     n92611 , n92612 , n92613 , n92614 , n92615 , n92616 , n92617 , n92618 , n92619 , n92620 , 
     n92621 , n92622 , n92623 , n92624 , n92625 , n92626 , n92627 , n92628 , n92629 , n92630 , 
     n92631 , n92632 , n92633 , n92634 , n92635 , n92636 , n92637 , n92638 , n92639 , n92640 , 
     n92641 , n92642 , n92643 , n92644 , n92645 , n92646 , n92647 , n92648 , n92649 , n92650 , 
     n92651 , n92652 , n92653 , n92654 , n92655 , n92656 , n92657 , n92658 , n92659 , n92660 , 
     n92661 , n92662 , n92663 , n92664 , n92665 , n92666 , n92667 , n92668 , n92669 , n92670 , 
     n92671 , n92672 , n92673 , n92674 , n92675 , n92676 , n92677 , n92678 , n92679 , n92680 , 
     n92681 , n92682 , n92683 , n92684 , n92685 , n92686 , n92687 , n92688 , n92689 , n92690 , 
     n92691 , n92692 , n92693 , n92694 , n92695 , n92696 , n92697 , n92698 , n92699 , n92700 , 
     n92701 , n92702 , n92703 , n92704 , n92705 , n92706 , n92707 , n92708 , n92709 , n92710 , 
     n92711 , n92712 , n92713 , n92714 , n92715 , n92716 , n92717 , n92718 , n92719 , n92720 , 
     n92721 , n92722 , n92723 , n92724 , n92725 , n92726 , n92727 , n92728 , n92729 , n92730 , 
     n92731 , n92732 , n92733 , n92734 , n92735 , n92736 , n92737 , n92738 , n92739 , n92740 , 
     n92741 , n92742 , n92743 , n92744 , n92745 , n92746 , n92747 , n92748 , n92749 , n92750 , 
     n92751 , n92752 , n92753 , n92754 , n92755 , n92756 , n92757 , n92758 , n92759 , n92760 , 
     n92761 , n92762 , n92763 , n92764 , n92765 , n92766 , n92767 , n92768 , n92769 , n92770 , 
     n92771 , n92772 , n92773 , n92774 , n92775 , n92776 , n92777 , n92778 , n92779 , n92780 , 
     n92781 , n92782 , n92783 , n92784 , n92785 , n92786 , n92787 , n92788 , n92789 , n92790 , 
     n92791 , n92792 , n92793 , n92794 , n92795 , n92796 , n92797 , n92798 , n92799 , n92800 , 
     n92801 , n92802 , n92803 , n92804 , n92805 , n92806 , n92807 , n92808 , n92809 , n92810 , 
     n92811 , n92812 , n92813 , n92814 , n92815 , n92816 , n92817 , n92818 , n92819 , n92820 , 
     n92821 , n92822 , n92823 , n92824 , n92825 , n92826 , n92827 , n92828 , n92829 , n92830 , 
     n92831 , n92832 , n92833 , n92834 , n92835 , n92836 , n92837 , n92838 , n92839 , n92840 , 
     n92841 , n92842 , n92843 , n92844 , n92845 , n92846 , n92847 , n92848 , n92849 , n92850 , 
     n92851 , n92852 , n92853 , n92854 , n92855 , n92856 , n92857 , n92858 , n92859 , n92860 , 
     n92861 , n92862 , n92863 , n92864 , n92865 , n92866 , n92867 , n92868 , n92869 , n92870 , 
     n92871 , n92872 , n92873 , n92874 , n92875 , n92876 , n92877 , n92878 , n92879 , n92880 , 
     n92881 , n92882 , n92883 , n92884 , n92885 , n92886 , n92887 , n92888 , n92889 , n92890 , 
     n92891 , n92892 , n92893 , n92894 , n92895 , n92896 , n92897 , n92898 , n92899 , n92900 , 
     n92901 , n92902 , n92903 , n92904 , n92905 , n92906 , n92907 , n92908 , n92909 , n92910 , 
     n92911 , n92912 , n92913 , n92914 , n92915 , n92916 , n92917 , n92918 , n92919 , n92920 , 
     n92921 , n92922 , n92923 , n92924 , n92925 , n92926 , n92927 , n92928 , n92929 , n92930 , 
     n92931 , n92932 , n92933 , n92934 , n92935 , n92936 , n92937 , n92938 , n92939 , n92940 , 
     n92941 , n92942 , n92943 , n92944 , n92945 , n92946 , n92947 , n92948 , n92949 , n92950 , 
     n92951 , n92952 , n92953 , n92954 , n92955 , n92956 , n92957 , n92958 , n92959 , n92960 , 
     n92961 , n92962 , n92963 , n92964 , n92965 , n92966 , n92967 , n92968 , n92969 , n92970 , 
     n92971 , n92972 , n92973 , n92974 , n92975 , n92976 , n92977 , n92978 , n92979 , n92980 , 
     n92981 , n92982 , n92983 , n92984 , n92985 , n92986 , n92987 , n92988 , n92989 , n92990 , 
     n92991 , n92992 , n92993 , n92994 , n92995 , n92996 , n92997 , n92998 , n92999 , n93000 , 
     n93001 , n93002 , n93003 , n93004 , n93005 , n93006 , n93007 , n93008 , n93009 , n93010 , 
     n93011 , n93012 , n93013 , n93014 , n93015 , n93016 , n93017 , n93018 , n93019 , n93020 , 
     n93021 , n93022 , n93023 , n93024 , n93025 , n93026 , n93027 , n93028 , n93029 , n93030 , 
     n93031 , n93032 , n93033 , n93034 , n93035 , n93036 , n93037 , n93038 , n93039 , n93040 , 
     n93041 , n93042 , n93043 , n93044 , n93045 , n93046 , n93047 , n93048 , n93049 , n93050 , 
     n93051 , n93052 , n93053 , n93054 , n93055 , n93056 , n93057 , n93058 , n93059 , n93060 , 
     n93061 , n93062 , n93063 , n93064 , n93065 , n93066 , n93067 , n93068 , n93069 , n93070 , 
     n93071 , n93072 , n93073 , n93074 , n93075 , n93076 , n93077 , n93078 , n93079 , n93080 , 
     n93081 , n93082 , n93083 , n93084 , n93085 , n93086 , n93087 , n93088 , n93089 , n93090 , 
     n93091 , n93092 , n93093 , n93094 , n93095 , n93096 , n93097 , n93098 , n93099 , n93100 , 
     n93101 , n93102 , n93103 , n93104 , n93105 , n93106 , n93107 , n93108 , n93109 , n93110 , 
     n93111 , n93112 , n93113 , n93114 , n93115 , n93116 , n93117 , n93118 , n93119 , n93120 , 
     n93121 , n93122 , n93123 , n93124 , n93125 , n93126 , n93127 , n93128 , n93129 , n93130 , 
     n93131 , n93132 , n93133 , n93134 , n93135 , n93136 , n93137 , n93138 , n93139 , n93140 , 
     n93141 , n93142 , n93143 , n93144 , n93145 , n93146 , n93147 , n93148 , n93149 , n93150 , 
     n93151 , n93152 , n93153 , n93154 , n93155 , n93156 , n93157 , n93158 , n93159 , n93160 , 
     n93161 , n93162 , n93163 , n93164 , n93165 , n93166 , n93167 , n93168 , n93169 , n93170 , 
     n93171 , n93172 , n93173 , n93174 , n93175 , n93176 , n93177 , n93178 , n93179 , n93180 , 
     n93181 , n93182 , n93183 , n93184 , n93185 , n93186 , n93187 , n93188 , n93189 , n93190 , 
     n93191 , n93192 , n93193 , n93194 , n93195 , n93196 , n93197 , n93198 , n93199 , n93200 , 
     n93201 , n93202 , n93203 , n93204 , n93205 , n93206 , n93207 , n93208 , n93209 , n93210 , 
     n93211 , n93212 , n93213 , n93214 , n93215 , n93216 , n93217 , n93218 , n93219 , n93220 , 
     n93221 , n93222 , n93223 , n93224 , n93225 , n93226 , n93227 , n93228 , n93229 , n93230 , 
     n93231 , n93232 , n93233 , n93234 , n93235 , n93236 , n93237 , n93238 , n93239 , n93240 , 
     n93241 , n93242 , n93243 , n93244 , n93245 , n93246 , n93247 , n93248 , n93249 , n93250 , 
     n93251 , n93252 , n93253 , n93254 , n93255 , n93256 , n93257 , n93258 , n93259 , n93260 , 
     n93261 , n93262 , n93263 , n93264 , n93265 , n93266 , n93267 , n93268 , n93269 , n93270 , 
     n93271 , n93272 , n93273 , n93274 , n93275 , n93276 , n93277 , n93278 , n93279 , n93280 , 
     n93281 , n93282 , n93283 , n93284 , n93285 , n93286 , n93287 , n93288 , n93289 , n93290 , 
     n93291 , n93292 , n93293 , n93294 , n93295 , n93296 , n93297 , n93298 , n93299 , n93300 , 
     n93301 , n93302 , n93303 , n93304 , n93305 , n93306 , n93307 , n93308 , n93309 , n93310 , 
     n93311 , n93312 , n93313 , n93314 , n93315 , n93316 , n93317 , n93318 , n93319 , n93320 , 
     n93321 , n93322 , n93323 , n93324 , n93325 , n93326 , n93327 , n93328 , n93329 , n93330 , 
     n93331 , n93332 , n93333 , n93334 , n93335 , n93336 , n93337 , n93338 , n93339 , n93340 , 
     n93341 , n93342 , n93343 , n93344 , n93345 , n93346 , n93347 , n93348 , n93349 , n93350 , 
     n93351 , n93352 , n93353 , n93354 , n93355 , n93356 , n93357 , n93358 , n93359 , n93360 , 
     n93361 , n93362 , n93363 , n93364 , n93365 , n93366 , n93367 , n93368 , n93369 , n93370 , 
     n93371 , n93372 , n93373 , n93374 , n93375 , n93376 , n93377 , n93378 , n93379 , n93380 , 
     n93381 , n93382 , n93383 , n93384 , n93385 , n93386 , n93387 , n93388 , n93389 , n93390 , 
     n93391 , n93392 , n93393 , n93394 , n93395 , n93396 , n93397 , n93398 , n93399 , n93400 , 
     n93401 , n93402 , n93403 , n93404 , n93405 , n93406 , n93407 , n93408 , n93409 , n93410 , 
     n93411 , n93412 , n93413 , n93414 , n93415 , n93416 , n93417 , n93418 , n93419 , n93420 , 
     n93421 , n93422 , n93423 , n93424 , n93425 , n93426 , n93427 , n93428 , n93429 , n93430 , 
     n93431 , n93432 , n93433 , n93434 , n93435 , n93436 , n93437 , n93438 , n93439 , n93440 , 
     n93441 , n93442 , n93443 , n93444 , n93445 , n93446 , n93447 , n93448 , n93449 , n93450 , 
     n93451 , n93452 , n93453 , n93454 , n93455 , n93456 , n93457 , n93458 , n93459 , n93460 , 
     n93461 , n93462 , n93463 , n93464 , n93465 , n93466 , n93467 , n93468 , n93469 , n93470 , 
     n93471 , n93472 , n93473 , n93474 , n93475 , n93476 , n93477 , n93478 , n93479 , n93480 , 
     n93481 , n93482 , n93483 , n93484 , n93485 , n93486 , n93487 , n93488 , n93489 , n93490 , 
     n93491 , n93492 , n93493 , n93494 , n93495 , n93496 , n93497 , n93498 , n93499 , n93500 , 
     n93501 , n93502 , n93503 , n93504 , n93505 , n93506 , n93507 , n93508 , n93509 , n93510 , 
     n93511 , n93512 , n93513 , n93514 , n93515 , n93516 , n93517 , n93518 , n93519 , n93520 , 
     n93521 , n93522 , n93523 , n93524 , n93525 , n93526 , n93527 , n93528 , n93529 , n93530 , 
     n93531 , n93532 , n93533 , n93534 , n93535 , n93536 , n93537 , n93538 , n93539 , n93540 , 
     n93541 , n93542 , n93543 , n93544 , n93545 , n93546 , n93547 , n93548 , n93549 , n93550 , 
     n93551 , n93552 , n93553 , n93554 , n93555 , n93556 , n93557 , n93558 , n93559 , n93560 , 
     n93561 , n93562 , n93563 , n93564 , n93565 , n93566 , n93567 , n93568 , n93569 , n93570 , 
     n93571 , n93572 , n93573 , n93574 , n93575 , n93576 , n93577 , n93578 , n93579 , n93580 , 
     n93581 , n93582 , n93583 , n93584 , n93585 , n93586 , n93587 , n93588 , n93589 , n93590 , 
     n93591 , n93592 , n93593 , n93594 , n93595 , n93596 , n93597 , n93598 , n93599 , n93600 , 
     n93601 , n93602 , n93603 , n93604 , n93605 , n93606 , n93607 , n93608 , n93609 , n93610 , 
     n93611 , n93612 , n93613 , n93614 , n93615 , n93616 , n93617 , n93618 , n93619 , n93620 , 
     n93621 , n93622 , n93623 , n93624 , n93625 , n93626 , n93627 , n93628 , n93629 , n93630 , 
     n93631 , n93632 , n93633 , n93634 , n93635 , n93636 , n93637 , n93638 , n93639 , n93640 , 
     n93641 , n93642 , n93643 , n93644 , n93645 , n93646 , n93647 , n93648 , n93649 , n93650 , 
     n93651 , n93652 , n93653 , n93654 , n93655 , n93656 , n93657 , n93658 , n93659 , n93660 , 
     n93661 , n93662 , n93663 , n93664 , n93665 , n93666 , n93667 , n93668 , n93669 , n93670 , 
     n93671 , n93672 , n93673 , n93674 , n93675 , n93676 , n93677 , n93678 , n93679 , n93680 , 
     n93681 , n93682 , n93683 , n93684 , n93685 , n93686 , n93687 , n93688 , n93689 , n93690 , 
     n93691 , n93692 , n93693 , n93694 , n93695 , n93696 , n93697 , n93698 , n93699 , n93700 , 
     n93701 , n93702 , n93703 , n93704 , n93705 , n93706 , n93707 , n93708 , n93709 , n93710 , 
     n93711 , n93712 , n93713 , n93714 , n93715 , n93716 , n93717 , n93718 , n93719 , n93720 , 
     n93721 , n93722 , n93723 , n93724 , n93725 , n93726 , n93727 , n93728 , n93729 , n93730 , 
     n93731 , n93732 , n93733 , n93734 , n93735 , n93736 , n93737 , n93738 , n93739 , n93740 , 
     n93741 , n93742 , n93743 , n93744 , n93745 , n93746 , n93747 , n93748 , n93749 , n93750 , 
     n93751 , n93752 , n93753 , n93754 , n93755 , n93756 , n93757 , n93758 , n93759 , n93760 , 
     n93761 , n93762 , n93763 , n93764 , n93765 , n93766 , n93767 , n93768 , n93769 , n93770 , 
     n93771 , n93772 , n93773 , n93774 , n93775 , n93776 , n93777 , n93778 , n93779 , n93780 , 
     n93781 , n93782 , n93783 , n93784 , n93785 , n93786 , n93787 , n93788 , n93789 , n93790 , 
     n93791 , n93792 , n93793 , n93794 , n93795 , n93796 , n93797 , n93798 , n93799 , n93800 , 
     n93801 , n93802 , n93803 , n93804 , n93805 , n93806 , n93807 , n93808 , n93809 , n93810 , 
     n93811 , n93812 , n93813 , n93814 , n93815 , n93816 , n93817 , n93818 , n93819 , n93820 , 
     n93821 , n93822 , n93823 , n93824 , n93825 , n93826 , n93827 , n93828 , n93829 , n93830 , 
     n93831 , n93832 , n93833 , n93834 , n93835 , n93836 , n93837 , n93838 , n93839 , n93840 , 
     n93841 , n93842 , n93843 , n93844 , n93845 , n93846 , n93847 , n93848 , n93849 , n93850 , 
     n93851 , n93852 , n93853 , n93854 , n93855 , n93856 , n93857 , n93858 , n93859 , n93860 , 
     n93861 , n93862 , n93863 , n93864 , n93865 , n93866 , n93867 , n93868 , n93869 , n93870 , 
     n93871 , n93872 , n93873 , n93874 , n93875 , n93876 , n93877 , n93878 , n93879 , n93880 , 
     n93881 , n93882 , n93883 , n93884 , n93885 , n93886 , n93887 , n93888 , n93889 , n93890 , 
     n93891 , n93892 , n93893 , n93894 , n93895 , n93896 , n93897 , n93898 , n93899 , n93900 , 
     n93901 , n93902 , n93903 , n93904 , n93905 , n93906 , n93907 , n93908 , n93909 , n93910 , 
     n93911 , n93912 , n93913 , n93914 , n93915 , n93916 , n93917 , n93918 , n93919 , n93920 , 
     n93921 , n93922 , n93923 , n93924 , n93925 , n93926 , n93927 , n93928 , n93929 , n93930 , 
     n93931 , n93932 , n93933 , n93934 , n93935 , n93936 , n93937 , n93938 , n93939 , n93940 , 
     n93941 , n93942 , n93943 , n93944 , n93945 , n93946 , n93947 , n93948 , n93949 , n93950 , 
     n93951 , n93952 , n93953 , n93954 , n93955 , n93956 , n93957 , n93958 , n93959 , n93960 , 
     n93961 , n93962 , n93963 , n93964 , n93965 , n93966 , n93967 , n93968 , n93969 , n93970 , 
     n93971 , n93972 , n93973 , n93974 , n93975 , n93976 , n93977 , n93978 , n93979 , n93980 , 
     n93981 , n93982 , n93983 , n93984 , n93985 , n93986 , n93987 , n93988 , n93989 , n93990 , 
     n93991 , n93992 , n93993 , n93994 , n93995 , n93996 , n93997 , n93998 , n93999 , n94000 , 
     n94001 , n94002 , n94003 , n94004 , n94005 , n94006 , n94007 , n94008 , n94009 , n94010 , 
     n94011 , n94012 , n94013 , n94014 , n94015 , n94016 , n94017 , n94018 , n94019 , n94020 , 
     n94021 , n94022 , n94023 , n94024 , n94025 , n94026 , n94027 , n94028 , n94029 , n94030 , 
     n94031 , n94032 , n94033 , n94034 , n94035 , n94036 , n94037 , n94038 , n94039 , n94040 , 
     n94041 , n94042 , n94043 , n94044 , n94045 , n94046 , n94047 , n94048 , n94049 , n94050 , 
     n94051 , n94052 , n94053 , n94054 , n94055 , n94056 , n94057 , n94058 , n94059 , n94060 , 
     n94061 , n94062 , n94063 , n94064 , n94065 , n94066 , n94067 , n94068 , n94069 , n94070 , 
     n94071 , n94072 , n94073 , n94074 , n94075 , n94076 , n94077 , n94078 , n94079 , n94080 , 
     n94081 , n94082 , n94083 , n94084 , n94085 , n94086 , n94087 , n94088 , n94089 , n94090 , 
     n94091 , n94092 , n94093 , n94094 , n94095 , n94096 , n94097 , n94098 , n94099 , n94100 , 
     n94101 , n94102 , n94103 , n94104 , n94105 , n94106 , n94107 , n94108 , n94109 , n94110 , 
     n94111 , n94112 , n94113 , n94114 , n94115 , n94116 , n94117 , n94118 , n94119 , n94120 , 
     n94121 , n94122 , n94123 , n94124 , n94125 , n94126 , n94127 , n94128 , n94129 , n94130 , 
     n94131 , n94132 , n94133 , n94134 , n94135 , n94136 , n94137 , n94138 , n94139 , n94140 , 
     n94141 , n94142 , n94143 , n94144 , n94145 , n94146 , n94147 , n94148 , n94149 , n94150 , 
     n94151 , n94152 , n94153 , n94154 , n94155 , n94156 , n94157 , n94158 , n94159 , n94160 , 
     n94161 , n94162 , n94163 , n94164 , n94165 , n94166 , n94167 , n94168 , n94169 , n94170 , 
     n94171 , n94172 , n94173 , n94174 , n94175 , n94176 , n94177 , n94178 , n94179 , n94180 , 
     n94181 , n94182 , n94183 , n94184 , n94185 , n94186 , n94187 , n94188 , n94189 , n94190 , 
     n94191 , n94192 , n94193 , n94194 , n94195 , n94196 , n94197 , n94198 , n94199 , n94200 , 
     n94201 , n94202 , n94203 , n94204 , n94205 , n94206 , n94207 , n94208 , n94209 , n94210 , 
     n94211 , n94212 , n94213 , n94214 , n94215 , n94216 , n94217 , n94218 , n94219 , n94220 , 
     n94221 , n94222 , n94223 , n94224 , n94225 , n94226 , n94227 , n94228 , n94229 , n94230 , 
     n94231 , n94232 , n94233 , n94234 , n94235 , n94236 , n94237 , n94238 , n94239 , n94240 , 
     n94241 , n94242 , n94243 , n94244 , n94245 , n94246 , n94247 , n94248 , n94249 , n94250 , 
     n94251 , n94252 , n94253 , n94254 , n94255 , n94256 , n94257 , n94258 , n94259 , n94260 , 
     n94261 , n94262 , n94263 , n94264 , n94265 , n94266 , n94267 , n94268 , n94269 , n94270 , 
     n94271 , n94272 , n94273 , n94274 , n94275 , n94276 , n94277 , n94278 , n94279 , n94280 , 
     n94281 , n94282 , n94283 , n94284 , n94285 , n94286 , n94287 , n94288 , n94289 , n94290 , 
     n94291 , n94292 , n94293 , n94294 , n94295 , n94296 , n94297 , n94298 , n94299 , n94300 , 
     n94301 , n94302 , n94303 , n94304 , n94305 , n94306 , n94307 , n94308 , n94309 , n94310 , 
     n94311 , n94312 , n94313 , n94314 , n94315 , n94316 , n94317 , n94318 , n94319 , n94320 , 
     n94321 , n94322 , n94323 , n94324 , n94325 , n94326 , n94327 , n94328 , n94329 , n94330 , 
     n94331 , n94332 , n94333 , n94334 , n94335 , n94336 , n94337 , n94338 , n94339 , n94340 , 
     n94341 , n94342 , n94343 , n94344 , n94345 , n94346 , n94347 , n94348 , n94349 , n94350 , 
     n94351 , n94352 , n94353 , n94354 , n94355 , n94356 , n94357 , n94358 , n94359 , n94360 , 
     n94361 , n94362 , n94363 , n94364 , n94365 , n94366 , n94367 , n94368 , n94369 , n94370 , 
     n94371 , n94372 , n94373 , n94374 , n94375 , n94376 , n94377 , n94378 , n94379 , n94380 , 
     n94381 , n94382 , n94383 , n94384 , n94385 , n94386 , n94387 , n94388 , n94389 , n94390 , 
     n94391 , n94392 , n94393 , n94394 , n94395 , n94396 , n94397 , n94398 , n94399 , n94400 , 
     n94401 , n94402 , n94403 , n94404 , n94405 , n94406 , n94407 , n94408 , n94409 , n94410 , 
     n94411 , n94412 , n94413 , n94414 , n94415 , n94416 , n94417 , n94418 , n94419 , n94420 , 
     n94421 , n94422 , n94423 , n94424 , n94425 , n94426 , n94427 , n94428 , n94429 , n94430 , 
     n94431 , n94432 , n94433 , n94434 , n94435 , n94436 , n94437 , n94438 , n94439 , n94440 , 
     n94441 , n94442 , n94443 , n94444 , n94445 , n94446 , n94447 , n94448 , n94449 , n94450 , 
     n94451 , n94452 , n94453 , n94454 , n94455 , n94456 , n94457 , n94458 , n94459 , n94460 , 
     n94461 , n94462 , n94463 , n94464 , n94465 , n94466 , n94467 , n94468 , n94469 , n94470 , 
     n94471 , n94472 , n94473 , n94474 , n94475 , n94476 , n94477 , n94478 , n94479 , n94480 , 
     n94481 , n94482 , n94483 , n94484 , n94485 , n94486 , n94487 , n94488 , n94489 , n94490 , 
     n94491 , n94492 , n94493 , n94494 , n94495 , n94496 , n94497 , n94498 , n94499 , n94500 , 
     n94501 , n94502 , n94503 , n94504 , n94505 , n94506 , n94507 , n94508 , n94509 , n94510 , 
     n94511 , n94512 , n94513 , n94514 , n94515 , n94516 , n94517 , n94518 , n94519 , n94520 , 
     n94521 , n94522 , n94523 , n94524 , n94525 , n94526 , n94527 , n94528 , n94529 , n94530 , 
     n94531 , n94532 , n94533 , n94534 , n94535 , n94536 , n94537 , n94538 , n94539 , n94540 , 
     n94541 , n94542 , n94543 , n94544 , n94545 , n94546 , n94547 , n94548 , n94549 , n94550 , 
     n94551 , n94552 , n94553 , n94554 , n94555 , n94556 , n94557 , n94558 , n94559 , n94560 , 
     n94561 , n94562 , n94563 , n94564 , n94565 , n94566 , n94567 , n94568 , n94569 , n94570 , 
     n94571 , n94572 , n94573 , n94574 , n94575 , n94576 , n94577 , n94578 , n94579 , n94580 , 
     n94581 , n94582 , n94583 , n94584 , n94585 , n94586 , n94587 , n94588 , n94589 , n94590 , 
     n94591 , n94592 , n94593 , n94594 , n94595 , n94596 , n94597 , n94598 , n94599 , n94600 , 
     n94601 , n94602 , n94603 , n94604 , n94605 , n94606 , n94607 , n94608 , n94609 , n94610 , 
     n94611 , n94612 , n94613 , n94614 , n94615 , n94616 , n94617 , n94618 , n94619 , n94620 , 
     n94621 , n94622 , n94623 , n94624 , n94625 , n94626 , n94627 , n94628 , n94629 , n94630 , 
     n94631 , n94632 , n94633 , n94634 , n94635 , n94636 , n94637 , n94638 , n94639 , n94640 , 
     n94641 , n94642 , n94643 , n94644 , n94645 , n94646 , n94647 , n94648 , n94649 , n94650 , 
     n94651 , n94652 , n94653 , n94654 , n94655 , n94656 , n94657 , n94658 , n94659 , n94660 , 
     n94661 , n94662 , n94663 , n94664 , n94665 , n94666 , n94667 , n94668 , n94669 , n94670 , 
     n94671 , n94672 , n94673 , n94674 , n94675 , n94676 , n94677 , n94678 , n94679 , n94680 , 
     n94681 , n94682 , n94683 , n94684 , n94685 , n94686 , n94687 , n94688 , n94689 , n94690 , 
     n94691 , n94692 , n94693 , n94694 , n94695 , n94696 , n94697 , n94698 , n94699 , n94700 , 
     n94701 , n94702 , n94703 , n94704 , n94705 , n94706 , n94707 , n94708 , n94709 , n94710 , 
     n94711 , n94712 , n94713 , n94714 , n94715 , n94716 , n94717 , n94718 , n94719 , n94720 , 
     n94721 , n94722 , n94723 , n94724 , n94725 , n94726 , n94727 , n94728 , n94729 , n94730 , 
     n94731 , n94732 , n94733 , n94734 , n94735 , n94736 , n94737 , n94738 , n94739 , n94740 , 
     n94741 , n94742 , n94743 , n94744 , n94745 , n94746 , n94747 , n94748 , n94749 , n94750 , 
     n94751 , n94752 , n94753 , n94754 , n94755 , n94756 , n94757 , n94758 , n94759 , n94760 , 
     n94761 , n94762 , n94763 , n94764 , n94765 , n94766 , n94767 , n94768 , n94769 , n94770 , 
     n94771 , n94772 , n94773 , n94774 , n94775 , n94776 , n94777 , n94778 , n94779 , n94780 , 
     n94781 , n94782 , n94783 , n94784 , n94785 , n94786 , n94787 , n94788 , n94789 , n94790 , 
     n94791 , n94792 , n94793 , n94794 , n94795 , n94796 , n94797 , n94798 , n94799 , n94800 , 
     n94801 , n94802 , n94803 , n94804 , n94805 , n94806 , n94807 , n94808 , n94809 , n94810 , 
     n94811 , n94812 , n94813 , n94814 , n94815 , n94816 , n94817 , n94818 , n94819 , n94820 , 
     n94821 , n94822 , n94823 , n94824 , n94825 , n94826 , n94827 , n94828 , n94829 , n94830 , 
     n94831 , n94832 , n94833 , n94834 , n94835 , n94836 , n94837 , n94838 , n94839 , n94840 , 
     n94841 , n94842 , n94843 , n94844 , n94845 , n94846 , n94847 , n94848 , n94849 , n94850 , 
     n94851 , n94852 , n94853 , n94854 , n94855 , n94856 , n94857 , n94858 , n94859 , n94860 , 
     n94861 , n94862 , n94863 , n94864 , n94865 , n94866 , n94867 , n94868 , n94869 , n94870 , 
     n94871 , n94872 , n94873 , n94874 , n94875 , n94876 , n94877 , n94878 , n94879 , n94880 , 
     n94881 , n94882 , n94883 , n94884 , n94885 , n94886 , n94887 , n94888 , n94889 , n94890 , 
     n94891 , n94892 , n94893 , n94894 , n94895 , n94896 , n94897 , n94898 , n94899 , n94900 , 
     n94901 , n94902 , n94903 , n94904 , n94905 , n94906 , n94907 , n94908 , n94909 , n94910 , 
     n94911 , n94912 , n94913 , n94914 , n94915 , n94916 , n94917 , n94918 , n94919 , n94920 , 
     n94921 , n94922 , n94923 , n94924 , n94925 , n94926 , n94927 , n94928 , n94929 , n94930 , 
     n94931 , n94932 , n94933 , n94934 , n94935 , n94936 , n94937 , n94938 , n94939 , n94940 , 
     n94941 , n94942 , n94943 , n94944 , n94945 , n94946 , n94947 , n94948 , n94949 , n94950 , 
     n94951 , n94952 , n94953 , n94954 , n94955 , n94956 , n94957 , n94958 , n94959 , n94960 , 
     n94961 , n94962 , n94963 , n94964 , n94965 , n94966 , n94967 , n94968 , n94969 , n94970 , 
     n94971 , n94972 , n94973 , n94974 , n94975 , n94976 , n94977 , n94978 , n94979 , n94980 , 
     n94981 , n94982 , n94983 , n94984 , n94985 , n94986 , n94987 , n94988 , n94989 , n94990 , 
     n94991 , n94992 , n94993 , n94994 , n94995 , n94996 , n94997 , n94998 , n94999 , n95000 , 
     n95001 , n95002 , n95003 , n95004 , n95005 , n95006 , n95007 , n95008 , n95009 , n95010 , 
     n95011 , n95012 , n95013 , n95014 , n95015 , n95016 , n95017 , n95018 , n95019 , n95020 , 
     n95021 , n95022 , n95023 , n95024 , n95025 , n95026 , n95027 , n95028 , n95029 , n95030 , 
     n95031 , n95032 , n95033 , n95034 , n95035 , n95036 , n95037 , n95038 , n95039 , n95040 , 
     n95041 , n95042 , n95043 , n95044 , n95045 , n95046 , n95047 , n95048 , n95049 , n95050 , 
     n95051 , n95052 , n95053 , n95054 , n95055 , n95056 , n95057 , n95058 , n95059 , n95060 , 
     n95061 , n95062 , n95063 , n95064 , n95065 , n95066 , n95067 , n95068 , n95069 , n95070 , 
     n95071 , n95072 , n95073 , n95074 , n95075 , n95076 , n95077 , n95078 , n95079 , n95080 , 
     n95081 , n95082 , n95083 , n95084 , n95085 , n95086 , n95087 , n95088 , n95089 , n95090 , 
     n95091 , n95092 , n95093 , n95094 , n95095 , n95096 , n95097 , n95098 , n95099 , n95100 , 
     n95101 , n95102 , n95103 , n95104 , n95105 , n95106 , n95107 , n95108 , n95109 , n95110 , 
     n95111 , n95112 , n95113 , n95114 , n95115 , n95116 , n95117 , n95118 , n95119 , n95120 , 
     n95121 , n95122 , n95123 , n95124 , n95125 , n95126 , n95127 , n95128 , n95129 , n95130 , 
     n95131 , n95132 , n95133 , n95134 , n95135 , n95136 , n95137 , n95138 , n95139 , n95140 , 
     n95141 , n95142 , n95143 , n95144 , n95145 , n95146 , n95147 , n95148 , n95149 , n95150 , 
     n95151 , n95152 , n95153 , n95154 , n95155 , n95156 , n95157 , n95158 , n95159 , n95160 , 
     n95161 , n95162 , n95163 , n95164 , n95165 , n95166 , n95167 , n95168 , n95169 , n95170 , 
     n95171 , n95172 , n95173 , n95174 , n95175 , n95176 , n95177 , n95178 , n95179 , n95180 , 
     n95181 , n95182 , n95183 , n95184 , n95185 , n95186 , n95187 , n95188 , n95189 , n95190 , 
     n95191 , n95192 , n95193 , n95194 , n95195 , n95196 , n95197 , n95198 , n95199 , n95200 , 
     n95201 , n95202 , n95203 , n95204 , n95205 , n95206 , n95207 , n95208 , n95209 , n95210 , 
     n95211 , n95212 , n95213 , n95214 , n95215 , n95216 , n95217 , n95218 , n95219 , n95220 , 
     n95221 , n95222 , n95223 , n95224 , n95225 , n95226 , n95227 , n95228 , n95229 , n95230 , 
     n95231 , n95232 , n95233 , n95234 , n95235 , n95236 , n95237 , n95238 , n95239 , n95240 , 
     n95241 , n95242 , n95243 , n95244 , n95245 , n95246 , n95247 , n95248 , n95249 , n95250 , 
     n95251 , n95252 , n95253 , n95254 , n95255 , n95256 , n95257 , n95258 , n95259 , n95260 , 
     n95261 , n95262 , n95263 , n95264 , n95265 , n95266 , n95267 , n95268 , n95269 , n95270 , 
     n95271 , n95272 , n95273 , n95274 , n95275 , n95276 , n95277 , n95278 , n95279 , n95280 , 
     n95281 , n95282 , n95283 , n95284 , n95285 , n95286 , n95287 , n95288 , n95289 , n95290 , 
     n95291 , n95292 , n95293 , n95294 , n95295 , n95296 , n95297 , n95298 , n95299 , n95300 , 
     n95301 , n95302 , n95303 , n95304 , n95305 , n95306 , n95307 , n95308 , n95309 , n95310 , 
     n95311 , n95312 , n95313 , n95314 , n95315 , n95316 , n95317 , n95318 , n95319 , n95320 , 
     n95321 , n95322 , n95323 , n95324 , n95325 , n95326 , n95327 , n95328 , n95329 , n95330 , 
     n95331 , n95332 , n95333 , n95334 , n95335 , n95336 , n95337 , n95338 , n95339 , n95340 , 
     n95341 , n95342 , n95343 , n95344 , n95345 , n95346 , n95347 , n95348 , n95349 , n95350 , 
     n95351 , n95352 , n95353 , n95354 , n95355 , n95356 , n95357 , n95358 , n95359 , n95360 , 
     n95361 , n95362 , n95363 , n95364 , n95365 , n95366 , n95367 , n95368 , n95369 , n95370 , 
     n95371 , n95372 , n95373 , n95374 , n95375 , n95376 , n95377 , n95378 , n95379 , n95380 , 
     n95381 , n95382 , n95383 , n95384 , n95385 , n95386 , n95387 , n95388 , n95389 , n95390 , 
     n95391 , n95392 , n95393 , n95394 , n95395 , n95396 , n95397 , n95398 , n95399 , n95400 , 
     n95401 , n95402 , n95403 , n95404 , n95405 , n95406 , n95407 , n95408 , n95409 , n95410 , 
     n95411 , n95412 , n95413 , n95414 , n95415 , n95416 , n95417 , n95418 , n95419 , n95420 , 
     n95421 , n95422 , n95423 , n95424 , n95425 , n95426 , n95427 , n95428 , n95429 , n95430 , 
     n95431 , n95432 , n95433 , n95434 , n95435 , n95436 , n95437 , n95438 , n95439 , n95440 , 
     n95441 , n95442 , n95443 , n95444 , n95445 , n95446 , n95447 , n95448 , n95449 , n95450 , 
     n95451 , n95452 , n95453 , n95454 , n95455 , n95456 , n95457 , n95458 , n95459 , n95460 , 
     n95461 , n95462 , n95463 , n95464 , n95465 , n95466 , n95467 , n95468 , n95469 , n95470 , 
     n95471 , n95472 , n95473 , n95474 , n95475 , n95476 , n95477 , n95478 , n95479 , n95480 , 
     n95481 , n95482 , n95483 , n95484 , n95485 , n95486 , n95487 , n95488 , n95489 , n95490 , 
     n95491 , n95492 , n95493 , n95494 , n95495 , n95496 , n95497 , n95498 , n95499 , n95500 , 
     n95501 , n95502 , n95503 , n95504 , n95505 , n95506 , n95507 , n95508 , n95509 , n95510 , 
     n95511 , n95512 , n95513 , n95514 , n95515 , n95516 , n95517 , n95518 , n95519 , n95520 , 
     n95521 , n95522 , n95523 , n95524 , n95525 , n95526 , n95527 , n95528 , n95529 , n95530 , 
     n95531 , n95532 , n95533 , n95534 , n95535 , n95536 , n95537 , n95538 , n95539 , n95540 , 
     n95541 , n95542 , n95543 , n95544 , n95545 , n95546 , n95547 , n95548 , n95549 , n95550 , 
     n95551 , n95552 , n95553 , n95554 , n95555 , n95556 , n95557 , n95558 , n95559 , n95560 , 
     n95561 , n95562 , n95563 , n95564 , n95565 , n95566 , n95567 , n95568 , n95569 , n95570 , 
     n95571 , n95572 , n95573 , n95574 , n95575 , n95576 , n95577 , n95578 , n95579 , n95580 , 
     n95581 , n95582 , n95583 , n95584 , n95585 , n95586 , n95587 , n95588 , n95589 , n95590 , 
     n95591 , n95592 , n95593 , n95594 , n95595 , n95596 , n95597 , n95598 , n95599 , n95600 , 
     n95601 , n95602 , n95603 , n95604 , n95605 , n95606 , n95607 , n95608 , n95609 , n95610 , 
     n95611 , n95612 , n95613 , n95614 , n95615 , n95616 , n95617 , n95618 , n95619 , n95620 , 
     n95621 , n95622 , n95623 , n95624 , n95625 , n95626 , n95627 , n95628 , n95629 , n95630 , 
     n95631 , n95632 , n95633 , n95634 , n95635 , n95636 , n95637 , n95638 , n95639 , n95640 , 
     n95641 , n95642 , n95643 , n95644 , n95645 , n95646 , n95647 , n95648 , n95649 , n95650 , 
     n95651 , n95652 , n95653 , n95654 , n95655 , n95656 , n95657 , n95658 , n95659 , n95660 , 
     n95661 , n95662 , n95663 , n95664 , n95665 , n95666 , n95667 , n95668 , n95669 , n95670 , 
     n95671 , n95672 , n95673 , n95674 , n95675 , n95676 , n95677 , n95678 , n95679 , n95680 , 
     n95681 , n95682 , n95683 , n95684 , n95685 , n95686 , n95687 , n95688 , n95689 , n95690 , 
     n95691 , n95692 , n95693 , n95694 , n95695 , n95696 , n95697 , n95698 , n95699 , n95700 , 
     n95701 , n95702 , n95703 , n95704 , n95705 , n95706 , n95707 , n95708 , n95709 , n95710 , 
     n95711 , n95712 , n95713 , n95714 , n95715 , n95716 , n95717 , n95718 , n95719 , n95720 , 
     n95721 , n95722 , n95723 , n95724 , n95725 , n95726 , n95727 , n95728 , n95729 , n95730 , 
     n95731 , n95732 , n95733 , n95734 , n95735 , n95736 , n95737 , n95738 , n95739 , n95740 , 
     n95741 , n95742 , n95743 , n95744 , n95745 , n95746 , n95747 , n95748 , n95749 , n95750 , 
     n95751 , n95752 , n95753 , n95754 , n95755 , n95756 , n95757 , n95758 , n95759 , n95760 , 
     n95761 , n95762 , n95763 , n95764 , n95765 , n95766 , n95767 , n95768 , n95769 , n95770 , 
     n95771 , n95772 , n95773 , n95774 , n95775 , n95776 , n95777 , n95778 , n95779 , n95780 , 
     n95781 , n95782 , n95783 , n95784 , n95785 , n95786 , n95787 , n95788 , n95789 , n95790 , 
     n95791 , n95792 , n95793 , n95794 , n95795 , n95796 , n95797 , n95798 , n95799 , n95800 , 
     n95801 , n95802 , n95803 , n95804 , n95805 , n95806 , n95807 , n95808 , n95809 , n95810 , 
     n95811 , n95812 , n95813 , n95814 , n95815 , n95816 , n95817 , n95818 , n95819 , n95820 , 
     n95821 , n95822 , n95823 , n95824 , n95825 , n95826 , n95827 , n95828 , n95829 , n95830 , 
     n95831 , n95832 , n95833 , n95834 , n95835 , n95836 , n95837 , n95838 , n95839 , n95840 , 
     n95841 , n95842 , n95843 , n95844 , n95845 , n95846 , n95847 , n95848 , n95849 , n95850 , 
     n95851 , n95852 , n95853 , n95854 , n95855 , n95856 , n95857 , n95858 , n95859 , n95860 , 
     n95861 , n95862 , n95863 , n95864 , n95865 , n95866 , n95867 , n95868 , n95869 , n95870 , 
     n95871 , n95872 , n95873 , n95874 , n95875 , n95876 , n95877 , n95878 , n95879 , n95880 , 
     n95881 , n95882 , n95883 , n95884 , n95885 , n95886 , n95887 , n95888 , n95889 , n95890 , 
     n95891 , n95892 , n95893 , n95894 , n95895 , n95896 , n95897 , n95898 , n95899 , n95900 , 
     n95901 , n95902 , n95903 , n95904 , n95905 , n95906 , n95907 , n95908 , n95909 , n95910 , 
     n95911 , n95912 , n95913 , n95914 , n95915 , n95916 , n95917 , n95918 , n95919 , n95920 , 
     n95921 , n95922 , n95923 , n95924 , n95925 , n95926 , n95927 , n95928 , n95929 , n95930 , 
     n95931 , n95932 , n95933 , n95934 , n95935 , n95936 , n95937 , n95938 , n95939 , n95940 , 
     n95941 , n95942 , n95943 , n95944 , n95945 , n95946 , n95947 , n95948 , n95949 , n95950 , 
     n95951 , n95952 , n95953 , n95954 , n95955 , n95956 , n95957 , n95958 , n95959 , n95960 , 
     n95961 , n95962 , n95963 , n95964 , n95965 , n95966 , n95967 , n95968 , n95969 , n95970 , 
     n95971 , n95972 , n95973 , n95974 , n95975 , n95976 , n95977 , n95978 , n95979 , n95980 , 
     n95981 , n95982 , n95983 , n95984 , n95985 , n95986 , n95987 , n95988 , n95989 , n95990 , 
     n95991 , n95992 , n95993 , n95994 , n95995 , n95996 , n95997 , n95998 , n95999 , n96000 , 
     n96001 , n96002 , n96003 , n96004 , n96005 , n96006 , n96007 , n96008 , n96009 , n96010 , 
     n96011 , n96012 , n96013 , n96014 , n96015 , n96016 , n96017 , n96018 , n96019 , n96020 , 
     n96021 , n96022 , n96023 , n96024 , n96025 , n96026 , n96027 , n96028 , n96029 , n96030 , 
     n96031 , n96032 , n96033 , n96034 , n96035 , n96036 , n96037 , n96038 , n96039 , n96040 , 
     n96041 , n96042 , n96043 , n96044 , n96045 , n96046 , n96047 , n96048 , n96049 , n96050 , 
     n96051 , n96052 , n96053 , n96054 , n96055 , n96056 , n96057 , n96058 , n96059 , n96060 , 
     n96061 , n96062 , n96063 , n96064 , n96065 , n96066 , n96067 , n96068 , n96069 , n96070 , 
     n96071 , n96072 , n96073 , n96074 , n96075 , n96076 , n96077 , n96078 , n96079 , n96080 , 
     n96081 , n96082 , n96083 , n96084 , n96085 , n96086 , n96087 , n96088 , n96089 , n96090 , 
     n96091 , n96092 , n96093 , n96094 , n96095 , n96096 , n96097 , n96098 , n96099 , n96100 , 
     n96101 , n96102 , n96103 , n96104 , n96105 , n96106 , n96107 , n96108 , n96109 , n96110 , 
     n96111 , n96112 , n96113 , n96114 , n96115 , n96116 , n96117 , n96118 , n96119 , n96120 , 
     n96121 , n96122 , n96123 , n96124 , n96125 , n96126 , n96127 , n96128 , n96129 , n96130 , 
     n96131 , n96132 , n96133 , n96134 , n96135 , n96136 , n96137 , n96138 , n96139 , n96140 , 
     n96141 , n96142 , n96143 , n96144 , n96145 , n96146 , n96147 , n96148 , n96149 , n96150 , 
     n96151 , n96152 , n96153 , n96154 , n96155 , n96156 , n96157 , n96158 , n96159 , n96160 , 
     n96161 , n96162 , n96163 , n96164 , n96165 , n96166 , n96167 , n96168 , n96169 , n96170 , 
     n96171 , n96172 , n96173 , n96174 , n96175 , n96176 , n96177 , n96178 , n96179 , n96180 , 
     n96181 , n96182 , n96183 , n96184 , n96185 , n96186 , n96187 , n96188 , n96189 , n96190 , 
     n96191 , n96192 , n96193 , n96194 , n96195 , n96196 , n96197 , n96198 , n96199 , n96200 , 
     n96201 , n96202 , n96203 , n96204 , n96205 , n96206 , n96207 , n96208 , n96209 , n96210 , 
     n96211 , n96212 , n96213 , n96214 , n96215 , n96216 , n96217 , n96218 , n96219 , n96220 , 
     n96221 , n96222 , n96223 , n96224 , n96225 , n96226 , n96227 , n96228 , n96229 , n96230 , 
     n96231 , n96232 , n96233 , n96234 , n96235 , n96236 , n96237 , n96238 , n96239 , n96240 , 
     n96241 , n96242 , n96243 , n96244 , n96245 , n96246 , n96247 , n96248 , n96249 , n96250 , 
     n96251 , n96252 , n96253 , n96254 , n96255 , n96256 , n96257 , n96258 , n96259 , n96260 , 
     n96261 , n96262 , n96263 , n96264 , n96265 , n96266 , n96267 , n96268 , n96269 , n96270 , 
     n96271 , n96272 , n96273 , n96274 , n96275 , n96276 , n96277 , n96278 , n96279 , n96280 , 
     n96281 , n96282 , n96283 , n96284 , n96285 , n96286 , n96287 , n96288 , n96289 , n96290 , 
     n96291 , n96292 , n96293 , n96294 , n96295 , n96296 , n96297 , n96298 , n96299 , n96300 , 
     n96301 , n96302 , n96303 , n96304 , n96305 , n96306 , n96307 , n96308 , n96309 , n96310 , 
     n96311 , n96312 , n96313 , n96314 , n96315 , n96316 , n96317 , n96318 , n96319 , n96320 , 
     n96321 , n96322 , n96323 , n96324 , n96325 , n96326 , n96327 , n96328 , n96329 , n96330 , 
     n96331 , n96332 , n96333 , n96334 , n96335 , n96336 , n96337 , n96338 , n96339 , n96340 , 
     n96341 , n96342 , n96343 , n96344 , n96345 , n96346 , n96347 , n96348 , n96349 , n96350 , 
     n96351 , n96352 , n96353 , n96354 , n96355 , n96356 , n96357 , n96358 , n96359 , n96360 , 
     n96361 , n96362 , n96363 , n96364 , n96365 , n96366 , n96367 , n96368 , n96369 , n96370 , 
     n96371 , n96372 , n96373 , n96374 , n96375 , n96376 , n96377 , n96378 , n96379 , n96380 , 
     n96381 , n96382 , n96383 , n96384 , n96385 , n96386 , n96387 , n96388 , n96389 , n96390 , 
     n96391 , n96392 , n96393 , n96394 , n96395 , n96396 , n96397 , n96398 , n96399 , n96400 , 
     n96401 , n96402 , n96403 , n96404 , n96405 , n96406 , n96407 , n96408 , n96409 , n96410 , 
     n96411 , n96412 , n96413 , n96414 , n96415 , n96416 , n96417 , n96418 , n96419 , n96420 , 
     n96421 , n96422 , n96423 , n96424 , n96425 , n96426 , n96427 , n96428 , n96429 , n96430 , 
     n96431 , n96432 , n96433 , n96434 , n96435 , n96436 , n96437 , n96438 , n96439 , n96440 , 
     n96441 , n96442 , n96443 , n96444 , n96445 , n96446 , n96447 , n96448 , n96449 , n96450 , 
     n96451 , n96452 , n96453 , n96454 , n96455 , n96456 , n96457 , n96458 , n96459 , n96460 , 
     n96461 , n96462 , n96463 , n96464 , n96465 , n96466 , n96467 , n96468 , n96469 , n96470 , 
     n96471 , n96472 , n96473 , n96474 , n96475 , n96476 , n96477 , n96478 , n96479 , n96480 , 
     n96481 , n96482 , n96483 , n96484 , n96485 , n96486 , n96487 , n96488 , n96489 , n96490 , 
     n96491 , n96492 , n96493 , n96494 , n96495 , n96496 , n96497 , n96498 , n96499 , n96500 , 
     n96501 , n96502 , n96503 , n96504 , n96505 , n96506 , n96507 , n96508 , n96509 , n96510 , 
     n96511 , n96512 , n96513 , n96514 , n96515 , n96516 , n96517 , n96518 , n96519 , n96520 , 
     n96521 , n96522 , n96523 , n96524 , n96525 , n96526 , n96527 , n96528 , n96529 , n96530 , 
     n96531 , n96532 , n96533 , n96534 , n96535 , n96536 , n96537 , n96538 , n96539 , n96540 , 
     n96541 , n96542 , n96543 , n96544 , n96545 , n96546 , n96547 , n96548 , n96549 , n96550 , 
     n96551 , n96552 , n96553 , n96554 , n96555 , n96556 , n96557 , n96558 , n96559 , n96560 , 
     n96561 , n96562 , n96563 , n96564 , n96565 , n96566 , n96567 , n96568 , n96569 , n96570 , 
     n96571 , n96572 , n96573 , n96574 , n96575 , n96576 , n96577 , n96578 , n96579 , n96580 , 
     n96581 , n96582 , n96583 , n96584 , n96585 , n96586 , n96587 , n96588 , n96589 , n96590 , 
     n96591 , n96592 , n96593 , n96594 , n96595 , n96596 , n96597 , n96598 , n96599 , n96600 , 
     n96601 , n96602 , n96603 , n96604 , n96605 , n96606 , n96607 , n96608 , n96609 , n96610 , 
     n96611 , n96612 , n96613 , n96614 , n96615 , n96616 , n96617 , n96618 , n96619 , n96620 , 
     n96621 , n96622 , n96623 , n96624 , n96625 , n96626 , n96627 , n96628 , n96629 , n96630 , 
     n96631 , n96632 , n96633 , n96634 , n96635 , n96636 , n96637 , n96638 , n96639 , n96640 , 
     n96641 , n96642 , n96643 , n96644 , n96645 , n96646 , n96647 , n96648 , n96649 , n96650 , 
     n96651 , n96652 , n96653 , n96654 , n96655 , n96656 , n96657 , n96658 , n96659 , n96660 , 
     n96661 , n96662 , n96663 , n96664 , n96665 , n96666 , n96667 , n96668 , n96669 , n96670 , 
     n96671 , n96672 , n96673 , n96674 , n96675 , n96676 , n96677 , n96678 , n96679 , n96680 , 
     n96681 , n96682 , n96683 , n96684 , n96685 , n96686 , n96687 , n96688 , n96689 , n96690 , 
     n96691 , n96692 , n96693 , n96694 , n96695 , n96696 , n96697 , n96698 , n96699 , n96700 , 
     n96701 , n96702 , n96703 , n96704 , n96705 , n96706 , n96707 , n96708 , n96709 , n96710 , 
     n96711 , n96712 , n96713 , n96714 , n96715 , n96716 , n96717 , n96718 , n96719 , n96720 , 
     n96721 , n96722 , n96723 , n96724 , n96725 , n96726 , n96727 , n96728 , n96729 , n96730 , 
     n96731 , n96732 , n96733 , n96734 , n96735 , n96736 , n96737 , n96738 , n96739 , n96740 , 
     n96741 , n96742 , n96743 , n96744 , n96745 , n96746 , n96747 , n96748 , n96749 , n96750 , 
     n96751 , n96752 , n96753 , n96754 , n96755 , n96756 , n96757 , n96758 , n96759 , n96760 , 
     n96761 , n96762 , n96763 , n96764 , n96765 , n96766 , n96767 , n96768 , n96769 , n96770 , 
     n96771 , n96772 , n96773 , n96774 , n96775 , n96776 , n96777 , n96778 , n96779 , n96780 , 
     n96781 , n96782 , n96783 , n96784 , n96785 , n96786 , n96787 , n96788 , n96789 , n96790 , 
     n96791 , n96792 , n96793 , n96794 , n96795 , n96796 , n96797 , n96798 , n96799 , n96800 , 
     n96801 , n96802 , n96803 , n96804 , n96805 , n96806 , n96807 , n96808 , n96809 , n96810 , 
     n96811 , n96812 , n96813 , n96814 , n96815 , n96816 , n96817 , n96818 , n96819 , n96820 , 
     n96821 , n96822 , n96823 , n96824 , n96825 , n96826 , n96827 , n96828 , n96829 , n96830 , 
     n96831 , n96832 , n96833 , n96834 , n96835 , n96836 , n96837 , n96838 , n96839 , n96840 , 
     n96841 , n96842 , n96843 , n96844 , n96845 , n96846 , n96847 , n96848 , n96849 , n96850 , 
     n96851 , n96852 , n96853 , n96854 , n96855 , n96856 , n96857 , n96858 , n96859 , n96860 , 
     n96861 , n96862 , n96863 , n96864 , n96865 , n96866 , n96867 , n96868 , n96869 , n96870 , 
     n96871 , n96872 , n96873 , n96874 , n96875 , n96876 , n96877 , n96878 , n96879 , n96880 , 
     n96881 , n96882 , n96883 , n96884 , n96885 , n96886 , n96887 , n96888 , n96889 , n96890 , 
     n96891 , n96892 , n96893 , n96894 , n96895 , n96896 , n96897 , n96898 , n96899 , n96900 , 
     n96901 , n96902 , n96903 , n96904 , n96905 , n96906 , n96907 , n96908 , n96909 , n96910 , 
     n96911 , n96912 , n96913 , n96914 , n96915 , n96916 , n96917 , n96918 , n96919 , n96920 , 
     n96921 , n96922 , n96923 , n96924 , n96925 , n96926 , n96927 , n96928 , n96929 , n96930 , 
     n96931 , n96932 , n96933 , n96934 , n96935 , n96936 , n96937 , n96938 , n96939 , n96940 , 
     n96941 , n96942 , n96943 , n96944 , n96945 , n96946 , n96947 , n96948 , n96949 , n96950 , 
     n96951 , n96952 , n96953 , n96954 , n96955 , n96956 , n96957 , n96958 , n96959 , n96960 , 
     n96961 , n96962 , n96963 , n96964 , n96965 , n96966 , n96967 , n96968 , n96969 , n96970 , 
     n96971 , n96972 , n96973 , n96974 , n96975 , n96976 , n96977 , n96978 , n96979 , n96980 , 
     n96981 , n96982 , n96983 , n96984 , n96985 , n96986 , n96987 , n96988 , n96989 , n96990 , 
     n96991 , n96992 , n96993 , n96994 , n96995 ;
buf ( RI15b3e9d0_1 , n0 );
buf ( RI15b56850_817 , n1 );
buf ( RI15b51120_631 , n2 );
buf ( RI15b51288_634 , n3 );
buf ( RI15b51198_632 , n4 );
buf ( RI15b51210_633 , n5 );
buf ( RI15b4c2d8_464 , n6 );
buf ( RI15b51030_629 , n7 );
buf ( RI15b4c260_463 , n8 );
buf ( RI15b50fb8_628 , n9 );
buf ( RI15b4c1e8_462 , n10 );
buf ( RI15b50f40_627 , n11 );
buf ( RI15b4c170_461 , n12 );
buf ( RI15b50ec8_626 , n13 );
buf ( RI15b4c0f8_460 , n14 );
buf ( RI15b50e50_625 , n15 );
buf ( RI15b57750_849 , n16 );
buf ( RI15b4fb90_585 , n17 );
buf ( RI15b4f7d0_577 , n18 );
buf ( RI15b4f410_569 , n19 );
buf ( RI15b4f050_561 , n20 );
buf ( RI15b4ec90_553 , n21 );
buf ( RI15b4e8d0_545 , n22 );
buf ( RI15b4e510_537 , n23 );
buf ( RI15b4e150_529 , n24 );
buf ( RI15b4dd90_521 , n25 );
buf ( RI15b4d9d0_513 , n26 );
buf ( RI15b4d610_505 , n27 );
buf ( RI15b4d250_497 , n28 );
buf ( RI15b4ce90_489 , n29 );
buf ( RI15b4cad0_481 , n30 );
buf ( RI15b4c710_473 , n31 );
buf ( RI15b4c350_465 , n32 );
buf ( RI15b4fc08_586 , n33 );
buf ( RI15b4f848_578 , n34 );
buf ( RI15b4f488_570 , n35 );
buf ( RI15b4f0c8_562 , n36 );
buf ( RI15b4ed08_554 , n37 );
buf ( RI15b4e948_546 , n38 );
buf ( RI15b4e588_538 , n39 );
buf ( RI15b4e1c8_530 , n40 );
buf ( RI15b4de08_522 , n41 );
buf ( RI15b4da48_514 , n42 );
buf ( RI15b4d688_506 , n43 );
buf ( RI15b4d2c8_498 , n44 );
buf ( RI15b4cf08_490 , n45 );
buf ( RI15b4cb48_482 , n46 );
buf ( RI15b4c788_474 , n47 );
buf ( RI15b4c3c8_466 , n48 );
buf ( RI15b4fc80_587 , n49 );
buf ( RI15b4f8c0_579 , n50 );
buf ( RI15b4f500_571 , n51 );
buf ( RI15b4f140_563 , n52 );
buf ( RI15b4ed80_555 , n53 );
buf ( RI15b4e9c0_547 , n54 );
buf ( RI15b4e600_539 , n55 );
buf ( RI15b4e240_531 , n56 );
buf ( RI15b4de80_523 , n57 );
buf ( RI15b4dac0_515 , n58 );
buf ( RI15b4d700_507 , n59 );
buf ( RI15b4d340_499 , n60 );
buf ( RI15b4cf80_491 , n61 );
buf ( RI15b4cbc0_483 , n62 );
buf ( RI15b4c800_475 , n63 );
buf ( RI15b4c440_467 , n64 );
buf ( RI15b4fcf8_588 , n65 );
buf ( RI15b4f938_580 , n66 );
buf ( RI15b4f578_572 , n67 );
buf ( RI15b4f1b8_564 , n68 );
buf ( RI15b4edf8_556 , n69 );
buf ( RI15b4ea38_548 , n70 );
buf ( RI15b4e678_540 , n71 );
buf ( RI15b4e2b8_532 , n72 );
buf ( RI15b4def8_524 , n73 );
buf ( RI15b4db38_516 , n74 );
buf ( RI15b4d778_508 , n75 );
buf ( RI15b4d3b8_500 , n76 );
buf ( RI15b4cff8_492 , n77 );
buf ( RI15b4cc38_484 , n78 );
buf ( RI15b4c878_476 , n79 );
buf ( RI15b4c4b8_468 , n80 );
buf ( RI15b4fd70_589 , n81 );
buf ( RI15b4f9b0_581 , n82 );
buf ( RI15b4f5f0_573 , n83 );
buf ( RI15b4f230_565 , n84 );
buf ( RI15b4ee70_557 , n85 );
buf ( RI15b4eab0_549 , n86 );
buf ( RI15b4e6f0_541 , n87 );
buf ( RI15b4e330_533 , n88 );
buf ( RI15b4df70_525 , n89 );
buf ( RI15b4dbb0_517 , n90 );
buf ( RI15b4d7f0_509 , n91 );
buf ( RI15b4d430_501 , n92 );
buf ( RI15b4d070_493 , n93 );
buf ( RI15b4ccb0_485 , n94 );
buf ( RI15b4c8f0_477 , n95 );
buf ( RI15b4c530_469 , n96 );
buf ( RI15b4fde8_590 , n97 );
buf ( RI15b4fa28_582 , n98 );
buf ( RI15b4f668_574 , n99 );
buf ( RI15b4f2a8_566 , n100 );
buf ( RI15b4eee8_558 , n101 );
buf ( RI15b4eb28_550 , n102 );
buf ( RI15b4e768_542 , n103 );
buf ( RI15b4e3a8_534 , n104 );
buf ( RI15b4dfe8_526 , n105 );
buf ( RI15b4dc28_518 , n106 );
buf ( RI15b4d868_510 , n107 );
buf ( RI15b4d4a8_502 , n108 );
buf ( RI15b4d0e8_494 , n109 );
buf ( RI15b4cd28_486 , n110 );
buf ( RI15b4c968_478 , n111 );
buf ( RI15b4c5a8_470 , n112 );
buf ( RI15b4fe60_591 , n113 );
buf ( RI15b4faa0_583 , n114 );
buf ( RI15b4f6e0_575 , n115 );
buf ( RI15b4f320_567 , n116 );
buf ( RI15b4ef60_559 , n117 );
buf ( RI15b4eba0_551 , n118 );
buf ( RI15b4e7e0_543 , n119 );
buf ( RI15b4e420_535 , n120 );
buf ( RI15b4e060_527 , n121 );
buf ( RI15b4dca0_519 , n122 );
buf ( RI15b4d8e0_511 , n123 );
buf ( RI15b4d520_503 , n124 );
buf ( RI15b4d160_495 , n125 );
buf ( RI15b4cda0_487 , n126 );
buf ( RI15b4c9e0_479 , n127 );
buf ( RI15b4c620_471 , n128 );
buf ( RI15b4fed8_592 , n129 );
buf ( RI15b4fb18_584 , n130 );
buf ( RI15b4f758_576 , n131 );
buf ( RI15b4f398_568 , n132 );
buf ( RI15b4efd8_560 , n133 );
buf ( RI15b4ec18_552 , n134 );
buf ( RI15b4e858_544 , n135 );
buf ( RI15b4e498_536 , n136 );
buf ( RI15b4e0d8_528 , n137 );
buf ( RI15b4dd18_520 , n138 );
buf ( RI15b4d958_512 , n139 );
buf ( RI15b4d598_504 , n140 );
buf ( RI15b4d1d8_496 , n141 );
buf ( RI15b4ce18_488 , n142 );
buf ( RI15b4ca58_480 , n143 );
buf ( RI15b4c698_472 , n144 );
buf ( RI15b54780_747 , n145 );
buf ( RI15b547f8_748 , n146 );
buf ( RI15b54870_749 , n147 );
buf ( RI15b667c8_1362 , n148 );
buf ( RI15b66840_1363 , n149 );
buf ( RI15b54690_745 , n150 );
buf ( RI15b55950_785 , n151 );
buf ( RI15b576d8_848 , n152 );
buf ( RI15b57660_847 , n153 );
buf ( RI15b56670_813 , n154 );
buf ( RI15b558d8_784 , n155 );
buf ( RI15b55860_783 , n156 );
buf ( RI15b557e8_782 , n157 );
buf ( RI15b57570_845 , n158 );
buf ( RI15b574f8_844 , n159 );
buf ( RI15b57480_843 , n160 );
buf ( RI15b57408_842 , n161 );
buf ( RI15b57390_841 , n162 );
buf ( RI15b57318_840 , n163 );
buf ( RI15b572a0_839 , n164 );
buf ( RI15b57228_838 , n165 );
buf ( RI15b571b0_837 , n166 );
buf ( RI15b57138_836 , n167 );
buf ( RI15b570c0_835 , n168 );
buf ( RI15b57048_834 , n169 );
buf ( RI15b56fd0_833 , n170 );
buf ( RI15b56f58_832 , n171 );
buf ( RI15b56ee0_831 , n172 );
buf ( RI15b56e68_830 , n173 );
buf ( RI15b56df0_829 , n174 );
buf ( RI15b56d78_828 , n175 );
buf ( RI15b56d00_827 , n176 );
buf ( RI15b56c88_826 , n177 );
buf ( RI15b56c10_825 , n178 );
buf ( RI15b56b98_824 , n179 );
buf ( RI15b56b20_823 , n180 );
buf ( RI15b56aa8_822 , n181 );
buf ( RI15b56a30_821 , n182 );
buf ( RI15b569b8_820 , n183 );
buf ( RI15b56940_819 , n184 );
buf ( RI15b568c8_818 , n185 );
buf ( RI15b567d8_816 , n186 );
buf ( RI15b56760_815 , n187 );
buf ( RI15b566e8_814 , n188 );
buf ( RI15b3ea48_2 , n189 );
buf ( RI15b58740_883 , n190 );
buf ( RI15b5d498_1048 , n191 );
buf ( RI15b586c8_882 , n192 );
buf ( RI15b5d420_1047 , n193 );
buf ( RI15b58650_881 , n194 );
buf ( RI15b5d3a8_1046 , n195 );
buf ( RI15b585d8_880 , n196 );
buf ( RI15b5d330_1045 , n197 );
buf ( RI15b58560_879 , n198 );
buf ( RI15b5d2b8_1044 , n199 );
buf ( RI15b62f10_1241 , n200 );
buf ( RI15b5c778_1020 , n201 );
buf ( RI15b5c700_1019 , n202 );
buf ( RI15b5c688_1018 , n203 );
buf ( RI15b5c610_1017 , n204 );
buf ( RI15b5c598_1016 , n205 );
buf ( RI15b5c520_1015 , n206 );
buf ( RI15b5c4a8_1014 , n207 );
buf ( RI15b5c430_1013 , n208 );
buf ( RI15b5c3b8_1012 , n209 );
buf ( RI15b5c340_1011 , n210 );
buf ( RI15b5bf80_1003 , n211 );
buf ( RI15b5bbc0_995 , n212 );
buf ( RI15b5b800_987 , n213 );
buf ( RI15b5b440_979 , n214 );
buf ( RI15b5b080_971 , n215 );
buf ( RI15b5acc0_963 , n216 );
buf ( RI15b5a900_955 , n217 );
buf ( RI15b5a540_947 , n218 );
buf ( RI15b5a180_939 , n219 );
buf ( RI15b59dc0_931 , n220 );
buf ( RI15b59a00_923 , n221 );
buf ( RI15b59640_915 , n222 );
buf ( RI15b59280_907 , n223 );
buf ( RI15b58ec0_899 , n224 );
buf ( RI15b58b00_891 , n225 );
buf ( RI15b5c2c8_1010 , n226 );
buf ( RI15b5bf08_1002 , n227 );
buf ( RI15b5bb48_994 , n228 );
buf ( RI15b5b788_986 , n229 );
buf ( RI15b5b3c8_978 , n230 );
buf ( RI15b5b008_970 , n231 );
buf ( RI15b5ac48_962 , n232 );
buf ( RI15b5a888_954 , n233 );
buf ( RI15b5a4c8_946 , n234 );
buf ( RI15b5a108_938 , n235 );
buf ( RI15b59d48_930 , n236 );
buf ( RI15b59988_922 , n237 );
buf ( RI15b595c8_914 , n238 );
buf ( RI15b59208_906 , n239 );
buf ( RI15b58e48_898 , n240 );
buf ( RI15b58a88_890 , n241 );
buf ( RI15b5c250_1009 , n242 );
buf ( RI15b5be90_1001 , n243 );
buf ( RI15b5bad0_993 , n244 );
buf ( RI15b5b710_985 , n245 );
buf ( RI15b5b350_977 , n246 );
buf ( RI15b5af90_969 , n247 );
buf ( RI15b5abd0_961 , n248 );
buf ( RI15b5a810_953 , n249 );
buf ( RI15b5a450_945 , n250 );
buf ( RI15b5a090_937 , n251 );
buf ( RI15b59cd0_929 , n252 );
buf ( RI15b59910_921 , n253 );
buf ( RI15b59550_913 , n254 );
buf ( RI15b59190_905 , n255 );
buf ( RI15b58dd0_897 , n256 );
buf ( RI15b58a10_889 , n257 );
buf ( RI15b5c1d8_1008 , n258 );
buf ( RI15b5be18_1000 , n259 );
buf ( RI15b5ba58_992 , n260 );
buf ( RI15b5b698_984 , n261 );
buf ( RI15b5b2d8_976 , n262 );
buf ( RI15b5af18_968 , n263 );
buf ( RI15b5ab58_960 , n264 );
buf ( RI15b5a798_952 , n265 );
buf ( RI15b5a3d8_944 , n266 );
buf ( RI15b5a018_936 , n267 );
buf ( RI15b59c58_928 , n268 );
buf ( RI15b59898_920 , n269 );
buf ( RI15b594d8_912 , n270 );
buf ( RI15b59118_904 , n271 );
buf ( RI15b58d58_896 , n272 );
buf ( RI15b58998_888 , n273 );
buf ( RI15b5c160_1007 , n274 );
buf ( RI15b5bda0_999 , n275 );
buf ( RI15b5b9e0_991 , n276 );
buf ( RI15b5b620_983 , n277 );
buf ( RI15b5b260_975 , n278 );
buf ( RI15b5aea0_967 , n279 );
buf ( RI15b5aae0_959 , n280 );
buf ( RI15b5a720_951 , n281 );
buf ( RI15b5a360_943 , n282 );
buf ( RI15b59fa0_935 , n283 );
buf ( RI15b59be0_927 , n284 );
buf ( RI15b59820_919 , n285 );
buf ( RI15b59460_911 , n286 );
buf ( RI15b590a0_903 , n287 );
buf ( RI15b58ce0_895 , n288 );
buf ( RI15b58920_887 , n289 );
buf ( RI15b5c0e8_1006 , n290 );
buf ( RI15b5bd28_998 , n291 );
buf ( RI15b5b968_990 , n292 );
buf ( RI15b5b5a8_982 , n293 );
buf ( RI15b5b1e8_974 , n294 );
buf ( RI15b5ae28_966 , n295 );
buf ( RI15b5aa68_958 , n296 );
buf ( RI15b5a6a8_950 , n297 );
buf ( RI15b5a2e8_942 , n298 );
buf ( RI15b59f28_934 , n299 );
buf ( RI15b59b68_926 , n300 );
buf ( RI15b597a8_918 , n301 );
buf ( RI15b593e8_910 , n302 );
buf ( RI15b59028_902 , n303 );
buf ( RI15b58c68_894 , n304 );
buf ( RI15b588a8_886 , n305 );
buf ( RI15b5c070_1005 , n306 );
buf ( RI15b5bcb0_997 , n307 );
buf ( RI15b5b8f0_989 , n308 );
buf ( RI15b5b530_981 , n309 );
buf ( RI15b5b170_973 , n310 );
buf ( RI15b5adb0_965 , n311 );
buf ( RI15b5a9f0_957 , n312 );
buf ( RI15b5a630_949 , n313 );
buf ( RI15b5a270_941 , n314 );
buf ( RI15b59eb0_933 , n315 );
buf ( RI15b59af0_925 , n316 );
buf ( RI15b59730_917 , n317 );
buf ( RI15b59370_909 , n318 );
buf ( RI15b58fb0_901 , n319 );
buf ( RI15b58bf0_893 , n320 );
buf ( RI15b58830_885 , n321 );
buf ( RI15b5bff8_1004 , n322 );
buf ( RI15b5bc38_996 , n323 );
buf ( RI15b5b878_988 , n324 );
buf ( RI15b5b4b8_980 , n325 );
buf ( RI15b5b0f8_972 , n326 );
buf ( RI15b5ad38_964 , n327 );
buf ( RI15b5a978_956 , n328 );
buf ( RI15b5a5b8_948 , n329 );
buf ( RI15b5a1f8_940 , n330 );
buf ( RI15b59e38_932 , n331 );
buf ( RI15b59a78_924 , n332 );
buf ( RI15b596b8_916 , n333 );
buf ( RI15b592f8_908 , n334 );
buf ( RI15b58f38_900 , n335 );
buf ( RI15b58b78_892 , n336 );
buf ( RI15b587b8_884 , n337 );
buf ( RI15b5d588_1050 , n338 );
buf ( RI15b5d6f0_1053 , n339 );
buf ( RI15b5d600_1051 , n340 );
buf ( RI15b5d678_1052 , n341 );
buf ( RI15b62e98_1240 , n342 );
buf ( RI15b62e20_1239 , n343 );
buf ( RI15b62da8_1238 , n344 );
buf ( RI15b62d30_1237 , n345 );
buf ( RI15b62cb8_1236 , n346 );
buf ( RI15b62c40_1235 , n347 );
buf ( RI15b62bc8_1234 , n348 );
buf ( RI15b606c0_1155 , n349 );
buf ( RI15b63e10_1273 , n350 );
buf ( RI15b4b090_425 , n351 );
buf ( RI15b44cb8_212 , n352 );
buf ( RI15b44e20_215 , n353 );
buf ( RI15b44d30_213 , n354 );
buf ( RI15b44da8_214 , n355 );
buf ( RI15b3fe70_45 , n356 );
buf ( RI15b44bc8_210 , n357 );
buf ( RI15b3fdf8_44 , n358 );
buf ( RI15b44b50_209 , n359 );
buf ( RI15b3fd80_43 , n360 );
buf ( RI15b44ad8_208 , n361 );
buf ( RI15b3fd08_42 , n362 );
buf ( RI15b44a60_207 , n363 );
buf ( RI15b3fc90_41 , n364 );
buf ( RI15b449e8_206 , n365 );
buf ( RI15b4bf90_457 , n366 );
buf ( RI15b43728_166 , n367 );
buf ( RI15b43368_158 , n368 );
buf ( RI15b42fa8_150 , n369 );
buf ( RI15b42be8_142 , n370 );
buf ( RI15b42828_134 , n371 );
buf ( RI15b42468_126 , n372 );
buf ( RI15b420a8_118 , n373 );
buf ( RI15b41ce8_110 , n374 );
buf ( RI15b41928_102 , n375 );
buf ( RI15b41568_94 , n376 );
buf ( RI15b411a8_86 , n377 );
buf ( RI15b40de8_78 , n378 );
buf ( RI15b40a28_70 , n379 );
buf ( RI15b40668_62 , n380 );
buf ( RI15b402a8_54 , n381 );
buf ( RI15b3fee8_46 , n382 );
buf ( RI15b437a0_167 , n383 );
buf ( RI15b433e0_159 , n384 );
buf ( RI15b43020_151 , n385 );
buf ( RI15b42c60_143 , n386 );
buf ( RI15b428a0_135 , n387 );
buf ( RI15b424e0_127 , n388 );
buf ( RI15b42120_119 , n389 );
buf ( RI15b41d60_111 , n390 );
buf ( RI15b419a0_103 , n391 );
buf ( RI15b415e0_95 , n392 );
buf ( RI15b41220_87 , n393 );
buf ( RI15b40e60_79 , n394 );
buf ( RI15b40aa0_71 , n395 );
buf ( RI15b406e0_63 , n396 );
buf ( RI15b40320_55 , n397 );
buf ( RI15b3ff60_47 , n398 );
buf ( RI15b43818_168 , n399 );
buf ( RI15b43458_160 , n400 );
buf ( RI15b43098_152 , n401 );
buf ( RI15b42cd8_144 , n402 );
buf ( RI15b42918_136 , n403 );
buf ( RI15b42558_128 , n404 );
buf ( RI15b42198_120 , n405 );
buf ( RI15b41dd8_112 , n406 );
buf ( RI15b41a18_104 , n407 );
buf ( RI15b41658_96 , n408 );
buf ( RI15b41298_88 , n409 );
buf ( RI15b40ed8_80 , n410 );
buf ( RI15b40b18_72 , n411 );
buf ( RI15b40758_64 , n412 );
buf ( RI15b40398_56 , n413 );
buf ( RI15b3ffd8_48 , n414 );
buf ( RI15b43890_169 , n415 );
buf ( RI15b434d0_161 , n416 );
buf ( RI15b43110_153 , n417 );
buf ( RI15b42d50_145 , n418 );
buf ( RI15b42990_137 , n419 );
buf ( RI15b425d0_129 , n420 );
buf ( RI15b42210_121 , n421 );
buf ( RI15b41e50_113 , n422 );
buf ( RI15b41a90_105 , n423 );
buf ( RI15b416d0_97 , n424 );
buf ( RI15b41310_89 , n425 );
buf ( RI15b40f50_81 , n426 );
buf ( RI15b40b90_73 , n427 );
buf ( RI15b407d0_65 , n428 );
buf ( RI15b40410_57 , n429 );
buf ( RI15b40050_49 , n430 );
buf ( RI15b43908_170 , n431 );
buf ( RI15b43548_162 , n432 );
buf ( RI15b43188_154 , n433 );
buf ( RI15b42dc8_146 , n434 );
buf ( RI15b42a08_138 , n435 );
buf ( RI15b42648_130 , n436 );
buf ( RI15b42288_122 , n437 );
buf ( RI15b41ec8_114 , n438 );
buf ( RI15b41b08_106 , n439 );
buf ( RI15b41748_98 , n440 );
buf ( RI15b41388_90 , n441 );
buf ( RI15b40fc8_82 , n442 );
buf ( RI15b40c08_74 , n443 );
buf ( RI15b40848_66 , n444 );
buf ( RI15b40488_58 , n445 );
buf ( RI15b400c8_50 , n446 );
buf ( RI15b43980_171 , n447 );
buf ( RI15b435c0_163 , n448 );
buf ( RI15b43200_155 , n449 );
buf ( RI15b42e40_147 , n450 );
buf ( RI15b42a80_139 , n451 );
buf ( RI15b426c0_131 , n452 );
buf ( RI15b42300_123 , n453 );
buf ( RI15b41f40_115 , n454 );
buf ( RI15b41b80_107 , n455 );
buf ( RI15b417c0_99 , n456 );
buf ( RI15b41400_91 , n457 );
buf ( RI15b41040_83 , n458 );
buf ( RI15b40c80_75 , n459 );
buf ( RI15b408c0_67 , n460 );
buf ( RI15b40500_59 , n461 );
buf ( RI15b40140_51 , n462 );
buf ( RI15b439f8_172 , n463 );
buf ( RI15b43638_164 , n464 );
buf ( RI15b43278_156 , n465 );
buf ( RI15b42eb8_148 , n466 );
buf ( RI15b42af8_140 , n467 );
buf ( RI15b42738_132 , n468 );
buf ( RI15b42378_124 , n469 );
buf ( RI15b41fb8_116 , n470 );
buf ( RI15b41bf8_108 , n471 );
buf ( RI15b41838_100 , n472 );
buf ( RI15b41478_92 , n473 );
buf ( RI15b410b8_84 , n474 );
buf ( RI15b40cf8_76 , n475 );
buf ( RI15b40938_68 , n476 );
buf ( RI15b40578_60 , n477 );
buf ( RI15b401b8_52 , n478 );
buf ( RI15b43a70_173 , n479 );
buf ( RI15b436b0_165 , n480 );
buf ( RI15b432f0_157 , n481 );
buf ( RI15b42f30_149 , n482 );
buf ( RI15b42b70_141 , n483 );
buf ( RI15b427b0_133 , n484 );
buf ( RI15b423f0_125 , n485 );
buf ( RI15b42030_117 , n486 );
buf ( RI15b41c70_109 , n487 );
buf ( RI15b418b0_101 , n488 );
buf ( RI15b414f0_93 , n489 );
buf ( RI15b41130_85 , n490 );
buf ( RI15b40d70_77 , n491 );
buf ( RI15b409b0_69 , n492 );
buf ( RI15b405f0_61 , n493 );
buf ( RI15b40230_53 , n494 );
buf ( RI15b48318_328 , n495 );
buf ( RI15b48390_329 , n496 );
buf ( RI15b48408_330 , n497 );
buf ( RI15b668b8_1364 , n498 );
buf ( RI15b3fba0_39 , n499 );
buf ( RI15b47df0_317 , n500 );
buf ( RI15b4a190_393 , n501 );
buf ( RI15b4bf18_456 , n502 );
buf ( RI15b4bea0_455 , n503 );
buf ( RI15b4be28_454 , n504 );
buf ( RI15b4bdb0_453 , n505 );
buf ( RI15b4bd38_452 , n506 );
buf ( RI15b4bcc0_451 , n507 );
buf ( RI15b4bc48_450 , n508 );
buf ( RI15b4bbd0_449 , n509 );
buf ( RI15b4bb58_448 , n510 );
buf ( RI15b4bae0_447 , n511 );
buf ( RI15b4ba68_446 , n512 );
buf ( RI15b4b9f0_445 , n513 );
buf ( RI15b4b978_444 , n514 );
buf ( RI15b4b900_443 , n515 );
buf ( RI15b4b888_442 , n516 );
buf ( RI15b4b810_441 , n517 );
buf ( RI15b4b798_440 , n518 );
buf ( RI15b4b720_439 , n519 );
buf ( RI15b4b6a8_438 , n520 );
buf ( RI15b4b630_437 , n521 );
buf ( RI15b4b5b8_436 , n522 );
buf ( RI15b4b540_435 , n523 );
buf ( RI15b4b4c8_434 , n524 );
buf ( RI15b4b450_433 , n525 );
buf ( RI15b4b3d8_432 , n526 );
buf ( RI15b4b360_431 , n527 );
buf ( RI15b4b2e8_430 , n528 );
buf ( RI15b4b270_429 , n529 );
buf ( RI15b4b1f8_428 , n530 );
buf ( RI15b4a208_394 , n531 );
buf ( RI15b4a118_392 , n532 );
buf ( RI15b4a0a0_391 , n533 );
buf ( RI15b4a028_390 , n534 );
buf ( RI15b49fb0_389 , n535 );
buf ( RI15b49f38_388 , n536 );
buf ( RI15b49ec0_387 , n537 );
buf ( RI15b49e48_386 , n538 );
buf ( RI15b49dd0_385 , n539 );
buf ( RI15b49d58_384 , n540 );
buf ( RI15b49ce0_383 , n541 );
buf ( RI15b49c68_382 , n542 );
buf ( RI15b49bf0_381 , n543 );
buf ( RI15b49b78_380 , n544 );
buf ( RI15b49b00_379 , n545 );
buf ( RI15b49a88_378 , n546 );
buf ( RI15b49a10_377 , n547 );
buf ( RI15b49998_376 , n548 );
buf ( RI15b49920_375 , n549 );
buf ( RI15b498a8_374 , n550 );
buf ( RI15b49830_373 , n551 );
buf ( RI15b497b8_372 , n552 );
buf ( RI15b49740_371 , n553 );
buf ( RI15b496c8_370 , n554 );
buf ( RI15b49650_369 , n555 );
buf ( RI15b495d8_368 , n556 );
buf ( RI15b49560_367 , n557 );
buf ( RI15b494e8_366 , n558 );
buf ( RI15b49470_365 , n559 );
buf ( RI15b493f8_364 , n560 );
buf ( RI15b49380_363 , n561 );
buf ( RI15b4b108_426 , n562 );
buf ( RI15b4b018_424 , n563 );
buf ( RI15b4afa0_423 , n564 );
buf ( RI15b4af28_422 , n565 );
buf ( RI15b4aeb0_421 , n566 );
buf ( RI15b4ae38_420 , n567 );
buf ( RI15b4adc0_419 , n568 );
buf ( RI15b4ad48_418 , n569 );
buf ( RI15b4acd0_417 , n570 );
buf ( RI15b4ac58_416 , n571 );
buf ( RI15b4abe0_415 , n572 );
buf ( RI15b4ab68_414 , n573 );
buf ( RI15b4aaf0_413 , n574 );
buf ( RI15b4aa78_412 , n575 );
buf ( RI15b4aa00_411 , n576 );
buf ( RI15b4a988_410 , n577 );
buf ( RI15b4a910_409 , n578 );
buf ( RI15b4a898_408 , n579 );
buf ( RI15b4a820_407 , n580 );
buf ( RI15b4a7a8_406 , n581 );
buf ( RI15b4a730_405 , n582 );
buf ( RI15b4a6b8_404 , n583 );
buf ( RI15b4a640_403 , n584 );
buf ( RI15b4a5c8_402 , n585 );
buf ( RI15b4a550_401 , n586 );
buf ( RI15b4a4d8_400 , n587 );
buf ( RI15b4a460_399 , n588 );
buf ( RI15b4a3e8_398 , n589 );
buf ( RI15b4a370_397 , n590 );
buf ( RI15b4a2f8_396 , n591 );
buf ( RI15b4a280_395 , n592 );
buf ( RI15b50928_614 , n593 );
buf ( RI15b508b0_613 , n594 );
buf ( RI15b50838_612 , n595 );
buf ( RI15b507c0_611 , n596 );
buf ( RI15b50748_610 , n597 );
buf ( RI15b506d0_609 , n598 );
buf ( RI15b50658_608 , n599 );
buf ( RI15b505e0_607 , n600 );
buf ( RI15b50568_606 , n601 );
buf ( RI15b504f0_605 , n602 );
buf ( RI15b50478_604 , n603 );
buf ( RI15b50400_603 , n604 );
buf ( RI15b50388_602 , n605 );
buf ( RI15b50310_601 , n606 );
buf ( RI15b50298_600 , n607 );
buf ( RI15b50220_599 , n608 );
buf ( RI15b501a8_598 , n609 );
buf ( RI15b50130_597 , n610 );
buf ( RI15b500b8_596 , n611 );
buf ( RI15b50040_595 , n612 );
buf ( RI15b4ffc8_594 , n613 );
buf ( RI15b4ff50_593 , n614 );
buf ( RI15b57fc0_867 , n615 );
buf ( RI15b57de0_863 , n616 );
buf ( RI15b55fe0_799 , n617 );
buf ( RI15b57d68_862 , n618 );
buf ( RI15b57cf0_861 , n619 );
buf ( RI15b57c78_860 , n620 );
buf ( RI15b57c00_859 , n621 );
buf ( RI15b57b88_858 , n622 );
buf ( RI15b57b10_857 , n623 );
buf ( RI15b57a98_856 , n624 );
buf ( RI15b57a20_855 , n625 );
buf ( RI15b579a8_854 , n626 );
buf ( RI15b57930_853 , n627 );
buf ( RI15b578b8_852 , n628 );
buf ( RI15b57840_851 , n629 );
buf ( RI15b577c8_850 , n630 );
buf ( RI15b55f68_798 , n631 );
buf ( RI15b55ef0_797 , n632 );
buf ( RI15b55e78_796 , n633 );
buf ( RI15b55e00_795 , n634 );
buf ( RI15b55d88_794 , n635 );
buf ( RI15b55d10_793 , n636 );
buf ( RI15b55c98_792 , n637 );
buf ( RI15b55c20_791 , n638 );
buf ( RI15b55ba8_790 , n639 );
buf ( RI15b55b30_789 , n640 );
buf ( RI15b55ab8_788 , n641 );
buf ( RI15b55a40_787 , n642 );
buf ( RI15b559c8_786 , n643 );
buf ( RI15b65850_1329 , n644 );
buf ( RI15b666d8_1360 , n645 );
buf ( RI15b658c8_1330 , n646 );
buf ( RI15b65940_1331 , n647 );
buf ( RI15b659b8_1332 , n648 );
buf ( RI15b65a30_1333 , n649 );
buf ( RI15b65aa8_1334 , n650 );
buf ( RI15b65b20_1335 , n651 );
buf ( RI15b65b98_1336 , n652 );
buf ( RI15b65fd0_1345 , n653 );
buf ( RI15b65f58_1344 , n654 );
buf ( RI15b65ee0_1343 , n655 );
buf ( RI15b65e68_1342 , n656 );
buf ( RI15b65df0_1341 , n657 );
buf ( RI15b65d78_1340 , n658 );
buf ( RI15b65d00_1339 , n659 );
buf ( RI15b65c88_1338 , n660 );
buf ( RI15b65c10_1337 , n661 );
buf ( RI15b66660_1359 , n662 );
buf ( RI15b665e8_1358 , n663 );
buf ( RI15b66570_1357 , n664 );
buf ( RI15b664f8_1356 , n665 );
buf ( RI15b66480_1355 , n666 );
buf ( RI15b66408_1354 , n667 );
buf ( RI15b66390_1353 , n668 );
buf ( RI15b66318_1352 , n669 );
buf ( RI15b662a0_1351 , n670 );
buf ( RI15b66228_1350 , n671 );
buf ( RI15b661b0_1349 , n672 );
buf ( RI15b66138_1348 , n673 );
buf ( RI15b660c0_1347 , n674 );
buf ( RI15b66048_1346 , n675 );
buf ( RI15b62b50_1233 , n676 );
buf ( RI15b63a50_1265 , n677 );
buf ( RI15b60be8_1166 , n678 );
buf ( RI15b60c60_1167 , n679 );
buf ( RI15b60cd8_1168 , n680 );
buf ( RI15b66750_1361 , n681 );
buf ( RI15b3fb28_38 , n682 );
buf ( RI15b61c50_1201 , n683 );
buf ( RI15b58470_877 , n684 );
buf ( RI15b583f8_876 , n685 );
buf ( RI15b58380_875 , n686 );
buf ( RI15b58308_874 , n687 );
buf ( RI15b58290_873 , n688 );
buf ( RI15b58218_872 , n689 );
buf ( RI15b581a0_871 , n690 );
buf ( RI15b58128_870 , n691 );
buf ( RI15b580b0_869 , n692 );
buf ( RI15b58038_868 , n693 );
buf ( RI15b57f48_866 , n694 );
buf ( RI15b57ed0_865 , n695 );
buf ( RI15b57e58_864 , n696 );
buf ( RI15b565f8_812 , n697 );
buf ( RI15b56580_811 , n698 );
buf ( RI15b56508_810 , n699 );
buf ( RI15b56490_809 , n700 );
buf ( RI15b56418_808 , n701 );
buf ( RI15b563a0_807 , n702 );
buf ( RI15b56328_806 , n703 );
buf ( RI15b562b0_805 , n704 );
buf ( RI15b56238_804 , n705 );
buf ( RI15b561c0_803 , n706 );
buf ( RI15b56148_802 , n707 );
buf ( RI15b560d0_801 , n708 );
buf ( RI15b56058_800 , n709 );
buf ( RI15b605d0_1153 , n710 );
buf ( RI15b60648_1154 , n711 );
buf ( RI15b54168_734 , n712 );
buf ( RI15b541e0_735 , n713 );
buf ( RI15b47d00_315 , n714 );
buf ( RI15b47d78_316 , n715 );
buf ( RI15b51558_640 , n716 );
buf ( RI15b450f0_221 , n717 );
buf ( RI15b4c008_458 , n718 );
buf ( RI15b63d98_1272 , n719 );
buf ( RI15b575e8_846 , n720 );
buf ( RI15b648d8_1296 , n721 );
buf ( RI15b63ac8_1266 , n722 );
buf ( RI15b64860_1295 , n723 );
buf ( RI15b647e8_1294 , n724 );
buf ( RI15b64770_1293 , n725 );
buf ( RI15b646f8_1292 , n726 );
buf ( RI15b64680_1291 , n727 );
buf ( RI15b64608_1290 , n728 );
buf ( RI15b64590_1289 , n729 );
buf ( RI15b64518_1288 , n730 );
buf ( RI15b644a0_1287 , n731 );
buf ( RI15b64428_1286 , n732 );
buf ( RI15b643b0_1285 , n733 );
buf ( RI15b64338_1284 , n734 );
buf ( RI15b642c0_1283 , n735 );
buf ( RI15b64248_1282 , n736 );
buf ( RI15b641d0_1281 , n737 );
buf ( RI15b64158_1280 , n738 );
buf ( RI15b640e0_1279 , n739 );
buf ( RI15b64068_1278 , n740 );
buf ( RI15b63ff0_1277 , n741 );
buf ( RI15b63f78_1276 , n742 );
buf ( RI15b63f00_1275 , n743 );
buf ( RI15b63e88_1274 , n744 );
buf ( RI15b63d20_1271 , n745 );
buf ( RI15b63ca8_1270 , n746 );
buf ( RI15b63c30_1269 , n747 );
buf ( RI15b63bb8_1268 , n748 );
buf ( RI15b63b40_1267 , n749 );
buf ( RI15b5d948_1058 , n750 );
buf ( RI15b467e8_270 , n751 );
buf ( RI15b48480_331 , n752 );
buf ( RI15b49308_362 , n753 );
buf ( RI15b484f8_332 , n754 );
buf ( RI15b48570_333 , n755 );
buf ( RI15b485e8_334 , n756 );
buf ( RI15b48660_335 , n757 );
buf ( RI15b486d8_336 , n758 );
buf ( RI15b48750_337 , n759 );
buf ( RI15b487c8_338 , n760 );
buf ( RI15b48840_339 , n761 );
buf ( RI15b488b8_340 , n762 );
buf ( RI15b48930_341 , n763 );
buf ( RI15b489a8_342 , n764 );
buf ( RI15b48a20_343 , n765 );
buf ( RI15b48a98_344 , n766 );
buf ( RI15b48b10_345 , n767 );
buf ( RI15b48b88_346 , n768 );
buf ( RI15b5e5f0_1085 , n769 );
buf ( RI15b5e6e0_1087 , n770 );
buf ( RI15b5d9c0_1059 , n771 );
buf ( RI15b5da38_1060 , n772 );
buf ( RI15b5dab0_1061 , n773 );
buf ( RI15b5db28_1062 , n774 );
buf ( RI15b5dba0_1063 , n775 );
buf ( RI15b5dc18_1064 , n776 );
buf ( RI15b5dc90_1065 , n777 );
buf ( RI15b5dd08_1066 , n778 );
buf ( RI15b5dd80_1067 , n779 );
buf ( RI15b5ddf8_1068 , n780 );
buf ( RI15b5de70_1069 , n781 );
buf ( RI15b5dee8_1070 , n782 );
buf ( RI15b5df60_1071 , n783 );
buf ( RI15b5dfd8_1072 , n784 );
buf ( RI15b5e050_1073 , n785 );
buf ( RI15b5e0c8_1074 , n786 );
buf ( RI15b5e140_1075 , n787 );
buf ( RI15b5e1b8_1076 , n788 );
buf ( RI15b5e230_1077 , n789 );
buf ( RI15b5e2a8_1078 , n790 );
buf ( RI15b5e320_1079 , n791 );
buf ( RI15b5e398_1080 , n792 );
buf ( RI15b5e410_1081 , n793 );
buf ( RI15b5e488_1082 , n794 );
buf ( RI15b5e500_1083 , n795 );
buf ( RI15b5e578_1084 , n796 );
buf ( RI15b5e668_1086 , n797 );
buf ( RI15b3f948_34 , n798 );
buf ( RI15b64950_1297 , n799 );
buf ( RI15b3eac0_3 , n800 );
buf ( RI15b657d8_1328 , n801 );
buf ( RI15b3f8d0_33 , n802 );
buf ( RI15b649c8_1298 , n803 );
buf ( RI15b3f858_32 , n804 );
buf ( RI15b64a40_1299 , n805 );
buf ( RI15b3f7e0_31 , n806 );
buf ( RI15b64ab8_1300 , n807 );
buf ( RI15b3f768_30 , n808 );
buf ( RI15b64b30_1301 , n809 );
buf ( RI15b3f6f0_29 , n810 );
buf ( RI15b64ba8_1302 , n811 );
buf ( RI15b3f678_28 , n812 );
buf ( RI15b64c20_1303 , n813 );
buf ( RI15b3f600_27 , n814 );
buf ( RI15b64c98_1304 , n815 );
buf ( RI15b3f1c8_18 , n816 );
buf ( RI15b650d0_1313 , n817 );
buf ( RI15b3f240_19 , n818 );
buf ( RI15b65058_1312 , n819 );
buf ( RI15b3f2b8_20 , n820 );
buf ( RI15b64fe0_1311 , n821 );
buf ( RI15b3f330_21 , n822 );
buf ( RI15b64f68_1310 , n823 );
buf ( RI15b3f3a8_22 , n824 );
buf ( RI15b64ef0_1309 , n825 );
buf ( RI15b3f420_23 , n826 );
buf ( RI15b64e78_1308 , n827 );
buf ( RI15b3f498_24 , n828 );
buf ( RI15b64e00_1307 , n829 );
buf ( RI15b3f510_25 , n830 );
buf ( RI15b64d88_1306 , n831 );
buf ( RI15b3f588_26 , n832 );
buf ( RI15b64d10_1305 , n833 );
buf ( RI15b3eb38_4 , n834 );
buf ( RI15b65760_1327 , n835 );
buf ( RI15b3ebb0_5 , n836 );
buf ( RI15b656e8_1326 , n837 );
buf ( RI15b3ec28_6 , n838 );
buf ( RI15b65670_1325 , n839 );
buf ( RI15b3eca0_7 , n840 );
buf ( RI15b655f8_1324 , n841 );
buf ( RI15b3ed18_8 , n842 );
buf ( RI15b65580_1323 , n843 );
buf ( RI15b3ed90_9 , n844 );
buf ( RI15b65508_1322 , n845 );
buf ( RI15b3ee08_10 , n846 );
buf ( RI15b65490_1321 , n847 );
buf ( RI15b3ee80_11 , n848 );
buf ( RI15b65418_1320 , n849 );
buf ( RI15b3eef8_12 , n850 );
buf ( RI15b653a0_1319 , n851 );
buf ( RI15b3ef70_13 , n852 );
buf ( RI15b65328_1318 , n853 );
buf ( RI15b3efe8_14 , n854 );
buf ( RI15b652b0_1317 , n855 );
buf ( RI15b3f060_15 , n856 );
buf ( RI15b65238_1316 , n857 );
buf ( RI15b3f0d8_16 , n858 );
buf ( RI15b651c0_1315 , n859 );
buf ( RI15b3f150_17 , n860 );
buf ( RI15b65148_1314 , n861 );
buf ( RI15b62f88_1242 , n862 );
buf ( RI15b5c7f0_1021 , n863 );
buf ( RI15b479b8_308 , n864 );
buf ( RI15b47b98_312 , n865 );
buf ( RI15b52278_668 , n866 );
buf ( RI15b52458_672 , n867 );
buf ( RI15b523e0_671 , n868 );
buf ( RI15b52368_670 , n869 );
buf ( RI15b522f0_669 , n870 );
buf ( RI15b51300_635 , n871 );
buf ( RI15b51378_636 , n872 );
buf ( RI15b513f0_637 , n873 );
buf ( RI15b51468_638 , n874 );
buf ( RI15b534c0_707 , n875 );
buf ( RI15b52f98_696 , n876 );
buf ( RI15b548e8_750 , n877 );
buf ( RI15b55770_781 , n878 );
buf ( RI15b54960_751 , n879 );
buf ( RI15b549d8_752 , n880 );
buf ( RI15b54a50_753 , n881 );
buf ( RI15b54ac8_754 , n882 );
buf ( RI15b54b40_755 , n883 );
buf ( RI15b54bb8_756 , n884 );
buf ( RI15b54c30_757 , n885 );
buf ( RI15b54ca8_758 , n886 );
buf ( RI15b54d20_759 , n887 );
buf ( RI15b54d98_760 , n888 );
buf ( RI15b54e10_761 , n889 );
buf ( RI15b54e88_762 , n890 );
buf ( RI15b54f00_763 , n891 );
buf ( RI15b54f78_764 , n892 );
buf ( RI15b54ff0_765 , n893 );
buf ( RI15b514e0_639 , n894 );
buf ( RI15b515d0_641 , n895 );
buf ( RI15b51648_642 , n896 );
buf ( RI15b516c0_643 , n897 );
buf ( RI15b51738_644 , n898 );
buf ( RI15b517b0_645 , n899 );
buf ( RI15b51828_646 , n900 );
buf ( RI15b518a0_647 , n901 );
buf ( RI15b51918_648 , n902 );
buf ( RI15b51990_649 , n903 );
buf ( RI15b51a08_650 , n904 );
buf ( RI15b51a80_651 , n905 );
buf ( RI15b51af8_652 , n906 );
buf ( RI15b51b70_653 , n907 );
buf ( RI15b51be8_654 , n908 );
buf ( RI15b51c60_655 , n909 );
buf ( RI15b51cd8_656 , n910 );
buf ( RI15b51d50_657 , n911 );
buf ( RI15b51dc8_658 , n912 );
buf ( RI15b51e40_659 , n913 );
buf ( RI15b51eb8_660 , n914 );
buf ( RI15b51f30_661 , n915 );
buf ( RI15b51fa8_662 , n916 );
buf ( RI15b52020_663 , n917 );
buf ( RI15b52098_664 , n918 );
buf ( RI15b52110_665 , n919 );
buf ( RI15b52188_666 , n920 );
buf ( RI15b52200_667 , n921 );
buf ( RI15b50b08_618 , n922 );
buf ( RI15b50a90_617 , n923 );
buf ( RI15b50a18_616 , n924 );
buf ( RI15b509a0_615 , n925 );
buf ( RI15b46e00_283 , n926 );
buf ( RI15b4b180_427 , n927 );
buf ( RI15b48228_326 , n928 );
buf ( RI15b482a0_327 , n929 );
buf ( RI15b45348_226 , n930 );
buf ( RI15b4c080_459 , n931 );
buf ( RI15b55680_779 , n932 );
buf ( RI15b55608_778 , n933 );
buf ( RI15b55590_777 , n934 );
buf ( RI15b55518_776 , n935 );
buf ( RI15b554a0_775 , n936 );
buf ( RI15b55428_774 , n937 );
buf ( RI15b553b0_773 , n938 );
buf ( RI15b55338_772 , n939 );
buf ( RI15b552c0_771 , n940 );
buf ( RI15b55248_770 , n941 );
buf ( RI15b551d0_769 , n942 );
buf ( RI15b55158_768 , n943 );
buf ( RI15b550e0_767 , n944 );
buf ( RI15b55068_766 , n945 );
buf ( RI15b52908_682 , n946 );
buf ( RI15b53f10_729 , n947 );
buf ( RI15b556f8_780 , n948 );
buf ( RI15b52b60_687 , n949 );
buf ( RI15b61d40_1203 , n950 );
buf ( RI15b62ad8_1232 , n951 );
buf ( RI15b61cc8_1202 , n952 );
buf ( RI15b639d8_1264 , n953 );
buf ( RI15b63960_1263 , n954 );
buf ( RI15b638e8_1262 , n955 );
buf ( RI15b63870_1261 , n956 );
buf ( RI15b637f8_1260 , n957 );
buf ( RI15b63780_1259 , n958 );
buf ( RI15b63708_1258 , n959 );
buf ( RI15b63690_1257 , n960 );
buf ( RI15b63618_1256 , n961 );
buf ( RI15b635a0_1255 , n962 );
buf ( RI15b63528_1254 , n963 );
buf ( RI15b634b0_1253 , n964 );
buf ( RI15b63438_1252 , n965 );
buf ( RI15b633c0_1251 , n966 );
buf ( RI15b63348_1250 , n967 );
buf ( RI15b632d0_1249 , n968 );
buf ( RI15b63258_1248 , n969 );
buf ( RI15b631e0_1247 , n970 );
buf ( RI15b63168_1246 , n971 );
buf ( RI15b630f0_1245 , n972 );
buf ( RI15b63078_1244 , n973 );
buf ( RI15b63000_1243 , n974 );
buf ( RI15b5f658_1120 , n975 );
buf ( RI15b5fdd8_1136 , n976 );
buf ( RI15b60d50_1169 , n977 );
buf ( RI15b61bd8_1200 , n978 );
buf ( RI15b60dc8_1170 , n979 );
buf ( RI15b60e40_1171 , n980 );
buf ( RI15b60eb8_1172 , n981 );
buf ( RI15b60f30_1173 , n982 );
buf ( RI15b60fa8_1174 , n983 );
buf ( RI15b61020_1175 , n984 );
buf ( RI15b61098_1176 , n985 );
buf ( RI15b61110_1177 , n986 );
buf ( RI15b61188_1178 , n987 );
buf ( RI15b61200_1179 , n988 );
buf ( RI15b61278_1180 , n989 );
buf ( RI15b612f0_1181 , n990 );
buf ( RI15b61368_1182 , n991 );
buf ( RI15b613e0_1183 , n992 );
buf ( RI15b61458_1184 , n993 );
buf ( RI15b62100_1211 , n994 );
buf ( RI15b62088_1210 , n995 );
buf ( RI15b62010_1209 , n996 );
buf ( RI15b61f98_1208 , n997 );
buf ( RI15b61f20_1207 , n998 );
buf ( RI15b61ea8_1206 , n999 );
buf ( RI15b61e30_1205 , n1000 );
buf ( RI15b61db8_1204 , n1001 );
buf ( RI15b45438_228 , n1002 );
buf ( RI15b477d8_304 , n1003 );
buf ( RI15b5cf70_1037 , n1004 );
buf ( RI15b5cef8_1036 , n1005 );
buf ( RI15b5ce80_1035 , n1006 );
buf ( RI15b5ce08_1034 , n1007 );
buf ( RI15b5cd90_1033 , n1008 );
buf ( RI15b5cd18_1032 , n1009 );
buf ( RI15b5cca0_1031 , n1010 );
buf ( RI15b5cc28_1030 , n1011 );
buf ( RI15b5cbb0_1029 , n1012 );
buf ( RI15b5cb38_1028 , n1013 );
buf ( RI15b5cac0_1027 , n1014 );
buf ( RI15b5ca48_1026 , n1015 );
buf ( RI15b5c9d0_1025 , n1016 );
buf ( RI15b5c958_1024 , n1017 );
buf ( RI15b5c8e0_1023 , n1018 );
buf ( RI15b5c868_1022 , n1019 );
buf ( RI15b5f388_1114 , n1020 );
buf ( RI15b60738_1156 , n1021 );
buf ( RI15b3f9c0_35 , n1022 );
buf ( RI15b3fa38_36 , n1023 );
buf ( RI15b60828_1158 , n1024 );
buf ( RI15b5e848_1090 , n1025 );
buf ( RI15b46950_273 , n1026 );
buf ( RI15b470d0_289 , n1027 );
buf ( RI15b44880_203 , n1028 );
buf ( RI15b44808_202 , n1029 );
buf ( RI15b44790_201 , n1030 );
buf ( RI15b44718_200 , n1031 );
buf ( RI15b446a0_199 , n1032 );
buf ( RI15b44628_198 , n1033 );
buf ( RI15b445b0_197 , n1034 );
buf ( RI15b44538_196 , n1035 );
buf ( RI15b444c0_195 , n1036 );
buf ( RI15b44448_194 , n1037 );
buf ( RI15b443d0_193 , n1038 );
buf ( RI15b44358_192 , n1039 );
buf ( RI15b442e0_191 , n1040 );
buf ( RI15b44268_190 , n1041 );
buf ( RI15b441f0_189 , n1042 );
buf ( RI15b44178_188 , n1043 );
buf ( RI15b44100_187 , n1044 );
buf ( RI15b44088_186 , n1045 );
buf ( RI15b44010_185 , n1046 );
buf ( RI15b43f98_184 , n1047 );
buf ( RI15b43f20_183 , n1048 );
buf ( RI15b43ea8_182 , n1049 );
buf ( RI15b43e30_181 , n1050 );
buf ( RI15b43db8_180 , n1051 );
buf ( RI15b43d40_179 , n1052 );
buf ( RI15b43cc8_178 , n1053 );
buf ( RI15b43c50_177 , n1054 );
buf ( RI15b43bd8_176 , n1055 );
buf ( RI15b43b60_175 , n1056 );
buf ( RI15b43ae8_174 , n1057 );
buf ( RI15b532e0_703 , n1058 );
buf ( RI15b62a60_1231 , n1059 );
buf ( RI15b629e8_1230 , n1060 );
buf ( RI15b62970_1229 , n1061 );
buf ( RI15b628f8_1228 , n1062 );
buf ( RI15b62880_1227 , n1063 );
buf ( RI15b62808_1226 , n1064 );
buf ( RI15b62790_1225 , n1065 );
buf ( RI15b62718_1224 , n1066 );
buf ( RI15b626a0_1223 , n1067 );
buf ( RI15b62628_1222 , n1068 );
buf ( RI15b625b0_1221 , n1069 );
buf ( RI15b62538_1220 , n1070 );
buf ( RI15b624c0_1219 , n1071 );
buf ( RI15b62448_1218 , n1072 );
buf ( RI15b623d0_1217 , n1073 );
buf ( RI15b62358_1216 , n1074 );
buf ( RI15b622e0_1215 , n1075 );
buf ( RI15b62268_1214 , n1076 );
buf ( RI15b621f0_1213 , n1077 );
buf ( RI15b62178_1212 , n1078 );
buf ( RI15b5f6d0_1121 , n1079 );
buf ( RI15b5d1c8_1042 , n1080 );
buf ( RI15b5d150_1041 , n1081 );
buf ( RI15b5d0d8_1040 , n1082 );
buf ( RI15b5d060_1039 , n1083 );
buf ( RI15b5cfe8_1038 , n1084 );
buf ( RI15b45618_232 , n1085 );
buf ( RI15b52c50_689 , n1086 );
buf ( RI15b5e8c0_1091 , n1087 );
buf ( RI15b5e7d0_1089 , n1088 );
buf ( RI15b5e758_1088 , n1089 );
buf ( RI15b5d768_1054 , n1090 );
buf ( RI15b5d7e0_1055 , n1091 );
buf ( RI15b5d858_1056 , n1092 );
buf ( RI15b5d8d0_1057 , n1093 );
buf ( RI15b53538_708 , n1094 );
buf ( RI15b5f9a0_1127 , n1095 );
buf ( RI15b5ec08_1098 , n1096 );
buf ( RI15b614d0_1185 , n1097 );
buf ( RI15b61b60_1199 , n1098 );
buf ( RI15b61ae8_1198 , n1099 );
buf ( RI15b61a70_1197 , n1100 );
buf ( RI15b619f8_1196 , n1101 );
buf ( RI15b61980_1195 , n1102 );
buf ( RI15b61908_1194 , n1103 );
buf ( RI15b61890_1193 , n1104 );
buf ( RI15b61818_1192 , n1105 );
buf ( RI15b617a0_1191 , n1106 );
buf ( RI15b61728_1190 , n1107 );
buf ( RI15b616b0_1189 , n1108 );
buf ( RI15b61638_1188 , n1109 );
buf ( RI15b615c0_1187 , n1110 );
buf ( RI15b61548_1186 , n1111 );
buf ( RI15b526b0_677 , n1112 );
buf ( RI15b53100_699 , n1113 );
buf ( RI15b52cc8_690 , n1114 );
buf ( RI15b46ba8_278 , n1115 );
buf ( RI15b52bd8_688 , n1116 );
buf ( RI15b53f88_730 , n1117 );
buf ( RI15b603f0_1149 , n1118 );
buf ( RI15b45d98_248 , n1119 );
buf ( RI15b50dd8_624 , n1120 );
buf ( RI15b50d60_623 , n1121 );
buf ( RI15b50ce8_622 , n1122 );
buf ( RI15b50c70_621 , n1123 );
buf ( RI15b50bf8_620 , n1124 );
buf ( RI15b50b80_619 , n1125 );
buf ( RI15b475f8_300 , n1126 );
buf ( RI15b3fab0_37 , n1127 );
buf ( RI15b45168_222 , n1128 );
buf ( RI15b542d0_737 , n1129 );
buf ( RI15b45ac8_242 , n1130 );
buf ( RI15b527a0_679 , n1131 );
buf ( RI15b53088_698 , n1132 );
buf ( RI15b53808_714 , n1133 );
buf ( RI15b5ee60_1103 , n1134 );
buf ( RI15b60468_1150 , n1135 );
buf ( RI15b54618_744 , n1136 );
buf ( RI15b54708_746 , n1137 );
buf ( RI15b46fe0_287 , n1138 );
buf ( RI15b60918_1160 , n1139 );
buf ( RI15b52d40_691 , n1140 );
buf ( RI15b460e0_255 , n1141 );
buf ( RI15b476e8_302 , n1142 );
buf ( RI15b48c00_347 , n1143 );
buf ( RI15b49290_361 , n1144 );
buf ( RI15b49218_360 , n1145 );
buf ( RI15b491a0_359 , n1146 );
buf ( RI15b49128_358 , n1147 );
buf ( RI15b490b0_357 , n1148 );
buf ( RI15b49038_356 , n1149 );
buf ( RI15b48fc0_355 , n1150 );
buf ( RI15b48f48_354 , n1151 );
buf ( RI15b48ed0_353 , n1152 );
buf ( RI15b48e58_352 , n1153 );
buf ( RI15b48de0_351 , n1154 );
buf ( RI15b48d68_350 , n1155 );
buf ( RI15b48cf0_349 , n1156 );
buf ( RI15b48c78_348 , n1157 );
buf ( RI15b52638_676 , n1158 );
buf ( RI15b53c40_723 , n1159 );
buf ( RI15b468d8_272 , n1160 );
buf ( RI15b45ff0_253 , n1161 );
buf ( RI15b45f78_252 , n1162 );
buf ( RI15b45f00_251 , n1163 );
buf ( RI15b45e88_250 , n1164 );
buf ( RI15b44e98_216 , n1165 );
buf ( RI15b44f10_217 , n1166 );
buf ( RI15b44f88_218 , n1167 );
buf ( RI15b45000_219 , n1168 );
buf ( RI15b54258_736 , n1169 );
buf ( RI15b53b50_721 , n1170 );
buf ( RI15b5f0b8_1108 , n1171 );
buf ( RI15b53da8_726 , n1172 );
buf ( RI15b469c8_274 , n1173 );
buf ( RI15b5f220_1111 , n1174 );
buf ( RI15b47328_294 , n1175 );
buf ( RI15b45a50_241 , n1176 );
buf ( RI15b584e8_878 , n1177 );
buf ( RI15b5d240_1043 , n1178 );
buf ( RI15b52e30_693 , n1179 );
buf ( RI15b535b0_709 , n1180 );
buf ( RI15b53e20_727 , n1181 );
buf ( RI15b60288_1146 , n1182 );
buf ( RI15b3fc18_40 , n1183 );
buf ( RI15b44970_205 , n1184 );
buf ( RI15b448f8_204 , n1185 );
buf ( RI15b608a0_1159 , n1186 );
buf ( RI15b45780_235 , n1187 );
buf ( RI15b525c0_675 , n1188 );
buf ( RI15b47418_296 , n1189 );
buf ( RI15b5f310_1113 , n1190 );
buf ( RI15b44c40_211 , n1191 );
buf ( RI15b46a40_275 , n1192 );
buf ( RI15b60af8_1164 , n1193 );
buf ( RI15b47f58_320 , n1194 );
buf ( RI15b53718_712 , n1195 );
buf ( RI15b5fb80_1131 , n1196 );
buf ( RI15b52db8_692 , n1197 );
buf ( RI15b45d20_247 , n1198 );
buf ( RI15b52f20_695 , n1199 );
buf ( RI15b47ee0_319 , n1200 );
buf ( RI15b543c0_739 , n1201 );
buf ( RI15b5ef50_1105 , n1202 );
buf ( RI15b5ec80_1099 , n1203 );
buf ( RI15b53448_706 , n1204 );
buf ( RI15b529f8_684 , n1205 );
buf ( RI15b54000_731 , n1206 );
buf ( RI15b5f838_1124 , n1207 );
buf ( RI15b53880_715 , n1208 );
buf ( RI15b5fce8_1134 , n1209 );
buf ( RI15b46d10_281 , n1210 );
buf ( RI15b52890_681 , n1211 );
buf ( RI15b5f5e0_1119 , n1212 );
buf ( RI15b5fd60_1135 , n1213 );
buf ( RI15b454b0_229 , n1214 );
buf ( RI15b46860_271 , n1215 );
buf ( RI15b46ab8_276 , n1216 );
buf ( RI15b5f478_1116 , n1217 );
buf ( RI15b540f0_733 , n1218 );
buf ( RI15b60558_1152 , n1219 );
buf ( RI15b47490_297 , n1220 );
buf ( RI15b471c0_291 , n1221 );
buf ( RI15b47238_292 , n1222 );
buf ( RI15b53268_702 , n1223 );
buf ( RI15b539e8_718 , n1224 );
buf ( RI15b5f130_1109 , n1225 );
buf ( RI15b5fb08_1130 , n1226 );
buf ( RI15b607b0_1157 , n1227 );
buf ( RI15b544b0_741 , n1228 );
buf ( RI15b5eed8_1104 , n1229 );
buf ( RI15b604e0_1151 , n1230 );
buf ( RI15b510a8_630 , n1231 );
buf ( RI15b463b0_261 , n1232 );
buf ( RI15b46428_262 , n1233 );
buf ( RI15b5f298_1112 , n1234 );
buf ( RI15b5f1a8_1110 , n1235 );
buf ( RI15b47a30_309 , n1236 );
buf ( RI15b53bc8_722 , n1237 );
buf ( RI15b46338_260 , n1238 );
buf ( RI15b47c10_313 , n1239 );
buf ( RI15b48048_322 , n1240 );
buf ( RI15b464a0_263 , n1241 );
buf ( RI15b5ecf8_1100 , n1242 );
buf ( RI15b52ea8_694 , n1243 );
buf ( RI15b53628_710 , n1244 );
buf ( RI15b47850_305 , n1245 );
buf ( RI15b46068_254 , n1246 );
buf ( RI15b47670_301 , n1247 );
buf ( RI15b524d0_673 , n1248 );
buf ( RI15b53178_700 , n1249 );
buf ( RI15b52ae8_686 , n1250 );
buf ( RI15b451e0_223 , n1251 );
buf ( RI15b52548_674 , n1252 );
buf ( RI15b60030_1141 , n1253 );
buf ( RI15b457f8_236 , n1254 );
buf ( RI15b60990_1161 , n1255 );
buf ( RI15b53ad8_720 , n1256 );
buf ( RI15b5ff40_1139 , n1257 );
buf ( RI15b45528_230 , n1258 );
buf ( RI15b5fa18_1128 , n1259 );
buf ( RI15b53358_704 , n1260 );
buf ( RI15b5f7c0_1123 , n1261 );
buf ( RI15b462c0_259 , n1262 );
buf ( RI15b453c0_227 , n1263 );
buf ( RI15b45870_237 , n1264 );
buf ( RI15b46518_264 , n1265 );
buf ( RI15b47058_288 , n1266 );
buf ( RI15b60b70_1165 , n1267 );
buf ( RI15b45bb8_244 , n1268 );
buf ( RI15b533d0_705 , n1269 );
buf ( RI15b47e68_318 , n1270 );
buf ( RI15b47fd0_321 , n1271 );
buf ( RI15b5f568_1118 , n1272 );
buf ( RI15b480c0_323 , n1273 );
buf ( RI15b45960_239 , n1274 );
buf ( RI15b52980_683 , n1275 );
buf ( RI15b53cb8_724 , n1276 );
buf ( RI15b60120_1143 , n1277 );
buf ( RI15b5f4f0_1117 , n1278 );
buf ( RI15b46248_258 , n1279 );
buf ( RI15b46e78_284 , n1280 );
buf ( RI15b46590_265 , n1281 );
buf ( RI15b5fe50_1137 , n1282 );
buf ( RI15b47aa8_310 , n1283 );
buf ( RI15b47b20_311 , n1284 );
buf ( RI15b5efc8_1106 , n1285 );
buf ( RI15b60378_1148 , n1286 );
buf ( RI15b5ed70_1101 , n1287 );
buf ( RI15b46c20_279 , n1288 );
buf ( RI15b5d510_1049 , n1289 );
buf ( RI15b45258_224 , n1290 );
buf ( RI15b46f68_286 , n1291 );
buf ( RI15b461d0_257 , n1292 );
buf ( RI15b472b0_293 , n1293 );
buf ( RI15b5f928_1126 , n1294 );
buf ( RI15b536a0_711 , n1295 );
buf ( RI15b45b40_243 , n1296 );
buf ( RI15b48138_324 , n1297 );
buf ( RI15b5f400_1115 , n1298 );
buf ( RI15b46b30_277 , n1299 );
buf ( RI15b46608_266 , n1300 );
buf ( RI15b45690_233 , n1301 );
buf ( RI15b53790_713 , n1302 );
buf ( RI15b5fbf8_1132 , n1303 );
buf ( RI15b54078_732 , n1304 );
buf ( RI15b46c98_280 , n1305 );
buf ( RI15b53e98_728 , n1306 );
buf ( RI15b455a0_231 , n1307 );
buf ( RI15b47940_307 , n1308 );
buf ( RI15b45e10_249 , n1309 );
buf ( RI15b5fa90_1129 , n1310 );
buf ( RI15b54348_738 , n1311 );
buf ( RI15b60a08_1162 , n1312 );
buf ( RI15b531f0_701 , n1313 );
buf ( RI15b60210_1145 , n1314 );
buf ( RI15b478c8_306 , n1315 );
buf ( RI15b47c88_314 , n1316 );
buf ( RI15b46680_267 , n1317 );
buf ( RI15b46158_256 , n1318 );
buf ( RI15b5fc70_1133 , n1319 );
buf ( RI15b53a60_719 , n1320 );
buf ( RI15b538f8_716 , n1321 );
buf ( RI15b5eb18_1096 , n1322 );
buf ( RI15b5f040_1107 , n1323 );
buf ( RI15b52728_678 , n1324 );
buf ( RI15b5eaa0_1095 , n1325 );
buf ( RI15b600a8_1142 , n1326 );
buf ( RI15b5ede8_1102 , n1327 );
buf ( RI15b5eb90_1097 , n1328 );
buf ( RI15b60198_1144 , n1329 );
buf ( RI15b481b0_325 , n1330 );
buf ( RI15b545a0_743 , n1331 );
buf ( RI15b452d0_225 , n1332 );
buf ( RI15b46d88_282 , n1333 );
buf ( RI15b5ea28_1094 , n1334 );
buf ( RI15b54438_740 , n1335 );
buf ( RI15b47508_298 , n1336 );
buf ( RI15b466f8_268 , n1337 );
buf ( RI15b47148_290 , n1338 );
buf ( RI15b458e8_238 , n1339 );
buf ( RI15b52a70_685 , n1340 );
buf ( RI15b52818_680 , n1341 );
buf ( RI15b5e9b0_1093 , n1342 );
buf ( RI15b5ffb8_1140 , n1343 );
buf ( RI15b5f8b0_1125 , n1344 );
buf ( RI15b46ef0_285 , n1345 );
buf ( RI15b45ca8_246 , n1346 );
buf ( RI15b53970_717 , n1347 );
buf ( RI15b47580_299 , n1348 );
buf ( RI15b53010_697 , n1349 );
buf ( RI15b5e938_1092 , n1350 );
buf ( RI15b45078_220 , n1351 );
buf ( RI15b60300_1147 , n1352 );
buf ( RI15b46770_269 , n1353 );
buf ( RI15b60a80_1163 , n1354 );
buf ( RI15b473a0_295 , n1355 );
buf ( RI15b47760_303 , n1356 );
buf ( RI15b5f748_1122 , n1357 );
buf ( RI15b5fec8_1138 , n1358 );
buf ( RI15b45c30_245 , n1359 );
buf ( RI15b53d30_725 , n1360 );
buf ( RI15b45708_234 , n1361 );
buf ( RI15b54528_742 , n1362 );
buf ( RI15b459d8_240 , n1363 );
buf ( n1364 , R_187c_13cca558 );
buf ( n1365 , R_125d_156aaaf8 );
buf ( n1366 , R_c3e_13d2c178 );
buf ( n1367 , R_61f_117eb278 );
buf ( n1368 , R_187d_117f5b38 );
buf ( n1369 , R_125e_13b8fe18 );
buf ( n1370 , R_c3f_123b4358 );
buf ( n1371 , R_187b_13ccb278 );
buf ( n1372 , R_620_13dfb518 );
buf ( n1373 , R_125c_15816b78 );
buf ( n1374 , R_c3d_13c22918 );
buf ( n1375 , R_61e_14a0c538 );
buf ( n1376 , R_5e7_10080958 );
buf ( n1377 , R_c06_170189e8 );
buf ( n1378 , R_18b4_1162f978 );
buf ( n1379 , R_1225_13c08298 );
buf ( n1380 , R_1844_117ef378 );
buf ( n1381 , R_1295_123bcf58 );
buf ( n1382 , R_c76_15ff42e8 );
buf ( n1383 , R_657_13bf5c78 );
buf ( n1384 , R_187e_140ac0d8 );
buf ( n1385 , R_125f_13c0f638 );
buf ( n1386 , R_c40_1580a9b8 );
buf ( n1387 , R_621_11c70318 );
buf ( n1388 , R_187a_13ddd2d8 );
buf ( n1389 , R_61d_123b84f8 );
buf ( n1390 , R_125b_1162bf58 );
buf ( n1391 , R_c3c_15ff9928 );
buf ( n1392 , R_12be_13ccf378 );
buf ( n1393 , R_5be_11c6a738 );
buf ( n1394 , R_bdd_17016508 );
buf ( n1395 , R_c9f_11636598 );
buf ( n1396 , R_11fc_13ddf7b8 );
buf ( n1397 , R_680_10085638 );
buf ( n1398 , R_181b_13d430d8 );
buf ( n1399 , R_18dd_13c062b8 );
buf ( n1400 , R_180c_156b4eb8 );
buf ( n1401 , R_12cd_13d535d8 );
buf ( n1402 , R_5af_1700c3c8 );
buf ( n1403 , R_cae_14a14ff8 );
buf ( n1404 , R_bce_15ff4608 );
buf ( n1405 , R_68f_13befcd8 );
buf ( n1406 , R_18ec_13d204b8 );
buf ( n1407 , R_11ed_116361d8 );
buf ( n1408 , R_187f_15811038 );
buf ( n1409 , R_1260_13d3b6f8 );
buf ( n1410 , R_c41_14a0bef8 );
buf ( n1411 , R_622_123b3bd8 );
buf ( n1412 , R_61c_13d56378 );
buf ( n1413 , R_c3b_150e7c58 );
buf ( n1414 , R_1879_15ff5c88 );
buf ( n1415 , R_125a_13bf58b8 );
buf ( n1416 , R_f82_13c1cd38 );
buf ( n1417 , R_963_13c209d8 );
buf ( n1418 , R_8fa_117ec678 );
buf ( n1419 , R_f19_15ff0648 );
buf ( n1420 , R_1538_13d29bf8 );
buf ( n1421 , R_15a1_150e22f8 );
buf ( n1422 , R_158f_13cd9058 );
buf ( n1423 , R_f70_17015608 );
buf ( n1424 , R_951_156b2578 );
buf ( n1425 , R_90c_13c0e0f8 );
buf ( n1426 , R_f2b_140b8838 );
buf ( n1427 , R_154a_1587f278 );
buf ( n1428 , R_1880_13c22738 );
buf ( n1429 , R_1261_13ccc0d8 );
buf ( n1430 , R_c42_117eb818 );
buf ( n1431 , R_623_140b3158 );
buf ( n1432 , R_61b_11c70458 );
buf ( n1433 , R_c3a_13b96218 );
buf ( n1434 , R_1259_13d23578 );
buf ( n1435 , R_1878_1162da38 );
buf ( n1436 , R_ce6_14875d78 );
buf ( n1437 , R_1924_13d1df38 );
buf ( n1438 , R_11b5_13d56f58 );
buf ( n1439 , R_577_1162c818 );
buf ( n1440 , R_6c7_10082438 );
buf ( n1441 , R_17d4_13cda278 );
buf ( n1442 , R_1305_10081fd8 );
buf ( n1443 , R_b96_15812b18 );
buf ( n1444 , R_1881_156b0638 );
buf ( n1445 , R_1262_12fc1698 );
buf ( n1446 , R_c43_140b0138 );
buf ( n1447 , R_624_13d421d8 );
buf ( n1448 , R_61a_14b2a318 );
buf ( n1449 , R_c39_117eaeb8 );
buf ( n1450 , R_1258_117e8618 );
buf ( n1451 , R_1877_1162cdb8 );
buf ( n1452 , R_119b_15ffa3c8 );
buf ( n1453 , R_55d_13b8e5b8 );
buf ( n1454 , R_131f_158106d8 );
buf ( n1455 , R_6e1_13c0fb38 );
buf ( n1456 , R_17ba_15fed6c8 );
buf ( n1457 , R_b7c_13b96e98 );
buf ( n1458 , R_193e_123b6018 );
buf ( n1459 , R_d00_117ec358 );
buf ( n1460 , R_1323_13d5b878 );
buf ( n1461 , R_6e5_15ff5328 );
buf ( n1462 , R_559_13c024d8 );
buf ( n1463 , R_1197_13bf4918 );
buf ( n1464 , R_1942_11c6dd98 );
buf ( n1465 , R_d04_14a16df8 );
buf ( n1466 , R_17b6_13dec158 );
buf ( n1467 , R_b78_13c10c18 );
buf ( n1468 , R_13ca_13d2c718 );
buf ( n1469 , R_19e9_13bf62b8 );
buf ( n1470 , R_170f_150defb8 );
buf ( n1471 , R_10f0_140b1ad8 );
buf ( n1472 , R_ad1_11c6ac38 );
buf ( n1473 , R_78c_13d5d3f8 );
buf ( n1474 , R_dab_140b3dd8 );
buf ( n1475 , R_883_13b936f8 );
buf ( n1476 , R_ff9_11631958 );
buf ( n1477 , R_ea2_150dd758 );
buf ( n1478 , R_9da_13cd8018 );
buf ( n1479 , R_1618_117f3658 );
buf ( n1480 , R_14c1_123ba4d8 );
buf ( n1481 , R_b5e_14a0f918 );
buf ( n1482 , R_179c_123bb018 );
buf ( n1483 , R_133d_13cd4e18 );
buf ( n1484 , R_6ff_14a0a918 );
buf ( n1485 , R_195c_150ddf78 );
buf ( n1486 , R_117d_123b8c78 );
buf ( n1487 , R_d1e_124c2cd8 );
buf ( n1488 , R_5f7_12fbf758 );
buf ( n1489 , R_c16_13df9858 );
buf ( n1490 , R_1235_15880cb8 );
buf ( n1491 , R_1854_1580fd78 );
buf ( n1492 , R_18a4_13bf2d98 );
buf ( n1493 , R_1285_100890f8 );
buf ( n1494 , R_c66_13bed2f8 );
buf ( n1495 , R_647_13d51af8 );
buf ( n1496 , R_1882_13d1fbf8 );
buf ( n1497 , R_1263_123be498 );
buf ( n1498 , R_c44_13c229b8 );
buf ( n1499 , R_625_13c1e638 );
buf ( n1500 , R_619_156b6718 );
buf ( n1501 , R_c38_117efd78 );
buf ( n1502 , R_1257_14a0f0f8 );
buf ( n1503 , R_1876_15ffcb28 );
buf ( n1504 , R_985_1587c4d8 );
buf ( n1505 , R_1516_12fc1eb8 );
buf ( n1506 , R_15c3_13c02078 );
buf ( n1507 , R_8d8_13d22fd8 );
buf ( n1508 , R_fa4_13d1e898 );
buf ( n1509 , R_ef7_1162bd78 );
buf ( n1510 , R_1663_124c2698 );
buf ( n1511 , R_838_1580b8b8 );
buf ( n1512 , R_a25_13bf4ff8 );
buf ( n1513 , R_1476_1486bd78 );
buf ( n1514 , R_1044_13d57818 );
buf ( n1515 , R_e57_13b8f738 );
buf ( n1516 , R_15fa_13c0bb78 );
buf ( n1517 , R_ec0_13c1bf78 );
buf ( n1518 , R_fdb_15ff7308 );
buf ( n1519 , R_14df_14a0cdf8 );
buf ( n1520 , R_9bc_15812758 );
buf ( n1521 , R_8a1_13d21818 );
buf ( n1522 , R_1883_13d41058 );
buf ( n1523 , R_1264_13c02758 );
buf ( n1524 , R_c45_13d24c98 );
buf ( n1525 , R_626_123b86d8 );
buf ( n1526 , R_618_1587ea58 );
buf ( n1527 , R_c37_13c0bfd8 );
buf ( n1528 , R_1256_13d54258 );
buf ( n1529 , R_1875_158179d8 );
buf ( n1530 , R_1145_13b98658 );
buf ( n1531 , R_737_116313b8 );
buf ( n1532 , R_b26_1486a518 );
buf ( n1533 , R_d56_117e9d38 );
buf ( n1534 , R_1764_13ccf7d8 );
buf ( n1535 , R_1375_13c275f8 );
buf ( n1536 , R_1994_123bac58 );
buf ( n1537 , R_143d_13bf2258 );
buf ( n1538 , R_a5e_1587ed78 );
buf ( n1539 , R_e1e_13c1bbb8 );
buf ( n1540 , R_107d_15888418 );
buf ( n1541 , R_7ff_13cd45f8 );
buf ( n1542 , R_169c_15885fd8 );
buf ( n1543 , R_1a5c_13de04d8 );
buf ( n1544 , R_1a48_13c1ff38 );
buf ( n1545 , R_a72_1486d358 );
buf ( n1546 , R_1429_13d23438 );
buf ( n1547 , R_1091_14a11d58 );
buf ( n1548 , R_e0a_13bfa3b8 );
buf ( n1549 , R_16b0_140aae18 );
buf ( n1550 , R_7eb_123b8278 );
buf ( n1551 , R_12c6_13cd49b8 );
buf ( n1552 , R_5b6_117f1f38 );
buf ( n1553 , R_ca7_140b4418 );
buf ( n1554 , R_bd5_13d51698 );
buf ( n1555 , R_688_13b99af8 );
buf ( n1556 , R_11f4_13d1e6b8 );
buf ( n1557 , R_18e5_13d45658 );
buf ( n1558 , R_1813_13d29c98 );
buf ( n1559 , R_16d9_14a17cf8 );
buf ( n1560 , R_1a1f_11c70958 );
buf ( n1561 , R_1400_14b29b98 );
buf ( n1562 , R_de1_13cd0638 );
buf ( n1563 , R_7c2_15ffa508 );
buf ( n1564 , R_a9b_100865d8 );
buf ( n1565 , R_10ba_15881938 );
buf ( n1566 , R_1805_14b271b8 );
buf ( n1567 , R_5a8_123b8318 );
buf ( n1568 , R_cb5_170107e8 );
buf ( n1569 , R_bc7_13c2a758 );
buf ( n1570 , R_696_10082ed8 );
buf ( n1571 , R_18f3_15ffc628 );
buf ( n1572 , R_11e6_14b222f8 );
buf ( n1573 , R_12d4_11634d38 );
buf ( n1574 , R_119f_156b4738 );
buf ( n1575 , R_561_1162a658 );
buf ( n1576 , R_6dd_117f36f8 );
buf ( n1577 , R_131b_15ff76c8 );
buf ( n1578 , R_17be_15816538 );
buf ( n1579 , R_b80_13cd8338 );
buf ( n1580 , R_cfc_1700d2c8 );
buf ( n1581 , R_193a_15885718 );
buf ( n1582 , R_5da_13df70f8 );
buf ( n1583 , R_18c1_11c6f738 );
buf ( n1584 , R_bf9_13d28ed8 );
buf ( n1585 , R_12a2_13bf2578 );
buf ( n1586 , R_1218_13d28078 );
buf ( n1587 , R_c83_13d59f78 );
buf ( n1588 , R_1837_13deb9d8 );
buf ( n1589 , R_664_123b47b8 );
buf ( n1590 , R_e39_156b3518 );
buf ( n1591 , R_a43_14b1feb8 );
buf ( n1592 , R_81a_13cceb58 );
buf ( n1593 , R_1062_117eedd8 );
buf ( n1594 , R_1458_13df07f8 );
buf ( n1595 , R_1681_140b99b8 );
buf ( n1596 , R_1327_124c2b98 );
buf ( n1597 , R_6e9_156b3158 );
buf ( n1598 , R_555_13d59b18 );
buf ( n1599 , R_1193_13b97438 );
buf ( n1600 , R_1946_14a16858 );
buf ( n1601 , R_d08_13d59938 );
buf ( n1602 , R_b74_123c0478 );
buf ( n1603 , R_17b2_13cd6498 );
buf ( n1604 , R_113a_117eb458 );
buf ( n1605 , R_742_14a129d8 );
buf ( n1606 , R_b1b_11629758 );
buf ( n1607 , R_d61_11633618 );
buf ( n1608 , R_1380_15887338 );
buf ( n1609 , R_1759_14874518 );
buf ( n1610 , R_199f_13d3c9b8 );
buf ( n1611 , R_1884_13cd1c18 );
buf ( n1612 , R_1265_156b0818 );
buf ( n1613 , R_c46_1580b598 );
buf ( n1614 , R_627_117efb98 );
buf ( n1615 , R_617_158807b8 );
buf ( n1616 , R_c36_156b63f8 );
buf ( n1617 , R_1255_1580dbb8 );
buf ( n1618 , R_1874_13df9c18 );
buf ( n1619 , R_87a_13c286d8 );
buf ( n1620 , R_1002_14a17938 );
buf ( n1621 , R_e99_123ba258 );
buf ( n1622 , R_9e3_170110a8 );
buf ( n1623 , R_1621_117eacd8 );
buf ( n1624 , R_14b8_123b31d8 );
buf ( n1625 , R_edf_117f5bd8 );
buf ( n1626 , R_14fe_13d55518 );
buf ( n1627 , R_15db_117f7258 );
buf ( n1628 , R_fbc_13beb9f8 );
buf ( n1629 , R_8c0_11631ef8 );
buf ( n1630 , R_99d_13cd4d78 );
buf ( n1631 , R_845_15888918 );
buf ( n1632 , R_1656_117f4af8 );
buf ( n1633 , R_1483_13d53d58 );
buf ( n1634 , R_a18_12fbdef8 );
buf ( n1635 , R_e64_14875058 );
buf ( n1636 , R_1037_15815098 );
buf ( n1637 , R_d8e_11630878 );
buf ( n1638 , R_172c_13d39d58 );
buf ( n1639 , R_13ad_14a12618 );
buf ( n1640 , R_19cc_13cda1d8 );
buf ( n1641 , R_110d_13dd5cb8 );
buf ( n1642 , R_aee_117e9478 );
buf ( n1643 , R_76f_117f4378 );
buf ( n1644 , R_ccd_13b8c8f8 );
buf ( n1645 , R_590_13dd64d8 );
buf ( n1646 , R_17ed_156b36f8 );
buf ( n1647 , R_190b_14872038 );
buf ( n1648 , R_6ae_156ab958 );
buf ( n1649 , R_baf_1700cd28 );
buf ( n1650 , R_12ec_124c3778 );
buf ( n1651 , R_11ce_11c6cad8 );
buf ( n1652 , R_17a3_150e7398 );
buf ( n1653 , R_1336_148754b8 );
buf ( n1654 , R_6f8_13c1c018 );
buf ( n1655 , R_1184_150e6498 );
buf ( n1656 , R_1955_14b235b8 );
buf ( n1657 , R_d17_14b27398 );
buf ( n1658 , R_b65_13dde318 );
buf ( n1659 , R_1885_1486cdb8 );
buf ( n1660 , R_1266_14a12438 );
buf ( n1661 , R_c47_100803b8 );
buf ( n1662 , R_628_117eb098 );
buf ( n1663 , R_616_170152e8 );
buf ( n1664 , R_c35_123b88b8 );
buf ( n1665 , R_1254_150e59f8 );
buf ( n1666 , R_1873_12fc2278 );
buf ( n1667 , R_74a_1008cb18 );
buf ( n1668 , R_1132_15880e98 );
buf ( n1669 , R_d69_14b23158 );
buf ( n1670 , R_b13_140b3d38 );
buf ( n1671 , R_1388_140aaf58 );
buf ( n1672 , R_19a7_140b9b98 );
buf ( n1673 , R_1751_1007feb8 );
buf ( n1674 , R_b57_13ccd6b8 );
buf ( n1675 , R_1344_117f3018 );
buf ( n1676 , R_1795_1008b678 );
buf ( n1677 , R_706_1580bd18 );
buf ( n1678 , R_1963_13d1f478 );
buf ( n1679 , R_1176_17015b08 );
buf ( n1680 , R_d25_15882298 );
buf ( n1681 , R_1590_150e4b98 );
buf ( n1682 , R_f71_124c4998 );
buf ( n1683 , R_952_14b26e98 );
buf ( n1684 , R_90b_13d41af8 );
buf ( n1685 , R_f2a_1162a158 );
buf ( n1686 , R_1549_1587ff98 );
buf ( n1687 , R_5c6_15816218 );
buf ( n1688 , R_12b6_1587db58 );
buf ( n1689 , R_be5_140b5818 );
buf ( n1690 , R_c97_156b09f8 );
buf ( n1691 , R_1204_13c23b38 );
buf ( n1692 , R_678_15884ef8 );
buf ( n1693 , R_1823_13d53df8 );
buf ( n1694 , R_18d5_11636098 );
buf ( n1695 , R_ed8_117e9c98 );
buf ( n1696 , R_15e2_14a140f8 );
buf ( n1697 , R_14f7_13b965d8 );
buf ( n1698 , R_fc3_14b27e38 );
buf ( n1699 , R_8b9_14875e18 );
buf ( n1700 , R_9a4_117ee018 );
buf ( n1701 , R_1a04_13c22b98 );
buf ( n1702 , R_13e5_13de07f8 );
buf ( n1703 , R_16f4_123b9fd8 );
buf ( n1704 , R_dc6_14873f78 );
buf ( n1705 , R_10d5_13b94a58 );
buf ( n1706 , R_7a7_116355f8 );
buf ( n1707 , R_ab6_15814e18 );
buf ( n1708 , R_1886_11638c58 );
buf ( n1709 , R_1267_14b23f18 );
buf ( n1710 , R_c48_13bf5e58 );
buf ( n1711 , R_629_150e7e38 );
buf ( n1712 , R_615_13c1d7d8 );
buf ( n1713 , R_c34_15ff1228 );
buf ( n1714 , R_1253_13d222b8 );
buf ( n1715 , R_1872_13ccb4f8 );
buf ( n1716 , R_16f6_116389d8 );
buf ( n1717 , R_10d7_156b5778 );
buf ( n1718 , R_ab8_156ac8f8 );
buf ( n1719 , R_1a02_13cd8298 );
buf ( n1720 , R_13e3_14a0a7d8 );
buf ( n1721 , R_7a5_13d456f8 );
buf ( n1722 , R_dc4_11634b58 );
buf ( n1723 , R_b4d_1700f208 );
buf ( n1724 , R_710_156ac718 );
buf ( n1725 , R_178b_1580ca38 );
buf ( n1726 , R_196d_117eb8b8 );
buf ( n1727 , R_d2f_13dedf58 );
buf ( n1728 , R_116c_140b8338 );
buf ( n1729 , R_134e_13d282f8 );
buf ( n1730 , R_1a06_1486e1b8 );
buf ( n1731 , R_13e7_116377b8 );
buf ( n1732 , R_dc8_1162b058 );
buf ( n1733 , R_7a9_123bd458 );
buf ( n1734 , R_16f2_158857b8 );
buf ( n1735 , R_ab4_12fbed58 );
buf ( n1736 , R_10d3_158899f8 );
buf ( n1737 , R_85a_156b1a38 );
buf ( n1738 , R_1498_15811c18 );
buf ( n1739 , R_1641_150db8b8 );
buf ( n1740 , R_a03_123bd818 );
buf ( n1741 , R_e79_13cd8658 );
buf ( n1742 , R_1022_11c6cf38 );
buf ( n1743 , R_150d_14b21678 );
buf ( n1744 , R_15cc_14a0ba98 );
buf ( n1745 , R_8cf_13ded9b8 );
buf ( n1746 , R_fad_140ac038 );
buf ( n1747 , R_eee_11632e98 );
buf ( n1748 , R_98e_12fbecb8 );
buf ( n1749 , R_13bd_13df6c98 );
buf ( n1750 , R_19dc_156b6858 );
buf ( n1751 , R_171c_117ecb78 );
buf ( n1752 , R_10fd_117eef18 );
buf ( n1753 , R_ade_13dd7658 );
buf ( n1754 , R_77f_117f4558 );
buf ( n1755 , R_d9e_13ddc3d8 );
buf ( n1756 , R_16f8_14a0e018 );
buf ( n1757 , R_10d9_123b9538 );
buf ( n1758 , R_aba_13c29678 );
buf ( n1759 , R_7a3_13ccb138 );
buf ( n1760 , R_dc2_158108b8 );
buf ( n1761 , R_13e1_156b8478 );
buf ( n1762 , R_1a00_123b7f58 );
buf ( n1763 , R_971_13df5618 );
buf ( n1764 , R_8ec_123bbd38 );
buf ( n1765 , R_15af_14866eb8 );
buf ( n1766 , R_f0b_13cd72f8 );
buf ( n1767 , R_f90_15812438 );
buf ( n1768 , R_152a_13df8818 );
buf ( n1769 , R_c15_15fee528 );
buf ( n1770 , R_1234_15ff9e28 );
buf ( n1771 , R_1853_13dd8738 );
buf ( n1772 , R_18a5_170177c8 );
buf ( n1773 , R_1286_124c4858 );
buf ( n1774 , R_c67_13ccba98 );
buf ( n1775 , R_648_15814058 );
buf ( n1776 , R_5f6_13cce018 );
buf ( n1777 , R_c05_14866d78 );
buf ( n1778 , R_18b5_10087cf8 );
buf ( n1779 , R_1224_13ccff58 );
buf ( n1780 , R_1296_13dda7b8 );
buf ( n1781 , R_1843_1580a878 );
buf ( n1782 , R_c77_13d523b8 );
buf ( n1783 , R_658_140ae1f8 );
buf ( n1784 , R_5e6_13d46698 );
buf ( n1785 , R_1a08_14b1b958 );
buf ( n1786 , R_13e9_13d22358 );
buf ( n1787 , R_dca_14b297d8 );
buf ( n1788 , R_7ab_15887ab8 );
buf ( n1789 , R_ab2_13df75f8 );
buf ( n1790 , R_10d1_13d55d38 );
buf ( n1791 , R_16f0_14b1e978 );
buf ( n1792 , R_d87_123bae38 );
buf ( n1793 , R_1733_15ff79e8 );
buf ( n1794 , R_13a6_156b1718 );
buf ( n1795 , R_1114_13d46ff8 );
buf ( n1796 , R_19c5_13bf6ad8 );
buf ( n1797 , R_af5_13c1b6b8 );
buf ( n1798 , R_768_158896d8 );
buf ( n1799 , R_964_123c1f58 );
buf ( n1800 , R_8f9_117ee658 );
buf ( n1801 , R_f18_14a19d78 );
buf ( n1802 , R_1537_117e9b58 );
buf ( n1803 , R_15a2_13ccce98 );
buf ( n1804 , R_f83_14a0e978 );
buf ( n1805 , R_1887_17018da8 );
buf ( n1806 , R_1268_13d38278 );
buf ( n1807 , R_c49_123b36d8 );
buf ( n1808 , R_62a_13d42278 );
buf ( n1809 , R_614_13c2a258 );
buf ( n1810 , R_c33_150e7bb8 );
buf ( n1811 , R_1252_116378f8 );
buf ( n1812 , R_1871_13defad8 );
buf ( n1813 , R_11a3_13c1be38 );
buf ( n1814 , R_565_13ddbb18 );
buf ( n1815 , R_6d9_11636818 );
buf ( n1816 , R_1317_1580c5d8 );
buf ( n1817 , R_17c2_13c03518 );
buf ( n1818 , R_b84_156b5278 );
buf ( n1819 , R_cf8_15881a78 );
buf ( n1820 , R_1936_13d2a558 );
buf ( n1821 , R_13b4_156abb38 );
buf ( n1822 , R_19d3_13bf92d8 );
buf ( n1823 , R_1725_13cd9a58 );
buf ( n1824 , R_1106_14b1c718 );
buf ( n1825 , R_ae7_13cd22f8 );
buf ( n1826 , R_776_14873bb8 );
buf ( n1827 , R_d95_15815778 );
buf ( n1828 , R_feb_1486c818 );
buf ( n1829 , R_eb0_13d53498 );
buf ( n1830 , R_14cf_14b1bd18 );
buf ( n1831 , R_9cc_158172f8 );
buf ( n1832 , R_160a_17010ce8 );
buf ( n1833 , R_891_13b8ab98 );
buf ( n1834 , R_132b_1007f7d8 );
buf ( n1835 , R_6ed_140b6538 );
buf ( n1836 , R_118f_14b1ee78 );
buf ( n1837 , R_194a_13d2ae18 );
buf ( n1838 , R_d0c_13dee8b8 );
buf ( n1839 , R_b70_13d20f58 );
buf ( n1840 , R_17ae_13d29a18 );
buf ( n1841 , R_1a3c_13b95278 );
buf ( n1842 , R_109d_10084878 );
buf ( n1843 , R_141d_13d441b8 );
buf ( n1844 , R_16bc_14a0bdb8 );
buf ( n1845 , R_dfe_15ff38e8 );
buf ( n1846 , R_7df_1587d338 );
buf ( n1847 , R_a7e_14a0bb38 );
buf ( n1848 , R_151f_12fbe998 );
buf ( n1849 , R_97c_13d528b8 );
buf ( n1850 , R_15ba_1008b0d8 );
buf ( n1851 , R_8e1_15889818 );
buf ( n1852 , R_f00_17017ae8 );
buf ( n1853 , R_f9b_13b974d8 );
buf ( n1854 , R_16fa_14b299b8 );
buf ( n1855 , R_10db_13cd6cb8 );
buf ( n1856 , R_abc_15882b58 );
buf ( n1857 , R_7a1_15ffcd08 );
buf ( n1858 , R_dc0_117f53b8 );
buf ( n1859 , R_13df_156b9238 );
buf ( n1860 , R_19fe_13c01fd8 );
buf ( n1861 , R_5cf_124c4678 );
buf ( n1862 , R_12ad_13cca878 );
buf ( n1863 , R_bee_156ac498 );
buf ( n1864 , R_c8e_156b6cb8 );
buf ( n1865 , R_120d_123be218 );
buf ( n1866 , R_66f_13df8d18 );
buf ( n1867 , R_182c_13b90598 );
buf ( n1868 , R_18cc_170190c8 );
buf ( n1869 , R_1505_13d27858 );
buf ( n1870 , R_15d4_13d3a078 );
buf ( n1871 , R_fb5_13c265b8 );
buf ( n1872 , R_8c7_13ccf738 );
buf ( n1873 , R_996_13cd1498 );
buf ( n1874 , R_ee6_156ae158 );
buf ( n1875 , R_1a0a_140b9238 );
buf ( n1876 , R_13eb_150e7438 );
buf ( n1877 , R_dcc_15815c78 );
buf ( n1878 , R_7ad_1008c078 );
buf ( n1879 , R_ab0_11629618 );
buf ( n1880 , R_10cf_1580df78 );
buf ( n1881 , R_16ee_123bf758 );
buf ( n1882 , R_1660_13dd6258 );
buf ( n1883 , R_83b_117f03b8 );
buf ( n1884 , R_a22_156b92d8 );
buf ( n1885 , R_1479_13ddc518 );
buf ( n1886 , R_1041_14a0db18 );
buf ( n1887 , R_e5a_11633118 );
buf ( n1888 , R_1711_11c69d38 );
buf ( n1889 , R_10f2_1486ad38 );
buf ( n1890 , R_ad3_13d5a5b8 );
buf ( n1891 , R_78a_13dfa2f8 );
buf ( n1892 , R_da9_123bc9b8 );
buf ( n1893 , R_13c8_11628e98 );
buf ( n1894 , R_19e7_14a10098 );
buf ( n1895 , R_eb5_13cd9cd8 );
buf ( n1896 , R_fe6_13df1d38 );
buf ( n1897 , R_14d4_13c27a58 );
buf ( n1898 , R_9c7_140af5f8 );
buf ( n1899 , R_896_123b6658 );
buf ( n1900 , R_1605_156b1b78 );
buf ( n1901 , R_1888_1580c858 );
buf ( n1902 , R_1269_13b99c38 );
buf ( n1903 , R_c4a_14a0cb78 );
buf ( n1904 , R_62b_1162a1f8 );
buf ( n1905 , R_613_124c47b8 );
buf ( n1906 , R_c32_14b23518 );
buf ( n1907 , R_1251_13d3fed8 );
buf ( n1908 , R_1870_13b92bb8 );
buf ( n1909 , R_16cc_156ba318 );
buf ( n1910 , R_1a2c_156b08b8 );
buf ( n1911 , R_140d_11638258 );
buf ( n1912 , R_dee_13c0e058 );
buf ( n1913 , R_7cf_123bbe78 );
buf ( n1914 , R_a8e_170160a8 );
buf ( n1915 , R_10ad_10082618 );
buf ( n1916 , R_11b0_13b99f58 );
buf ( n1917 , R_572_140ab458 );
buf ( n1918 , R_6cc_117e8a78 );
buf ( n1919 , R_130a_13dda498 );
buf ( n1920 , R_17cf_13d389f8 );
buf ( n1921 , R_b91_14b1f418 );
buf ( n1922 , R_ceb_13d56d78 );
buf ( n1923 , R_1929_13cd4af8 );
buf ( n1924 , R_f72_13c2a1b8 );
buf ( n1925 , R_953_14b20a98 );
buf ( n1926 , R_90a_156ae658 );
buf ( n1927 , R_f29_11630698 );
buf ( n1928 , R_1548_140ac538 );
buf ( n1929 , R_1591_13c25618 );
buf ( n1930 , R_16fc_156b9a58 );
buf ( n1931 , R_10dd_13d551f8 );
buf ( n1932 , R_abe_14a15958 );
buf ( n1933 , R_79f_140af7d8 );
buf ( n1934 , R_dbe_13cd4c38 );
buf ( n1935 , R_13dd_15884b38 );
buf ( n1936 , R_19fc_13b96fd8 );
buf ( n1937 , R_ff0_123b3b38 );
buf ( n1938 , R_eab_11634518 );
buf ( n1939 , R_9d1_13d4ed58 );
buf ( n1940 , R_14ca_11631e58 );
buf ( n1941 , R_160f_170102e8 );
buf ( n1942 , R_88c_116319f8 );
buf ( n1943 , R_e36_13c05b38 );
buf ( n1944 , R_a46_11637e98 );
buf ( n1945 , R_817_116294d8 );
buf ( n1946 , R_1065_13c0b218 );
buf ( n1947 , R_1455_117ef238 );
buf ( n1948 , R_1684_13dd5ad8 );
buf ( n1949 , R_e2b_13d28578 );
buf ( n1950 , R_a51_11630ff8 );
buf ( n1951 , R_80c_13d2acd8 );
buf ( n1952 , R_1070_150e2d98 );
buf ( n1953 , R_1a69_11c6fe18 );
buf ( n1954 , R_168f_13d295b8 );
buf ( n1955 , R_144a_1580c678 );
buf ( n1956 , R_1a0c_13ccacd8 );
buf ( n1957 , R_13ed_13cd4ff8 );
buf ( n1958 , R_dce_14871f98 );
buf ( n1959 , R_7af_11633578 );
buf ( n1960 , R_aae_15814238 );
buf ( n1961 , R_10cd_13d20878 );
buf ( n1962 , R_16ec_13df6a18 );
buf ( n1963 , R_1889_13bf9c38 );
buf ( n1964 , R_126a_15886a78 );
buf ( n1965 , R_c4b_13cd76b8 );
buf ( n1966 , R_62c_10086038 );
buf ( n1967 , R_612_10088dd8 );
buf ( n1968 , R_c31_13b90778 );
buf ( n1969 , R_1250_13d58c18 );
buf ( n1970 , R_186f_1162dcb8 );
buf ( n1971 , R_1a21_150e5598 );
buf ( n1972 , R_1402_140b1cb8 );
buf ( n1973 , R_de3_140b0778 );
buf ( n1974 , R_7c4_13cd5138 );
buf ( n1975 , R_a99_13cd0a98 );
buf ( n1976 , R_10b8_13bea7d8 );
buf ( n1977 , R_16d7_15888a58 );
buf ( n1978 , R_b23_1587bc18 );
buf ( n1979 , R_d59_14868cb8 );
buf ( n1980 , R_1378_14b28158 );
buf ( n1981 , R_1761_11631f98 );
buf ( n1982 , R_1997_13d45158 );
buf ( n1983 , R_1142_117f06d8 );
buf ( n1984 , R_73a_13de1158 );
buf ( n1985 , R_1a35_1486d7b8 );
buf ( n1986 , R_16c3_13c01498 );
buf ( n1987 , R_1416_1162ee38 );
buf ( n1988 , R_df7_117f35b8 );
buf ( n1989 , R_7d8_156abc78 );
buf ( n1990 , R_a85_17014168 );
buf ( n1991 , R_10a4_1486b0f8 );
buf ( n1992 , R_a59_14a1a1d8 );
buf ( n1993 , R_e23_13df5f78 );
buf ( n1994 , R_1078_1580f558 );
buf ( n1995 , R_804_156b6f38 );
buf ( n1996 , R_1697_13d59d98 );
buf ( n1997 , R_1a61_14a195f8 );
buf ( n1998 , R_1442_14a18c98 );
buf ( n1999 , R_1096_13dd6f78 );
buf ( n2000 , R_1424_13b906d8 );
buf ( n2001 , R_16b5_13c045f8 );
buf ( n2002 , R_e05_140ad938 );
buf ( n2003 , R_7e6_1486dd58 );
buf ( n2004 , R_a77_100895f8 );
buf ( n2005 , R_1a43_170104c8 );
buf ( n2006 , R_15ef_15889318 );
buf ( n2007 , R_ecb_13df7198 );
buf ( n2008 , R_14ea_13cd2078 );
buf ( n2009 , R_fd0_13cd59f8 );
buf ( n2010 , R_8ac_15889278 );
buf ( n2011 , R_9b1_1008a3b8 );
buf ( n2012 , R_cc2_14a11218 );
buf ( n2013 , R_17f8_13c28d18 );
buf ( n2014 , R_59b_15812bb8 );
buf ( n2015 , R_1900_1486c318 );
buf ( n2016 , R_6a3_11c69658 );
buf ( n2017 , R_bba_13deb7f8 );
buf ( n2018 , R_12e1_123bbf18 );
buf ( n2019 , R_11d9_14a18518 );
buf ( n2020 , R_1125_124c3e58 );
buf ( n2021 , R_d76_156b6218 );
buf ( n2022 , R_b06_14b24af8 );
buf ( n2023 , R_1395_13c0d978 );
buf ( n2024 , R_19b4_14a10598 );
buf ( n2025 , R_1744_11c6e3d8 );
buf ( n2026 , R_757_13d3ceb8 );
buf ( n2027 , R_16fe_123b51b8 );
buf ( n2028 , R_10df_156b31f8 );
buf ( n2029 , R_ac0_123c19b8 );
buf ( n2030 , R_79d_13ddd698 );
buf ( n2031 , R_dbc_13d207d8 );
buf ( n2032 , R_13db_13d412d8 );
buf ( n2033 , R_19fa_140afeb8 );
buf ( n2034 , R_188a_14a0dd98 );
buf ( n2035 , R_126b_170193e8 );
buf ( n2036 , R_c4c_14874a18 );
buf ( n2037 , R_62d_123c23b8 );
buf ( n2038 , R_611_156aa558 );
buf ( n2039 , R_c30_13cd8158 );
buf ( n2040 , R_124f_13cd9418 );
buf ( n2041 , R_186e_1162cb38 );
buf ( n2042 , R_1233_13d5c318 );
buf ( n2043 , R_1852_11635698 );
buf ( n2044 , R_18a6_15885218 );
buf ( n2045 , R_1287_13c29e98 );
buf ( n2046 , R_c68_12fc1cd8 );
buf ( n2047 , R_649_150e1f38 );
buf ( n2048 , R_5f5_13bf7398 );
buf ( n2049 , R_c14_13defe98 );
buf ( n2050 , R_18c2_13d5d998 );
buf ( n2051 , R_bf8_13bf77f8 );
buf ( n2052 , R_12a3_14b20278 );
buf ( n2053 , R_1217_123bdd18 );
buf ( n2054 , R_c84_123bee98 );
buf ( n2055 , R_1836_14a16038 );
buf ( n2056 , R_665_117eefb8 );
buf ( n2057 , R_5d9_15fed588 );
buf ( n2058 , R_84f_1587bdf8 );
buf ( n2059 , R_148d_156b2d98 );
buf ( n2060 , R_164c_156b65d8 );
buf ( n2061 , R_a0e_13cd5098 );
buf ( n2062 , R_e6e_13c1e818 );
buf ( n2063 , R_102d_14a14878 );
buf ( n2064 , R_d7b_1007dbb8 );
buf ( n2065 , R_1120_13cd3158 );
buf ( n2066 , R_139a_12fbf398 );
buf ( n2067 , R_b01_1587af98 );
buf ( n2068 , R_19b9_116327b8 );
buf ( n2069 , R_75c_13d54b18 );
buf ( n2070 , R_173f_14a0d1b8 );
buf ( n2071 , R_ca0_117f3978 );
buf ( n2072 , R_bdc_14867a98 );
buf ( n2073 , R_11fb_13d26638 );
buf ( n2074 , R_681_13c02c58 );
buf ( n2075 , R_18de_1162c638 );
buf ( n2076 , R_181a_15887fb8 );
buf ( n2077 , R_12bf_12fbe3f8 );
buf ( n2078 , R_5bd_123b9678 );
buf ( n2079 , R_1a0e_1486b698 );
buf ( n2080 , R_13ef_156ba1d8 );
buf ( n2081 , R_dd0_12fc0798 );
buf ( n2082 , R_7b1_14a13478 );
buf ( n2083 , R_aac_116311d8 );
buf ( n2084 , R_10cb_150dccb8 );
buf ( n2085 , R_16ea_140b6cb8 );
buf ( n2086 , R_ffe_13ccf198 );
buf ( n2087 , R_e9d_13d27038 );
buf ( n2088 , R_9df_14a17398 );
buf ( n2089 , R_161d_13b962b8 );
buf ( n2090 , R_14bc_117f0598 );
buf ( n2091 , R_87e_140b08b8 );
buf ( n2092 , R_5a1_13d446b8 );
buf ( n2093 , R_cbc_12fc1b98 );
buf ( n2094 , R_bc0_13dfb338 );
buf ( n2095 , R_69d_11c69798 );
buf ( n2096 , R_18fa_140b5098 );
buf ( n2097 , R_11df_15880998 );
buf ( n2098 , R_12db_156b4af8 );
buf ( n2099 , R_17fe_1580f5f8 );
buf ( n2100 , R_191b_13c25f78 );
buf ( n2101 , R_580_1162b4b8 );
buf ( n2102 , R_6be_158101d8 );
buf ( n2103 , R_17dd_14872358 );
buf ( n2104 , R_12fc_15813dd8 );
buf ( n2105 , R_b9f_140b49b8 );
buf ( n2106 , R_cdd_13bf42d8 );
buf ( n2107 , R_11be_150e4378 );
buf ( n2108 , R_eba_13d29158 );
buf ( n2109 , R_fe1_13d2bef8 );
buf ( n2110 , R_14d9_13c21338 );
buf ( n2111 , R_9c2_116297f8 );
buf ( n2112 , R_89b_117ed118 );
buf ( n2113 , R_1600_117e96f8 );
buf ( n2114 , R_585_14a19b98 );
buf ( n2115 , R_1916_150e99b8 );
buf ( n2116 , R_17e2_123c1d78 );
buf ( n2117 , R_6b9_150dc998 );
buf ( n2118 , R_ba4_13c04d78 );
buf ( n2119 , R_12f7_117f4ff8 );
buf ( n2120 , R_11c3_117ee158 );
buf ( n2121 , R_cd8_150deab8 );
buf ( n2122 , R_15c4_13d46e18 );
buf ( n2123 , R_8d7_13de10b8 );
buf ( n2124 , R_fa5_13df4858 );
buf ( n2125 , R_ef6_13c1f358 );
buf ( n2126 , R_986_11631278 );
buf ( n2127 , R_1515_13ccb8b8 );
buf ( n2128 , R_11a7_123b9b78 );
buf ( n2129 , R_569_12fbfd98 );
buf ( n2130 , R_6d5_14b25958 );
buf ( n2131 , R_1313_1587dab8 );
buf ( n2132 , R_17c6_13d290b8 );
buf ( n2133 , R_b88_14a0d9d8 );
buf ( n2134 , R_cf4_13bea558 );
buf ( n2135 , R_1932_13cd1538 );
buf ( n2136 , R_1778_11631598 );
buf ( n2137 , R_d42_1580f918 );
buf ( n2138 , R_1159_148722b8 );
buf ( n2139 , R_1361_14a18658 );
buf ( n2140 , R_b3a_11637678 );
buf ( n2141 , R_1980_15883a58 );
buf ( n2142 , R_723_14a0aeb8 );
buf ( n2143 , R_ec5_123c1eb8 );
buf ( n2144 , R_fd6_15ff7448 );
buf ( n2145 , R_14e4_14a121b8 );
buf ( n2146 , R_9b7_117eaaf8 );
buf ( n2147 , R_8a6_156b3018 );
buf ( n2148 , R_15f5_140ade38 );
buf ( n2149 , R_d45_117f4418 );
buf ( n2150 , R_1775_140b5d18 );
buf ( n2151 , R_1364_13c1d918 );
buf ( n2152 , R_1156_15ff6fe8 );
buf ( n2153 , R_1983_100863f8 );
buf ( n2154 , R_726_13d39498 );
buf ( n2155 , R_b37_10089b98 );
buf ( n2156 , R_15e9_11636db8 );
buf ( n2157 , R_14f0_13b92398 );
buf ( n2158 , R_fca_156b44b8 );
buf ( n2159 , R_8b2_11629078 );
buf ( n2160 , R_9ab_14866698 );
buf ( n2161 , R_ed1_158870b8 );
buf ( n2162 , R_1632_117f1178 );
buf ( n2163 , R_9f4_1486d2b8 );
buf ( n2164 , R_e88_124c4498 );
buf ( n2165 , R_1013_14a135b8 );
buf ( n2166 , R_14a7_15814af8 );
buf ( n2167 , R_869_14a19e18 );
buf ( n2168 , R_132f_13c0b8f8 );
buf ( n2169 , R_6f1_150df878 );
buf ( n2170 , R_118b_14b27618 );
buf ( n2171 , R_194e_14b236f8 );
buf ( n2172 , R_d10_123b2d78 );
buf ( n2173 , R_b6c_123b8138 );
buf ( n2174 , R_17aa_13dfac58 );
buf ( n2175 , R_188b_117e9978 );
buf ( n2176 , R_126c_1580edd8 );
buf ( n2177 , R_c4d_13d24b58 );
buf ( n2178 , R_62e_13bf7438 );
buf ( n2179 , R_610_14a186f8 );
buf ( n2180 , R_c2f_14a0c038 );
buf ( n2181 , R_124e_117ee338 );
buf ( n2182 , R_186d_15fee348 );
buf ( n2183 , R_e8c_1587e738 );
buf ( n2184 , R_162e_123b25f8 );
buf ( n2185 , R_9f0_140abe58 );
buf ( n2186 , R_14ab_13dd50d8 );
buf ( n2187 , R_86d_14a18dd8 );
buf ( n2188 , R_100f_13d5dad8 );
buf ( n2189 , R_8f8_15ff8668 );
buf ( n2190 , R_f17_14a18e78 );
buf ( n2191 , R_1536_14a0dc58 );
buf ( n2192 , R_15a3_12fc08d8 );
buf ( n2193 , R_f84_117e8d98 );
buf ( n2194 , R_965_140b2578 );
buf ( n2195 , R_d71_14b23018 );
buf ( n2196 , R_b0b_13c21e78 );
buf ( n2197 , R_1390_17016a08 );
buf ( n2198 , R_19af_11636458 );
buf ( n2199 , R_1749_117ec178 );
buf ( n2200 , R_752_15ff64a8 );
buf ( n2201 , R_112a_1587e0f8 );
buf ( n2202 , R_18b6_13bf3018 );
buf ( n2203 , R_1223_13dd8418 );
buf ( n2204 , R_1297_13b99738 );
buf ( n2205 , R_1842_123b43f8 );
buf ( n2206 , R_c78_15887018 );
buf ( n2207 , R_659_123b34f8 );
buf ( n2208 , R_5e5_13df0578 );
buf ( n2209 , R_c04_13cd6f38 );
buf ( n2210 , R_954_17014988 );
buf ( n2211 , R_909_13d3efd8 );
buf ( n2212 , R_f28_13bf6fd8 );
buf ( n2213 , R_1547_13df7b98 );
buf ( n2214 , R_1592_156b9918 );
buf ( n2215 , R_f73_13d22a38 );
buf ( n2216 , R_70d_13beb098 );
buf ( n2217 , R_178e_13c1cb58 );
buf ( n2218 , R_196a_156b6d58 );
buf ( n2219 , R_d2c_14a0ec98 );
buf ( n2220 , R_116f_13d3e7b8 );
buf ( n2221 , R_134b_15ff6cc8 );
buf ( n2222 , R_b50_15815598 );
buf ( n2223 , R_caf_156adc58 );
buf ( n2224 , R_bcd_1162baf8 );
buf ( n2225 , R_690_13c1e098 );
buf ( n2226 , R_18ed_124c3278 );
buf ( n2227 , R_11ec_1008d0b8 );
buf ( n2228 , R_12ce_13c071b8 );
buf ( n2229 , R_180b_1008abd8 );
buf ( n2230 , R_5ae_13cd7ed8 );
buf ( n2231 , R_177b_1007d6b8 );
buf ( n2232 , R_d3f_13cd10d8 );
buf ( n2233 , R_115c_150e8f18 );
buf ( n2234 , R_135e_11c696f8 );
buf ( n2235 , R_b3d_13dddeb8 );
buf ( n2236 , R_720_13d395d8 );
buf ( n2237 , R_197d_14a15458 );
buf ( n2238 , R_1700_140ae8d8 );
buf ( n2239 , R_10e1_13c07758 );
buf ( n2240 , R_ac2_156ad2f8 );
buf ( n2241 , R_79b_15886398 );
buf ( n2242 , R_dba_116373f8 );
buf ( n2243 , R_13d9_14a14378 );
buf ( n2244 , R_19f8_117ef558 );
buf ( n2245 , R_595_13def178 );
buf ( n2246 , R_17f2_1580c998 );
buf ( n2247 , R_1906_13ccad78 );
buf ( n2248 , R_6a9_15ff4ba8 );
buf ( n2249 , R_bb4_117f4d78 );
buf ( n2250 , R_12e7_13cd42d8 );
buf ( n2251 , R_11d3_1162b0f8 );
buf ( n2252 , R_cc8_123b7738 );
buf ( n2253 , R_d48_13c21c98 );
buf ( n2254 , R_1772_14a16998 );
buf ( n2255 , R_1367_15880858 );
buf ( n2256 , R_1153_117f1678 );
buf ( n2257 , R_1986_11c6c038 );
buf ( n2258 , R_729_117f72f8 );
buf ( n2259 , R_b34_158825b8 );
buf ( n2260 , R_ff5_13c2a618 );
buf ( n2261 , R_ea6_150dd7f8 );
buf ( n2262 , R_9d6_13c01f38 );
buf ( n2263 , R_14c5_14a0e518 );
buf ( n2264 , R_1614_156b2b18 );
buf ( n2265 , R_887_14a18298 );
buf ( n2266 , R_848_13ddf218 );
buf ( n2267 , R_1653_14869438 );
buf ( n2268 , R_1486_156afe18 );
buf ( n2269 , R_a15_1700ed08 );
buf ( n2270 , R_e67_117f4e18 );
buf ( n2271 , R_1034_156ac5d8 );
buf ( n2272 , R_8eb_150db1d8 );
buf ( n2273 , R_15b0_1580bdb8 );
buf ( n2274 , R_f0a_14a0ce98 );
buf ( n2275 , R_f91_117f6f38 );
buf ( n2276 , R_1529_123bca58 );
buf ( n2277 , R_972_13ccc038 );
buf ( n2278 , R_1a10_123b4718 );
buf ( n2279 , R_13f1_13d24298 );
buf ( n2280 , R_dd2_14a19198 );
buf ( n2281 , R_7b3_13c07938 );
buf ( n2282 , R_aaa_13b8cfd8 );
buf ( n2283 , R_10c9_15812a78 );
buf ( n2284 , R_16e8_13cd8d38 );
buf ( n2285 , R_d64_15ff5968 );
buf ( n2286 , R_b18_117f40f8 );
buf ( n2287 , R_1383_13c2a438 );
buf ( n2288 , R_19a2_117f01d8 );
buf ( n2289 , R_1756_123c0f18 );
buf ( n2290 , R_1137_13d20ff8 );
buf ( n2291 , R_745_13c1d5f8 );
buf ( n2292 , R_1636_14b22618 );
buf ( n2293 , R_9f8_13decdd8 );
buf ( n2294 , R_e84_14875b98 );
buf ( n2295 , R_1017_13d3bbf8 );
buf ( n2296 , R_865_13d4e7b8 );
buf ( n2297 , R_14a3_11c6d078 );
buf ( n2298 , R_83e_13d43ad8 );
buf ( n2299 , R_a1f_13d22d58 );
buf ( n2300 , R_147c_1580d398 );
buf ( n2301 , R_103e_13d57958 );
buf ( n2302 , R_e5d_1486ddf8 );
buf ( n2303 , R_165d_13bec038 );
buf ( n2304 , R_1494_117f6718 );
buf ( n2305 , R_1645_11c6c178 );
buf ( n2306 , R_a07_14b251d8 );
buf ( n2307 , R_e75_1580a5f8 );
buf ( n2308 , R_1026_158103b8 );
buf ( n2309 , R_856_13cd2a78 );
buf ( n2310 , R_188c_13d39ad8 );
buf ( n2311 , R_126d_11636638 );
buf ( n2312 , R_c4e_13c0fe58 );
buf ( n2313 , R_62f_116305f8 );
buf ( n2314 , R_60f_13bf44b8 );
buf ( n2315 , R_c2e_156b6c18 );
buf ( n2316 , R_124d_123b5438 );
buf ( n2317 , R_186c_15817758 );
buf ( n2318 , R_57b_12fc1f58 );
buf ( n2319 , R_6c3_14a11718 );
buf ( n2320 , R_17d8_13bf24d8 );
buf ( n2321 , R_1301_13ccee78 );
buf ( n2322 , R_b9a_140b40f8 );
buf ( n2323 , R_ce2_156b49b8 );
buf ( n2324 , R_11b9_13d5d5d8 );
buf ( n2325 , R_1920_117ea198 );
buf ( n2326 , R_1713_14a0f878 );
buf ( n2327 , R_10f4_13de4c18 );
buf ( n2328 , R_ad5_117ed1b8 );
buf ( n2329 , R_788_117e8ed8 );
buf ( n2330 , R_da7_11635ff8 );
buf ( n2331 , R_13c6_123c10f8 );
buf ( n2332 , R_19e5_1580eb58 );
buf ( n2333 , R_e90_11637038 );
buf ( n2334 , R_9ec_117eb958 );
buf ( n2335 , R_162a_117ec0d8 );
buf ( n2336 , R_14af_156abdb8 );
buf ( n2337 , R_871_1587f138 );
buf ( n2338 , R_100b_11631d18 );
buf ( n2339 , R_111b_1580faf8 );
buf ( n2340 , R_139f_150df058 );
buf ( n2341 , R_afc_117f8158 );
buf ( n2342 , R_19be_13ccfff8 );
buf ( n2343 , R_761_12fbf078 );
buf ( n2344 , R_173a_156b5a98 );
buf ( n2345 , R_d80_13c1d418 );
buf ( n2346 , R_58a_13ddaf38 );
buf ( n2347 , R_1911_124c4038 );
buf ( n2348 , R_17e7_15883198 );
buf ( n2349 , R_6b4_15881bb8 );
buf ( n2350 , R_ba9_13d5c958 );
buf ( n2351 , R_12f2_17013c68 );
buf ( n2352 , R_11c8_11634fb8 );
buf ( n2353 , R_cd3_13c06178 );
buf ( n2354 , R_6fc_13de34f8 );
buf ( n2355 , R_1180_13ddc298 );
buf ( n2356 , R_1959_14a14698 );
buf ( n2357 , R_d1b_13cd9558 );
buf ( n2358 , R_b61_13d22538 );
buf ( n2359 , R_179f_150e5818 );
buf ( n2360 , R_133a_13d57138 );
buf ( n2361 , R_be4_15817bb8 );
buf ( n2362 , R_c98_13dec298 );
buf ( n2363 , R_1203_1587d978 );
buf ( n2364 , R_679_123b7918 );
buf ( n2365 , R_1822_117e9018 );
buf ( n2366 , R_18d6_13c2ad98 );
buf ( n2367 , R_5c5_1162b5f8 );
buf ( n2368 , R_12b7_117f83d8 );
buf ( n2369 , R_ca8_14a11038 );
buf ( n2370 , R_bd4_11637ad8 );
buf ( n2371 , R_689_158869d8 );
buf ( n2372 , R_11f3_116300f8 );
buf ( n2373 , R_18e6_156b1678 );
buf ( n2374 , R_1812_11c6f558 );
buf ( n2375 , R_12c7_13b97c58 );
buf ( n2376 , R_5b5_11637fd8 );
buf ( n2377 , R_177e_14b1a738 );
buf ( n2378 , R_d3c_13b8b278 );
buf ( n2379 , R_115f_156ac7b8 );
buf ( n2380 , R_135b_13d38b38 );
buf ( n2381 , R_b40_158142d8 );
buf ( n2382 , R_71d_13c1ea98 );
buf ( n2383 , R_197a_13c0a318 );
buf ( n2384 , R_e16_17018088 );
buf ( n2385 , R_1085_13c03e78 );
buf ( n2386 , R_7f7_15888b98 );
buf ( n2387 , R_16a4_158821f8 );
buf ( n2388 , R_1a54_13de0438 );
buf ( n2389 , R_1435_10082258 );
buf ( n2390 , R_a66_15882838 );
buf ( n2391 , R_703_14867bd8 );
buf ( n2392 , R_1960_1162c958 );
buf ( n2393 , R_1179_13d3c7d8 );
buf ( n2394 , R_d22_13d599d8 );
buf ( n2395 , R_b5a_13bf68f8 );
buf ( n2396 , R_1341_13d458d8 );
buf ( n2397 , R_1798_1700e9e8 );
buf ( n2398 , R_171e_13df60b8 );
buf ( n2399 , R_10ff_13ddcab8 );
buf ( n2400 , R_ae0_14a11f38 );
buf ( n2401 , R_77d_13d27df8 );
buf ( n2402 , R_d9c_13ccd4d8 );
buf ( n2403 , R_13bb_1587d478 );
buf ( n2404 , R_19da_13dd5a38 );
buf ( n2405 , R_108a_1486e938 );
buf ( n2406 , R_e11_13cd8c98 );
buf ( n2407 , R_16a9_14a130b8 );
buf ( n2408 , R_7f2_156b2938 );
buf ( n2409 , R_1a4f_13d3a618 );
buf ( n2410 , R_a6b_13b8e1f8 );
buf ( n2411 , R_1430_13dd84b8 );
buf ( n2412 , R_d4b_117f6178 );
buf ( n2413 , R_176f_13d447f8 );
buf ( n2414 , R_136a_13c26838 );
buf ( n2415 , R_1150_15ff71c8 );
buf ( n2416 , R_1989_13ccbc78 );
buf ( n2417 , R_72c_10083c98 );
buf ( n2418 , R_b31_13d44c58 );
buf ( n2419 , R_814_13d51eb8 );
buf ( n2420 , R_1068_1580ea18 );
buf ( n2421 , R_1687_123b81d8 );
buf ( n2422 , R_1452_13df0938 );
buf ( n2423 , R_e33_14a0c3f8 );
buf ( n2424 , R_a49_14a0eb58 );
buf ( n2425 , R_1851_13d5b058 );
buf ( n2426 , R_18a7_13b96858 );
buf ( n2427 , R_1288_13c1daf8 );
buf ( n2428 , R_c69_156af738 );
buf ( n2429 , R_64a_11629438 );
buf ( n2430 , R_5f4_140b13f8 );
buf ( n2431 , R_c13_1162db78 );
buf ( n2432 , R_1232_156aaa58 );
buf ( n2433 , R_15bb_117f3338 );
buf ( n2434 , R_8e0_14a0f698 );
buf ( n2435 , R_f9c_14a104f8 );
buf ( n2436 , R_eff_13d381d8 );
buf ( n2437 , R_151e_15883af8 );
buf ( n2438 , R_97d_14a16178 );
buf ( n2439 , R_1702_13cd9198 );
buf ( n2440 , R_10e3_117f2f78 );
buf ( n2441 , R_ac4_1700f028 );
buf ( n2442 , R_799_13d5a018 );
buf ( n2443 , R_db8_150e6998 );
buf ( n2444 , R_13d7_14b1d1b8 );
buf ( n2445 , R_19f6_1580aa58 );
buf ( n2446 , R_14fd_156b56d8 );
buf ( n2447 , R_15dc_123bfd98 );
buf ( n2448 , R_fbd_14a0b098 );
buf ( n2449 , R_8bf_14875f58 );
buf ( n2450 , R_99e_15ff9388 );
buf ( n2451 , R_ede_11634338 );
buf ( n2452 , R_188d_17018e48 );
buf ( n2453 , R_126e_150e04f8 );
buf ( n2454 , R_c4f_15814918 );
buf ( n2455 , R_630_13d25558 );
buf ( n2456 , R_60e_13cd3d38 );
buf ( n2457 , R_c2d_1580aaf8 );
buf ( n2458 , R_124c_13d40018 );
buf ( n2459 , R_186b_13d42bd8 );
buf ( n2460 , R_1a23_13d52458 );
buf ( n2461 , R_1404_1486a8d8 );
buf ( n2462 , R_de5_11633a78 );
buf ( n2463 , R_7c6_156b9738 );
buf ( n2464 , R_a97_13c05e58 );
buf ( n2465 , R_10b6_124c3638 );
buf ( n2466 , R_16d5_123bc4b8 );
buf ( n2467 , R_bed_13b90db8 );
buf ( n2468 , R_c8f_117ef4b8 );
buf ( n2469 , R_120c_13ddcd38 );
buf ( n2470 , R_670_13ccfaf8 );
buf ( n2471 , R_182b_13cd80b8 );
buf ( n2472 , R_18cd_13c1ca18 );
buf ( n2473 , R_5ce_14b1ded8 );
buf ( n2474 , R_12ae_13c1f178 );
buf ( n2475 , R_bc6_13cd7bb8 );
buf ( n2476 , R_697_13bf83d8 );
buf ( n2477 , R_18f4_15881cf8 );
buf ( n2478 , R_11e5_1162add8 );
buf ( n2479 , R_12d5_17015928 );
buf ( n2480 , R_1804_150e44b8 );
buf ( n2481 , R_5a7_12fbe178 );
buf ( n2482 , R_cb6_1162e398 );
buf ( n2483 , R_110f_15887518 );
buf ( n2484 , R_19ca_156b8a18 );
buf ( n2485 , R_af0_17012a48 );
buf ( n2486 , R_76d_156b1df8 );
buf ( n2487 , R_d8c_15814b98 );
buf ( n2488 , R_172e_117ed438 );
buf ( n2489 , R_13ab_13b99878 );
buf ( n2490 , R_1a12_13d52ef8 );
buf ( n2491 , R_13f3_156b74d8 );
buf ( n2492 , R_dd4_140ac5d8 );
buf ( n2493 , R_7b5_13c1f718 );
buf ( n2494 , R_aa8_14a0ea18 );
buf ( n2495 , R_10c7_13df2c38 );
buf ( n2496 , R_16e6_156b9eb8 );
buf ( n2497 , R_15cd_13cd86f8 );
buf ( n2498 , R_8ce_13d1e2f8 );
buf ( n2499 , R_fae_13bf6df8 );
buf ( n2500 , R_eed_15812578 );
buf ( n2501 , R_98f_117f62b8 );
buf ( n2502 , R_150c_15ff3848 );
buf ( n2503 , R_908_123c0658 );
buf ( n2504 , R_f27_13cd08b8 );
buf ( n2505 , R_1546_14a18f18 );
buf ( n2506 , R_1593_13d58e98 );
buf ( n2507 , R_f74_158805d8 );
buf ( n2508 , R_955_1580f0f8 );
buf ( n2509 , R_d5c_1580ed38 );
buf ( n2510 , R_137b_13d5cc78 );
buf ( n2511 , R_175e_15813478 );
buf ( n2512 , R_199a_117e8b18 );
buf ( n2513 , R_113f_123b3098 );
buf ( n2514 , R_73d_13c220f8 );
buf ( n2515 , R_b20_13c06c18 );
buf ( n2516 , R_163a_13d3ddb8 );
buf ( n2517 , R_9fc_14a0b818 );
buf ( n2518 , R_e80_11633ed8 );
buf ( n2519 , R_101b_123b6518 );
buf ( n2520 , R_861_124c3bd8 );
buf ( n2521 , R_149f_123b5e38 );
buf ( n2522 , R_1080_14a149b8 );
buf ( n2523 , R_7fc_13d3f258 );
buf ( n2524 , R_169f_124c2d78 );
buf ( n2525 , R_1a59_117eded8 );
buf ( n2526 , R_143a_14a0edd8 );
buf ( n2527 , R_a61_1700dd68 );
buf ( n2528 , R_e1b_13cd1178 );
buf ( n2529 , R_140f_117f1cb8 );
buf ( n2530 , R_df0_13c09cd8 );
buf ( n2531 , R_7d1_14b28978 );
buf ( n2532 , R_a8c_123c0338 );
buf ( n2533 , R_10ab_13df0398 );
buf ( n2534 , R_16ca_13d52f98 );
buf ( n2535 , R_1a2e_13c22698 );
buf ( n2536 , R_b10_14b21fd8 );
buf ( n2537 , R_138b_156b0318 );
buf ( n2538 , R_19aa_14a194b8 );
buf ( n2539 , R_174e_15811a38 );
buf ( n2540 , R_74d_117f0e58 );
buf ( n2541 , R_112f_156aac38 );
buf ( n2542 , R_d6c_156b62b8 );
buf ( n2543 , R_1781_1162d5d8 );
buf ( n2544 , R_d39_15811b78 );
buf ( n2545 , R_1162_124c2558 );
buf ( n2546 , R_1358_156b8e78 );
buf ( n2547 , R_b43_13c06858 );
buf ( n2548 , R_71a_117ee798 );
buf ( n2549 , R_1977_15880b78 );
buf ( n2550 , R_1108_13ccfb98 );
buf ( n2551 , R_ae9_1580cd58 );
buf ( n2552 , R_774_1700a7a8 );
buf ( n2553 , R_d93_13cce0b8 );
buf ( n2554 , R_13b2_15886898 );
buf ( n2555 , R_1727_14870e18 );
buf ( n2556 , R_19d1_123b5b18 );
buf ( n2557 , R_188e_11c6a698 );
buf ( n2558 , R_126f_14b23c98 );
buf ( n2559 , R_c50_13d471d8 );
buf ( n2560 , R_631_13ddd7d8 );
buf ( n2561 , R_60d_117f3a18 );
buf ( n2562 , R_c2c_13d2c498 );
buf ( n2563 , R_124b_156b97d8 );
buf ( n2564 , R_186a_13ddb118 );
buf ( n2565 , R_fdc_1162ca98 );
buf ( n2566 , R_14de_13c202f8 );
buf ( n2567 , R_9bd_11632cb8 );
buf ( n2568 , R_8a0_13bf81f8 );
buf ( n2569 , R_15fb_123ba078 );
buf ( n2570 , R_ebf_13b91678 );
buf ( n2571 , R_e94_148719f8 );
buf ( n2572 , R_9e8_15ff97e8 );
buf ( n2573 , R_1626_13de2918 );
buf ( n2574 , R_14b3_13dde9f8 );
buf ( n2575 , R_875_156aea18 );
buf ( n2576 , R_1007_15881578 );
buf ( n2577 , R_14f6_11638938 );
buf ( n2578 , R_fc4_1580d578 );
buf ( n2579 , R_8b8_123ba2f8 );
buf ( n2580 , R_9a5_117ecc18 );
buf ( n2581 , R_ed7_14a0da78 );
buf ( n2582 , R_15e3_123c0158 );
buf ( n2583 , R_e0c_1700d0e8 );
buf ( n2584 , R_16ae_123b38b8 );
buf ( n2585 , R_7ed_117ef738 );
buf ( n2586 , R_1a4a_12fc1c38 );
buf ( n2587 , R_a70_150dbc78 );
buf ( n2588 , R_142b_15889bd8 );
buf ( n2589 , R_108f_13de36d8 );
buf ( n2590 , R_d4e_11c6b6d8 );
buf ( n2591 , R_176c_13ddfcb8 );
buf ( n2592 , R_136d_11634dd8 );
buf ( n2593 , R_114d_158861b8 );
buf ( n2594 , R_198c_13d53a38 );
buf ( n2595 , R_72f_11637498 );
buf ( n2596 , R_b2e_170098a8 );
buf ( n2597 , R_8f7_13b8e298 );
buf ( n2598 , R_f16_1587d838 );
buf ( n2599 , R_1535_13ded2d8 );
buf ( n2600 , R_15a4_1162bcd8 );
buf ( n2601 , R_f85_170174a8 );
buf ( n2602 , R_966_156acd58 );
buf ( n2603 , R_12a4_13cd0db8 );
buf ( n2604 , R_1216_13c26518 );
buf ( n2605 , R_c85_13d505b8 );
buf ( n2606 , R_1835_13b8eb58 );
buf ( n2607 , R_666_13cd8798 );
buf ( n2608 , R_5d8_14a11fd8 );
buf ( n2609 , R_18c3_156b8c98 );
buf ( n2610 , R_bf7_156b4418 );
buf ( n2611 , R_15d5_117ed898 );
buf ( n2612 , R_fb6_14b24558 );
buf ( n2613 , R_8c6_13d442f8 );
buf ( n2614 , R_997_123bb478 );
buf ( n2615 , R_ee5_14a14af8 );
buf ( n2616 , R_1504_13d553d8 );
buf ( n2617 , R_6d1_158167b8 );
buf ( n2618 , R_130f_156ab4f8 );
buf ( n2619 , R_17ca_150df9b8 );
buf ( n2620 , R_b8c_124c3ef8 );
buf ( n2621 , R_cf0_11c6a878 );
buf ( n2622 , R_192e_150e8a18 );
buf ( n2623 , R_11ab_13d29d38 );
buf ( n2624 , R_56d_156b76b8 );
buf ( n2625 , R_1704_13bf4238 );
buf ( n2626 , R_10e5_14871778 );
buf ( n2627 , R_ac6_1587bcb8 );
buf ( n2628 , R_797_14b1c178 );
buf ( n2629 , R_db6_13ddd058 );
buf ( n2630 , R_13d5_1587c618 );
buf ( n2631 , R_19f4_150e3ab8 );
buf ( n2632 , R_1298_156b1d58 );
buf ( n2633 , R_1841_13d2c538 );
buf ( n2634 , R_c79_156b5598 );
buf ( n2635 , R_65a_14874ab8 );
buf ( n2636 , R_5e4_13bf0278 );
buf ( n2637 , R_c03_14a0d2f8 );
buf ( n2638 , R_18b7_13ccd1b8 );
buf ( n2639 , R_1222_14b1acd8 );
buf ( n2640 , R_1073_14b20f98 );
buf ( n2641 , R_809_13d3e678 );
buf ( n2642 , R_1a66_123b6158 );
buf ( n2643 , R_1692_117f31f8 );
buf ( n2644 , R_1447_13b93338 );
buf ( n2645 , R_e28_156abbd8 );
buf ( n2646 , R_a54_13cce838 );
buf ( n2647 , R_1054_13bf8ab8 );
buf ( n2648 , R_1466_13d5abf8 );
buf ( n2649 , R_1673_1580e798 );
buf ( n2650 , R_e47_1587b178 );
buf ( n2651 , R_a35_117f5db8 );
buf ( n2652 , R_828_10081f38 );
buf ( n2653 , R_1469_1587ee18 );
buf ( n2654 , R_1051_11635c38 );
buf ( n2655 , R_e4a_11629118 );
buf ( n2656 , R_1670_1007f238 );
buf ( n2657 , R_82b_13cd7258 );
buf ( n2658 , R_a32_1486afb8 );
buf ( n2659 , R_1187_117f4198 );
buf ( n2660 , R_1952_14a0c0d8 );
buf ( n2661 , R_d14_13dee778 );
buf ( n2662 , R_b68_10089d78 );
buf ( n2663 , R_17a6_15811f38 );
buf ( n2664 , R_1333_117f21b8 );
buf ( n2665 , R_6f5_13d43678 );
buf ( n2666 , R_6c8_1580d758 );
buf ( n2667 , R_1306_1580d938 );
buf ( n2668 , R_17d3_13d3a578 );
buf ( n2669 , R_b95_117f7618 );
buf ( n2670 , R_ce7_13d27218 );
buf ( n2671 , R_1925_15ff0328 );
buf ( n2672 , R_11b4_13b8ec98 );
buf ( n2673 , R_576_13d2bf98 );
buf ( n2674 , R_e00_13cd8bf8 );
buf ( n2675 , R_7e1_150e4058 );
buf ( n2676 , R_a7c_156b7118 );
buf ( n2677 , R_1a3e_14a0b278 );
buf ( n2678 , R_109b_123bd4f8 );
buf ( n2679 , R_141f_1008c578 );
buf ( n2680 , R_16ba_156b6e98 );
buf ( n2681 , R_188f_156b5458 );
buf ( n2682 , R_1270_14a103b8 );
buf ( n2683 , R_c51_11630af8 );
buf ( n2684 , R_632_13ccde38 );
buf ( n2685 , R_60c_13dd9c78 );
buf ( n2686 , R_c2b_14b23478 );
buf ( n2687 , R_124a_140b7898 );
buf ( n2688 , R_1869_14b29cd8 );
buf ( n2689 , R_1a14_117ebbd8 );
buf ( n2690 , R_13f5_13cd8a18 );
buf ( n2691 , R_dd6_13de0d98 );
buf ( n2692 , R_7b7_15816a38 );
buf ( n2693 , R_aa6_13d28c58 );
buf ( n2694 , R_10c5_11632998 );
buf ( n2695 , R_16e4_10087078 );
buf ( n2696 , R_190c_13d1d998 );
buf ( n2697 , R_6af_124c33b8 );
buf ( n2698 , R_bae_1587b5d8 );
buf ( n2699 , R_12ed_14a176b8 );
buf ( n2700 , R_11cd_13cd27f8 );
buf ( n2701 , R_cce_116331b8 );
buf ( n2702 , R_58f_156b9558 );
buf ( n2703 , R_17ec_13dd7fb8 );
buf ( n2704 , R_1057_123bd278 );
buf ( n2705 , R_1463_124c4b78 );
buf ( n2706 , R_1676_140ae6f8 );
buf ( n2707 , R_e44_148741f8 );
buf ( n2708 , R_a38_150dc3f8 );
buf ( n2709 , R_825_123b3278 );
buf ( n2710 , R_18a8_1580c8f8 );
buf ( n2711 , R_1289_13c09738 );
buf ( n2712 , R_c6a_15811fd8 );
buf ( n2713 , R_64b_1007d938 );
buf ( n2714 , R_5f3_116307d8 );
buf ( n2715 , R_c12_1162cc78 );
buf ( n2716 , R_1231_13dee9f8 );
buf ( n2717 , R_1850_1587f778 );
buf ( n2718 , R_146c_14872f38 );
buf ( n2719 , R_104e_1580f7d8 );
buf ( n2720 , R_e4d_14b20d18 );
buf ( n2721 , R_166d_13d20058 );
buf ( n2722 , R_82e_1580f2d8 );
buf ( n2723 , R_a2f_123b3db8 );
buf ( n2724 , R_19c3_116340b8 );
buf ( n2725 , R_af7_13cd2d98 );
buf ( n2726 , R_766_13c07618 );
buf ( n2727 , R_1735_13bf9f58 );
buf ( n2728 , R_d85_13dd7518 );
buf ( n2729 , R_13a4_150ea138 );
buf ( n2730 , R_1116_13c02438 );
buf ( n2731 , R_df9_13dd9458 );
buf ( n2732 , R_7da_14a16fd8 );
buf ( n2733 , R_a83_13b9a278 );
buf ( n2734 , R_10a2_123b3d18 );
buf ( n2735 , R_1a37_1587f958 );
buf ( n2736 , R_16c1_13d3d458 );
buf ( n2737 , R_1418_13d2b1d8 );
buf ( n2738 , R_ea1_156b5c78 );
buf ( n2739 , R_9db_13c05bd8 );
buf ( n2740 , R_1619_15888d78 );
buf ( n2741 , R_14c0_17012fe8 );
buf ( n2742 , R_882_13dee458 );
buf ( n2743 , R_ffa_11c68f78 );
buf ( n2744 , R_1967_15ff9608 );
buf ( n2745 , R_1172_170122c8 );
buf ( n2746 , R_d29_13bed898 );
buf ( n2747 , R_1348_156b1178 );
buf ( n2748 , R_b53_1162fe78 );
buf ( n2749 , R_1791_15ff73a8 );
buf ( n2750 , R_70a_13dee818 );
buf ( n2751 , R_8ea_13b91c18 );
buf ( n2752 , R_15b1_140b0d18 );
buf ( n2753 , R_f09_13d4f9d8 );
buf ( n2754 , R_f92_13b99238 );
buf ( n2755 , R_1528_13cca918 );
buf ( n2756 , R_973_12fc1738 );
buf ( n2757 , R_907_13d1cef8 );
buf ( n2758 , R_f26_13d51378 );
buf ( n2759 , R_1545_13ddab78 );
buf ( n2760 , R_1594_123b52f8 );
buf ( n2761 , R_f75_1587ec38 );
buf ( n2762 , R_956_117f3bf8 );
buf ( n2763 , R_a1c_13d42098 );
buf ( n2764 , R_147f_15ffd208 );
buf ( n2765 , R_103b_12fbfbb8 );
buf ( n2766 , R_e60_13b98dd8 );
buf ( n2767 , R_165a_156b9418 );
buf ( n2768 , R_841_13de1e78 );
buf ( n2769 , R_1715_13c03ab8 );
buf ( n2770 , R_10f6_1587fc78 );
buf ( n2771 , R_ad7_11c6aaf8 );
buf ( n2772 , R_786_13bf7938 );
buf ( n2773 , R_da5_13c24c18 );
buf ( n2774 , R_13c4_156adbb8 );
buf ( n2775 , R_19e3_13b8b4f8 );
buf ( n2776 , R_15c5_13cce478 );
buf ( n2777 , R_8d6_14a156d8 );
buf ( n2778 , R_fa6_13ccd7f8 );
buf ( n2779 , R_ef5_13c0f8b8 );
buf ( n2780 , R_987_148737f8 );
buf ( n2781 , R_1514_13d4ea38 );
buf ( n2782 , R_d36_13cd2938 );
buf ( n2783 , R_1165_1700dae8 );
buf ( n2784 , R_1355_13c0e2d8 );
buf ( n2785 , R_b46_12fbedf8 );
buf ( n2786 , R_717_13c1ebd8 );
buf ( n2787 , R_1974_13b938d8 );
buf ( n2788 , R_1784_14b1b3b8 );
buf ( n2789 , R_156d_13b91d58 );
buf ( n2790 , R_f4e_13d2bb38 );
buf ( n2791 , R_156c_1486f8d8 );
buf ( n2792 , R_92f_1587e418 );
buf ( n2793 , R_f4d_158174d8 );
buf ( n2794 , R_92e_15880df8 );
buf ( n2795 , R_156e_13bee0b8 );
buf ( n2796 , R_f4f_13d1f298 );
buf ( n2797 , R_930_117f5818 );
buf ( n2798 , R_156b_13cd6a38 );
buf ( n2799 , R_f4c_13d4edf8 );
buf ( n2800 , R_92d_13b93838 );
buf ( n2801 , R_156f_1700c828 );
buf ( n2802 , R_f50_13d5d038 );
buf ( n2803 , R_931_1007f198 );
buf ( n2804 , R_92c_13bef238 );
buf ( n2805 , R_156a_14a0d7f8 );
buf ( n2806 , R_f4b_1162df38 );
buf ( n2807 , R_682_13dd6a78 );
buf ( n2808 , R_11fa_12fbfe38 );
buf ( n2809 , R_18df_1162e1b8 );
buf ( n2810 , R_1819_117f44b8 );
buf ( n2811 , R_12c0_156b3478 );
buf ( n2812 , R_5bc_150db098 );
buf ( n2813 , R_ca1_15888af8 );
buf ( n2814 , R_bdb_123b9178 );
buf ( n2815 , R_1890_13c0a4f8 );
buf ( n2816 , R_1271_13cd3e78 );
buf ( n2817 , R_c52_11629cf8 );
buf ( n2818 , R_633_1587c6b8 );
buf ( n2819 , R_60b_17014c08 );
buf ( n2820 , R_c2a_13c01d58 );
buf ( n2821 , R_1249_150de798 );
buf ( n2822 , R_1868_13cd62b8 );
buf ( n2823 , R_105a_14a112b8 );
buf ( n2824 , R_1460_158862f8 );
buf ( n2825 , R_1679_13cd44b8 );
buf ( n2826 , R_e41_14a14e18 );
buf ( n2827 , R_a3b_13cd1998 );
buf ( n2828 , R_822_117e9158 );
buf ( n2829 , R_1570_13d44118 );
buf ( n2830 , R_f51_13ccb778 );
buf ( n2831 , R_932_15810d18 );
buf ( n2832 , R_92b_14a180b8 );
buf ( n2833 , R_f4a_1162c8b8 );
buf ( n2834 , R_1569_13bede38 );
buf ( n2835 , R_163e_12fc0338 );
buf ( n2836 , R_a00_13df4df8 );
buf ( n2837 , R_e7c_13c08798 );
buf ( n2838 , R_101f_117ed9d8 );
buf ( n2839 , R_85d_117f4738 );
buf ( n2840 , R_149b_13cd1038 );
buf ( n2841 , R_146f_117f47d8 );
buf ( n2842 , R_104b_158885f8 );
buf ( n2843 , R_e50_12fbe858 );
buf ( n2844 , R_166a_1587c938 );
buf ( n2845 , R_831_156b2398 );
buf ( n2846 , R_a2c_11c701d8 );
buf ( n2847 , R_801_150e6e98 );
buf ( n2848 , R_169a_13b94878 );
buf ( n2849 , R_1a5e_1162d3f8 );
buf ( n2850 , R_143f_13b8c218 );
buf ( n2851 , R_a5c_13b8c178 );
buf ( n2852 , R_e20_13ddd0f8 );
buf ( n2853 , R_107b_156b2118 );
buf ( n2854 , R_d51_13df3b38 );
buf ( n2855 , R_1769_14b21038 );
buf ( n2856 , R_1370_13cd2618 );
buf ( n2857 , R_114a_13c218d8 );
buf ( n2858 , R_198f_13d28bb8 );
buf ( n2859 , R_732_13d55fb8 );
buf ( n2860 , R_b2b_13ccd2f8 );
buf ( n2861 , R_1571_1580af58 );
buf ( n2862 , R_f52_12fc1ff8 );
buf ( n2863 , R_933_14868718 );
buf ( n2864 , R_92a_13c01a38 );
buf ( n2865 , R_f49_13d4f4d8 );
buf ( n2866 , R_1568_1580c218 );
buf ( n2867 , R_1706_15814eb8 );
buf ( n2868 , R_10e7_14a160d8 );
buf ( n2869 , R_ac8_156afa58 );
buf ( n2870 , R_795_14a12b18 );
buf ( n2871 , R_db4_117edd98 );
buf ( n2872 , R_13d3_13b90f98 );
buf ( n2873 , R_19f2_12fbf258 );
buf ( n2874 , R_17b9_156b0b38 );
buf ( n2875 , R_193f_13d3aa78 );
buf ( n2876 , R_b7b_13befeb8 );
buf ( n2877 , R_d01_140ab318 );
buf ( n2878 , R_119a_13b8a5f8 );
buf ( n2879 , R_1320_14b27f78 );
buf ( n2880 , R_55c_11630e18 );
buf ( n2881 , R_6e2_158149b8 );
buf ( n2882 , R_106b_117f3518 );
buf ( n2883 , R_168a_117eb598 );
buf ( n2884 , R_144f_14b26718 );
buf ( n2885 , R_e30_123b3e58 );
buf ( n2886 , R_a4c_170172c8 );
buf ( n2887 , R_811_15882478 );
buf ( n2888 , R_1406_148665f8 );
buf ( n2889 , R_de7_1007fcd8 );
buf ( n2890 , R_7c8_156b7f78 );
buf ( n2891 , R_a95_117f6cb8 );
buf ( n2892 , R_10b4_13d3d598 );
buf ( n2893 , R_16d3_1700be28 );
buf ( n2894 , R_1a25_13b9a318 );
buf ( n2895 , R_1572_156b67b8 );
buf ( n2896 , R_f53_123c01f8 );
buf ( n2897 , R_934_156b0958 );
buf ( n2898 , R_929_13d5bf58 );
buf ( n2899 , R_f48_13c256b8 );
buf ( n2900 , R_1567_13b91e98 );
buf ( n2901 , R_1943_11c70598 );
buf ( n2902 , R_d05_13c0cd98 );
buf ( n2903 , R_b77_13d415f8 );
buf ( n2904 , R_17b5_14a12118 );
buf ( n2905 , R_1324_15887298 );
buf ( n2906 , R_6e6_13becb78 );
buf ( n2907 , R_558_116299d8 );
buf ( n2908 , R_1196_13d4f398 );
buf ( n2909 , R_e98_13d433f8 );
buf ( n2910 , R_9e4_13cccdf8 );
buf ( n2911 , R_1622_13c044b8 );
buf ( n2912 , R_14b7_13d21318 );
buf ( n2913 , R_879_15884c78 );
buf ( n2914 , R_1003_124c39f8 );
buf ( n2915 , R_1a16_1486b418 );
buf ( n2916 , R_13f7_13d24338 );
buf ( n2917 , R_dd8_1587fd18 );
buf ( n2918 , R_7b9_13c0f458 );
buf ( n2919 , R_aa4_13c1d0f8 );
buf ( n2920 , R_10c3_13ccbef8 );
buf ( n2921 , R_16e2_140b6df8 );
buf ( n2922 , R_1573_14a0c498 );
buf ( n2923 , R_f54_11632858 );
buf ( n2924 , R_935_150e5318 );
buf ( n2925 , R_928_156aab98 );
buf ( n2926 , R_f47_13cd9238 );
buf ( n2927 , R_1566_123b2a58 );
buf ( n2928 , R_a0b_11637858 );
buf ( n2929 , R_e71_14b21a38 );
buf ( n2930 , R_102a_11c6ccb8 );
buf ( n2931 , R_852_14b1d938 );
buf ( n2932 , R_1490_13bf8158 );
buf ( n2933 , R_1649_13dd4f98 );
buf ( n2934 , R_a12_1008b358 );
buf ( n2935 , R_e6a_156b7a78 );
buf ( n2936 , R_1031_14b25778 );
buf ( n2937 , R_84b_156ad1b8 );
buf ( n2938 , R_1650_13dd4e58 );
buf ( n2939 , R_1489_13c21978 );
buf ( n2940 , R_7e8_1486a0b8 );
buf ( n2941 , R_1a45_1162e2f8 );
buf ( n2942 , R_a75_156b0778 );
buf ( n2943 , R_1426_11637718 );
buf ( n2944 , R_1094_13d28398 );
buf ( n2945 , R_16b3_117efeb8 );
buf ( n2946 , R_e07_13d453d8 );
buf ( n2947 , R_17bd_1162b918 );
buf ( n2948 , R_b7f_14a0be58 );
buf ( n2949 , R_cfd_13d1d038 );
buf ( n2950 , R_193b_13d39f38 );
buf ( n2951 , R_119e_13c1bcf8 );
buf ( n2952 , R_560_12fbf118 );
buf ( n2953 , R_6de_13cd4058 );
buf ( n2954 , R_131c_13c245d8 );
buf ( n2955 , R_1891_123b9858 );
buf ( n2956 , R_1272_13dd9ef8 );
buf ( n2957 , R_c53_15ff5148 );
buf ( n2958 , R_634_11631818 );
buf ( n2959 , R_60a_156b2758 );
buf ( n2960 , R_c29_13cd0598 );
buf ( n2961 , R_1248_12fbfcf8 );
buf ( n2962 , R_1867_14a0ded8 );
buf ( n2963 , R_9cd_13d1f518 );
buf ( n2964 , R_14ce_1008b5d8 );
buf ( n2965 , R_160b_14b24cd8 );
buf ( n2966 , R_890_11628df8 );
buf ( n2967 , R_fec_13ccc5d8 );
buf ( n2968 , R_eaf_13d5baf8 );
buf ( n2969 , R_15bc_15889138 );
buf ( n2970 , R_8df_11637358 );
buf ( n2971 , R_f9d_158889b8 );
buf ( n2972 , R_efe_11632b78 );
buf ( n2973 , R_97e_13c29718 );
buf ( n2974 , R_151d_1700bc48 );
buf ( n2975 , R_ae2_123bdef8 );
buf ( n2976 , R_77b_17011828 );
buf ( n2977 , R_d9a_13c047d8 );
buf ( n2978 , R_13b9_15ffc948 );
buf ( n2979 , R_19d8_14870b98 );
buf ( n2980 , R_1720_156b9198 );
buf ( n2981 , R_1101_140b7398 );
buf ( n2982 , R_1202_15881898 );
buf ( n2983 , R_67a_13de2878 );
buf ( n2984 , R_1821_117f1c18 );
buf ( n2985 , R_18d7_1580f378 );
buf ( n2986 , R_5c4_14868fd8 );
buf ( n2987 , R_12b8_11631b38 );
buf ( n2988 , R_be3_13de2198 );
buf ( n2989 , R_c99_13c029d8 );
buf ( n2990 , R_fd1_13c1d058 );
buf ( n2991 , R_14e9_14868538 );
buf ( n2992 , R_9b2_1580b6d8 );
buf ( n2993 , R_8ab_14a0fc38 );
buf ( n2994 , R_15f0_140ae3d8 );
buf ( n2995 , R_eca_14a11df8 );
buf ( n2996 , R_1574_13cd7cf8 );
buf ( n2997 , R_f55_14b1ac38 );
buf ( n2998 , R_936_140acf38 );
buf ( n2999 , R_927_124c4178 );
buf ( n3000 , R_f46_14a0af58 );
buf ( n3001 , R_1565_1700e808 );
buf ( n3002 , R_14d3_1580e5b8 );
buf ( n3003 , R_9c8_15fef248 );
buf ( n3004 , R_895_13d532b8 );
buf ( n3005 , R_1606_1007ef18 );
buf ( n3006 , R_eb4_117eda78 );
buf ( n3007 , R_fe7_1162ba58 );
buf ( n3008 , R_8f6_156b7b18 );
buf ( n3009 , R_f15_158819d8 );
buf ( n3010 , R_15a5_158168f8 );
buf ( n3011 , R_1534_123b9c18 );
buf ( n3012 , R_f86_13c1ce78 );
buf ( n3013 , R_967_11c68938 );
buf ( n3014 , R_1901_15817ed8 );
buf ( n3015 , R_6a4_1162c1d8 );
buf ( n3016 , R_bb9_156ab1d8 );
buf ( n3017 , R_12e2_11636a98 );
buf ( n3018 , R_11d8_156aa738 );
buf ( n3019 , R_cc3_15887c98 );
buf ( n3020 , R_59a_117f76b8 );
buf ( n3021 , R_17f7_117e9838 );
buf ( n3022 , R_105d_123b4998 );
buf ( n3023 , R_145d_123bec18 );
buf ( n3024 , R_167c_140b6178 );
buf ( n3025 , R_e3e_150da7d8 );
buf ( n3026 , R_a3e_11635cd8 );
buf ( n3027 , R_81f_156b45f8 );
buf ( n3028 , R_120b_13def358 );
buf ( n3029 , R_671_140b4058 );
buf ( n3030 , R_182a_117ef698 );
buf ( n3031 , R_18ce_156b4e18 );
buf ( n3032 , R_5cd_14a185b8 );
buf ( n3033 , R_12af_15ff69a8 );
buf ( n3034 , R_bec_124c2878 );
buf ( n3035 , R_c90_117eb778 );
buf ( n3036 , R_1386_14a0c7b8 );
buf ( n3037 , R_19a5_1008a598 );
buf ( n3038 , R_1753_13cd1218 );
buf ( n3039 , R_748_13d3b518 );
buf ( n3040 , R_1134_1580ad78 );
buf ( n3041 , R_d67_13d3caf8 );
buf ( n3042 , R_b15_156b2078 );
buf ( n3043 , R_128a_15880718 );
buf ( n3044 , R_c6b_14a13518 );
buf ( n3045 , R_64c_148739d8 );
buf ( n3046 , R_5f2_13dd5538 );
buf ( n3047 , R_c11_15ff5aa8 );
buf ( n3048 , R_1230_124c42b8 );
buf ( n3049 , R_184f_1587fa98 );
buf ( n3050 , R_18a9_11c6f918 );
buf ( n3051 , R_bbf_1587ddd8 );
buf ( n3052 , R_69e_123b5bb8 );
buf ( n3053 , R_18fb_13df16f8 );
buf ( n3054 , R_11de_10089058 );
buf ( n3055 , R_12dc_13c0bc18 );
buf ( n3056 , R_17fd_13d408d8 );
buf ( n3057 , R_5a0_11631db8 );
buf ( n3058 , R_cbd_14872df8 );
buf ( n3059 , R_691_15883378 );
buf ( n3060 , R_18ee_14a171b8 );
buf ( n3061 , R_11eb_13d4f078 );
buf ( n3062 , R_12cf_158850d8 );
buf ( n3063 , R_180a_13d3fc58 );
buf ( n3064 , R_5ad_14a0c2b8 );
buf ( n3065 , R_cb0_13de1658 );
buf ( n3066 , R_bcc_13df1f18 );
buf ( n3067 , R_1472_13d3c698 );
buf ( n3068 , R_1048_13df8bd8 );
buf ( n3069 , R_e53_10087b18 );
buf ( n3070 , R_1667_13beaf58 );
buf ( n3071 , R_834_15888698 );
buf ( n3072 , R_a29_13de0618 );
buf ( n3073 , R_1575_13d42598 );
buf ( n3074 , R_f56_13c0c578 );
buf ( n3075 , R_937_15886c58 );
buf ( n3076 , R_926_158846d8 );
buf ( n3077 , R_f45_13d4f438 );
buf ( n3078 , R_1564_1587b038 );
buf ( n3079 , R_906_14a145f8 );
buf ( n3080 , R_f25_13d24e78 );
buf ( n3081 , R_1544_124c4fd8 );
buf ( n3082 , R_1595_14b1f698 );
buf ( n3083 , R_f76_117f6fd8 );
buf ( n3084 , R_957_15888878 );
buf ( n3085 , R_c7a_140ac998 );
buf ( n3086 , R_65b_1580b778 );
buf ( n3087 , R_5e3_117eba98 );
buf ( n3088 , R_c02_123b2f58 );
buf ( n3089 , R_18b8_12fc05b8 );
buf ( n3090 , R_1221_15812cf8 );
buf ( n3091 , R_1299_14b1fc38 );
buf ( n3092 , R_1840_13d549d8 );
buf ( n3093 , R_1947_156ac3f8 );
buf ( n3094 , R_d09_150dd438 );
buf ( n3095 , R_b73_117f7938 );
buf ( n3096 , R_17b1_14a0dcf8 );
buf ( n3097 , R_1328_13d2aeb8 );
buf ( n3098 , R_6ea_123bbb58 );
buf ( n3099 , R_1192_1587dbf8 );
buf ( n3100 , R_137e_13c27738 );
buf ( n3101 , R_175b_15883ff8 );
buf ( n3102 , R_199d_1008a6d8 );
buf ( n3103 , R_113c_13d20eb8 );
buf ( n3104 , R_740_13bf6b78 );
buf ( n3105 , R_b1d_123c1918 );
buf ( n3106 , R_d5f_15888c38 );
buf ( n3107 , R_fcb_13def8f8 );
buf ( n3108 , R_8b1_170124a8 );
buf ( n3109 , R_9ac_14a190f8 );
buf ( n3110 , R_ed0_13d23d98 );
buf ( n3111 , R_15ea_1580e658 );
buf ( n3112 , R_14ef_123bead8 );
buf ( n3113 , R_d33_123bd8b8 );
buf ( n3114 , R_1168_156b6fd8 );
buf ( n3115 , R_1352_13c10b78 );
buf ( n3116 , R_b49_14a158b8 );
buf ( n3117 , R_714_1587c898 );
buf ( n3118 , R_1971_13ddfe98 );
buf ( n3119 , R_1787_1486e2f8 );
buf ( n3120 , R_68a_14a15b38 );
buf ( n3121 , R_11f2_1162a6f8 );
buf ( n3122 , R_18e7_13c08c98 );
buf ( n3123 , R_1811_117e9a18 );
buf ( n3124 , R_12c8_140aa878 );
buf ( n3125 , R_5b4_140b2a78 );
buf ( n3126 , R_ca9_15887e78 );
buf ( n3127 , R_bd3_13c0e9b8 );
buf ( n3128 , R_195d_15884818 );
buf ( n3129 , R_117c_14874838 );
buf ( n3130 , R_d1f_1007f698 );
buf ( n3131 , R_b5d_123bb8d8 );
buf ( n3132 , R_133e_13d55dd8 );
buf ( n3133 , R_179b_12fbde58 );
buf ( n3134 , R_700_13cd9878 );
buf ( n3135 , R_1576_1700c6e8 );
buf ( n3136 , R_f57_14a14198 );
buf ( n3137 , R_938_13bedc58 );
buf ( n3138 , R_925_13df1338 );
buf ( n3139 , R_f44_156b99b8 );
buf ( n3140 , R_1563_158841d8 );
buf ( n3141 , R_c86_14a12e38 );
buf ( n3142 , R_1834_13cd3f18 );
buf ( n3143 , R_667_1486b558 );
buf ( n3144 , R_5d7_156b0c78 );
buf ( n3145 , R_18c4_11c709f8 );
buf ( n3146 , R_bf6_11c6f378 );
buf ( n3147 , R_12a5_1162d718 );
buf ( n3148 , R_1215_117f51d8 );
buf ( n3149 , R_1892_13d3b1f8 );
buf ( n3150 , R_1273_13dd5c18 );
buf ( n3151 , R_c54_13becd58 );
buf ( n3152 , R_635_13d2c678 );
buf ( n3153 , R_609_1580ef18 );
buf ( n3154 , R_c28_140ba098 );
buf ( n3155 , R_1247_13ccda78 );
buf ( n3156 , R_1866_13bf9eb8 );
buf ( n3157 , R_9d2_13ccb958 );
buf ( n3158 , R_14c9_117f80b8 );
buf ( n3159 , R_1610_1700a988 );
buf ( n3160 , R_88b_1587e5f8 );
buf ( n3161 , R_ff1_13b8bd18 );
buf ( n3162 , R_eaa_13dd6618 );
buf ( n3163 , R_1708_11630558 );
buf ( n3164 , R_10e9_123c2138 );
buf ( n3165 , R_aca_14a131f8 );
buf ( n3166 , R_793_12fc2138 );
buf ( n3167 , R_db2_123b68d8 );
buf ( n3168 , R_13d1_156ac998 );
buf ( n3169 , R_19f0_13d47138 );
buf ( n3170 , R_7d3_13dd99f8 );
buf ( n3171 , R_a8a_150e0ef8 );
buf ( n3172 , R_10a9_1486ae78 );
buf ( n3173 , R_16c8_13dfaed8 );
buf ( n3174 , R_1a30_14a19698 );
buf ( n3175 , R_1411_13dfa438 );
buf ( n3176 , R_df2_150e09f8 );
buf ( n3177 , R_14e3_11634838 );
buf ( n3178 , R_9b8_13d43b78 );
buf ( n3179 , R_8a5_13bee798 );
buf ( n3180 , R_15f6_117f0458 );
buf ( n3181 , R_ec4_11c68a78 );
buf ( n3182 , R_fd7_116387f8 );
buf ( n3183 , R_17c1_13d57d18 );
buf ( n3184 , R_b83_13bedd98 );
buf ( n3185 , R_cf9_1587d798 );
buf ( n3186 , R_1937_150e3c98 );
buf ( n3187 , R_11a2_13c05138 );
buf ( n3188 , R_564_15815278 );
buf ( n3189 , R_6da_13c00f98 );
buf ( n3190 , R_1318_1008a9f8 );
buf ( n3191 , R_faf_158866b8 );
buf ( n3192 , R_8cd_15ff2ee8 );
buf ( n3193 , R_eec_117f7078 );
buf ( n3194 , R_990_11633c58 );
buf ( n3195 , R_150b_13cd8dd8 );
buf ( n3196 , R_15ce_13df0898 );
buf ( n3197 , R_1766_116318b8 );
buf ( n3198 , R_1373_15810598 );
buf ( n3199 , R_1147_13b8d438 );
buf ( n3200 , R_1992_13b8d1b8 );
buf ( n3201 , R_735_13cd4cd8 );
buf ( n3202 , R_b28_1162fab8 );
buf ( n3203 , R_d54_150e15d8 );
buf ( n3204 , R_1577_13d44ed8 );
buf ( n3205 , R_f58_13d3e178 );
buf ( n3206 , R_939_123b2878 );
buf ( n3207 , R_924_140b7118 );
buf ( n3208 , R_f43_140aeab8 );
buf ( n3209 , R_1562_100874d8 );
buf ( n3210 , R_17ce_13d50b58 );
buf ( n3211 , R_b90_14a17e38 );
buf ( n3212 , R_cec_156b8fb8 );
buf ( n3213 , R_192a_13df93f8 );
buf ( n3214 , R_11af_156b2a78 );
buf ( n3215 , R_571_13b96ad8 );
buf ( n3216 , R_6cd_150dc5d8 );
buf ( n3217 , R_130b_14b1eab8 );
buf ( n3218 , R_19b7_117f7758 );
buf ( n3219 , R_75a_150de5b8 );
buf ( n3220 , R_1741_100824d8 );
buf ( n3221 , R_d79_1008a638 );
buf ( n3222 , R_1122_150e9a58 );
buf ( n3223 , R_1398_10083978 );
buf ( n3224 , R_b03_158129d8 );
buf ( n3225 , R_14d8_13cd4698 );
buf ( n3226 , R_9c3_13befa58 );
buf ( n3227 , R_89a_117edb18 );
buf ( n3228 , R_1601_13d272b8 );
buf ( n3229 , R_eb9_11638438 );
buf ( n3230 , R_fe2_13defdf8 );
buf ( n3231 , R_13f9_1580cb78 );
buf ( n3232 , R_dda_117f7118 );
buf ( n3233 , R_7bb_13bf54f8 );
buf ( n3234 , R_aa2_12fc1a58 );
buf ( n3235 , R_10c1_13b901d8 );
buf ( n3236 , R_16e0_158811b8 );
buf ( n3237 , R_1a18_156b8bf8 );
buf ( n3238 , R_fbe_13cd90f8 );
buf ( n3239 , R_8be_13df3278 );
buf ( n3240 , R_99f_123b6b58 );
buf ( n3241 , R_edd_13b99cd8 );
buf ( n3242 , R_15dd_156aef18 );
buf ( n3243 , R_14fc_140b09f8 );
buf ( n3244 , R_19b2_150e0318 );
buf ( n3245 , R_1746_123b75f8 );
buf ( n3246 , R_755_14a13338 );
buf ( n3247 , R_1127_13de3318 );
buf ( n3248 , R_d74_17011d28 );
buf ( n3249 , R_b08_150dce98 );
buf ( n3250 , R_1393_11c68c58 );
buf ( n3251 , R_1956_15813158 );
buf ( n3252 , R_d18_156b9698 );
buf ( n3253 , R_b64_156b3a18 );
buf ( n3254 , R_17a2_117e8758 );
buf ( n3255 , R_1337_13d20af8 );
buf ( n3256 , R_6f9_17012b88 );
buf ( n3257 , R_1183_1580f698 );
buf ( n3258 , R_bb3_17013d08 );
buf ( n3259 , R_12e8_14b1e158 );
buf ( n3260 , R_11d2_124c3318 );
buf ( n3261 , R_cc9_11c6e018 );
buf ( n3262 , R_594_13cd9698 );
buf ( n3263 , R_17f1_13c0bdf8 );
buf ( n3264 , R_1907_13ccaa58 );
buf ( n3265 , R_6aa_13de4038 );
buf ( n3266 , R_ba3_13cd5bd8 );
buf ( n3267 , R_12f8_13cd2758 );
buf ( n3268 , R_11c2_13c1fc18 );
buf ( n3269 , R_cd9_14b1f878 );
buf ( n3270 , R_584_12fc0bf8 );
buf ( n3271 , R_1917_13d21f98 );
buf ( n3272 , R_17e1_13d37878 );
buf ( n3273 , R_6ba_11637b78 );
buf ( n3274 , R_8e9_13cd6b78 );
buf ( n3275 , R_15b2_117f08b8 );
buf ( n3276 , R_f08_156b5db8 );
buf ( n3277 , R_f93_13b92758 );
buf ( n3278 , R_1527_13ccaeb8 );
buf ( n3279 , R_974_13c0c2f8 );
buf ( n3280 , R_ad9_150e2a78 );
buf ( n3281 , R_784_13dfa4d8 );
buf ( n3282 , R_da3_14a0cd58 );
buf ( n3283 , R_13c2_13d2a4b8 );
buf ( n3284 , R_19e1_1700c5a8 );
buf ( n3285 , R_1717_13df61f8 );
buf ( n3286 , R_10f8_156b7258 );
buf ( n3287 , R_1578_123bab18 );
buf ( n3288 , R_f59_13c10358 );
buf ( n3289 , R_93a_1486f978 );
buf ( n3290 , R_923_11632178 );
buf ( n3291 , R_f42_14b1f9b8 );
buf ( n3292 , R_1561_13bf4a58 );
buf ( n3293 , R_1060_13c0b358 );
buf ( n3294 , R_145a_14a12bb8 );
buf ( n3295 , R_167f_14a19378 );
buf ( n3296 , R_e3b_13dd7f18 );
buf ( n3297 , R_a41_14a10d18 );
buf ( n3298 , R_81c_13bf79d8 );
buf ( n3299 , R_12fd_1007d9d8 );
buf ( n3300 , R_b9e_123ba618 );
buf ( n3301 , R_cde_13d39218 );
buf ( n3302 , R_11bd_11c6dcf8 );
buf ( n3303 , R_191c_1580c038 );
buf ( n3304 , R_57f_158160d8 );
buf ( n3305 , R_6bf_13df4e98 );
buf ( n3306 , R_17dc_15ff5508 );
buf ( n3307 , R_1893_117f0d18 );
buf ( n3308 , R_1274_156b1218 );
buf ( n3309 , R_c55_13cce338 );
buf ( n3310 , R_636_123c1238 );
buf ( n3311 , R_608_13d58678 );
buf ( n3312 , R_c27_13bf2a78 );
buf ( n3313 , R_1246_14b229d8 );
buf ( n3314 , R_1865_156b4d78 );
buf ( n3315 , R_772_11634a18 );
buf ( n3316 , R_d91_13c0fdb8 );
buf ( n3317 , R_13b0_1486d0d8 );
buf ( n3318 , R_1729_123b6338 );
buf ( n3319 , R_19cf_11c70c78 );
buf ( n3320 , R_110a_156b12b8 );
buf ( n3321 , R_aeb_11638758 );
buf ( n3322 , R_e78_117ef0f8 );
buf ( n3323 , R_1023_15ff3ac8 );
buf ( n3324 , R_859_13c0f098 );
buf ( n3325 , R_1497_116337f8 );
buf ( n3326 , R_1642_1162e578 );
buf ( n3327 , R_a04_13c22e18 );
buf ( n3328 , R_76b_13ddaad8 );
buf ( n3329 , R_d8a_10085458 );
buf ( n3330 , R_1730_11c6fd78 );
buf ( n3331 , R_13a9_15887978 );
buf ( n3332 , R_1111_11629c58 );
buf ( n3333 , R_19c8_123b61f8 );
buf ( n3334 , R_af2_11635558 );
buf ( n3335 , R_1045_13c2abb8 );
buf ( n3336 , R_e56_13c1f0d8 );
buf ( n3337 , R_1664_1700d9a8 );
buf ( n3338 , R_837_13d43c18 );
buf ( n3339 , R_a26_13c28c78 );
buf ( n3340 , R_1475_123b8bd8 );
buf ( n3341 , R_e63_156b1358 );
buf ( n3342 , R_1038_10085f98 );
buf ( n3343 , R_1657_13cd2c58 );
buf ( n3344 , R_844_117f3ab8 );
buf ( n3345 , R_1482_140b29d8 );
buf ( n3346 , R_a19_156ad4d8 );
buf ( n3347 , R_18f5_1587d518 );
buf ( n3348 , R_11e4_158159f8 );
buf ( n3349 , R_12d6_11c6c5d8 );
buf ( n3350 , R_1803_123b54d8 );
buf ( n3351 , R_5a6_13ccf5f8 );
buf ( n3352 , R_cb7_1162c458 );
buf ( n3353 , R_bc5_14a0c5d8 );
buf ( n3354 , R_698_14a0feb8 );
buf ( n3355 , R_194b_15882658 );
buf ( n3356 , R_d0d_1580bef8 );
buf ( n3357 , R_b6f_117eb638 );
buf ( n3358 , R_17ad_156b4f58 );
buf ( n3359 , R_132c_158823d8 );
buf ( n3360 , R_6ee_14a0faf8 );
buf ( n3361 , R_118e_156ab3b8 );
buf ( n3362 , R_75f_14870918 );
buf ( n3363 , R_173c_123b9218 );
buf ( n3364 , R_d7e_11634018 );
buf ( n3365 , R_111d_13beeb58 );
buf ( n3366 , R_139d_100868f8 );
buf ( n3367 , R_afe_15ff7ee8 );
buf ( n3368 , R_19bc_17010248 );
buf ( n3369 , R_1175_11634c98 );
buf ( n3370 , R_d26_1587cf78 );
buf ( n3371 , R_b56_13c236d8 );
buf ( n3372 , R_1345_13cd4738 );
buf ( n3373 , R_1794_15813338 );
buf ( n3374 , R_707_13d580d8 );
buf ( n3375 , R_1964_13d42b38 );
buf ( n3376 , R_f24_13b92938 );
buf ( n3377 , R_1543_15ff0828 );
buf ( n3378 , R_1596_15ff8a28 );
buf ( n3379 , R_f77_158124d8 );
buf ( n3380 , R_958_13df5bb8 );
buf ( n3381 , R_905_13d4f758 );
buf ( n3382 , R_1579_13b8d078 );
buf ( n3383 , R_f5a_15884d18 );
buf ( n3384 , R_93b_1580c3f8 );
buf ( n3385 , R_922_140af198 );
buf ( n3386 , R_f41_156b7cf8 );
buf ( n3387 , R_1560_14a14cd8 );
buf ( n3388 , R_c6c_14b20318 );
buf ( n3389 , R_64d_13ccebf8 );
buf ( n3390 , R_5f1_15814c38 );
buf ( n3391 , R_c10_15817898 );
buf ( n3392 , R_122f_13d22038 );
buf ( n3393 , R_184e_14b1b8b8 );
buf ( n3394 , R_18aa_11638b18 );
buf ( n3395 , R_128b_1587eaf8 );
buf ( n3396 , R_1695_14a12ed8 );
buf ( n3397 , R_1a63_1486ec58 );
buf ( n3398 , R_1444_15ff0788 );
buf ( n3399 , R_a57_13d5aa18 );
buf ( n3400 , R_e25_14a17078 );
buf ( n3401 , R_1076_1587b678 );
buf ( n3402 , R_806_14a0bd18 );
buf ( n3403 , R_fb7_15887158 );
buf ( n3404 , R_8c5_1008b2b8 );
buf ( n3405 , R_998_13d573b8 );
buf ( n3406 , R_ee4_15ff7da8 );
buf ( n3407 , R_1503_150daf58 );
buf ( n3408 , R_15d6_117ed398 );
buf ( n3409 , R_7ca_150de978 );
buf ( n3410 , R_a93_156af4b8 );
buf ( n3411 , R_10b2_100826b8 );
buf ( n3412 , R_16d1_156b27f8 );
buf ( n3413 , R_1a27_13cd2118 );
buf ( n3414 , R_1408_1587fbd8 );
buf ( n3415 , R_de9_13cd12b8 );
buf ( n3416 , R_9e0_15ffc9e8 );
buf ( n3417 , R_161e_123b8a98 );
buf ( n3418 , R_14bb_10081cb8 );
buf ( n3419 , R_87d_123b9498 );
buf ( n3420 , R_fff_12fbe5d8 );
buf ( n3421 , R_e9c_13df34f8 );
buf ( n3422 , R_ba8_123c12d8 );
buf ( n3423 , R_12f3_11634f18 );
buf ( n3424 , R_11c7_17013b28 );
buf ( n3425 , R_cd4_13c2b018 );
buf ( n3426 , R_589_14a19058 );
buf ( n3427 , R_1912_156aacd8 );
buf ( n3428 , R_17e6_140b2758 );
buf ( n3429 , R_6b5_1587d658 );
buf ( n3430 , R_f14_13d26458 );
buf ( n3431 , R_15a6_1162eb18 );
buf ( n3432 , R_1533_14b268f8 );
buf ( n3433 , R_f87_11637998 );
buf ( n3434 , R_968_13d2b958 );
buf ( n3435 , R_8f5_13bebe58 );
buf ( n3436 , R_8d5_150e1c18 );
buf ( n3437 , R_fa7_12fbff78 );
buf ( n3438 , R_ef4_1162ea78 );
buf ( n3439 , R_988_15814198 );
buf ( n3440 , R_1513_13c06498 );
buf ( n3441 , R_15c6_12fbf2f8 );
buf ( n3442 , R_8b7_15ffa468 );
buf ( n3443 , R_9a6_13d46058 );
buf ( n3444 , R_ed6_13d57598 );
buf ( n3445 , R_15e4_156aeb58 );
buf ( n3446 , R_14f5_13c29178 );
buf ( n3447 , R_fc5_13b8d258 );
buf ( n3448 , R_acc_13df8638 );
buf ( n3449 , R_791_13d42818 );
buf ( n3450 , R_db0_13bf9418 );
buf ( n3451 , R_13cf_123c2318 );
buf ( n3452 , R_19ee_11630cd8 );
buf ( n3453 , R_170a_13d25698 );
buf ( n3454 , R_10eb_13debbb8 );
buf ( n3455 , R_19ad_1587f9f8 );
buf ( n3456 , R_174b_15ff3528 );
buf ( n3457 , R_750_1008c9d8 );
buf ( n3458 , R_112c_13c015d8 );
buf ( n3459 , R_d6f_117eae18 );
buf ( n3460 , R_b0d_13d41c38 );
buf ( n3461 , R_138e_158113f8 );
buf ( n3462 , R_168d_156b2f78 );
buf ( n3463 , R_144c_14a0dbb8 );
buf ( n3464 , R_e2d_1587d3d8 );
buf ( n3465 , R_a4f_15814418 );
buf ( n3466 , R_80e_156ac218 );
buf ( n3467 , R_106e_14a15318 );
buf ( n3468 , R_157a_156b4198 );
buf ( n3469 , R_f5b_1162d7b8 );
buf ( n3470 , R_93c_13b933d8 );
buf ( n3471 , R_921_15813298 );
buf ( n3472 , R_f40_13cd1fd8 );
buf ( n3473 , R_155f_148745b8 );
buf ( n3474 , R_1275_13d26bd8 );
buf ( n3475 , R_c56_12fbf438 );
buf ( n3476 , R_637_14b20db8 );
buf ( n3477 , R_607_15886258 );
buf ( n3478 , R_c26_13d3ac58 );
buf ( n3479 , R_1245_13d261d8 );
buf ( n3480 , R_1864_13ddb2f8 );
buf ( n3481 , R_1894_13cd6998 );
buf ( n3482 , R_9d7_1580ac38 );
buf ( n3483 , R_1615_150e0598 );
buf ( n3484 , R_14c4_15ffa148 );
buf ( n3485 , R_886_156aa9b8 );
buf ( n3486 , R_ff6_13d424f8 );
buf ( n3487 , R_ea5_13d23b18 );
buf ( n3488 , R_1a51_13cda098 );
buf ( n3489 , R_a69_123b4f38 );
buf ( n3490 , R_1432_14b1d258 );
buf ( n3491 , R_1088_13bec3f8 );
buf ( n3492 , R_e13_140ab1d8 );
buf ( n3493 , R_16a7_156afb98 );
buf ( n3494 , R_7f4_14b238d8 );
buf ( n3495 , R_17c5_12fc1058 );
buf ( n3496 , R_b87_140b0db8 );
buf ( n3497 , R_cf5_156ab818 );
buf ( n3498 , R_1933_11633258 );
buf ( n3499 , R_11a6_13c243f8 );
buf ( n3500 , R_568_13ccd9d8 );
buf ( n3501 , R_6d6_13ccc498 );
buf ( n3502 , R_1314_13b93158 );
buf ( n3503 , R_a81_11c6b098 );
buf ( n3504 , R_10a0_148694d8 );
buf ( n3505 , R_1a39_150e4cd8 );
buf ( n3506 , R_16bf_13d3e8f8 );
buf ( n3507 , R_141a_13ccc678 );
buf ( n3508 , R_dfb_123b4c18 );
buf ( n3509 , R_7dc_14b22578 );
buf ( n3510 , R_116b_13ddcb58 );
buf ( n3511 , R_134f_14b1c7b8 );
buf ( n3512 , R_b4c_13d41eb8 );
buf ( n3513 , R_711_140b8798 );
buf ( n3514 , R_178a_13b96538 );
buf ( n3515 , R_196e_150e3658 );
buf ( n3516 , R_d30_13df5118 );
buf ( n3517 , R_b99_13df2ff8 );
buf ( n3518 , R_ce3_10088b58 );
buf ( n3519 , R_11b8_156b8798 );
buf ( n3520 , R_1921_13b91df8 );
buf ( n3521 , R_57a_13ccb818 );
buf ( n3522 , R_6c4_15887798 );
buf ( n3523 , R_17d7_11c6faf8 );
buf ( n3524 , R_1302_12fbe8f8 );
buf ( n3525 , R_65c_117f0278 );
buf ( n3526 , R_5e2_117ef198 );
buf ( n3527 , R_c01_13df0118 );
buf ( n3528 , R_18b9_13ded058 );
buf ( n3529 , R_1220_117f77f8 );
buf ( n3530 , R_129a_14a10ef8 );
buf ( n3531 , R_183f_140b7f78 );
buf ( n3532 , R_c7b_1580c178 );
buf ( n3533 , R_7bd_12fc1558 );
buf ( n3534 , R_aa0_11c6be58 );
buf ( n3535 , R_10bf_13df54d8 );
buf ( n3536 , R_16de_13de3138 );
buf ( n3537 , R_1a1a_156b8ab8 );
buf ( n3538 , R_13fb_156b4b98 );
buf ( n3539 , R_ddc_11632df8 );
buf ( n3540 , R_a7a_11c6b1d8 );
buf ( n3541 , R_1a40_140b6d58 );
buf ( n3542 , R_1099_116354b8 );
buf ( n3543 , R_1421_117ef7d8 );
buf ( n3544 , R_16b8_13d3ea38 );
buf ( n3545 , R_e02_15ff37a8 );
buf ( n3546 , R_7e3_15812118 );
buf ( n3547 , R_1a56_13bf0818 );
buf ( n3548 , R_1437_123bad98 );
buf ( n3549 , R_a64_13beb318 );
buf ( n3550 , R_e18_156afc38 );
buf ( n3551 , R_1083_123c0a18 );
buf ( n3552 , R_7f9_156b30b8 );
buf ( n3553 , R_16a2_150e9418 );
buf ( n3554 , R_18e0_13c201b8 );
buf ( n3555 , R_1818_140b47d8 );
buf ( n3556 , R_12c1_123bb838 );
buf ( n3557 , R_5bb_156b5638 );
buf ( n3558 , R_ca2_13dd9d18 );
buf ( n3559 , R_bda_13b985b8 );
buf ( n3560 , R_683_11634478 );
buf ( n3561 , R_11f9_13ccd938 );
buf ( n3562 , R_157b_1486f0b8 );
buf ( n3563 , R_f5c_13de2378 );
buf ( n3564 , R_93d_117f0ef8 );
buf ( n3565 , R_920_13df90d8 );
buf ( n3566 , R_f3f_13bf1a38 );
buf ( n3567 , R_155e_123c0d38 );
buf ( n3568 , R_8de_13d4e0d8 );
buf ( n3569 , R_f9e_13b8a738 );
buf ( n3570 , R_efd_123bfed8 );
buf ( n3571 , R_97f_123c21d8 );
buf ( n3572 , R_151c_13d5c4f8 );
buf ( n3573 , R_15bd_13df43f8 );
buf ( n3574 , R_1763_13d44618 );
buf ( n3575 , R_1995_17017548 );
buf ( n3576 , R_1144_17018948 );
buf ( n3577 , R_738_1700bce8 );
buf ( n3578 , R_b25_1162ad38 );
buf ( n3579 , R_d57_13c242b8 );
buf ( n3580 , R_1376_117f5098 );
buf ( n3581 , R_9be_140aaaf8 );
buf ( n3582 , R_89f_156b2ed8 );
buf ( n3583 , R_15fc_13c28db8 );
buf ( n3584 , R_ebe_13cd5c78 );
buf ( n3585 , R_fdd_1162dd58 );
buf ( n3586 , R_14dd_123b8db8 );
buf ( n3587 , R_14aa_13c0f9f8 );
buf ( n3588 , R_86c_13df77d8 );
buf ( n3589 , R_1010_15884278 );
buf ( n3590 , R_e8b_15880ad8 );
buf ( n3591 , R_162f_15ff7808 );
buf ( n3592 , R_9f1_123be718 );
buf ( n3593 , R_1457_13d54758 );
buf ( n3594 , R_1682_1587fb38 );
buf ( n3595 , R_e38_150debf8 );
buf ( n3596 , R_a44_1580d618 );
buf ( n3597 , R_819_14873898 );
buf ( n3598 , R_1063_13cd8978 );
buf ( n3599 , R_1a4c_156b8b58 );
buf ( n3600 , R_a6e_117ec3f8 );
buf ( n3601 , R_142d_14b1c998 );
buf ( n3602 , R_108d_14a0a878 );
buf ( n3603 , R_e0e_156b9f58 );
buf ( n3604 , R_16ac_13bf1218 );
buf ( n3605 , R_7ef_1700c788 );
buf ( n3606 , R_1014_13c079d8 );
buf ( n3607 , R_868_1587de78 );
buf ( n3608 , R_14a6_10081998 );
buf ( n3609 , R_1633_117e9ab8 );
buf ( n3610 , R_9f5_13d25c38 );
buf ( n3611 , R_e87_15ff9ce8 );
buf ( n3612 , R_1829_123b40d8 );
buf ( n3613 , R_18cf_13ded238 );
buf ( n3614 , R_5cc_156aa698 );
buf ( n3615 , R_12b0_14a177f8 );
buf ( n3616 , R_beb_13cca738 );
buf ( n3617 , R_c91_15ff1cc8 );
buf ( n3618 , R_120a_13cd9738 );
buf ( n3619 , R_672_13c06fd8 );
buf ( n3620 , R_779_13cd2258 );
buf ( n3621 , R_d98_13b958b8 );
buf ( n3622 , R_13b7_1700e308 );
buf ( n3623 , R_19d6_117ecfd8 );
buf ( n3624 , R_1722_123b5a78 );
buf ( n3625 , R_1103_117f7bb8 );
buf ( n3626 , R_ae4_11634ab8 );
buf ( n3627 , R_c57_15814f58 );
buf ( n3628 , R_638_14a151d8 );
buf ( n3629 , R_606_13d50838 );
buf ( n3630 , R_c25_10083bf8 );
buf ( n3631 , R_1244_13ddb898 );
buf ( n3632 , R_1863_123b9f38 );
buf ( n3633 , R_1895_13df3a98 );
buf ( n3634 , R_1276_123bda98 );
buf ( n3635 , R_1042_13cd6718 );
buf ( n3636 , R_e59_1587dd38 );
buf ( n3637 , R_1661_13de0758 );
buf ( n3638 , R_83a_13d21598 );
buf ( n3639 , R_a23_14869cf8 );
buf ( n3640 , R_1478_13cd7618 );
buf ( n3641 , R_668_11c6aff8 );
buf ( n3642 , R_5d6_13d24158 );
buf ( n3643 , R_18c5_123b5f78 );
buf ( n3644 , R_bf5_123ba7f8 );
buf ( n3645 , R_12a6_148674f8 );
buf ( n3646 , R_1214_15886cf8 );
buf ( n3647 , R_c87_13c21bf8 );
buf ( n3648 , R_1833_117f3838 );
buf ( n3649 , R_1820_14872a38 );
buf ( n3650 , R_18d8_13b8ef18 );
buf ( n3651 , R_5c3_10080778 );
buf ( n3652 , R_12b9_140abb38 );
buf ( n3653 , R_be2_13b98338 );
buf ( n3654 , R_c9a_13cd1f38 );
buf ( n3655 , R_1201_15ff65e8 );
buf ( n3656 , R_67b_13c02bb8 );
buf ( n3657 , R_1542_14a19cd8 );
buf ( n3658 , R_1597_117ee478 );
buf ( n3659 , R_f78_156af198 );
buf ( n3660 , R_959_11631bd8 );
buf ( n3661 , R_904_13bebbd8 );
buf ( n3662 , R_f23_13c2b338 );
buf ( n3663 , R_157c_14a0eab8 );
buf ( n3664 , R_f5d_15817c58 );
buf ( n3665 , R_93e_13cd6858 );
buf ( n3666 , R_91f_117f7d98 );
buf ( n3667 , R_f3e_1700a708 );
buf ( n3668 , R_155d_1700fa28 );
buf ( n3669 , R_764_150dee78 );
buf ( n3670 , R_1737_13cd6538 );
buf ( n3671 , R_d83_150dc678 );
buf ( n3672 , R_1118_13cce3d8 );
buf ( n3673 , R_13a2_13df95d8 );
buf ( n3674 , R_af9_14b1bc78 );
buf ( n3675 , R_19c1_15811358 );
buf ( n3676 , R_14ae_14b22438 );
buf ( n3677 , R_870_158800d8 );
buf ( n3678 , R_100c_14b1bef8 );
buf ( n3679 , R_e8f_13c27cd8 );
buf ( n3680 , R_9ed_150e3a18 );
buf ( n3681 , R_162b_13d24478 );
buf ( n3682 , R_64e_12fbeb78 );
buf ( n3683 , R_5f0_13d25738 );
buf ( n3684 , R_c0f_1587ef58 );
buf ( n3685 , R_122e_14a181f8 );
buf ( n3686 , R_184d_1486ac98 );
buf ( n3687 , R_18ab_13bf9d78 );
buf ( n3688 , R_128c_11c6a378 );
buf ( n3689 , R_c6d_13d3be78 );
buf ( n3690 , R_d11_117f09f8 );
buf ( n3691 , R_b6b_13c0e878 );
buf ( n3692 , R_17a9_15ff62c8 );
buf ( n3693 , R_1330_1580d6b8 );
buf ( n3694 , R_6f2_123ba398 );
buf ( n3695 , R_118a_13c1eef8 );
buf ( n3696 , R_194f_13c0e738 );
buf ( n3697 , R_1758_14a14eb8 );
buf ( n3698 , R_19a0_13c204d8 );
buf ( n3699 , R_1139_117ef878 );
buf ( n3700 , R_743_13d5a478 );
buf ( n3701 , R_b1a_13c01038 );
buf ( n3702 , R_d62_15811df8 );
buf ( n3703 , R_1381_123b3a98 );
buf ( n3704 , R_e6d_123b7238 );
buf ( n3705 , R_102e_150ddd98 );
buf ( n3706 , R_84e_15883418 );
buf ( n3707 , R_164d_14a0c678 );
buf ( n3708 , R_148c_1580e8d8 );
buf ( n3709 , R_a0f_15ffbae8 );
buf ( n3710 , R_12ee_13d3d958 );
buf ( n3711 , R_11cc_14a11a38 );
buf ( n3712 , R_ccf_15812258 );
buf ( n3713 , R_58e_150e4558 );
buf ( n3714 , R_17eb_150e6538 );
buf ( n3715 , R_190d_14b294b8 );
buf ( n3716 , R_6b0_14a172f8 );
buf ( n3717 , R_bad_15883c38 );
buf ( n3718 , R_1018_13d2a878 );
buf ( n3719 , R_864_13c09238 );
buf ( n3720 , R_14a2_13cd9e18 );
buf ( n3721 , R_1637_1162fbf8 );
buf ( n3722 , R_9f9_156b7438 );
buf ( n3723 , R_e83_15886438 );
buf ( n3724 , R_1a5b_13df6158 );
buf ( n3725 , R_143c_15ff2a88 );
buf ( n3726 , R_a5f_13df1518 );
buf ( n3727 , R_e1d_13c288b8 );
buf ( n3728 , R_107e_13c1c298 );
buf ( n3729 , R_7fe_117f30b8 );
buf ( n3730 , R_169d_156abf98 );
buf ( n3731 , R_15b3_13cd6e98 );
buf ( n3732 , R_f07_13b953b8 );
buf ( n3733 , R_f94_13d25198 );
buf ( n3734 , R_1526_1486bf58 );
buf ( n3735 , R_975_13d529f8 );
buf ( n3736 , R_8e8_117f0bd8 );
buf ( n3737 , R_78f_1162c9f8 );
buf ( n3738 , R_dae_11c6d578 );
buf ( n3739 , R_13cd_14a162b8 );
buf ( n3740 , R_19ec_15814738 );
buf ( n3741 , R_170c_13ccdd98 );
buf ( n3742 , R_10ed_15882dd8 );
buf ( n3743 , R_ace_15885cb8 );
buf ( n3744 , R_157d_13cd56d8 );
buf ( n3745 , R_f5e_140b53b8 );
buf ( n3746 , R_93f_13d57778 );
buf ( n3747 , R_91e_15886f78 );
buf ( n3748 , R_f3d_11634798 );
buf ( n3749 , R_155c_156adf78 );
buf ( n3750 , R_782_15ffd168 );
buf ( n3751 , R_da1_14b290f8 );
buf ( n3752 , R_13c0_117f6b78 );
buf ( n3753 , R_19df_117eb318 );
buf ( n3754 , R_1719_13c1f8f8 );
buf ( n3755 , R_10fa_13decd38 );
buf ( n3756 , R_adb_17014708 );
buf ( n3757 , R_a88_13cd40f8 );
buf ( n3758 , R_10a7_117eb1d8 );
buf ( n3759 , R_16c6_158880f8 );
buf ( n3760 , R_1a32_15818018 );
buf ( n3761 , R_1413_13d57ef8 );
buf ( n3762 , R_df4_17013f88 );
buf ( n3763 , R_7d5_15889098 );
buf ( n3764 , R_639_13df0cf8 );
buf ( n3765 , R_605_14b1c3f8 );
buf ( n3766 , R_c24_11632d58 );
buf ( n3767 , R_1243_158151d8 );
buf ( n3768 , R_1862_140b94b8 );
buf ( n3769 , R_1896_13c0a598 );
buf ( n3770 , R_1277_13c27378 );
buf ( n3771 , R_c58_13dddc38 );
buf ( n3772 , R_15a7_17013448 );
buf ( n3773 , R_1532_156b4ff8 );
buf ( n3774 , R_f88_13d225d8 );
buf ( n3775 , R_969_13cce298 );
buf ( n3776 , R_8f4_156b9af8 );
buf ( n3777 , R_f13_13c2b478 );
buf ( n3778 , R_1750_14a13018 );
buf ( n3779 , R_74b_123b9998 );
buf ( n3780 , R_1131_13d21c78 );
buf ( n3781 , R_d6a_13c0c118 );
buf ( n3782 , R_b12_1587bb78 );
buf ( n3783 , R_1389_13c2a4d8 );
buf ( n3784 , R_19a8_124c5578 );
buf ( n3785 , R_a9e_13de43f8 );
buf ( n3786 , R_10bd_1162e6b8 );
buf ( n3787 , R_16dc_14b1f058 );
buf ( n3788 , R_1a1c_13cda138 );
buf ( n3789 , R_13fd_14a0e0b8 );
buf ( n3790 , R_dde_15ffc448 );
buf ( n3791 , R_7bf_123bb0b8 );
buf ( n3792 , R_1027_13c277d8 );
buf ( n3793 , R_855_14a117b8 );
buf ( n3794 , R_1493_13bee3d8 );
buf ( n3795 , R_1646_13ccbdb8 );
buf ( n3796 , R_a08_15ffa5a8 );
buf ( n3797 , R_e74_123b4678 );
buf ( n3798 , R_12d0_14a11cb8 );
buf ( n3799 , R_1809_13d4f7f8 );
buf ( n3800 , R_5ac_11c6e838 );
buf ( n3801 , R_cb1_13d2c998 );
buf ( n3802 , R_bcb_1007e3d8 );
buf ( n3803 , R_692_1587be98 );
buf ( n3804 , R_18ef_13d28758 );
buf ( n3805 , R_11ea_1580f238 );
buf ( n3806 , R_991_1007ff58 );
buf ( n3807 , R_eeb_12fbe0d8 );
buf ( n3808 , R_150a_14a0b3b8 );
buf ( n3809 , R_15cf_10085958 );
buf ( n3810 , R_fb0_117f5318 );
buf ( n3811 , R_8cc_13bf3338 );
buf ( n3812 , R_ce8_11c6a7d8 );
buf ( n3813 , R_1926_116372b8 );
buf ( n3814 , R_11b3_13cd3fb8 );
buf ( n3815 , R_575_15817438 );
buf ( n3816 , R_6c9_13dee318 );
buf ( n3817 , R_1307_15ff2da8 );
buf ( n3818 , R_17d2_156b8978 );
buf ( n3819 , R_b94_1587e198 );
buf ( n3820 , R_1810_117f12b8 );
buf ( n3821 , R_12c9_17017868 );
buf ( n3822 , R_5b3_123baa78 );
buf ( n3823 , R_caa_15fedbc8 );
buf ( n3824 , R_bd2_1580d9d8 );
buf ( n3825 , R_68b_13ddf038 );
buf ( n3826 , R_11f1_13c2a938 );
buf ( n3827 , R_18e8_123bd638 );
buf ( n3828 , R_157e_13dee278 );
buf ( n3829 , R_f5f_1162d038 );
buf ( n3830 , R_940_1486f838 );
buf ( n3831 , R_91d_14b1cdf8 );
buf ( n3832 , R_f3c_148682b8 );
buf ( n3833 , R_155b_12fc0158 );
buf ( n3834 , R_14b2_15ff2628 );
buf ( n3835 , R_874_123c0298 );
buf ( n3836 , R_1008_1587dc98 );
buf ( n3837 , R_e93_13cd4878 );
buf ( n3838 , R_9e9_123b4498 );
buf ( n3839 , R_1627_156b7578 );
buf ( n3840 , R_cf1_124c34f8 );
buf ( n3841 , R_192f_14a12cf8 );
buf ( n3842 , R_11aa_117e9bf8 );
buf ( n3843 , R_56c_140ab598 );
buf ( n3844 , R_6d2_1162ec58 );
buf ( n3845 , R_1310_13ddf538 );
buf ( n3846 , R_17c9_11638578 );
buf ( n3847 , R_b8b_13df36d8 );
buf ( n3848 , R_a91_13ccfeb8 );
buf ( n3849 , R_10b0_117ea418 );
buf ( n3850 , R_16cf_11c6b138 );
buf ( n3851 , R_1a29_13d384f8 );
buf ( n3852 , R_140a_140aa5f8 );
buf ( n3853 , R_deb_140b71b8 );
buf ( n3854 , R_7cc_13cd94b8 );
buf ( n3855 , R_1a47_100862b8 );
buf ( n3856 , R_a73_123be538 );
buf ( n3857 , R_1428_13dde3b8 );
buf ( n3858 , R_1092_15ff41a8 );
buf ( n3859 , R_e09_15887a18 );
buf ( n3860 , R_16b1_13c0c258 );
buf ( n3861 , R_7ea_11c6e518 );
buf ( n3862 , R_e66_170138a8 );
buf ( n3863 , R_1035_1162a478 );
buf ( n3864 , R_847_14a15a98 );
buf ( n3865 , R_1654_1580fff8 );
buf ( n3866 , R_1485_117f6358 );
buf ( n3867 , R_a16_14b25638 );
buf ( n3868 , R_b60_13b97b18 );
buf ( n3869 , R_179e_156b3c98 );
buf ( n3870 , R_133b_13ddde18 );
buf ( n3871 , R_6fd_156b8338 );
buf ( n3872 , R_117f_13cd7578 );
buf ( n3873 , R_195a_150e1218 );
buf ( n3874 , R_d1c_13d3fd98 );
buf ( n3875 , R_134c_14a11ad8 );
buf ( n3876 , R_b4f_12fbee98 );
buf ( n3877 , R_70e_124c25f8 );
buf ( n3878 , R_178d_11638a78 );
buf ( n3879 , R_196b_1580a918 );
buf ( n3880 , R_d2d_13cd54f8 );
buf ( n3881 , R_116e_117ebb38 );
buf ( n3882 , R_5e1_14b286f8 );
buf ( n3883 , R_c00_150df558 );
buf ( n3884 , R_18ba_11638bb8 );
buf ( n3885 , R_121f_13dfa1b8 );
buf ( n3886 , R_129b_13cd3298 );
buf ( n3887 , R_183e_1587c398 );
buf ( n3888 , R_c7c_11c6a558 );
buf ( n3889 , R_65d_13cd74d8 );
buf ( n3890 , R_9b3_13df8138 );
buf ( n3891 , R_8aa_13dd9a98 );
buf ( n3892 , R_15f1_156b5d18 );
buf ( n3893 , R_ec9_1587c1b8 );
buf ( n3894 , R_fd2_13c05098 );
buf ( n3895 , R_14e8_1700a528 );
buf ( n3896 , R_11dd_14875918 );
buf ( n3897 , R_12dd_14a0e158 );
buf ( n3898 , R_17fc_11635eb8 );
buf ( n3899 , R_59f_14a14c38 );
buf ( n3900 , R_cbe_116357d8 );
buf ( n3901 , R_bbe_15881438 );
buf ( n3902 , R_18fc_17009bc8 );
buf ( n3903 , R_69f_13d56b98 );
buf ( n3904 , R_1598_13cd92d8 );
buf ( n3905 , R_f79_13bf2e38 );
buf ( n3906 , R_95a_13d37698 );
buf ( n3907 , R_903_117ec7b8 );
buf ( n3908 , R_f22_14a13978 );
buf ( n3909 , R_1541_15886758 );
buf ( n3910 , R_12e3_17014028 );
buf ( n3911 , R_11d7_1587d5b8 );
buf ( n3912 , R_cc4_13bead78 );
buf ( n3913 , R_599_150dcf38 );
buf ( n3914 , R_17f6_117f1498 );
buf ( n3915 , R_1902_14b1af58 );
buf ( n3916 , R_6a5_13df56b8 );
buf ( n3917 , R_bb8_124c3b38 );
buf ( n3918 , R_14bf_150dd938 );
buf ( n3919 , R_881_150db278 );
buf ( n3920 , R_ffb_15813ab8 );
buf ( n3921 , R_ea0_13b95778 );
buf ( n3922 , R_9dc_15ff19a8 );
buf ( n3923 , R_161a_14b23bf8 );
buf ( n3924 , R_1454_123b4538 );
buf ( n3925 , R_e35_11c70098 );
buf ( n3926 , R_a47_1486f3d8 );
buf ( n3927 , R_816_13c06cb8 );
buf ( n3928 , R_1066_13bee838 );
buf ( n3929 , R_1685_15ff1d68 );
buf ( n3930 , R_8b0_15813c98 );
buf ( n3931 , R_9ad_13de0bb8 );
buf ( n3932 , R_ecf_13c26798 );
buf ( n3933 , R_15eb_140b6498 );
buf ( n3934 , R_14ee_13d5a298 );
buf ( n3935 , R_fcc_150e33d8 );
buf ( n3936 , R_101c_11c6ce98 );
buf ( n3937 , R_860_14a17b18 );
buf ( n3938 , R_149e_11c6edd8 );
buf ( n3939 , R_163b_13c04b98 );
buf ( n3940 , R_9fd_117ebf98 );
buf ( n3941 , R_e7f_117f6038 );
buf ( n3942 , R_604_15811718 );
buf ( n3943 , R_c23_123bfc58 );
buf ( n3944 , R_1242_10080c78 );
buf ( n3945 , R_1861_12fbf7f8 );
buf ( n3946 , R_1897_13d3d1d8 );
buf ( n3947 , R_1278_117f4f58 );
buf ( n3948 , R_c59_116304b8 );
buf ( n3949 , R_63a_13c0a278 );
buf ( n3950 , R_b59_15feff68 );
buf ( n3951 , R_1342_148716d8 );
buf ( n3952 , R_1797_117f7e38 );
buf ( n3953 , R_704_123b2ff8 );
buf ( n3954 , R_1961_1162de98 );
buf ( n3955 , R_1178_13cd24d8 );
buf ( n3956 , R_d23_11c68618 );
buf ( n3957 , R_157f_13b8ce98 );
buf ( n3958 , R_f60_140af9b8 );
buf ( n3959 , R_941_13df8b38 );
buf ( n3960 , R_91c_13df6d38 );
buf ( n3961 , R_f3b_15810c78 );
buf ( n3962 , R_155a_15882338 );
buf ( n3963 , R_e5c_117f6df8 );
buf ( n3964 , R_165e_117edf78 );
buf ( n3965 , R_83d_13c24ad8 );
buf ( n3966 , R_a20_15883738 );
buf ( n3967 , R_147b_1700f5c8 );
buf ( n3968 , R_103f_123b9ad8 );
buf ( n3969 , R_5ef_1162a018 );
buf ( n3970 , R_c0e_158802b8 );
buf ( n3971 , R_122d_150e4eb8 );
buf ( n3972 , R_184c_14a19418 );
buf ( n3973 , R_18ac_117f13f8 );
buf ( n3974 , R_128d_123b2af8 );
buf ( n3975 , R_c6e_15ff6408 );
buf ( n3976 , R_64f_13bf1ad8 );
buf ( n3977 , R_9a0_13dd6078 );
buf ( n3978 , R_edc_123be678 );
buf ( n3979 , R_15de_15ff2268 );
buf ( n3980 , R_14fb_13c29038 );
buf ( n3981 , R_fbf_150e4f58 );
buf ( n3982 , R_8bd_13cd5ef8 );
buf ( n3983 , R_1998_14b279d8 );
buf ( n3984 , R_1141_1580bbd8 );
buf ( n3985 , R_73b_14a15638 );
buf ( n3986 , R_b22_13cce8d8 );
buf ( n3987 , R_d5a_13bf6178 );
buf ( n3988 , R_1379_123bdbd8 );
buf ( n3989 , R_1760_117f7f78 );
buf ( n3990 , R_1981_1587b7b8 );
buf ( n3991 , R_b39_15ffae68 );
buf ( n3992 , R_724_117ec8f8 );
buf ( n3993 , R_1777_1587ccf8 );
buf ( n3994 , R_d43_13beedd8 );
buf ( n3995 , R_1362_150dfcd8 );
buf ( n3996 , R_1158_13bf0f98 );
buf ( n3997 , R_770_15888058 );
buf ( n3998 , R_d8f_11629f78 );
buf ( n3999 , R_13ae_13bf3478 );
buf ( n4000 , R_172b_156b88d8 );
buf ( n4001 , R_19cd_117ed578 );
buf ( n4002 , R_110c_15810458 );
buf ( n4003 , R_aed_14a0e298 );
buf ( n4004 , R_1449_14b26678 );
buf ( n4005 , R_e2a_13c29858 );
buf ( n4006 , R_a52_140af378 );
buf ( n4007 , R_80b_158154f8 );
buf ( n4008 , R_1071_123c1378 );
buf ( n4009 , R_1a68_117ed618 );
buf ( n4010 , R_1690_13c216f8 );
buf ( n4011 , R_ef3_13cd06d8 );
buf ( n4012 , R_989_13c068f8 );
buf ( n4013 , R_1512_1162e078 );
buf ( n4014 , R_15c7_13d3c4b8 );
buf ( n4015 , R_8d4_123c1738 );
buf ( n4016 , R_fa8_123be858 );
buf ( n4017 , R_1984_1162e438 );
buf ( n4018 , R_727_1700aca8 );
buf ( n4019 , R_b36_123bb338 );
buf ( n4020 , R_d46_13cd3338 );
buf ( n4021 , R_1774_13c26c98 );
buf ( n4022 , R_1365_150db818 );
buf ( n4023 , R_1155_17012868 );
buf ( n4024 , R_b3c_13cd4eb8 );
buf ( n4025 , R_721_156b7d98 );
buf ( n4026 , R_197e_13d5c8b8 );
buf ( n4027 , R_177a_123c1418 );
buf ( n4028 , R_d40_11635af8 );
buf ( n4029 , R_115b_123bf2f8 );
buf ( n4030 , R_135f_11c6da78 );
buf ( n4031 , R_894_1587b2b8 );
buf ( n4032 , R_1607_123bd138 );
buf ( n4033 , R_eb3_123b5cf8 );
buf ( n4034 , R_fe8_15816678 );
buf ( n4035 , R_14d2_11636e58 );
buf ( n4036 , R_9c9_13cce798 );
buf ( n4037 , R_160c_117f74d8 );
buf ( n4038 , R_88f_13c0d338 );
buf ( n4039 , R_fed_12fc1198 );
buf ( n4040 , R_eae_13cd1d58 );
buf ( n4041 , R_9ce_1162c6d8 );
buf ( n4042 , R_14cd_10081178 );
buf ( n4043 , R_dac_14a109f8 );
buf ( n4044 , R_13cb_13ccf0f8 );
buf ( n4045 , R_19ea_11629b18 );
buf ( n4046 , R_170e_1580e338 );
buf ( n4047 , R_10ef_14a199b8 );
buf ( n4048 , R_ad0_123b65b8 );
buf ( n4049 , R_78d_15817618 );
buf ( n4050 , R_999_1008a138 );
buf ( n4051 , R_ee3_158135b8 );
buf ( n4052 , R_1502_117ea238 );
buf ( n4053 , R_15d7_11c6ab98 );
buf ( n4054 , R_fb8_156b7bb8 );
buf ( n4055 , R_8c4_117f8018 );
buf ( n4056 , R_efc_12fc14b8 );
buf ( n4057 , R_980_13d2b9f8 );
buf ( n4058 , R_151b_14a153b8 );
buf ( n4059 , R_15be_11629bb8 );
buf ( n4060 , R_8dd_13d1dcb8 );
buf ( n4061 , R_f9f_13bf1858 );
buf ( n4062 , R_8a4_13cd4418 );
buf ( n4063 , R_15f7_117ea878 );
buf ( n4064 , R_ec3_14a15e58 );
buf ( n4065 , R_fd8_117f1718 );
buf ( n4066 , R_14e2_13ddc478 );
buf ( n4067 , R_9b9_1008a458 );
buf ( n4068 , R_1580_123b3958 );
buf ( n4069 , R_f61_14867318 );
buf ( n4070 , R_942_140b3a18 );
buf ( n4071 , R_91b_156b0d18 );
buf ( n4072 , R_f3a_1007f4b8 );
buf ( n4073 , R_1559_13c234f8 );
buf ( n4074 , R_1441_13ded378 );
buf ( n4075 , R_a5a_13c097d8 );
buf ( n4076 , R_e22_117eccb8 );
buf ( n4077 , R_1079_13beb6d8 );
buf ( n4078 , R_803_140b8158 );
buf ( n4079 , R_1698_15811998 );
buf ( n4080 , R_1a60_14b1b778 );
buf ( n4081 , R_1987_140b7cf8 );
buf ( n4082 , R_72a_158127f8 );
buf ( n4083 , R_b33_13d2aaf8 );
buf ( n4084 , R_d49_15811678 );
buf ( n4085 , R_1771_17009c68 );
buf ( n4086 , R_1368_1587e9b8 );
buf ( n4087 , R_1152_13c0bd58 );
buf ( n4088 , R_5d5_123be038 );
buf ( n4089 , R_18c6_13d3a1b8 );
buf ( n4090 , R_bf4_1587cb18 );
buf ( n4091 , R_12a7_15817cf8 );
buf ( n4092 , R_1213_140ad078 );
buf ( n4093 , R_c88_17017cc8 );
buf ( n4094 , R_1832_123bc2d8 );
buf ( n4095 , R_669_116322b8 );
buf ( n4096 , R_769_150da558 );
buf ( n4097 , R_d88_117f22f8 );
buf ( n4098 , R_1732_123b2558 );
buf ( n4099 , R_13a7_13c08ab8 );
buf ( n4100 , R_1113_123c1e18 );
buf ( n4101 , R_19c6_13cd18f8 );
buf ( n4102 , R_af4_1580feb8 );
buf ( n4103 , R_b3f_13c22198 );
buf ( n4104 , R_71e_140aec98 );
buf ( n4105 , R_197b_123c14b8 );
buf ( n4106 , R_177d_17012728 );
buf ( n4107 , R_d3d_13c053b8 );
buf ( n4108 , R_115e_15885c18 );
buf ( n4109 , R_135c_13cda3b8 );
buf ( n4110 , R_12d7_13cd2578 );
buf ( n4111 , R_1802_13d3fbb8 );
buf ( n4112 , R_5a5_13d375f8 );
buf ( n4113 , R_cb8_11c6c218 );
buf ( n4114 , R_bc4_14b2a138 );
buf ( n4115 , R_699_15888ff8 );
buf ( n4116 , R_18f6_124c27d8 );
buf ( n4117 , R_11e3_1162fa18 );
buf ( n4118 , R_b67_13cd4f58 );
buf ( n4119 , R_17a5_116334d8 );
buf ( n4120 , R_1334_13cd5598 );
buf ( n4121 , R_6f6_117f1858 );
buf ( n4122 , R_1186_11635d78 );
buf ( n4123 , R_1953_117eb6d8 );
buf ( n4124 , R_d15_123b5578 );
buf ( n4125 , R_603_13ddbe38 );
buf ( n4126 , R_c22_117f71b8 );
buf ( n4127 , R_1241_1162a5b8 );
buf ( n4128 , R_1860_13ccdf78 );
buf ( n4129 , R_1898_11c6bb38 );
buf ( n4130 , R_1279_15887478 );
buf ( n4131 , R_c5a_14a16538 );
buf ( n4132 , R_63b_15883cd8 );
buf ( n4133 , R_10bb_1587d8d8 );
buf ( n4134 , R_16da_124c3db8 );
buf ( n4135 , R_1a1e_11c6ed38 );
buf ( n4136 , R_13ff_17012c28 );
buf ( n4137 , R_de0_13d3abb8 );
buf ( n4138 , R_7c1_156b3bf8 );
buf ( n4139 , R_a9c_1162e4d8 );
buf ( n4140 , R_18d0_117f1358 );
buf ( n4141 , R_5cb_12fc0d38 );
buf ( n4142 , R_12b1_124c38b8 );
buf ( n4143 , R_bea_13ccb098 );
buf ( n4144 , R_c92_150e3838 );
buf ( n4145 , R_1209_14a0aa58 );
buf ( n4146 , R_673_14a13fb8 );
buf ( n4147 , R_1828_1580ab98 );
buf ( n4148 , R_14b6_1587d1f8 );
buf ( n4149 , R_878_13c100d8 );
buf ( n4150 , R_1004_156ab318 );
buf ( n4151 , R_e97_14866918 );
buf ( n4152 , R_9e5_1587d6f8 );
buf ( n4153 , R_1623_13b96178 );
buf ( n4154 , R_11d1_1162f6f8 );
buf ( n4155 , R_cca_117eebf8 );
buf ( n4156 , R_593_117ee0b8 );
buf ( n4157 , R_17f0_100833d8 );
buf ( n4158 , R_1908_1162f5b8 );
buf ( n4159 , R_6ab_13ccbe58 );
buf ( n4160 , R_bb2_15810278 );
buf ( n4161 , R_12e9_13d26818 );
buf ( n4162 , R_f89_13d51738 );
buf ( n4163 , R_96a_1587c258 );
buf ( n4164 , R_8f3_10082b18 );
buf ( n4165 , R_f12_1162b2d8 );
buf ( n4166 , R_15a8_14b25db8 );
buf ( n4167 , R_1531_13c0ac78 );
buf ( n4168 , R_12c2_13d4e2b8 );
buf ( n4169 , R_5ba_13b94d78 );
buf ( n4170 , R_ca3_13ddaa38 );
buf ( n4171 , R_bd9_13d54398 );
buf ( n4172 , R_684_117f5a98 );
buf ( n4173 , R_11f8_13bf1538 );
buf ( n4174 , R_18e1_17010388 );
buf ( n4175 , R_1817_1580f9b8 );
buf ( n4176 , R_a7f_117ebc78 );
buf ( n4177 , R_1a3b_13d275d8 );
buf ( n4178 , R_109e_14a11538 );
buf ( n4179 , R_16bd_117eb9f8 );
buf ( n4180 , R_141c_123b3f98 );
buf ( n4181 , R_dfd_1700cf08 );
buf ( n4182 , R_7de_15881ed8 );
buf ( n4183 , R_f95_13d51058 );
buf ( n4184 , R_1525_140b5598 );
buf ( n4185 , R_976_140b2f78 );
buf ( n4186 , R_8e7_13dd8ff8 );
buf ( n4187 , R_15b4_13dee598 );
buf ( n4188 , R_f06_14b29238 );
buf ( n4189 , R_899_13d5a8d8 );
buf ( n4190 , R_1602_13c28ef8 );
buf ( n4191 , R_eb8_13c1c0b8 );
buf ( n4192 , R_fe3_13ccb598 );
buf ( n4193 , R_14d7_14a0fb98 );
buf ( n4194 , R_9c4_123c1a58 );
buf ( n4195 , R_1599_13bf40f8 );
buf ( n4196 , R_f7a_13d510f8 );
buf ( n4197 , R_95b_15813838 );
buf ( n4198 , R_902_14a0aff8 );
buf ( n4199 , R_f21_15812398 );
buf ( n4200 , R_1540_14871458 );
buf ( n4201 , R_1321_156b1038 );
buf ( n4202 , R_1199_13cd3bf8 );
buf ( n4203 , R_6e3_140b27f8 );
buf ( n4204 , R_55b_13d54f78 );
buf ( n4205 , R_1940_117ed758 );
buf ( n4206 , R_17b8_14b1ca38 );
buf ( n4207 , R_d02_14b21998 );
buf ( n4208 , R_b7a_140b8298 );
buf ( n4209 , R_ed5_123b27d8 );
buf ( n4210 , R_15e5_13d3e0d8 );
buf ( n4211 , R_14f4_1580cad8 );
buf ( n4212 , R_fc6_117f2078 );
buf ( n4213 , R_8b6_12fbe7b8 );
buf ( n4214 , R_9a7_13dd6118 );
buf ( n4215 , R_d96_13c23778 );
buf ( n4216 , R_13b5_124c31d8 );
buf ( n4217 , R_19d4_123b6798 );
buf ( n4218 , R_1724_117edcf8 );
buf ( n4219 , R_1105_158130b8 );
buf ( n4220 , R_ae6_14873e38 );
buf ( n4221 , R_777_17012228 );
buf ( n4222 , R_1581_10080458 );
buf ( n4223 , R_f62_13ccaff8 );
buf ( n4224 , R_943_156b21b8 );
buf ( n4225 , R_91a_13d23e38 );
buf ( n4226 , R_f39_117f5778 );
buf ( n4227 , R_1558_15ffb2c8 );
buf ( n4228 , R_88a_15880c18 );
buf ( n4229 , R_ff2_13d42638 );
buf ( n4230 , R_ea9_15810ef8 );
buf ( n4231 , R_9d3_12fc1e18 );
buf ( n4232 , R_14c8_13d50d38 );
buf ( n4233 , R_1611_13df2b98 );
buf ( n4234 , R_5c2_150db138 );
buf ( n4235 , R_12ba_158138d8 );
buf ( n4236 , R_be1_10082898 );
buf ( n4237 , R_c9b_13b977f8 );
buf ( n4238 , R_1200_13d3d778 );
buf ( n4239 , R_67c_13dec978 );
buf ( n4240 , R_181f_156b4558 );
buf ( n4241 , R_18d9_117f3e78 );
buf ( n4242 , R_1743_15ff3488 );
buf ( n4243 , R_758_13cd0ef8 );
buf ( n4244 , R_1124_14a17d98 );
buf ( n4245 , R_d77_14a0ca38 );
buf ( n4246 , R_1396_156ace98 );
buf ( n4247 , R_b05_13d37d78 );
buf ( n4248 , R_19b5_13cd3c98 );
buf ( n4249 , R_d9f_1580b818 );
buf ( n4250 , R_13be_156af5f8 );
buf ( n4251 , R_19dd_13d56238 );
buf ( n4252 , R_171b_14a0ac38 );
buf ( n4253 , R_10fc_13d52c78 );
buf ( n4254 , R_add_17015ce8 );
buf ( n4255 , R_780_13cd31f8 );
buf ( n4256 , R_198a_12fc1af8 );
buf ( n4257 , R_72d_13d467d8 );
buf ( n4258 , R_b30_156ac358 );
buf ( n4259 , R_d4c_11633d98 );
buf ( n4260 , R_176e_12fbe678 );
buf ( n4261 , R_136b_15810638 );
buf ( n4262 , R_114f_123ba1b8 );
buf ( n4263 , R_119d_123ba578 );
buf ( n4264 , R_55f_13cce658 );
buf ( n4265 , R_6df_13bf5ef8 );
buf ( n4266 , R_131d_14a11c18 );
buf ( n4267 , R_17bc_15886d98 );
buf ( n4268 , R_b7e_123b7eb8 );
buf ( n4269 , R_cfe_123b7418 );
buf ( n4270 , R_193c_123b6298 );
buf ( n4271 , R_b42_116296b8 );
buf ( n4272 , R_71b_13cd8fb8 );
buf ( n4273 , R_1978_1587e698 );
buf ( n4274 , R_1780_1587b718 );
buf ( n4275 , R_d3a_117f6678 );
buf ( n4276 , R_1161_13beb3b8 );
buf ( n4277 , R_1359_11c6d9d8 );
buf ( n4278 , R_1325_156ac178 );
buf ( n4279 , R_6e7_15882fb8 );
buf ( n4280 , R_557_15885f38 );
buf ( n4281 , R_1195_116363b8 );
buf ( n4282 , R_1944_124c2918 );
buf ( n4283 , R_d06_13dde818 );
buf ( n4284 , R_b76_13d41b98 );
buf ( n4285 , R_17b4_13d29ab8 );
buf ( n4286 , R_1020_117ed258 );
buf ( n4287 , R_85c_1580fc38 );
buf ( n4288 , R_149a_13bf0ef8 );
buf ( n4289 , R_163f_13de4218 );
buf ( n4290 , R_a01_156b1498 );
buf ( n4291 , R_e7b_1486b738 );
buf ( n4292 , R_11c1_123b5618 );
buf ( n4293 , R_cda_156b9878 );
buf ( n4294 , R_1918_15880f38 );
buf ( n4295 , R_583_13cccb78 );
buf ( n4296 , R_17e0_14a15d18 );
buf ( n4297 , R_6bb_117f2398 );
buf ( n4298 , R_ba2_14a0e5b8 );
buf ( n4299 , R_12f9_13d5c9f8 );
buf ( n4300 , R_5ee_12fc0c98 );
buf ( n4301 , R_c0d_13b93fb8 );
buf ( n4302 , R_122c_14b217b8 );
buf ( n4303 , R_18ad_13cd6358 );
buf ( n4304 , R_184b_1486d3f8 );
buf ( n4305 , R_128e_13b91a38 );
buf ( n4306 , R_c6f_150e83d8 );
buf ( n4307 , R_650_116346f8 );
buf ( n4308 , R_5e0_13df04d8 );
buf ( n4309 , R_bff_123b92b8 );
buf ( n4310 , R_18bb_11c6f698 );
buf ( n4311 , R_121e_14b1d438 );
buf ( n4312 , R_129c_1007ebf8 );
buf ( n4313 , R_183d_15882e78 );
buf ( n4314 , R_c7d_13c108f8 );
buf ( n4315 , R_65e_13d43998 );
buf ( n4316 , R_75d_156ad118 );
buf ( n4317 , R_173e_148678b8 );
buf ( n4318 , R_d7c_123be998 );
buf ( n4319 , R_111f_14a110d8 );
buf ( n4320 , R_139b_156b35b8 );
buf ( n4321 , R_b00_13ccf558 );
buf ( n4322 , R_19ba_17014d48 );
buf ( n4323 , R_a78_13cd1cb8 );
buf ( n4324 , R_1a42_15817118 );
buf ( n4325 , R_1097_13d240b8 );
buf ( n4326 , R_1423_13c05a98 );
buf ( n4327 , R_16b6_140aab98 );
buf ( n4328 , R_e04_156b17b8 );
buf ( n4329 , R_7e5_14b1e798 );
buf ( n4330 , R_746_170166e8 );
buf ( n4331 , R_1136_13d56558 );
buf ( n4332 , R_d65_1008bb78 );
buf ( n4333 , R_b17_123bcc38 );
buf ( n4334 , R_1384_140b3298 );
buf ( n4335 , R_19a3_117eaa58 );
buf ( n4336 , R_1755_10087258 );
buf ( n4337 , R_c21_1700d4a8 );
buf ( n4338 , R_1240_11630238 );
buf ( n4339 , R_185f_13bf7118 );
buf ( n4340 , R_1899_156b1fd8 );
buf ( n4341 , R_127a_14b28298 );
buf ( n4342 , R_c5b_13d26278 );
buf ( n4343 , R_63c_1587b538 );
buf ( n4344 , R_602_156afff8 );
buf ( n4345 , R_753_116336b8 );
buf ( n4346 , R_1129_13ccc3f8 );
buf ( n4347 , R_d72_13b95e58 );
buf ( n4348 , R_b0a_156ad438 );
buf ( n4349 , R_1391_15886578 );
buf ( n4350 , R_19b0_17014a28 );
buf ( n4351 , R_1748_117eeab8 );
buf ( n4352 , R_e32_13c05c78 );
buf ( n4353 , R_a4a_117e8bb8 );
buf ( n4354 , R_813_11631318 );
buf ( n4355 , R_1069_116369f8 );
buf ( n4356 , R_1688_156b6a38 );
buf ( n4357 , R_1451_150e6b78 );
buf ( n4358 , R_cdf_150dfa58 );
buf ( n4359 , R_11bc_11c6a9b8 );
buf ( n4360 , R_191d_13c10678 );
buf ( n4361 , R_57e_1162f338 );
buf ( n4362 , R_6c0_13b98c98 );
buf ( n4363 , R_17db_117f6858 );
buf ( n4364 , R_12fe_116291b8 );
buf ( n4365 , R_b9d_14872678 );
buf ( n4366 , R_1349_13d26db8 );
buf ( n4367 , R_b52_1162a978 );
buf ( n4368 , R_1790_117e9798 );
buf ( n4369 , R_70b_17018808 );
buf ( n4370 , R_1968_13bf0318 );
buf ( n4371 , R_d2a_15fef568 );
buf ( n4372 , R_1171_117f5278 );
buf ( n4373 , R_192b_11633cf8 );
buf ( n4374 , R_11ae_123bc238 );
buf ( n4375 , R_570_117ec218 );
buf ( n4376 , R_6ce_13dee1d8 );
buf ( n4377 , R_130c_15ff67c8 );
buf ( n4378 , R_17cd_13b91858 );
buf ( n4379 , R_b8f_14b25b38 );
buf ( n4380 , R_ced_14a0a558 );
buf ( n4381 , R_1582_150e7ed8 );
buf ( n4382 , R_f63_13cca7d8 );
buf ( n4383 , R_944_13d1fab8 );
buf ( n4384 , R_919_123bdf98 );
buf ( n4385 , R_f38_13d26958 );
buf ( n4386 , R_1557_14a16c18 );
buf ( n4387 , R_10ae_123b9358 );
buf ( n4388 , R_16cd_117eee78 );
buf ( n4389 , R_1a2b_140accb8 );
buf ( n4390 , R_140c_11c6f058 );
buf ( n4391 , R_ded_14a14738 );
buf ( n4392 , R_7ce_13d45d38 );
buf ( n4393 , R_a8f_17014de8 );
buf ( n4394 , R_10a5_13d564b8 );
buf ( n4395 , R_16c4_1580f878 );
buf ( n4396 , R_1a34_14a19558 );
buf ( n4397 , R_1415_158165d8 );
buf ( n4398 , R_df6_156b2bb8 );
buf ( n4399 , R_7d7_13c29998 );
buf ( n4400 , R_a86_123bc0f8 );
buf ( n4401 , R_165b_13de0898 );
buf ( n4402 , R_840_156b26b8 );
buf ( n4403 , R_a1d_14a15778 );
buf ( n4404 , R_147e_11638078 );
buf ( n4405 , R_103c_140b0ef8 );
buf ( n4406 , R_e5f_150e3d38 );
buf ( n4407 , R_11c6_13def038 );
buf ( n4408 , R_cd5_13cd09f8 );
buf ( n4409 , R_588_13de09d8 );
buf ( n4410 , R_1913_13beef18 );
buf ( n4411 , R_17e5_150de518 );
buf ( n4412 , R_6b6_13d519b8 );
buf ( n4413 , R_ba7_13d2ca38 );
buf ( n4414 , R_12f4_11c6ca38 );
buf ( n4415 , R_19e8_15888e18 );
buf ( n4416 , R_1710_13bf6718 );
buf ( n4417 , R_10f1_124c52f8 );
buf ( n4418 , R_ad2_156b8658 );
buf ( n4419 , R_78b_1162ddf8 );
buf ( n4420 , R_daa_1008ced8 );
buf ( n4421 , R_13c9_13de18d8 );
buf ( n4422 , R_11a1_117e91f8 );
buf ( n4423 , R_563_13d1ea78 );
buf ( n4424 , R_6db_13dd91d8 );
buf ( n4425 , R_1319_117f10d8 );
buf ( n4426 , R_17c0_15ff4888 );
buf ( n4427 , R_b82_13beff58 );
buf ( n4428 , R_cfa_14b21ad8 );
buf ( n4429 , R_1938_13df6ab8 );
buf ( n4430 , R_82a_14a0cfd8 );
buf ( n4431 , R_a33_11c70278 );
buf ( n4432 , R_1468_158803f8 );
buf ( n4433 , R_1052_117f42d8 );
buf ( n4434 , R_1671_13dd6898 );
buf ( n4435 , R_e49_15ff8f28 );
buf ( n4436 , R_1329_14a16ad8 );
buf ( n4437 , R_6eb_13d45b58 );
buf ( n4438 , R_1191_15881618 );
buf ( n4439 , R_1948_13c26a18 );
buf ( n4440 , R_d0a_158820b8 );
buf ( n4441 , R_b72_13c103f8 );
buf ( n4442 , R_17b0_13decf18 );
buf ( n4443 , R_a36_13b92438 );
buf ( n4444 , R_827_123b8f98 );
buf ( n4445 , R_1055_11635738 );
buf ( n4446 , R_1465_14a18ab8 );
buf ( n4447 , R_1674_11636c78 );
buf ( n4448 , R_e46_15884098 );
buf ( n4449 , R_851_11635238 );
buf ( n4450 , R_148f_13df4358 );
buf ( n4451 , R_164a_13c1e318 );
buf ( n4452 , R_a0c_100899b8 );
buf ( n4453 , R_e70_117ec538 );
buf ( n4454 , R_102b_13d38d18 );
buf ( n4455 , R_198d_156b4378 );
buf ( n4456 , R_730_123bb518 );
buf ( n4457 , R_b2d_124c29b8 );
buf ( n4458 , R_d4f_13cd15d8 );
buf ( n4459 , R_176b_150e5bd8 );
buf ( n4460 , R_136e_15ff6b88 );
buf ( n4461 , R_114c_140b06d8 );
buf ( n4462 , R_16f5_13d39b78 );
buf ( n4463 , R_1a03_14b23338 );
buf ( n4464 , R_10d6_150df4b8 );
buf ( n4465 , R_13e4_13cd99b8 );
buf ( n4466 , R_ab7_1700b748 );
buf ( n4467 , R_dc5_15ff3f28 );
buf ( n4468 , R_7a6_150dad78 );
buf ( n4469 , R_1a05_1162d498 );
buf ( n4470 , R_13e6_1486e578 );
buf ( n4471 , R_dc7_13cd2398 );
buf ( n4472 , R_16f3_10088bf8 );
buf ( n4473 , R_7a8_13beac38 );
buf ( n4474 , R_10d4_13d1de98 );
buf ( n4475 , R_ab5_13df25f8 );
buf ( n4476 , R_82d_13c24b78 );
buf ( n4477 , R_a30_117ef9b8 );
buf ( n4478 , R_146b_150da9b8 );
buf ( n4479 , R_104f_170118c8 );
buf ( n4480 , R_e4c_13ddfd58 );
buf ( n4481 , R_166e_123be3f8 );
buf ( n4482 , R_73e_15883878 );
buf ( n4483 , R_b1f_11631098 );
buf ( n4484 , R_d5d_11636778 );
buf ( n4485 , R_137c_11634e78 );
buf ( n4486 , R_175d_13df13d8 );
buf ( n4487 , R_199b_150dc8f8 );
buf ( n4488 , R_113e_10081ad8 );
buf ( n4489 , R_b45_13cce978 );
buf ( n4490 , R_718_123b4fd8 );
buf ( n4491 , R_1975_13deedb8 );
buf ( n4492 , R_1783_15817e38 );
buf ( n4493 , R_d37_13d26d18 );
buf ( n4494 , R_1164_13df29b8 );
buf ( n4495 , R_1356_15884958 );
buf ( n4496 , R_16f7_140b9558 );
buf ( n4497 , R_10d8_13d55158 );
buf ( n4498 , R_ab9_14a16358 );
buf ( n4499 , R_1a01_14a0bf98 );
buf ( n4500 , R_7a4_13cca698 );
buf ( n4501 , R_13e2_13d50338 );
buf ( n4502 , R_dc3_13d5b918 );
buf ( n4503 , R_1509_13c080b8 );
buf ( n4504 , R_15d0_13d5d7b8 );
buf ( n4505 , R_fb1_17011fa8 );
buf ( n4506 , R_8cb_1162afb8 );
buf ( n4507 , R_992_158117b8 );
buf ( n4508 , R_eea_158843b8 );
buf ( n4509 , R_1a07_15817f78 );
buf ( n4510 , R_13e8_13d57458 );
buf ( n4511 , R_dc9_13dedb98 );
buf ( n4512 , R_7aa_14a113f8 );
buf ( n4513 , R_ab3_13ccea18 );
buf ( n4514 , R_16f1_13c2b298 );
buf ( n4515 , R_10d2_14a0f4b8 );
buf ( n4516 , R_84a_1700eee8 );
buf ( n4517 , R_1651_100849b8 );
buf ( n4518 , R_1488_15811858 );
buf ( n4519 , R_a13_117f7ed8 );
buf ( n4520 , R_e69_14b24ff8 );
buf ( n4521 , R_1032_15884638 );
buf ( n4522 , R_1434_15884a98 );
buf ( n4523 , R_a67_1587c9d8 );
buf ( n4524 , R_e15_117f6538 );
buf ( n4525 , R_1086_158844f8 );
buf ( n4526 , R_16a5_1587d018 );
buf ( n4527 , R_7f6_14a10318 );
buf ( n4528 , R_1a53_11c70b38 );
buf ( n4529 , R_f7b_13c24f38 );
buf ( n4530 , R_95c_13b8ad78 );
buf ( n4531 , R_901_15ff0dc8 );
buf ( n4532 , R_f20_11633078 );
buf ( n4533 , R_153f_140abef8 );
buf ( n4534 , R_159a_13d58d58 );
buf ( n4535 , R_1a20_117f5638 );
buf ( n4536 , R_1401_14a19918 );
buf ( n4537 , R_de2_123bef38 );
buf ( n4538 , R_7c3_14a0f058 );
buf ( n4539 , R_a9a_15816f38 );
buf ( n4540 , R_10b9_15ff6908 );
buf ( n4541 , R_16d8_14b209f8 );
buf ( n4542 , R_1583_13b8ba98 );
buf ( n4543 , R_f64_123b9718 );
buf ( n4544 , R_945_123bcaf8 );
buf ( n4545 , R_918_13c20ed8 );
buf ( n4546 , R_f37_158875b8 );
buf ( n4547 , R_1556_140b5db8 );
buf ( n4548 , R_a39_17016d28 );
buf ( n4549 , R_824_140b4b98 );
buf ( n4550 , R_1058_13b8c7b8 );
buf ( n4551 , R_1462_13d228f8 );
buf ( n4552 , R_1677_1008aef8 );
buf ( n4553 , R_e43_140ab8b8 );
buf ( n4554 , R_123f_12fc2458 );
buf ( n4555 , R_185e_100815d8 );
buf ( n4556 , R_189a_15ff14a8 );
buf ( n4557 , R_127b_13de1a18 );
buf ( n4558 , R_c5c_140b8518 );
buf ( n4559 , R_63d_13df0438 );
buf ( n4560 , R_601_14a12c58 );
buf ( n4561 , R_c20_1486b7d8 );
buf ( n4562 , R_15fd_156b4c38 );
buf ( n4563 , R_ebd_117f1ad8 );
buf ( n4564 , R_fde_13d429f8 );
buf ( n4565 , R_14dc_13ddc5b8 );
buf ( n4566 , R_9bf_15ff2128 );
buf ( n4567 , R_89e_123bbdd8 );
buf ( n4568 , R_16f9_13cd6218 );
buf ( n4569 , R_10da_14a0d4d8 );
buf ( n4570 , R_abb_14b262b8 );
buf ( n4571 , R_7a2_13de1fb8 );
buf ( n4572 , R_dc1_13c211f8 );
buf ( n4573 , R_13e0_1486e4d8 );
buf ( n4574 , R_19ff_123b42b8 );
buf ( n4575 , R_1739_15ff78a8 );
buf ( n4576 , R_d81_140ad4d8 );
buf ( n4577 , R_111a_13d42ef8 );
buf ( n4578 , R_13a0_117f2bb8 );
buf ( n4579 , R_afb_13bf4af8 );
buf ( n4580 , R_19bf_117f5e58 );
buf ( n4581 , R_762_156b33d8 );
buf ( n4582 , R_1a09_1162d358 );
buf ( n4583 , R_13ea_1580dc58 );
buf ( n4584 , R_dcb_1162f798 );
buf ( n4585 , R_7ac_13c08838 );
buf ( n4586 , R_ab1_150e1b78 );
buf ( n4587 , R_10d0_150e7938 );
buf ( n4588 , R_16ef_14a136f8 );
buf ( n4589 , R_a6c_123b7378 );
buf ( n4590 , R_142f_117f79d8 );
buf ( n4591 , R_108b_156b83d8 );
buf ( n4592 , R_e10_14a0b4f8 );
buf ( n4593 , R_16aa_150e47d8 );
buf ( n4594 , R_7f1_123bc378 );
buf ( n4595 , R_1a4e_123b60b8 );
buf ( n4596 , R_5b2_1486f018 );
buf ( n4597 , R_cab_15fee028 );
buf ( n4598 , R_bd1_1587dfb8 );
buf ( n4599 , R_68c_123c1b98 );
buf ( n4600 , R_11f0_13cd3a18 );
buf ( n4601 , R_18e9_13b98a18 );
buf ( n4602 , R_180f_13c1cbf8 );
buf ( n4603 , R_12ca_14a13dd8 );
buf ( n4604 , R_1000_13d4e858 );
buf ( n4605 , R_e9b_13cd5f98 );
buf ( n4606 , R_9e1_13bea878 );
buf ( n4607 , R_161f_10080098 );
buf ( n4608 , R_14ba_1580ba98 );
buf ( n4609 , R_87c_13dee6d8 );
buf ( n4610 , R_830_1008cc58 );
buf ( n4611 , R_a2d_13d43f38 );
buf ( n4612 , R_146e_17010ba8 );
buf ( n4613 , R_104c_13d1f658 );
buf ( n4614 , R_e4f_13ccef18 );
buf ( n4615 , R_166b_116345b8 );
buf ( n4616 , R_ff7_13c0cf78 );
buf ( n4617 , R_ea4_117ea738 );
buf ( n4618 , R_9d8_156b6ad8 );
buf ( n4619 , R_1616_17009da8 );
buf ( n4620 , R_14c3_116384d8 );
buf ( n4621 , R_885_13de02f8 );
buf ( n4622 , R_11b7_11c6de38 );
buf ( n4623 , R_1922_13c26018 );
buf ( n4624 , R_579_13d5d358 );
buf ( n4625 , R_6c5_13d59398 );
buf ( n4626 , R_17d6_11c6d258 );
buf ( n4627 , R_1303_156b3d38 );
buf ( n4628 , R_b98_14b1aeb8 );
buf ( n4629 , R_ce4_117f17b8 );
buf ( n4630 , R_96b_15816c18 );
buf ( n4631 , R_8f2_158891d8 );
buf ( n4632 , R_f11_124c3598 );
buf ( n4633 , R_15a9_1007e0b8 );
buf ( n4634 , R_1530_13c1c5b8 );
buf ( n4635 , R_f8a_1580da78 );
buf ( n4636 , R_5ab_13d20b98 );
buf ( n4637 , R_cb2_15883eb8 );
buf ( n4638 , R_bca_1162ecf8 );
buf ( n4639 , R_693_1580e978 );
buf ( n4640 , R_18f0_14868178 );
buf ( n4641 , R_11e9_12fc0518 );
buf ( n4642 , R_12d1_15ff4388 );
buf ( n4643 , R_1808_117ec998 );
buf ( n4644 , R_112e_124c40d8 );
buf ( n4645 , R_d6d_10080278 );
buf ( n4646 , R_b0f_150e1e98 );
buf ( n4647 , R_138c_14a12938 );
buf ( n4648 , R_19ab_1486d5d8 );
buf ( n4649 , R_174d_13c05318 );
buf ( n4650 , R_74e_117e9dd8 );
buf ( n4651 , R_5d4_1587e918 );
buf ( n4652 , R_18c7_117ed7f8 );
buf ( n4653 , R_bf3_158826f8 );
buf ( n4654 , R_12a8_140b92d8 );
buf ( n4655 , R_1212_13debed8 );
buf ( n4656 , R_c89_15886078 );
buf ( n4657 , R_1831_13b99eb8 );
buf ( n4658 , R_66a_117f7c58 );
buf ( n4659 , R_16fb_13d39a38 );
buf ( n4660 , R_10dc_140acad8 );
buf ( n4661 , R_abd_12fbf938 );
buf ( n4662 , R_7a0_1162cef8 );
buf ( n4663 , R_dbf_13d1dd58 );
buf ( n4664 , R_13de_13bf51d8 );
buf ( n4665 , R_19fd_13c22cd8 );
buf ( n4666 , R_a62_11630378 );
buf ( n4667 , R_e1a_13d29f18 );
buf ( n4668 , R_1081_156ae298 );
buf ( n4669 , R_7fb_13c27c38 );
buf ( n4670 , R_16a0_1007f9b8 );
buf ( n4671 , R_1a58_123b6a18 );
buf ( n4672 , R_1439_11637c18 );
buf ( n4673 , R_1511_1162c778 );
buf ( n4674 , R_15c8_10085a98 );
buf ( n4675 , R_8d3_15fefba8 );
buf ( n4676 , R_fa9_150dc218 );
buf ( n4677 , R_ef2_13d3af78 );
buf ( n4678 , R_98a_11629578 );
buf ( n4679 , R_151a_15ff8d48 );
buf ( n4680 , R_15bf_15ff4f68 );
buf ( n4681 , R_8dc_13dd7b58 );
buf ( n4682 , R_fa0_1162a838 );
buf ( n4683 , R_efb_13ccc2b8 );
buf ( n4684 , R_981_156acad8 );
buf ( n4685 , R_133f_11636ef8 );
buf ( n4686 , R_179a_13ccf918 );
buf ( n4687 , R_701_13dd6438 );
buf ( n4688 , R_195e_15817578 );
buf ( n4689 , R_117b_156b5f98 );
buf ( n4690 , R_d20_1162aa18 );
buf ( n4691 , R_b5c_116370d8 );
buf ( n4692 , R_c0c_13d3f7f8 );
buf ( n4693 , R_122b_117ec498 );
buf ( n4694 , R_18ae_13d39998 );
buf ( n4695 , R_184a_124c54d8 );
buf ( n4696 , R_128f_123b97b8 );
buf ( n4697 , R_c70_15885998 );
buf ( n4698 , R_651_14a122f8 );
buf ( n4699 , R_5ed_13cccad8 );
buf ( n4700 , R_1a0b_1486ee38 );
buf ( n4701 , R_13ec_117f2758 );
buf ( n4702 , R_dcd_13d1e438 );
buf ( n4703 , R_7ae_13d3c058 );
buf ( n4704 , R_aaf_140af698 );
buf ( n4705 , R_10ce_11637538 );
buf ( n4706 , R_16ed_156af558 );
buf ( n4707 , R_a55_12fbef38 );
buf ( n4708 , R_e27_13d405b8 );
buf ( n4709 , R_1074_14b1a878 );
buf ( n4710 , R_808_13c22c38 );
buf ( n4711 , R_1693_13cd4558 );
buf ( n4712 , R_1a65_1587f8b8 );
buf ( n4713 , R_1446_1587eff8 );
buf ( n4714 , R_a3c_150e6038 );
buf ( n4715 , R_821_117f1b78 );
buf ( n4716 , R_105b_13cd2f78 );
buf ( n4717 , R_145f_13b8d398 );
buf ( n4718 , R_167a_13df45d8 );
buf ( n4719 , R_e40_13c26f18 );
buf ( n4720 , R_1584_1580b318 );
buf ( n4721 , R_f65_13d3b5b8 );
buf ( n4722 , R_946_14a10a98 );
buf ( n4723 , R_917_117f5458 );
buf ( n4724 , R_f36_14a118f8 );
buf ( n4725 , R_1555_15815638 );
buf ( n4726 , R_cd0_117f6d58 );
buf ( n4727 , R_58d_1587f3b8 );
buf ( n4728 , R_17ea_15ffadc8 );
buf ( n4729 , R_190e_13bf3d38 );
buf ( n4730 , R_6b1_15ffc808 );
buf ( n4731 , R_bac_13c0a098 );
buf ( n4732 , R_12ef_14b277f8 );
buf ( n4733 , R_11cb_15ff6f48 );
buf ( n4734 , R_977_1580b1d8 );
buf ( n4735 , R_8e6_1580c0d8 );
buf ( n4736 , R_15b5_14866f58 );
buf ( n4737 , R_f05_123b8ef8 );
buf ( n4738 , R_f96_15885538 );
buf ( n4739 , R_1524_1162d178 );
buf ( n4740 , R_11a5_156b5138 );
buf ( n4741 , R_567_13bf17b8 );
buf ( n4742 , R_6d7_12fc12d8 );
buf ( n4743 , R_1315_123b2698 );
buf ( n4744 , R_17c4_13ccc718 );
buf ( n4745 , R_b86_123b9a38 );
buf ( n4746 , R_cf6_14b29738 );
buf ( n4747 , R_1934_123bf7f8 );
buf ( n4748 , R_1338_116375d8 );
buf ( n4749 , R_6fa_13bec218 );
buf ( n4750 , R_1182_13c1c658 );
buf ( n4751 , R_1957_13d3ec18 );
buf ( n4752 , R_d19_13def3f8 );
buf ( n4753 , R_b63_15ffbb88 );
buf ( n4754 , R_17a1_117f24d8 );
buf ( n4755 , R_132d_1587ce38 );
buf ( n4756 , R_6ef_158893b8 );
buf ( n4757 , R_118d_124c3958 );
buf ( n4758 , R_194c_1587cbb8 );
buf ( n4759 , R_d0e_13c10998 );
buf ( n4760 , R_b6e_117ef5f8 );
buf ( n4761 , R_17ac_1486cb38 );
buf ( n4762 , R_12b2_156ab458 );
buf ( n4763 , R_be9_14867638 );
buf ( n4764 , R_c93_14a12258 );
buf ( n4765 , R_1208_13bec358 );
buf ( n4766 , R_674_123c0018 );
buf ( n4767 , R_1827_13c01b78 );
buf ( n4768 , R_18d1_117e98d8 );
buf ( n4769 , R_5ca_13ccca38 );
buf ( n4770 , R_16fd_13bf4378 );
buf ( n4771 , R_10de_140b68f8 );
buf ( n4772 , R_abf_13befd78 );
buf ( n4773 , R_79e_15817b18 );
buf ( n4774 , R_dbd_117f2b18 );
buf ( n4775 , R_13dc_13d1ce58 );
buf ( n4776 , R_19fb_150e3978 );
buf ( n4777 , R_858_150dae18 );
buf ( n4778 , R_1496_13b8b098 );
buf ( n4779 , R_1643_1162c278 );
buf ( n4780 , R_a05_117f4cd8 );
buf ( n4781 , R_e77_1486b878 );
buf ( n4782 , R_1024_11635058 );
buf ( n4783 , R_733_10086998 );
buf ( n4784 , R_b2a_150dd2f8 );
buf ( n4785 , R_d52_1580c498 );
buf ( n4786 , R_1768_15813b58 );
buf ( n4787 , R_1371_156b10d8 );
buf ( n4788 , R_1149_156aff58 );
buf ( n4789 , R_1990_117f1df8 );
buf ( n4790 , R_185d_1162a0b8 );
buf ( n4791 , R_189b_123bccd8 );
buf ( n4792 , R_127c_1580f198 );
buf ( n4793 , R_c5d_13bf88d8 );
buf ( n4794 , R_63e_170163c8 );
buf ( n4795 , R_600_150e8798 );
buf ( n4796 , R_c1f_117ebdb8 );
buf ( n4797 , R_123e_13ccb318 );
buf ( n4798 , R_bfe_17018b28 );
buf ( n4799 , R_18bc_123b9df8 );
buf ( n4800 , R_121d_11632718 );
buf ( n4801 , R_129d_117f6998 );
buf ( n4802 , R_183c_14b21498 );
buf ( n4803 , R_c7e_14a0d6b8 );
buf ( n4804 , R_65f_14874978 );
buf ( n4805 , R_5df_13c24178 );
buf ( n4806 , R_833_117f3dd8 );
buf ( n4807 , R_a2a_14869bb8 );
buf ( n4808 , R_1471_140adbb8 );
buf ( n4809 , R_1049_11636138 );
buf ( n4810 , R_e52_13d4e498 );
buf ( n4811 , R_1668_13b909f8 );
buf ( n4812 , R_15df_14b24c38 );
buf ( n4813 , R_14fa_15ff7128 );
buf ( n4814 , R_fc0_13beba98 );
buf ( n4815 , R_8bc_14a0e338 );
buf ( n4816 , R_9a1_123b5758 );
buf ( n4817 , R_edb_17017048 );
buf ( n4818 , R_1a0d_13ccaaf8 );
buf ( n4819 , R_13ee_13d23398 );
buf ( n4820 , R_dcf_13cccfd8 );
buf ( n4821 , R_7b0_123bf4d8 );
buf ( n4822 , R_aad_14873a78 );
buf ( n4823 , R_10cc_13cd01d8 );
buf ( n4824 , R_16eb_150e81f8 );
buf ( n4825 , R_172d_13cda318 );
buf ( n4826 , R_13ac_116343d8 );
buf ( n4827 , R_110e_14a11998 );
buf ( n4828 , R_19cb_13d3a758 );
buf ( n4829 , R_aef_13d50dd8 );
buf ( n4830 , R_76e_13bf8d38 );
buf ( n4831 , R_d8d_13dd52b8 );
buf ( n4832 , R_715_13b94ff8 );
buf ( n4833 , R_1972_156aa918 );
buf ( n4834 , R_1786_140b5778 );
buf ( n4835 , R_d34_15ff3b68 );
buf ( n4836 , R_1167_1587c7f8 );
buf ( n4837 , R_1353_123c05b8 );
buf ( n4838 , R_b48_15814378 );
buf ( n4839 , R_17fb_11c6bd18 );
buf ( n4840 , R_59e_13cd0098 );
buf ( n4841 , R_cbf_15fed948 );
buf ( n4842 , R_bbd_13b8f418 );
buf ( n4843 , R_18fd_15882798 );
buf ( n4844 , R_6a0_117edbb8 );
buf ( n4845 , R_11dc_150db458 );
buf ( n4846 , R_12de_117e9658 );
buf ( n4847 , R_19db_123b8458 );
buf ( n4848 , R_171d_13d45e78 );
buf ( n4849 , R_10fe_117ebd18 );
buf ( n4850 , R_adf_13ccfcd8 );
buf ( n4851 , R_77e_123bcff8 );
buf ( n4852 , R_d9d_12fc0298 );
buf ( n4853 , R_13bc_13c07cf8 );
buf ( n4854 , R_142a_14a0f2d8 );
buf ( n4855 , R_1090_1486e7f8 );
buf ( n4856 , R_e0b_156b7758 );
buf ( n4857 , R_16af_1486be18 );
buf ( n4858 , R_7ec_123b4038 );
buf ( n4859 , R_1a49_13ccbb38 );
buf ( n4860 , R_a71_117f59f8 );
buf ( n4861 , R_15f2_13d4fe38 );
buf ( n4862 , R_ec8_15883058 );
buf ( n4863 , R_fd3_10088798 );
buf ( n4864 , R_14e7_14b1ce98 );
buf ( n4865 , R_9b4_13bf5b38 );
buf ( n4866 , R_8a9_13c21298 );
buf ( n4867 , R_ece_11634bf8 );
buf ( n4868 , R_15ec_13d3f4d8 );
buf ( n4869 , R_14ed_117f5f98 );
buf ( n4870 , R_fcd_1580d258 );
buf ( n4871 , R_8af_13ddfb78 );
buf ( n4872 , R_9ae_140b18f8 );
buf ( n4873 , R_1501_117f0a98 );
buf ( n4874 , R_15d8_11c6ea18 );
buf ( n4875 , R_fb9_15ff0be8 );
buf ( n4876 , R_8c3_10081498 );
buf ( n4877 , R_99a_15ffaaa8 );
buf ( n4878 , R_ee2_13cd1b78 );
buf ( n4879 , R_1712_11637178 );
buf ( n4880 , R_10f3_14a19238 );
buf ( n4881 , R_ad4_14a0a5f8 );
buf ( n4882 , R_789_140b2cf8 );
buf ( n4883 , R_da8_140b3838 );
buf ( n4884 , R_13c7_13df0ed8 );
buf ( n4885 , R_19e6_11636958 );
buf ( n4886 , R_95d_117f8338 );
buf ( n4887 , R_900_140b74d8 );
buf ( n4888 , R_f1f_1587f1d8 );
buf ( n4889 , R_153e_13d410f8 );
buf ( n4890 , R_159b_1162f658 );
buf ( n4891 , R_f7c_15ffc268 );
buf ( n4892 , R_cc5_13b8c858 );
buf ( n4893 , R_598_17015108 );
buf ( n4894 , R_17f5_13c1c798 );
buf ( n4895 , R_1903_1162d2b8 );
buf ( n4896 , R_6a6_15816df8 );
buf ( n4897 , R_bb7_14a17a78 );
buf ( n4898 , R_12e4_13df4678 );
buf ( n4899 , R_11d6_13cccf38 );
buf ( n4900 , R_a4d_14a159f8 );
buf ( n4901 , R_810_1007f918 );
buf ( n4902 , R_106c_13cd4238 );
buf ( n4903 , R_168b_13d20d78 );
buf ( n4904 , R_144e_17019028 );
buf ( n4905 , R_e2f_123b83b8 );
buf ( n4906 , R_f66_1700e448 );
buf ( n4907 , R_947_13cd36f8 );
buf ( n4908 , R_916_12fbefd8 );
buf ( n4909 , R_f35_13dd5fd8 );
buf ( n4910 , R_1554_13c04918 );
buf ( n4911 , R_1585_117efe18 );
buf ( n4912 , R_16ff_13b95318 );
buf ( n4913 , R_10e0_1580e478 );
buf ( n4914 , R_ac1_13d23078 );
buf ( n4915 , R_79c_1162d8f8 );
buf ( n4916 , R_dbb_1580e018 );
buf ( n4917 , R_13da_123c03d8 );
buf ( n4918 , R_19f9_13cd81f8 );
buf ( n4919 , R_a3f_13c012b8 );
buf ( n4920 , R_81e_140b4cd8 );
buf ( n4921 , R_105e_156ba278 );
buf ( n4922 , R_145c_13ddc0b8 );
buf ( n4923 , R_167d_124c5438 );
buf ( n4924 , R_e3d_15889778 );
buf ( n4925 , R_be0_117ea5f8 );
buf ( n4926 , R_c9c_13b8ed38 );
buf ( n4927 , R_11ff_14a17618 );
buf ( n4928 , R_67d_156b7398 );
buf ( n4929 , R_181e_13c04e18 );
buf ( n4930 , R_18da_13cd38d8 );
buf ( n4931 , R_5c1_13c0a818 );
buf ( n4932 , R_12bb_13b8a918 );
buf ( n4933 , R_ca4_156b1c18 );
buf ( n4934 , R_bd8_117e87f8 );
buf ( n4935 , R_685_13bf38d8 );
buf ( n4936 , R_11f7_10080b38 );
buf ( n4937 , R_18e2_13becfd8 );
buf ( n4938 , R_1816_14b1ff58 );
buf ( n4939 , R_12c3_10083478 );
buf ( n4940 , R_5b9_140b2bb8 );
buf ( n4941 , R_1630_123b9cb8 );
buf ( n4942 , R_e8a_14b1db18 );
buf ( n4943 , R_9f2_10089418 );
buf ( n4944 , R_14a9_156acb78 );
buf ( n4945 , R_1011_12fbe218 );
buf ( n4946 , R_86b_124c4e98 );
buf ( n4947 , R_1726_14869a78 );
buf ( n4948 , R_19d2_13d533f8 );
buf ( n4949 , R_1107_13df9038 );
buf ( n4950 , R_ae8_13bef5f8 );
buf ( n4951 , R_775_158109f8 );
buf ( n4952 , R_d94_12fbf6b8 );
buf ( n4953 , R_13b3_13d40158 );
buf ( n4954 , R_1658_13bf9ff8 );
buf ( n4955 , R_843_150e0458 );
buf ( n4956 , R_1481_117e8e38 );
buf ( n4957 , R_a1a_15fefd88 );
buf ( n4958 , R_1039_13ddba78 );
buf ( n4959 , R_e62_13c23098 );
buf ( n4960 , R_1a0f_13c24038 );
buf ( n4961 , R_13f0_11c6e338 );
buf ( n4962 , R_dd1_13de4a38 );
buf ( n4963 , R_7b2_13bf2898 );
buf ( n4964 , R_aab_13c1cfb8 );
buf ( n4965 , R_10ca_1700ac08 );
buf ( n4966 , R_16e9_15ff3668 );
buf ( n4967 , R_1793_150de018 );
buf ( n4968 , R_708_14a0d258 );
buf ( n4969 , R_1965_13ccb6d8 );
buf ( n4970 , R_1174_11c6c358 );
buf ( n4971 , R_d27_13dee138 );
buf ( n4972 , R_b55_15ffb0e8 );
buf ( n4973 , R_1346_13d3f2f8 );
buf ( n4974 , R_e1f_123b6ab8 );
buf ( n4975 , R_107c_117f4058 );
buf ( n4976 , R_800_13d219f8 );
buf ( n4977 , R_169b_150e49b8 );
buf ( n4978 , R_1a5d_1486e398 );
buf ( n4979 , R_143e_14a19f58 );
buf ( n4980 , R_a5d_15880498 );
buf ( n4981 , R_1a22_15810b38 );
buf ( n4982 , R_1403_124c5398 );
buf ( n4983 , R_de4_117f6498 );
buf ( n4984 , R_7c5_15ffbe08 );
buf ( n4985 , R_a98_1486db78 );
buf ( n4986 , R_10b7_14a17578 );
buf ( n4987 , R_16d6_14a10458 );
buf ( n4988 , R_1a2d_13b8fcd8 );
buf ( n4989 , R_140e_13def718 );
buf ( n4990 , R_def_13d3eb78 );
buf ( n4991 , R_7d0_156b2e38 );
buf ( n4992 , R_a8d_11632678 );
buf ( n4993 , R_10ac_156b5958 );
buf ( n4994 , R_16cb_156b72f8 );
buf ( n4995 , R_1634_17018c68 );
buf ( n4996 , R_9f6_158867f8 );
buf ( n4997 , R_e86_14a183d8 );
buf ( n4998 , R_1015_14b1e6f8 );
buf ( n4999 , R_867_15881398 );
buf ( n5000 , R_14a5_11629ed8 );
buf ( n5001 , R_e8e_150da878 );
buf ( n5002 , R_9ee_13d54618 );
buf ( n5003 , R_162c_13b96c18 );
buf ( n5004 , R_14ad_12fbf618 );
buf ( n5005 , R_86f_15ff83e8 );
buf ( n5006 , R_100d_158136f8 );
buf ( n5007 , R_189c_14a10c78 );
buf ( n5008 , R_127d_11636318 );
buf ( n5009 , R_c5e_15882a18 );
buf ( n5010 , R_63f_156b5b38 );
buf ( n5011 , R_5ff_13d40ab8 );
buf ( n5012 , R_c1e_14a0b958 );
buf ( n5013 , R_123d_13ddd5f8 );
buf ( n5014 , R_185c_11630738 );
buf ( n5015 , R_141e_13b90818 );
buf ( n5016 , R_16bb_123b7d78 );
buf ( n5017 , R_dff_117eeb58 );
buf ( n5018 , R_7e0_13dfacf8 );
buf ( n5019 , R_a7d_123b7af8 );
buf ( n5020 , R_1a3d_156b9cd8 );
buf ( n5021 , R_109c_13b98d38 );
buf ( n5022 , R_cb9_150db638 );
buf ( n5023 , R_bc3_156b6678 );
buf ( n5024 , R_69a_13b8b6d8 );
buf ( n5025 , R_18f7_13b90bd8 );
buf ( n5026 , R_11e2_13d1e4d8 );
buf ( n5027 , R_12d8_13d43718 );
buf ( n5028 , R_1801_13c013f8 );
buf ( n5029 , R_5a4_15ff7d08 );
buf ( n5030 , R_13a5_13d45338 );
buf ( n5031 , R_1115_11630b98 );
buf ( n5032 , R_19c4_17016fa8 );
buf ( n5033 , R_af6_117f49b8 );
buf ( n5034 , R_767_117f2d98 );
buf ( n5035 , R_d86_15fef7e8 );
buf ( n5036 , R_1734_1580c718 );
buf ( n5037 , R_836_123b33b8 );
buf ( n5038 , R_a27_117ede38 );
buf ( n5039 , R_1474_13c042d8 );
buf ( n5040 , R_1046_123bc918 );
buf ( n5041 , R_e55_124c3a98 );
buf ( n5042 , R_1665_156ac678 );
buf ( n5043 , R_122a_14a0b318 );
buf ( n5044 , R_18af_11c6f7d8 );
buf ( n5045 , R_1849_140b6358 );
buf ( n5046 , R_1290_13dd8b98 );
buf ( n5047 , R_c71_14a11e98 );
buf ( n5048 , R_652_13d386d8 );
buf ( n5049 , R_5ec_14868df8 );
buf ( n5050 , R_c0b_13b8c038 );
buf ( n5051 , R_574_13d4ec18 );
buf ( n5052 , R_6ca_156b3f18 );
buf ( n5053 , R_1308_117f2438 );
buf ( n5054 , R_17d1_11c6fa58 );
buf ( n5055 , R_b93_15881078 );
buf ( n5056 , R_ce9_156b86f8 );
buf ( n5057 , R_1927_123bb6f8 );
buf ( n5058 , R_11b2_14a101d8 );
buf ( n5059 , R_8f1_14a0fcd8 );
buf ( n5060 , R_f10_156ab778 );
buf ( n5061 , R_15aa_13c1f498 );
buf ( n5062 , R_152f_158884b8 );
buf ( n5063 , R_f8b_13dda218 );
buf ( n5064 , R_96c_15ff4e28 );
buf ( n5065 , R_948_15ff1728 );
buf ( n5066 , R_915_158834b8 );
buf ( n5067 , R_f34_123bd958 );
buf ( n5068 , R_1553_1162fdd8 );
buf ( n5069 , R_1586_13cd7938 );
buf ( n5070 , R_f67_156b54f8 );
buf ( n5071 , R_1701_117ee5b8 );
buf ( n5072 , R_10e2_13b97cf8 );
buf ( n5073 , R_ac3_13d41ff8 );
buf ( n5074 , R_79a_13b8d758 );
buf ( n5075 , R_db9_13d4e358 );
buf ( n5076 , R_13d8_13c10178 );
buf ( n5077 , R_19f7_123b4218 );
buf ( n5078 , R_ec2_156acdf8 );
buf ( n5079 , R_fd9_13cd6038 );
buf ( n5080 , R_14e1_13d4fbb8 );
buf ( n5081 , R_9ba_13d3b018 );
buf ( n5082 , R_8a3_117f3298 );
buf ( n5083 , R_15f8_150dd618 );
buf ( n5084 , R_b1c_10084238 );
buf ( n5085 , R_d60_1700c1e8 );
buf ( n5086 , R_137f_13d27fd8 );
buf ( n5087 , R_175a_15fedda8 );
buf ( n5088 , R_199e_123b8d18 );
buf ( n5089 , R_113b_11c703b8 );
buf ( n5090 , R_741_156b0278 );
buf ( n5091 , R_15e6_140b4238 );
buf ( n5092 , R_14f3_10088a18 );
buf ( n5093 , R_fc7_117e8c58 );
buf ( n5094 , R_8b5_13ccefb8 );
buf ( n5095 , R_9a8_14a19af8 );
buf ( n5096 , R_ed4_150e1998 );
buf ( n5097 , R_d68_15885b78 );
buf ( n5098 , R_b14_11c6b8b8 );
buf ( n5099 , R_1387_117eaf58 );
buf ( n5100 , R_19a6_14a19738 );
buf ( n5101 , R_1752_150e4738 );
buf ( n5102 , R_749_123b2918 );
buf ( n5103 , R_1133_1587e378 );
buf ( n5104 , R_1417_15ff4428 );
buf ( n5105 , R_df8_15888eb8 );
buf ( n5106 , R_7d9_124c3098 );
buf ( n5107 , R_a84_13b8b778 );
buf ( n5108 , R_10a3_13c1e4f8 );
buf ( n5109 , R_1a36_14b1b318 );
buf ( n5110 , R_16c2_156b1e98 );
buf ( n5111 , R_1a11_123b7b98 );
buf ( n5112 , R_13f2_13de2738 );
buf ( n5113 , R_dd3_14a19a58 );
buf ( n5114 , R_7b4_15885a38 );
buf ( n5115 , R_aa9_13cd5818 );
buf ( n5116 , R_10c8_14a14058 );
buf ( n5117 , R_16e7_117eea18 );
buf ( n5118 , R_b27_10087e38 );
buf ( n5119 , R_d55_117f0f98 );
buf ( n5120 , R_1765_12fbdf98 );
buf ( n5121 , R_1374_17015888 );
buf ( n5122 , R_1146_123bed58 );
buf ( n5123 , R_1993_13d53b78 );
buf ( n5124 , R_736_15ff9108 );
buf ( n5125 , R_56b_123b7558 );
buf ( n5126 , R_6d3_1007e1f8 );
buf ( n5127 , R_1311_10087a78 );
buf ( n5128 , R_17c8_13d50a18 );
buf ( n5129 , R_b8a_14b26858 );
buf ( n5130 , R_cf2_14a17438 );
buf ( n5131 , R_1930_13c083d8 );
buf ( n5132 , R_11a9_117f1038 );
buf ( n5133 , R_1638_15815818 );
buf ( n5134 , R_9fa_123b77d8 );
buf ( n5135 , R_e82_13df3ef8 );
buf ( n5136 , R_1019_158858f8 );
buf ( n5137 , R_863_13d47318 );
buf ( n5138 , R_14a1_117ed938 );
buf ( n5139 , R_eb2_11c6d2f8 );
buf ( n5140 , R_fe9_1162ed98 );
buf ( n5141 , R_14d1_1587ae58 );
buf ( n5142 , R_9ca_1587bd58 );
buf ( n5143 , R_893_13ccf238 );
buf ( n5144 , R_1608_117f45f8 );
buf ( n5145 , R_6f3_17012cc8 );
buf ( n5146 , R_1189_13de2d78 );
buf ( n5147 , R_1950_123b8098 );
buf ( n5148 , R_d12_13cd6d58 );
buf ( n5149 , R_b6a_140afff8 );
buf ( n5150 , R_17a8_13d3cf58 );
buf ( n5151 , R_1331_148755f8 );
buf ( n5152 , R_e9f_17016288 );
buf ( n5153 , R_9dd_156ab8b8 );
buf ( n5154 , R_161b_13d3ca58 );
buf ( n5155 , R_14be_13b98478 );
buf ( n5156 , R_880_117ea2d8 );
buf ( n5157 , R_ffc_13b8acd8 );
buf ( n5158 , R_1789_13cca9b8 );
buf ( n5159 , R_196f_13bf01d8 );
buf ( n5160 , R_d31_156b13f8 );
buf ( n5161 , R_116a_13c23e58 );
buf ( n5162 , R_1350_11632498 );
buf ( n5163 , R_b4b_156ad398 );
buf ( n5164 , R_712_13b90d18 );
buf ( n5165 , R_e92_117f2ed8 );
buf ( n5166 , R_9ea_123b7e18 );
buf ( n5167 , R_1628_123b7698 );
buf ( n5168 , R_14b1_14a16e98 );
buf ( n5169 , R_873_14a14238 );
buf ( n5170 , R_1009_13b980b8 );
buf ( n5171 , R_bf2_170099e8 );
buf ( n5172 , R_12a9_1162d0d8 );
buf ( n5173 , R_1211_150e5278 );
buf ( n5174 , R_c8a_150e3798 );
buf ( n5175 , R_1830_13bf6358 );
buf ( n5176 , R_66b_150e1498 );
buf ( n5177 , R_5d3_158808f8 );
buf ( n5178 , R_18c8_13cd9f58 );
buf ( n5179 , R_a42_15888198 );
buf ( n5180 , R_81b_12fbec18 );
buf ( n5181 , R_1061_13d3c558 );
buf ( n5182 , R_1459_17016aa8 );
buf ( n5183 , R_1680_1486aab8 );
buf ( n5184 , R_e3a_123bb798 );
buf ( n5185 , R_17ef_15889958 );
buf ( n5186 , R_1909_15815e58 );
buf ( n5187 , R_6ac_12fc1918 );
buf ( n5188 , R_bb1_14874d38 );
buf ( n5189 , R_12ea_13ddf358 );
buf ( n5190 , R_11d0_170096c8 );
buf ( n5191 , R_ccb_117ec038 );
buf ( n5192 , R_592_13c23958 );
buf ( n5193 , R_fee_14b29f58 );
buf ( n5194 , R_ead_13c22378 );
buf ( n5195 , R_9cf_1162e118 );
buf ( n5196 , R_14cc_123c0b58 );
buf ( n5197 , R_160d_123bff78 );
buf ( n5198 , R_88e_123c0fb8 );
buf ( n5199 , R_8ff_156b7c58 );
buf ( n5200 , R_f1e_15880038 );
buf ( n5201 , R_153d_15811218 );
buf ( n5202 , R_159c_15815db8 );
buf ( n5203 , R_f7d_13cd0778 );
buf ( n5204 , R_95e_13b98018 );
buf ( n5205 , R_189d_13cd3518 );
buf ( n5206 , R_127e_13d4f118 );
buf ( n5207 , R_c5f_12fbfa78 );
buf ( n5208 , R_640_140b2258 );
buf ( n5209 , R_5fe_15888558 );
buf ( n5210 , R_c1d_13dfb1f8 );
buf ( n5211 , R_123c_15fee708 );
buf ( n5212 , R_185b_14b21538 );
buf ( n5213 , R_15d1_123b63d8 );
buf ( n5214 , R_fb2_15810818 );
buf ( n5215 , R_8ca_15815bd8 );
buf ( n5216 , R_993_11c6b598 );
buf ( n5217 , R_ee9_1700fca8 );
buf ( n5218 , R_1508_156b7898 );
buf ( n5219 , R_121c_158871f8 );
buf ( n5220 , R_129e_13d3cb98 );
buf ( n5221 , R_183b_13c20bb8 );
buf ( n5222 , R_c7f_13cd6ad8 );
buf ( n5223 , R_660_156ba458 );
buf ( n5224 , R_5de_123b7cd8 );
buf ( n5225 , R_18bd_140b9878 );
buf ( n5226 , R_bfd_11c6f238 );
buf ( n5227 , R_16b4_117ead78 );
buf ( n5228 , R_e06_1580ff58 );
buf ( n5229 , R_7e7_15885858 );
buf ( n5230 , R_1a44_1162c4f8 );
buf ( n5231 , R_a76_13d38638 );
buf ( n5232 , R_1095_156b0ef8 );
buf ( n5233 , R_1425_13d571d8 );
buf ( n5234 , R_8e5_150db318 );
buf ( n5235 , R_15b6_1580e838 );
buf ( n5236 , R_f04_15885038 );
buf ( n5237 , R_f97_1700c288 );
buf ( n5238 , R_1523_140b8e78 );
buf ( n5239 , R_978_156b6498 );
buf ( n5240 , R_914_13d54c58 );
buf ( n5241 , R_f33_13d59258 );
buf ( n5242 , R_1552_13ccfa58 );
buf ( n5243 , R_1587_140aacd8 );
buf ( n5244 , R_f68_140acb78 );
buf ( n5245 , R_949_14b26a38 );
buf ( n5246 , R_15c0_158147d8 );
buf ( n5247 , R_8db_1580e158 );
buf ( n5248 , R_fa1_1162ffb8 );
buf ( n5249 , R_efa_13bf5818 );
buf ( n5250 , R_982_13debcf8 );
buf ( n5251 , R_1519_15813e78 );
buf ( n5252 , R_164e_117eb138 );
buf ( n5253 , R_148b_15886118 );
buf ( n5254 , R_a10_13df0f78 );
buf ( n5255 , R_e6c_15ff0d28 );
buf ( n5256 , R_102f_123c08d8 );
buf ( n5257 , R_84d_15feee88 );
buf ( n5258 , R_1703_13c254d8 );
buf ( n5259 , R_10e4_158894f8 );
buf ( n5260 , R_ac5_15883558 );
buf ( n5261 , R_798_123beb78 );
buf ( n5262 , R_db7_14869938 );
buf ( n5263 , R_13d6_156ae8d8 );
buf ( n5264 , R_19f5_13d2c2b8 );
buf ( n5265 , R_eb7_11c6d1b8 );
buf ( n5266 , R_fe4_12fc21d8 );
buf ( n5267 , R_14d6_1008b178 );
buf ( n5268 , R_9c5_14b21d58 );
buf ( n5269 , R_898_123b5c58 );
buf ( n5270 , R_1603_14872fd8 );
buf ( n5271 , R_1714_15889638 );
buf ( n5272 , R_10f5_140b5f98 );
buf ( n5273 , R_ad6_14873258 );
buf ( n5274 , R_787_14a0e838 );
buf ( n5275 , R_da6_13ddc158 );
buf ( n5276 , R_13c5_15fee208 );
buf ( n5277 , R_19e4_13de3a98 );
buf ( n5278 , R_98b_13b8dcf8 );
buf ( n5279 , R_ef1_13b924d8 );
buf ( n5280 , R_8d2_156ad578 );
buf ( n5281 , R_faa_156b0458 );
buf ( n5282 , R_1510_13d1f0b8 );
buf ( n5283 , R_15c9_13bf0b38 );
buf ( n5284 , R_aa7_13d451f8 );
buf ( n5285 , R_7b6_14a18018 );
buf ( n5286 , R_dd5_124c5258 );
buf ( n5287 , R_10c6_1700ff28 );
buf ( n5288 , R_13f4_14a0b778 );
buf ( n5289 , R_16e5_13c07ed8 );
buf ( n5290 , R_1a13_117ef058 );
buf ( n5291 , R_839_14b28f18 );
buf ( n5292 , R_e58_158814d8 );
buf ( n5293 , R_a24_123b5938 );
buf ( n5294 , R_1043_14b26538 );
buf ( n5295 , R_1477_117f0098 );
buf ( n5296 , R_1662_13df1978 );
buf ( n5297 , R_854_15ff3e88 );
buf ( n5298 , R_e73_14b288d8 );
buf ( n5299 , R_a09_123bb158 );
buf ( n5300 , R_1028_117f4eb8 );
buf ( n5301 , R_1492_13cd4378 );
buf ( n5302 , R_1647_12fc19b8 );
buf ( n5303 , R_be8_15ffcee8 );
buf ( n5304 , R_5c9_14b27438 );
buf ( n5305 , R_675_156aec98 );
buf ( n5306 , R_c94_13b8fb98 );
buf ( n5307 , R_1207_156b81f8 );
buf ( n5308 , R_12b3_13ddf718 );
buf ( n5309 , R_1826_140b01d8 );
buf ( n5310 , R_18d2_13c290d8 );
buf ( n5311 , R_cac_123c1058 );
buf ( n5312 , R_5b1_13d28e38 );
buf ( n5313 , R_68d_1700f2a8 );
buf ( n5314 , R_bd0_13ccc538 );
buf ( n5315 , R_11ef_117f3d38 );
buf ( n5316 , R_12cb_123bfe38 );
buf ( n5317 , R_180e_1580c7b8 );
buf ( n5318 , R_18ea_14a115d8 );
buf ( n5319 , R_d75_1486bc38 );
buf ( n5320 , R_756_13b8ae18 );
buf ( n5321 , R_b07_140aaa58 );
buf ( n5322 , R_1126_156aaeb8 );
buf ( n5323 , R_1394_15814878 );
buf ( n5324 , R_1745_123b4cb8 );
buf ( n5325 , R_19b3_123bc558 );
buf ( n5326 , R_d7a_13b95ef8 );
buf ( n5327 , R_75b_15814558 );
buf ( n5328 , R_b02_14a13f18 );
buf ( n5329 , R_1121_150e9c38 );
buf ( n5330 , R_1399_158830f8 );
buf ( n5331 , R_1740_13cd6fd8 );
buf ( n5332 , R_19b8_15812c58 );
buf ( n5333 , R_c0a_14a19ff8 );
buf ( n5334 , R_5eb_15feeac8 );
buf ( n5335 , R_653_123be358 );
buf ( n5336 , R_c72_13df6fb8 );
buf ( n5337 , R_1229_156b7938 );
buf ( n5338 , R_1291_14a0d758 );
buf ( n5339 , R_1848_14a197d8 );
buf ( n5340 , R_18b0_15815a98 );
buf ( n5341 , R_a96_150e8478 );
buf ( n5342 , R_7c7_13d45c98 );
buf ( n5343 , R_de6_13c05778 );
buf ( n5344 , R_10b5_156ab6d8 );
buf ( n5345 , R_1405_14a192d8 );
buf ( n5346 , R_16d4_14868c18 );
buf ( n5347 , R_1a24_116348d8 );
buf ( n5348 , R_85f_13dd89b8 );
buf ( n5349 , R_e7e_140ad6b8 );
buf ( n5350 , R_9fe_13c02d98 );
buf ( n5351 , R_101d_123b5d98 );
buf ( n5352 , R_149d_156b8dd8 );
buf ( n5353 , R_163c_1486a6f8 );
buf ( n5354 , R_d9b_13d3dbd8 );
buf ( n5355 , R_77c_116359b8 );
buf ( n5356 , R_ae1_15fed768 );
buf ( n5357 , R_1100_10085818 );
buf ( n5358 , R_13ba_15881d98 );
buf ( n5359 , R_171f_13bf08b8 );
buf ( n5360 , R_19d9_1700c508 );
buf ( n5361 , R_889_15ff9b08 );
buf ( n5362 , R_9d4_11c6e6f8 );
buf ( n5363 , R_ea8_13d1fe78 );
buf ( n5364 , R_ff3_117efc38 );
buf ( n5365 , R_14c7_140b4918 );
buf ( n5366 , R_1612_13cd0278 );
buf ( n5367 , R_582_14869118 );
buf ( n5368 , R_cdb_14a0ae18 );
buf ( n5369 , R_ba1_13d29338 );
buf ( n5370 , R_6bc_13cd53b8 );
buf ( n5371 , R_11c0_13deef98 );
buf ( n5372 , R_12fa_11631638 );
buf ( n5373 , R_17df_13cd0e58 );
buf ( n5374 , R_1919_1587e2d8 );
buf ( n5375 , R_e24_13ddcfb8 );
buf ( n5376 , R_a58_14a18a18 );
buf ( n5377 , R_805_1580a7d8 );
buf ( n5378 , R_1077_11c6d898 );
buf ( n5379 , R_1443_13d3f9d8 );
buf ( n5380 , R_1696_156afd78 );
buf ( n5381 , R_1a62_14b1b138 );
buf ( n5382 , R_94a_156b24d8 );
buf ( n5383 , R_f32_116350f8 );
buf ( n5384 , R_913_100840f8 );
buf ( n5385 , R_f69_117f0c78 );
buf ( n5386 , R_1551_150dde38 );
buf ( n5387 , R_1588_150e7d98 );
buf ( n5388 , R_a50_13df7698 );
buf ( n5389 , R_e2c_15881e38 );
buf ( n5390 , R_80d_14a16a38 );
buf ( n5391 , R_106f_156ad938 );
buf ( n5392 , R_144b_1486ce58 );
buf ( n5393 , R_168e_123bbc98 );
buf ( n5394 , R_6fe_13bf5318 );
buf ( n5395 , R_b5f_13cd4918 );
buf ( n5396 , R_d1d_13def2b8 );
buf ( n5397 , R_117e_14a0ccb8 );
buf ( n5398 , R_133c_117f2938 );
buf ( n5399 , R_179d_10085138 );
buf ( n5400 , R_195b_14b1c8f8 );
buf ( n5401 , R_cb3_1587b358 );
buf ( n5402 , R_5aa_13dd5678 );
buf ( n5403 , R_694_11636b38 );
buf ( n5404 , R_bc9_124c3d18 );
buf ( n5405 , R_11e8_13ccd258 );
buf ( n5406 , R_12d2_123bdc78 );
buf ( n5407 , R_1807_117ee298 );
buf ( n5408 , R_18f1_156aba98 );
buf ( n5409 , R_c1c_156ba3b8 );
buf ( n5410 , R_5fd_14a10958 );
buf ( n5411 , R_641_123b90d8 );
buf ( n5412 , R_c60_158171b8 );
buf ( n5413 , R_123b_1162cd18 );
buf ( n5414 , R_127f_13b8a558 );
buf ( n5415 , R_185a_15814cd8 );
buf ( n5416 , R_189e_13bf8e78 );
buf ( n5417 , R_877_13d3e498 );
buf ( n5418 , R_9e6_14b28838 );
buf ( n5419 , R_e96_156b4a58 );
buf ( n5420 , R_1005_13c1edb8 );
buf ( n5421 , R_14b5_15882018 );
buf ( n5422 , R_1624_10086cb8 );
buf ( n5423 , R_db5_117ece98 );
buf ( n5424 , R_796_156b0138 );
buf ( n5425 , R_ac7_148725d8 );
buf ( n5426 , R_10e6_11630918 );
buf ( n5427 , R_13d4_15882bf8 );
buf ( n5428 , R_1705_10085db8 );
buf ( n5429 , R_19f3_1008c618 );
buf ( n5430 , R_96d_1162e7f8 );
buf ( n5431 , R_f0f_13d3d9f8 );
buf ( n5432 , R_8f0_13d29838 );
buf ( n5433 , R_f8c_117f2578 );
buf ( n5434 , R_152e_117f3f18 );
buf ( n5435 , R_15ab_13ccc358 );
buf ( n5436 , R_587_124c5118 );
buf ( n5437 , R_cd6_13d39178 );
buf ( n5438 , R_ba6_156ad9d8 );
buf ( n5439 , R_6b7_13c0b718 );
buf ( n5440 , R_11c5_13d39538 );
buf ( n5441 , R_12f5_158104f8 );
buf ( n5442 , R_17e4_156acf38 );
buf ( n5443 , R_1914_10084f58 );
buf ( n5444 , R_846_100885b8 );
buf ( n5445 , R_e65_15810318 );
buf ( n5446 , R_a17_13ccf878 );
buf ( n5447 , R_1036_140b5278 );
buf ( n5448 , R_1484_11c6b778 );
buf ( n5449 , R_1655_1700cdc8 );
buf ( n5450 , R_a45_17017188 );
buf ( n5451 , R_e37_10083018 );
buf ( n5452 , R_818_13b8dbb8 );
buf ( n5453 , R_1064_1700d5e8 );
buf ( n5454 , R_1456_13cd8518 );
buf ( n5455 , R_1683_1587f6d8 );
buf ( n5456 , R_57d_14b1ef18 );
buf ( n5457 , R_ce0_1580ccb8 );
buf ( n5458 , R_b9c_15884e58 );
buf ( n5459 , R_6c1_156b1538 );
buf ( n5460 , R_11bb_117ed2f8 );
buf ( n5461 , R_12ff_17012408 );
buf ( n5462 , R_17da_123bf398 );
buf ( n5463 , R_191e_140b0c78 );
buf ( n5464 , R_d58_13df39f8 );
buf ( n5465 , R_b24_15815958 );
buf ( n5466 , R_739_123c1698 );
buf ( n5467 , R_1143_13cd7078 );
buf ( n5468 , R_1377_158873d8 );
buf ( n5469 , R_1762_140aef18 );
buf ( n5470 , R_1996_156b4058 );
buf ( n5471 , R_95f_13bf9918 );
buf ( n5472 , R_f1d_15ff80c8 );
buf ( n5473 , R_8fe_13d4f898 );
buf ( n5474 , R_f7e_156b42d8 );
buf ( n5475 , R_153c_13c1d698 );
buf ( n5476 , R_159d_1162b198 );
buf ( n5477 , R_aa5_156b4238 );
buf ( n5478 , R_7b8_1162e9d8 );
buf ( n5479 , R_dd7_140b62b8 );
buf ( n5480 , R_10c4_12fc1878 );
buf ( n5481 , R_13f6_1700d728 );
buf ( n5482 , R_16e3_123b4d58 );
buf ( n5483 , R_1a15_13d3e998 );
buf ( n5484 , R_b0c_123c1878 );
buf ( n5485 , R_d70_13b96038 );
buf ( n5486 , R_751_13bf12b8 );
buf ( n5487 , R_112b_13d5c3b8 );
buf ( n5488 , R_138f_13df66f8 );
buf ( n5489 , R_174a_13d24658 );
buf ( n5490 , R_19ae_1587f818 );
buf ( n5491 , R_a8b_117f7898 );
buf ( n5492 , R_7d2_10082a78 );
buf ( n5493 , R_df1_15884778 );
buf ( n5494 , R_10aa_13c28458 );
buf ( n5495 , R_1410_13cd5a98 );
buf ( n5496 , R_16c9_13c03018 );
buf ( n5497 , R_1a2f_15886b18 );
buf ( n5498 , R_d7f_117f5ef8 );
buf ( n5499 , R_760_13cce6f8 );
buf ( n5500 , R_afd_156ae018 );
buf ( n5501 , R_111c_13c0f138 );
buf ( n5502 , R_139e_15ff9428 );
buf ( n5503 , R_173b_13d23758 );
buf ( n5504 , R_19bd_150e0c78 );
buf ( n5505 , R_70f_14b26038 );
buf ( n5506 , R_b4e_158835f8 );
buf ( n5507 , R_d2e_15ff2d08 );
buf ( n5508 , R_116d_14a0bc78 );
buf ( n5509 , R_134d_13cd26b8 );
buf ( n5510 , R_178c_13d39718 );
buf ( n5511 , R_196c_117ef418 );
buf ( n5512 , R_705_17018768 );
buf ( n5513 , R_b58_12fc00b8 );
buf ( n5514 , R_d24_13c0ca78 );
buf ( n5515 , R_1177_13d5b558 );
buf ( n5516 , R_1343_13d298d8 );
buf ( n5517 , R_1796_156ae338 );
buf ( n5518 , R_1962_13d5d218 );
buf ( n5519 , R_c9d_13c00ef8 );
buf ( n5520 , R_bdf_117f0638 );
buf ( n5521 , R_5c0_117ea0f8 );
buf ( n5522 , R_67e_14a0b8b8 );
buf ( n5523 , R_11fe_124c36d8 );
buf ( n5524 , R_12bc_13b981f8 );
buf ( n5525 , R_181d_123ba758 );
buf ( n5526 , R_18db_11c6d7f8 );
buf ( n5527 , R_ebc_1580cfd8 );
buf ( n5528 , R_89d_11c693d8 );
buf ( n5529 , R_9c0_13d46b98 );
buf ( n5530 , R_fdf_158176b8 );
buf ( n5531 , R_14db_156b5e58 );
buf ( n5532 , R_15fe_140b97d8 );
buf ( n5533 , R_ee1_13d40c98 );
buf ( n5534 , R_99b_156b3838 );
buf ( n5535 , R_8c2_15813518 );
buf ( n5536 , R_fba_140aebf8 );
buf ( n5537 , R_1500_1700e8a8 );
buf ( n5538 , R_15d9_13d53538 );
buf ( n5539 , R_eda_13d57638 );
buf ( n5540 , R_9a2_13c28bd8 );
buf ( n5541 , R_8bb_13d43498 );
buf ( n5542 , R_fc1_156b40f8 );
buf ( n5543 , R_14f9_13cd6178 );
buf ( n5544 , R_15e0_13cd0458 );
buf ( n5545 , R_d8b_150dc7b8 );
buf ( n5546 , R_76c_150e63f8 );
buf ( n5547 , R_af1_13b8c3f8 );
buf ( n5548 , R_1110_13d5cdb8 );
buf ( n5549 , R_13aa_14b1d898 );
buf ( n5550 , R_172f_11c6dbb8 );
buf ( n5551 , R_19c9_1509b4f8 );
buf ( n5552 , R_55a_158145f8 );
buf ( n5553 , R_6e4_11630a58 );
buf ( n5554 , R_b79_13ccfd78 );
buf ( n5555 , R_d03_124c2eb8 );
buf ( n5556 , R_1198_117f3b58 );
buf ( n5557 , R_1322_15ff6ea8 );
buf ( n5558 , R_17b7_15810bd8 );
buf ( n5559 , R_1941_117ed4d8 );
buf ( n5560 , R_6cf_1486c6d8 );
buf ( n5561 , R_56f_14a0b598 );
buf ( n5562 , R_cee_13cd9c38 );
buf ( n5563 , R_b8e_150e97d8 );
buf ( n5564 , R_11ad_13d569b8 );
buf ( n5565 , R_130d_124c3818 );
buf ( n5566 , R_17cc_117e9298 );
buf ( n5567 , R_192c_13b94918 );
buf ( n5568 , R_94b_100881f8 );
buf ( n5569 , R_f31_13c231d8 );
buf ( n5570 , R_912_11630f58 );
buf ( n5571 , R_f6a_117ea058 );
buf ( n5572 , R_1550_17014668 );
buf ( n5573 , R_1589_123b7198 );
buf ( n5574 , R_bd7_14a0ef18 );
buf ( n5575 , R_ca5_1007eb58 );
buf ( n5576 , R_5b8_170170e8 );
buf ( n5577 , R_686_15810f98 );
buf ( n5578 , R_11f6_14b22bb8 );
buf ( n5579 , R_12c4_15ff0008 );
buf ( n5580 , R_1815_156b1cb8 );
buf ( n5581 , R_18e3_13ccb9f8 );
buf ( n5582 , R_6e0_14a15f98 );
buf ( n5583 , R_55e_148707d8 );
buf ( n5584 , R_cff_14a0b458 );
buf ( n5585 , R_b7d_156b6df8 );
buf ( n5586 , R_119c_14872ad8 );
buf ( n5587 , R_131e_13dd6e38 );
buf ( n5588 , R_17bb_13bf1d58 );
buf ( n5589 , R_193d_11c70638 );
buf ( n5590 , R_d92_14b21358 );
buf ( n5591 , R_773_117f54f8 );
buf ( n5592 , R_aea_17012908 );
buf ( n5593 , R_1109_15ff3de8 );
buf ( n5594 , R_13b1_150dc358 );
buf ( n5595 , R_1728_13d5beb8 );
buf ( n5596 , R_19d0_14870af8 );
buf ( n5597 , R_e12_13b8cc18 );
buf ( n5598 , R_a6a_13d1d218 );
buf ( n5599 , R_7f3_148688f8 );
buf ( n5600 , R_1089_123b6838 );
buf ( n5601 , R_1431_15812ed8 );
buf ( n5602 , R_16a8_123bf118 );
buf ( n5603 , R_1a50_117ed6b8 );
buf ( n5604 , R_6f7_117e93d8 );
buf ( n5605 , R_b66_14a0f238 );
buf ( n5606 , R_d16_13c1b7f8 );
buf ( n5607 , R_1185_13d1ecf8 );
buf ( n5608 , R_1335_13bf1f38 );
buf ( n5609 , R_17a4_14b1ea18 );
buf ( n5610 , R_1954_15ff1ae8 );
buf ( n5611 , R_e17_13df86d8 );
buf ( n5612 , R_a65_14b22b18 );
buf ( n5613 , R_7f8_1700bec8 );
buf ( n5614 , R_1084_13d39038 );
buf ( n5615 , R_1436_15fef608 );
buf ( n5616 , R_16a3_15ff2768 );
buf ( n5617 , R_1a55_123b5898 );
buf ( n5618 , R_a21_1587bad8 );
buf ( n5619 , R_83c_13cd7398 );
buf ( n5620 , R_e5b_123bf898 );
buf ( n5621 , R_1040_1008ac78 );
buf ( n5622 , R_147a_13c04378 );
buf ( n5623 , R_165f_13cd97d8 );
buf ( n5624 , R_bfc_13d53cb8 );
buf ( n5625 , R_5dd_123b45d8 );
buf ( n5626 , R_661_13d3c2d8 );
buf ( n5627 , R_c80_1008ca78 );
buf ( n5628 , R_121b_14b24698 );
buf ( n5629 , R_129f_1008b7b8 );
buf ( n5630 , R_183a_156acc18 );
buf ( n5631 , R_18be_14a0de38 );
buf ( n5632 , R_c1b_123b48f8 );
buf ( n5633 , R_5fc_140b3518 );
buf ( n5634 , R_642_14a0d118 );
buf ( n5635 , R_c61_13c06718 );
buf ( n5636 , R_123a_15ffcf88 );
buf ( n5637 , R_1280_14a106d8 );
buf ( n5638 , R_1859_13d25378 );
buf ( n5639 , R_189f_14a13c98 );
buf ( n5640 , R_556_13d2a2d8 );
buf ( n5641 , R_6e8_12fbf4d8 );
buf ( n5642 , R_b75_156ae838 );
buf ( n5643 , R_d07_156abe58 );
buf ( n5644 , R_1194_1580f058 );
buf ( n5645 , R_1326_11c684d8 );
buf ( n5646 , R_17b3_13ddb4d8 );
buf ( n5647 , R_1945_14b22898 );
buf ( n5648 , R_bf1_13df18d8 );
buf ( n5649 , R_5d2_10088f18 );
buf ( n5650 , R_66c_123c06f8 );
buf ( n5651 , R_c8b_13c0e5f8 );
buf ( n5652 , R_1210_117f56d8 );
buf ( n5653 , R_12aa_140afb98 );
buf ( n5654 , R_182f_13d58998 );
buf ( n5655 , R_18c9_11c6eb58 );
buf ( n5656 , R_cc0_1580fcd8 );
buf ( n5657 , R_59d_13df9d58 );
buf ( n5658 , R_6a1_13cd9b98 );
buf ( n5659 , R_bbc_13d4e678 );
buf ( n5660 , R_11db_124c45d8 );
buf ( n5661 , R_12df_13d27178 );
buf ( n5662 , R_17fa_13beb8b8 );
buf ( n5663 , R_18fe_1587ca78 );
buf ( n5664 , R_d63_117f68f8 );
buf ( n5665 , R_b19_158882d8 );
buf ( n5666 , R_744_123bea38 );
buf ( n5667 , R_1138_14869ed8 );
buf ( n5668 , R_1382_13b8b958 );
buf ( n5669 , R_1757_13de1978 );
buf ( n5670 , R_19a1_123b3598 );
buf ( n5671 , R_db3_14869898 );
buf ( n5672 , R_794_17016788 );
buf ( n5673 , R_ac9_15811cb8 );
buf ( n5674 , R_10e8_140b1538 );
buf ( n5675 , R_13d2_13c292b8 );
buf ( n5676 , R_1707_13ddd9b8 );
buf ( n5677 , R_19f1_13cce518 );
buf ( n5678 , R_ecd_13d5b5f8 );
buf ( n5679 , R_9af_1587fdb8 );
buf ( n5680 , R_8ae_11631778 );
buf ( n5681 , R_fce_13c051d8 );
buf ( n5682 , R_14ec_156b01d8 );
buf ( n5683 , R_15ed_1008af98 );
buf ( n5684 , R_da4_13cd7438 );
buf ( n5685 , R_785_116381b8 );
buf ( n5686 , R_ad8_117f7a78 );
buf ( n5687 , R_10f7_1587f598 );
buf ( n5688 , R_13c3_13cd0b38 );
buf ( n5689 , R_1716_123b6bf8 );
buf ( n5690 , R_19e2_13d567d8 );
buf ( n5691 , R_58c_1587fe58 );
buf ( n5692 , R_cd1_1486dc18 );
buf ( n5693 , R_bab_13df0e38 );
buf ( n5694 , R_6b2_14867ef8 );
buf ( n5695 , R_11ca_123bd9f8 );
buf ( n5696 , R_12f0_158817f8 );
buf ( n5697 , R_17e9_123bb5b8 );
buf ( n5698 , R_190f_15881b18 );
buf ( n5699 , R_979_117efcd8 );
buf ( n5700 , R_f03_13c06f38 );
buf ( n5701 , R_8e4_123b2b98 );
buf ( n5702 , R_f98_13d588f8 );
buf ( n5703 , R_1522_15817d98 );
buf ( n5704 , R_15b7_11636bd8 );
buf ( n5705 , R_c09_14a18bf8 );
buf ( n5706 , R_5ea_1162b558 );
buf ( n5707 , R_654_150e54f8 );
buf ( n5708 , R_c73_15810958 );
buf ( n5709 , R_1228_150e4ff8 );
buf ( n5710 , R_1292_117e9fb8 );
buf ( n5711 , R_1847_13d54898 );
buf ( n5712 , R_18b1_1162ae78 );
buf ( n5713 , R_ec7_10083838 );
buf ( n5714 , R_8a8_140b6858 );
buf ( n5715 , R_9b5_156b6038 );
buf ( n5716 , R_fd4_13bef878 );
buf ( n5717 , R_14e6_123be178 );
buf ( n5718 , R_15f3_1580b958 );
buf ( n5719 , R_6dc_13d56738 );
buf ( n5720 , R_562_11630198 );
buf ( n5721 , R_cfb_156b77f8 );
buf ( n5722 , R_b81_14b23658 );
buf ( n5723 , R_11a0_117f1a38 );
buf ( n5724 , R_131a_13cd6678 );
buf ( n5725 , R_17bf_1162eed8 );
buf ( n5726 , R_1939_13b99198 );
buf ( n5727 , R_85b_150e9ff8 );
buf ( n5728 , R_e7a_13df06b8 );
buf ( n5729 , R_a02_13d20378 );
buf ( n5730 , R_1021_14873438 );
buf ( n5731 , R_1499_13c056d8 );
buf ( n5732 , R_1640_15816e98 );
buf ( n5733 , R_6c6_14b27a78 );
buf ( n5734 , R_578_13c06678 );
buf ( n5735 , R_ce5_117e9518 );
buf ( n5736 , R_b97_116328f8 );
buf ( n5737 , R_11b6_123b6478 );
buf ( n5738 , R_1304_150e5a98 );
buf ( n5739 , R_17d5_13cd9eb8 );
buf ( n5740 , R_1923_10086ad8 );
buf ( n5741 , R_aa3_123ba9d8 );
buf ( n5742 , R_7ba_17013308 );
buf ( n5743 , R_dd9_1587f4f8 );
buf ( n5744 , R_10c2_13de4358 );
buf ( n5745 , R_13f8_14866c38 );
buf ( n5746 , R_16e1_1587e058 );
buf ( n5747 , R_1a17_13d3a398 );
buf ( n5748 , R_ea3_117f04f8 );
buf ( n5749 , R_884_124c4358 );
buf ( n5750 , R_9d9_14a0c178 );
buf ( n5751 , R_ff8_14a15098 );
buf ( n5752 , R_14c2_13d50e78 );
buf ( n5753 , R_1617_13de3e58 );
buf ( n5754 , R_e0d_13c081f8 );
buf ( n5755 , R_a6f_140ab4f8 );
buf ( n5756 , R_7ee_117eb4f8 );
buf ( n5757 , R_108e_117ecf38 );
buf ( n5758 , R_142c_13d55f18 );
buf ( n5759 , R_16ad_15885df8 );
buf ( n5760 , R_1a4b_13d3a118 );
buf ( n5761 , R_e01_13b8ca38 );
buf ( n5762 , R_a7b_150e6f38 );
buf ( n5763 , R_7e2_116332f8 );
buf ( n5764 , R_109a_140adc58 );
buf ( n5765 , R_1420_1580acd8 );
buf ( n5766 , R_16b9_13b972f8 );
buf ( n5767 , R_1a3f_13cd8f18 );
buf ( n5768 , R_597_156aeab8 );
buf ( n5769 , R_cc6_1486fd38 );
buf ( n5770 , R_bb6_13d58fd8 );
buf ( n5771 , R_6a7_140b7938 );
buf ( n5772 , R_11d5_14871bd8 );
buf ( n5773 , R_12e5_14b28bf8 );
buf ( n5774 , R_17f4_156b4cd8 );
buf ( n5775 , R_1904_140b9058 );
buf ( n5776 , R_dfa_1486ff18 );
buf ( n5777 , R_a82_116368b8 );
buf ( n5778 , R_7db_150dd1b8 );
buf ( n5779 , R_10a1_123b8598 );
buf ( n5780 , R_1419_13df1b58 );
buf ( n5781 , R_16c0_13b994b8 );
buf ( n5782 , R_1a38_13ccab98 );
buf ( n5783 , R_911_14b22078 );
buf ( n5784 , R_94c_123bc7d8 );
buf ( n5785 , R_f30_12fbf898 );
buf ( n5786 , R_f6b_13c0a6d8 );
buf ( n5787 , R_154f_1700ea88 );
buf ( n5788 , R_158a_13c25758 );
buf ( n5789 , R_d44_13b99418 );
buf ( n5790 , R_b38_13d23618 );
buf ( n5791 , R_725_13d4f618 );
buf ( n5792 , R_1157_14a13298 );
buf ( n5793 , R_1363_124c4718 );
buf ( n5794 , R_1776_15882518 );
buf ( n5795 , R_1982_15816fd8 );
buf ( n5796 , R_983_1700b4c8 );
buf ( n5797 , R_ef9_1007e338 );
buf ( n5798 , R_8da_1587ba38 );
buf ( n5799 , R_fa2_15ffaf08 );
buf ( n5800 , R_1518_13c09ff8 );
buf ( n5801 , R_15c1_13c1e138 );
buf ( n5802 , R_d41_13bf8f18 );
buf ( n5803 , R_722_14b26fd8 );
buf ( n5804 , R_b3b_14a0f378 );
buf ( n5805 , R_115a_156af9b8 );
buf ( n5806 , R_1360_156aa5f8 );
buf ( n5807 , R_1779_13dec3d8 );
buf ( n5808 , R_197f_1700ba68 );
buf ( n5809 , R_7fd_13d29658 );
buf ( n5810 , R_e1c_156b8158 );
buf ( n5811 , R_a60_124c2738 );
buf ( n5812 , R_107f_13d55ab8 );
buf ( n5813 , R_143b_13cd5458 );
buf ( n5814 , R_169e_13d59618 );
buf ( n5815 , R_1a5a_117ecd58 );
buf ( n5816 , R_a94_158121b8 );
buf ( n5817 , R_7c9_13c1bb18 );
buf ( n5818 , R_de8_13df22d8 );
buf ( n5819 , R_10b3_17011328 );
buf ( n5820 , R_1407_140b9cd8 );
buf ( n5821 , R_16d2_150e0098 );
buf ( n5822 , R_1a26_14868678 );
buf ( n5823 , R_e9a_14a0e1f8 );
buf ( n5824 , R_87b_123b2e18 );
buf ( n5825 , R_9e2_148680d8 );
buf ( n5826 , R_1001_100877f8 );
buf ( n5827 , R_14b9_150dda78 );
buf ( n5828 , R_1620_117efff8 );
buf ( n5829 , R_bc2_1580b098 );
buf ( n5830 , R_cba_13c20118 );
buf ( n5831 , R_5a3_13b98298 );
buf ( n5832 , R_69b_13bf94b8 );
buf ( n5833 , R_11e1_1486a798 );
buf ( n5834 , R_12d9_123ba118 );
buf ( n5835 , R_1800_15888378 );
buf ( n5836 , R_18f8_156ac538 );
buf ( n5837 , R_960_13ccf418 );
buf ( n5838 , R_f1c_13df79b8 );
buf ( n5839 , R_8fd_123b6fb8 );
buf ( n5840 , R_f7f_140aa558 );
buf ( n5841 , R_153b_117f5d18 );
buf ( n5842 , R_159e_14871db8 );
buf ( n5843 , R_d47_13d27998 );
buf ( n5844 , R_b35_1587cc58 );
buf ( n5845 , R_728_140ba318 );
buf ( n5846 , R_1154_117e95b8 );
buf ( n5847 , R_1366_17015568 );
buf ( n5848 , R_1773_156ac2b8 );
buf ( n5849 , R_1985_1162c3b8 );
buf ( n5850 , R_b11_15883698 );
buf ( n5851 , R_d6b_123b8958 );
buf ( n5852 , R_74c_150e17b8 );
buf ( n5853 , R_1130_13bef0f8 );
buf ( n5854 , R_138a_13d25cd8 );
buf ( n5855 , R_174f_13df2058 );
buf ( n5856 , R_19a9_1486eed8 );
buf ( n5857 , R_6ec_13c03b58 );
buf ( n5858 , R_b71_140afd78 );
buf ( n5859 , R_d0b_1587d158 );
buf ( n5860 , R_1190_13c09198 );
buf ( n5861 , R_132a_13d44bb8 );
buf ( n5862 , R_17af_123b9d58 );
buf ( n5863 , R_1949_140b51d8 );
buf ( n5864 , R_815_158140f8 );
buf ( n5865 , R_a48_13bed6b8 );
buf ( n5866 , R_e34_13cd7e38 );
buf ( n5867 , R_1067_13b93ab8 );
buf ( n5868 , R_1453_15ff99c8 );
buf ( n5869 , R_1686_1008c258 );
buf ( n5870 , R_af8_148696b8 );
buf ( n5871 , R_d84_156b3e78 );
buf ( n5872 , R_765_13df9678 );
buf ( n5873 , R_1117_140b2398 );
buf ( n5874 , R_13a3_123bd598 );
buf ( n5875 , R_1736_117f1218 );
buf ( n5876 , R_19c2_14871098 );
buf ( n5877 , R_d3e_14870198 );
buf ( n5878 , R_71f_123b6e78 );
buf ( n5879 , R_b3e_11631138 );
buf ( n5880 , R_115d_1008bd58 );
buf ( n5881 , R_135d_13cd9d78 );
buf ( n5882 , R_177c_11629258 );
buf ( n5883 , R_197c_13bec8f8 );
buf ( n5884 , R_96e_1162bff8 );
buf ( n5885 , R_f0e_17010f68 );
buf ( n5886 , R_8ef_13dd96d8 );
buf ( n5887 , R_f8d_13cd51d8 );
buf ( n5888 , R_152d_13d1f8d8 );
buf ( n5889 , R_15ac_12fc1418 );
buf ( n5890 , R_ee8_13d55658 );
buf ( n5891 , R_994_13c086f8 );
buf ( n5892 , R_8c9_1162f838 );
buf ( n5893 , R_fb3_11c6c7b8 );
buf ( n5894 , R_1507_14b218f8 );
buf ( n5895 , R_15d2_11c6e978 );
buf ( n5896 , R_ed3_13b93018 );
buf ( n5897 , R_9a9_140ac3f8 );
buf ( n5898 , R_8b4_150e2e38 );
buf ( n5899 , R_fc8_14875238 );
buf ( n5900 , R_14f2_13cd1718 );
buf ( n5901 , R_15e7_150e0e58 );
buf ( n5902 , R_c1a_13d3c198 );
buf ( n5903 , R_5fb_156b22f8 );
buf ( n5904 , R_643_117ea698 );
buf ( n5905 , R_c62_1162c598 );
buf ( n5906 , R_1239_15817938 );
buf ( n5907 , R_1281_158887d8 );
buf ( n5908 , R_1858_13bea9b8 );
buf ( n5909 , R_18a0_123bfcf8 );
buf ( n5910 , R_98c_13c21f18 );
buf ( n5911 , R_ef0_13d51418 );
buf ( n5912 , R_8d1_12fc06f8 );
buf ( n5913 , R_fab_14a127f8 );
buf ( n5914 , R_150f_15817398 );
buf ( n5915 , R_15ca_156b71b8 );
buf ( n5916 , R_c95_123be2b8 );
buf ( n5917 , R_be7_1162d858 );
buf ( n5918 , R_5c8_15feeca8 );
buf ( n5919 , R_676_13d37e18 );
buf ( n5920 , R_1206_13ddcc98 );
buf ( n5921 , R_12b4_10087938 );
buf ( n5922 , R_1825_1486a298 );
buf ( n5923 , R_18d3_17018f88 );
buf ( n5924 , R_d5b_150e0958 );
buf ( n5925 , R_b21_14b21e98 );
buf ( n5926 , R_73c_13bec858 );
buf ( n5927 , R_1140_13b98798 );
buf ( n5928 , R_137a_13dd7018 );
buf ( n5929 , R_175f_15ff7f88 );
buf ( n5930 , R_1999_117f2118 );
buf ( n5931 , R_d4a_13df40d8 );
buf ( n5932 , R_b32_13c268d8 );
buf ( n5933 , R_72b_11632c18 );
buf ( n5934 , R_1151_11638898 );
buf ( n5935 , R_1369_117f5138 );
buf ( n5936 , R_1770_124c2a58 );
buf ( n5937 , R_1988_150dfaf8 );
buf ( n5938 , R_db1_13bf06d8 );
buf ( n5939 , R_792_13ccb638 );
buf ( n5940 , R_acb_13d2a378 );
buf ( n5941 , R_10ea_13d2b598 );
buf ( n5942 , R_13d0_1700b388 );
buf ( n5943 , R_1709_1162a298 );
buf ( n5944 , R_19ef_150de1f8 );
buf ( n5945 , R_ae3_14b24738 );
buf ( n5946 , R_d99_156abef8 );
buf ( n5947 , R_77a_13c0f3b8 );
buf ( n5948 , R_1102_11632358 );
buf ( n5949 , R_13b8_13c29c18 );
buf ( n5950 , R_1721_14870f58 );
buf ( n5951 , R_19d7_13de38b8 );
buf ( n5952 , R_6d8_1580ebf8 );
buf ( n5953 , R_566_140b4f58 );
buf ( n5954 , R_cf7_13d26778 );
buf ( n5955 , R_b85_13df3958 );
buf ( n5956 , R_11a4_140b1178 );
buf ( n5957 , R_1316_13c24718 );
buf ( n5958 , R_17c3_13df1e78 );
buf ( n5959 , R_1935_14a13798 );
buf ( n5960 , R_a0d_14a0f198 );
buf ( n5961 , R_850_1700cbe8 );
buf ( n5962 , R_e6f_117ee6f8 );
buf ( n5963 , R_102c_156ae3d8 );
buf ( n5964 , R_148e_17014208 );
buf ( n5965 , R_164b_123b8638 );
buf ( n5966 , R_f2f_13ccded8 );
buf ( n5967 , R_910_158144b8 );
buf ( n5968 , R_94d_13de1dd8 );
buf ( n5969 , R_f6c_140aca38 );
buf ( n5970 , R_154e_158131f8 );
buf ( n5971 , R_158b_123b5078 );
buf ( n5972 , R_70c_1162a338 );
buf ( n5973 , R_b51_13df4c18 );
buf ( n5974 , R_d2b_123bacf8 );
buf ( n5975 , R_1170_13ddca18 );
buf ( n5976 , R_134a_123bdb38 );
buf ( n5977 , R_178f_14a0df78 );
buf ( n5978 , R_1969_13c0e918 );
buf ( n5979 , R_ec1_13c0ddd8 );
buf ( n5980 , R_8a2_13dd9638 );
buf ( n5981 , R_9bb_14a13d38 );
buf ( n5982 , R_fda_14876098 );
buf ( n5983 , R_14e0_117ea9b8 );
buf ( n5984 , R_15f9_13d4fcf8 );
buf ( n5985 , R_d3b_150e4a58 );
buf ( n5986 , R_71c_150dba98 );
buf ( n5987 , R_b41_100844b8 );
buf ( n5988 , R_1160_14a16498 );
buf ( n5989 , R_135a_156b8838 );
buf ( n5990 , R_177f_13ccedd8 );
buf ( n5991 , R_1979_156ad7f8 );
buf ( n5992 , R_80a_11c686b8 );
buf ( n5993 , R_a53_13d54ed8 );
buf ( n5994 , R_e29_124c3138 );
buf ( n5995 , R_1072_13d5c598 );
buf ( n5996 , R_1448_156b5098 );
buf ( n5997 , R_1691_13bf8478 );
buf ( n5998 , R_1a67_13d3a898 );
buf ( n5999 , R_aa1_13ccbd18 );
buf ( n6000 , R_7bc_13ccc218 );
buf ( n6001 , R_ddb_15812618 );
buf ( n6002 , R_10c0_15816d58 );
buf ( n6003 , R_13fa_14b29a58 );
buf ( n6004 , R_16df_10084eb8 );
buf ( n6005 , R_1a19_11c70a98 );
buf ( n6006 , R_a1e_13de1338 );
buf ( n6007 , R_83f_123bc5f8 );
buf ( n6008 , R_e5e_13c25258 );
buf ( n6009 , R_103d_123b2738 );
buf ( n6010 , R_147d_13d53e98 );
buf ( n6011 , R_165c_123b57f8 );
buf ( n6012 , R_c74_14b242d8 );
buf ( n6013 , R_c08_13ded7d8 );
buf ( n6014 , R_5e9_15816178 );
buf ( n6015 , R_655_13c026b8 );
buf ( n6016 , R_1227_123b72d8 );
buf ( n6017 , R_1293_1008c6b8 );
buf ( n6018 , R_1846_13c22af8 );
buf ( n6019 , R_18b2_150dd4d8 );
buf ( n6020 , R_a14_11632038 );
buf ( n6021 , R_849_123c1af8 );
buf ( n6022 , R_e68_15887658 );
buf ( n6023 , R_1033_13bf8518 );
buf ( n6024 , R_1487_1007fc38 );
buf ( n6025 , R_1652_11635418 );
buf ( n6026 , R_68e_11630eb8 );
buf ( n6027 , R_bcf_1486c4f8 );
buf ( n6028 , R_cad_150e5c78 );
buf ( n6029 , R_5b0_13d20c38 );
buf ( n6030 , R_11ee_13df5938 );
buf ( n6031 , R_12cc_156aee78 );
buf ( n6032 , R_180d_13d29dd8 );
buf ( n6033 , R_18eb_13cd2bb8 );
buf ( n6034 , R_7e9_13b903b8 );
buf ( n6035 , R_e08_14a11498 );
buf ( n6036 , R_a74_13c02a78 );
buf ( n6037 , R_1093_123bddb8 );
buf ( n6038 , R_1427_1580dd98 );
buf ( n6039 , R_16b2_123b89f8 );
buf ( n6040 , R_1a46_150dff58 );
buf ( n6041 , R_c81_140ac718 );
buf ( n6042 , R_bfb_117e8f78 );
buf ( n6043 , R_5dc_13cd21b8 );
buf ( n6044 , R_662_11c6af58 );
buf ( n6045 , R_121a_13dd6bb8 );
buf ( n6046 , R_12a0_156af7d8 );
buf ( n6047 , R_1839_10083a18 );
buf ( n6048 , R_18bf_13cd63f8 );
buf ( n6049 , R_d4d_14b1c218 );
buf ( n6050 , R_b2f_14a168f8 );
buf ( n6051 , R_72e_15885178 );
buf ( n6052 , R_114e_14866878 );
buf ( n6053 , R_136c_13d5ce58 );
buf ( n6054 , R_176d_15883e18 );
buf ( n6055 , R_198b_123ba938 );
buf ( n6056 , R_bb0_11635198 );
buf ( n6057 , R_6ad_14b295f8 );
buf ( n6058 , R_591_123b56b8 );
buf ( n6059 , R_ccc_13c02f78 );
buf ( n6060 , R_11cf_13dedd78 );
buf ( n6061 , R_12eb_156ab598 );
buf ( n6062 , R_17ee_117f2a78 );
buf ( n6063 , R_190a_1162b238 );
buf ( n6064 , R_7d4_14a0fe18 );
buf ( n6065 , R_df3_14b1e478 );
buf ( n6066 , R_a89_13dd9278 );
buf ( n6067 , R_10a8_13d52958 );
buf ( n6068 , R_1412_11c6f198 );
buf ( n6069 , R_16c7_13d27d58 );
buf ( n6070 , R_1a31_140b9d78 );
buf ( n6071 , R_c19_1700d408 );
buf ( n6072 , R_5fa_13df88b8 );
buf ( n6073 , R_644_13d23938 );
buf ( n6074 , R_c63_1162e258 );
buf ( n6075 , R_1238_13df9a38 );
buf ( n6076 , R_1282_13c2acf8 );
buf ( n6077 , R_1857_13cd2ed8 );
buf ( n6078 , R_18a1_156aefb8 );
buf ( n6079 , R_6f0_140ae658 );
buf ( n6080 , R_b6d_123b4178 );
buf ( n6081 , R_d0f_150df0f8 );
buf ( n6082 , R_118c_14a17898 );
buf ( n6083 , R_132e_13bed758 );
buf ( n6084 , R_17ab_13cd0d18 );
buf ( n6085 , R_194d_1008c438 );
buf ( n6086 , R_802_13d3e5d8 );
buf ( n6087 , R_e21_14a0aaf8 );
buf ( n6088 , R_a5b_13bf7e38 );
buf ( n6089 , R_107a_13d1ed98 );
buf ( n6090 , R_1440_124c4d58 );
buf ( n6091 , R_1699_140b0318 );
buf ( n6092 , R_1a5f_124c5618 );
buf ( n6093 , R_8fc_13bebd18 );
buf ( n6094 , R_961_12fbe358 );
buf ( n6095 , R_f1b_13ddafd8 );
buf ( n6096 , R_f80_1486f478 );
buf ( n6097 , R_153a_116341f8 );
buf ( n6098 , R_159f_1008d338 );
buf ( n6099 , R_ada_15812f78 );
buf ( n6100 , R_da2_156b5ef8 );
buf ( n6101 , R_783_123ba898 );
buf ( n6102 , R_10f9_123b7a58 );
buf ( n6103 , R_13c1_13d3bfb8 );
buf ( n6104 , R_1718_156b8018 );
buf ( n6105 , R_19e0_13dd4ef8 );
buf ( n6106 , R_6cb_117f2258 );
buf ( n6107 , R_573_1162dfd8 );
buf ( n6108 , R_cea_13d5be18 );
buf ( n6109 , R_b92_13c01998 );
buf ( n6110 , R_11b1_1700a208 );
buf ( n6111 , R_1309_117e8898 );
buf ( n6112 , R_17d0_156b8d38 );
buf ( n6113 , R_1928_14a0f738 );
buf ( n6114 , R_eb1_156b8f18 );
buf ( n6115 , R_892_11c69018 );
buf ( n6116 , R_9cb_13bed1b8 );
buf ( n6117 , R_fea_13d2b3b8 );
buf ( n6118 , R_14d0_13ccf698 );
buf ( n6119 , R_1609_13cd30b8 );
buf ( n6120 , R_67f_13cd88d8 );
buf ( n6121 , R_c9e_1580ee78 );
buf ( n6122 , R_bde_123b3138 );
buf ( n6123 , R_5bf_117f0b38 );
buf ( n6124 , R_11fd_1162f3d8 );
buf ( n6125 , R_12bd_13bf9698 );
buf ( n6126 , R_181c_13bf7758 );
buf ( n6127 , R_18dc_15817258 );
buf ( n6128 , R_c8c_13b97258 );
buf ( n6129 , R_bf0_13c26d38 );
buf ( n6130 , R_5d1_14875af8 );
buf ( n6131 , R_66d_1700eda8 );
buf ( n6132 , R_120f_156b0a98 );
buf ( n6133 , R_12ab_1486c278 );
buf ( n6134 , R_182e_116366d8 );
buf ( n6135 , R_18ca_11c708b8 );
buf ( n6136 , R_f2e_13dddb98 );
buf ( n6137 , R_90f_13b8e3d8 );
buf ( n6138 , R_94e_117f3c98 );
buf ( n6139 , R_f6d_13bf7a78 );
buf ( n6140 , R_154d_13df8c78 );
buf ( n6141 , R_158c_13d278f8 );
buf ( n6142 , R_702_13de3598 );
buf ( n6143 , R_b5b_13d45bf8 );
buf ( n6144 , R_d21_156ac038 );
buf ( n6145 , R_117a_14b292d8 );
buf ( n6146 , R_1340_123bbab8 );
buf ( n6147 , R_1799_13df1018 );
buf ( n6148 , R_195f_13b92e38 );
buf ( n6149 , R_d38_156afaf8 );
buf ( n6150 , R_719_13d1d498 );
buf ( n6151 , R_b44_13df7238 );
buf ( n6152 , R_1163_13b91358 );
buf ( n6153 , R_1357_13d5bcd8 );
buf ( n6154 , R_1782_1486c138 );
buf ( n6155 , R_1976_14b1de38 );
buf ( n6156 , R_695_13b93b58 );
buf ( n6157 , R_bc8_13dfb3d8 );
buf ( n6158 , R_cb4_15817078 );
buf ( n6159 , R_5a9_156b6998 );
buf ( n6160 , R_11e7_13bf3298 );
buf ( n6161 , R_12d3_14b28338 );
buf ( n6162 , R_1806_123b6dd8 );
buf ( n6163 , R_18f2_13d40338 );
buf ( n6164 , R_a06_158876f8 );
buf ( n6165 , R_857_14874dd8 );
buf ( n6166 , R_e76_13bf0958 );
buf ( n6167 , R_1025_13d59438 );
buf ( n6168 , R_1495_14870238 );
buf ( n6169 , R_1644_15ff4d88 );
buf ( n6170 , R_6fb_156b9378 );
buf ( n6171 , R_b62_123bb298 );
buf ( n6172 , R_d1a_117ee1f8 );
buf ( n6173 , R_1181_148748d8 );
buf ( n6174 , R_1339_1580de38 );
buf ( n6175 , R_17a0_13dd7478 );
buf ( n6176 , R_1958_156ae5b8 );
buf ( n6177 , R_97a_117eaff8 );
buf ( n6178 , R_f02_13d538f8 );
buf ( n6179 , R_8e3_13c107b8 );
buf ( n6180 , R_f99_1580efb8 );
buf ( n6181 , R_1521_148676d8 );
buf ( n6182 , R_15b8_13b93e78 );
buf ( n6183 , R_829_13b954f8 );
buf ( n6184 , R_a34_156b03b8 );
buf ( n6185 , R_e48_15813d38 );
buf ( n6186 , R_1053_13cd3478 );
buf ( n6187 , R_1467_13b8be58 );
buf ( n6188 , R_1672_13cd1df8 );
buf ( n6189 , R_e89_13de0078 );
buf ( n6190 , R_9f3_156b0598 );
buf ( n6191 , R_86a_13b94378 );
buf ( n6192 , R_1012_123bf618 );
buf ( n6193 , R_14a8_13becdf8 );
buf ( n6194 , R_1631_1486c9f8 );
buf ( n6195 , R_acd_1008bfd8 );
buf ( n6196 , R_daf_123b59d8 );
buf ( n6197 , R_790_13d2bd18 );
buf ( n6198 , R_10ec_1700b6a8 );
buf ( n6199 , R_13ce_13df2a58 );
buf ( n6200 , R_170b_14b26178 );
buf ( n6201 , R_19ed_148709b8 );
buf ( n6202 , R_a31_13cd7d98 );
buf ( n6203 , R_82c_140b1e98 );
buf ( n6204 , R_e4b_116316d8 );
buf ( n6205 , R_1050_13d3d138 );
buf ( n6206 , R_146a_123bd318 );
buf ( n6207 , R_166f_140ad118 );
buf ( n6208 , R_eac_1007f418 );
buf ( n6209 , R_88d_13bf99b8 );
buf ( n6210 , R_9d0_17010748 );
buf ( n6211 , R_fef_1580b138 );
buf ( n6212 , R_14cb_13d44258 );
buf ( n6213 , R_160e_11632a38 );
buf ( n6214 , R_826_13c24cb8 );
buf ( n6215 , R_a37_158112b8 );
buf ( n6216 , R_e45_15fee168 );
buf ( n6217 , R_1056_15fedc68 );
buf ( n6218 , R_1464_13d3fa78 );
buf ( n6219 , R_1675_14b28dd8 );
buf ( n6220 , R_eb6_11c69518 );
buf ( n6221 , R_897_11c69338 );
buf ( n6222 , R_9c6_156ad258 );
buf ( n6223 , R_fe5_14b1f4b8 );
buf ( n6224 , R_14d5_14871a98 );
buf ( n6225 , R_1604_13beed38 );
buf ( n6226 , R_9ef_14a126b8 );
buf ( n6227 , R_e8d_13c07578 );
buf ( n6228 , R_86e_13ded738 );
buf ( n6229 , R_100e_100810d8 );
buf ( n6230 , R_14ac_13cce158 );
buf ( n6231 , R_162d_13c0adb8 );
buf ( n6232 , R_7cb_14a0acd8 );
buf ( n6233 , R_dea_123c0798 );
buf ( n6234 , R_a92_13d25238 );
buf ( n6235 , R_10b1_13d55478 );
buf ( n6236 , R_1409_1587f638 );
buf ( n6237 , R_16d0_13c02ed8 );
buf ( n6238 , R_1a28_14a12398 );
buf ( n6239 , R_ee0_13d1ffb8 );
buf ( n6240 , R_99c_14a0f418 );
buf ( n6241 , R_8c1_14b25818 );
buf ( n6242 , R_fbb_123b70f8 );
buf ( n6243 , R_14ff_1580bf98 );
buf ( n6244 , R_15da_140ba138 );
buf ( n6245 , R_687_14b23fb8 );
buf ( n6246 , R_bd6_13dd71f8 );
buf ( n6247 , R_ca6_123bd098 );
buf ( n6248 , R_5b7_117e8cf8 );
buf ( n6249 , R_11f5_15815318 );
buf ( n6250 , R_12c5_14a0f7d8 );
buf ( n6251 , R_1814_170116e8 );
buf ( n6252 , R_18e4_12fc1d78 );
buf ( n6253 , R_812_12fc0018 );
buf ( n6254 , R_a4b_13bf22f8 );
buf ( n6255 , R_e31_13bee338 );
buf ( n6256 , R_106a_13d56a58 );
buf ( n6257 , R_1450_1580a738 );
buf ( n6258 , R_1689_14a0c218 );
buf ( n6259 , R_e85_156aa878 );
buf ( n6260 , R_9f7_13d246f8 );
buf ( n6261 , R_866_15ffb868 );
buf ( n6262 , R_1016_156af698 );
buf ( n6263 , R_14a4_11c6ec98 );
buf ( n6264 , R_1635_15ff7588 );
buf ( n6265 , R_8ee_140ae338 );
buf ( n6266 , R_96f_13d3b8d8 );
buf ( n6267 , R_f0d_13d4fa78 );
buf ( n6268 , R_f8e_13d541b8 );
buf ( n6269 , R_152c_156b2258 );
buf ( n6270 , R_15ad_13d58218 );
buf ( n6271 , R_9de_124c3458 );
buf ( n6272 , R_e9e_123b9038 );
buf ( n6273 , R_87f_117f0958 );
buf ( n6274 , R_ffd_13c27f58 );
buf ( n6275 , R_14bd_13cd71b8 );
buf ( n6276 , R_161c_156b6178 );
buf ( n6277 , R_aec_14866b98 );
buf ( n6278 , R_d90_10081718 );
buf ( n6279 , R_771_1007ee78 );
buf ( n6280 , R_110b_14b24f58 );
buf ( n6281 , R_13af_158110d8 );
buf ( n6282 , R_172a_11c6feb8 );
buf ( n6283 , R_19ce_11c6fc38 );
buf ( n6284 , R_6d4_15ff47e8 );
buf ( n6285 , R_56a_17018268 );
buf ( n6286 , R_cf3_150e21b8 );
buf ( n6287 , R_b89_13cd67b8 );
buf ( n6288 , R_11a8_13c0ab38 );
buf ( n6289 , R_1312_15881758 );
buf ( n6290 , R_17c7_1580cf38 );
buf ( n6291 , R_1931_11c6b4f8 );
buf ( n6292 , R_7be_13d51918 );
buf ( n6293 , R_ddd_10083fb8 );
buf ( n6294 , R_a9f_140b7b18 );
buf ( n6295 , R_10be_1162c138 );
buf ( n6296 , R_13fc_13b967b8 );
buf ( n6297 , R_16dd_15ffb728 );
buf ( n6298 , R_1a1b_13d3ab18 );
buf ( n6299 , R_a2e_1580aeb8 );
buf ( n6300 , R_82f_14b26cb8 );
buf ( n6301 , R_e4e_13dec798 );
buf ( n6302 , R_104d_13de2af8 );
buf ( n6303 , R_146d_156b1998 );
buf ( n6304 , R_166c_117f5958 );
buf ( n6305 , R_d50_156b51d8 );
buf ( n6306 , R_b2c_12fc0478 );
buf ( n6307 , R_731_15ffaa08 );
buf ( n6308 , R_114b_13ddbed8 );
buf ( n6309 , R_136f_11c6c718 );
buf ( n6310 , R_176a_11628f38 );
buf ( n6311 , R_198e_150e3518 );
buf ( n6312 , R_ed9_15ff7948 );
buf ( n6313 , R_9a3_13c1fad8 );
buf ( n6314 , R_8ba_116386b8 );
buf ( n6315 , R_fc2_1700f7a8 );
buf ( n6316 , R_14f8_117f15d8 );
buf ( n6317 , R_15e1_150dcd58 );
buf ( n6318 , R_b16_13c1c1f8 );
buf ( n6319 , R_d66_13b8b1d8 );
buf ( n6320 , R_747_158864d8 );
buf ( n6321 , R_1135_156b68f8 );
buf ( n6322 , R_1385_1580b278 );
buf ( n6323 , R_1754_156add98 );
buf ( n6324 , R_19a4_13d4fd98 );
buf ( n6325 , R_823_11c6f2d8 );
buf ( n6326 , R_a3a_14871318 );
buf ( n6327 , R_e42_156ade38 );
buf ( n6328 , R_1059_13c0f318 );
buf ( n6329 , R_1461_14a1a138 );
buf ( n6330 , R_1678_14a0fd78 );
buf ( n6331 , R_8d9_158837d8 );
buf ( n6332 , R_984_15882d38 );
buf ( n6333 , R_ef8_15816998 );
buf ( n6334 , R_fa3_15815458 );
buf ( n6335 , R_1517_156ad898 );
buf ( n6336 , R_15c2_11630c38 );
buf ( n6337 , R_af3_13beae18 );
buf ( n6338 , R_d89_117e8938 );
buf ( n6339 , R_76a_123bceb8 );
buf ( n6340 , R_1112_13c20c58 );
buf ( n6341 , R_13a8_117f4a58 );
buf ( n6342 , R_1731_1008a818 );
buf ( n6343 , R_19c7_13d38bd8 );
buf ( n6344 , R_b04_156aed38 );
buf ( n6345 , R_d78_13cd7758 );
buf ( n6346 , R_759_11629938 );
buf ( n6347 , R_1123_15ffb908 );
buf ( n6348 , R_1397_13d37a58 );
buf ( n6349 , R_1742_13d237f8 );
buf ( n6350 , R_19b6_14b20778 );
buf ( n6351 , R_c64_13c1fdf8 );
buf ( n6352 , R_c18_12fc23b8 );
buf ( n6353 , R_5f9_13b8f238 );
buf ( n6354 , R_645_140b2118 );
buf ( n6355 , R_1237_1162dad8 );
buf ( n6356 , R_1283_14a18798 );
buf ( n6357 , R_1856_117f4878 );
buf ( n6358 , R_18a2_13d53998 );
buf ( n6359 , R_f2d_100818f8 );
buf ( n6360 , R_90e_11629898 );
buf ( n6361 , R_94f_15888738 );
buf ( n6362 , R_f6e_14a188d8 );
buf ( n6363 , R_154c_14a147d8 );
buf ( n6364 , R_158d_15ff0a08 );
buf ( n6365 , R_9eb_117ef2d8 );
buf ( n6366 , R_e91_1580e3d8 );
buf ( n6367 , R_872_13c0c7f8 );
buf ( n6368 , R_100a_117f81f8 );
buf ( n6369 , R_14b0_124c2f58 );
buf ( n6370 , R_1629_14a0b6d8 );
buf ( n6371 , R_656_15886bb8 );
buf ( n6372 , R_c75_156b0db8 );
buf ( n6373 , R_c07_124c4cb8 );
buf ( n6374 , R_5e8_1162f298 );
buf ( n6375 , R_1226_13b8e018 );
buf ( n6376 , R_1294_13b91ad8 );
buf ( n6377 , R_1845_13cd83d8 );
buf ( n6378 , R_18b3_13d1e118 );
buf ( n6379 , R_ba0_156b4698 );
buf ( n6380 , R_6bd_13c0ec38 );
buf ( n6381 , R_581_13d1d8f8 );
buf ( n6382 , R_cdc_13cd9378 );
buf ( n6383 , R_11bf_123b6c98 );
buf ( n6384 , R_12fb_150e3018 );
buf ( n6385 , R_17de_14b20458 );
buf ( n6386 , R_191a_123b2cd8 );
buf ( n6387 , R_d5e_14a10278 );
buf ( n6388 , R_b1e_13df7418 );
buf ( n6389 , R_73f_1587b998 );
buf ( n6390 , R_113d_13d58498 );
buf ( n6391 , R_137d_14a11b78 );
buf ( n6392 , R_175c_1587b218 );
buf ( n6393 , R_199c_17017408 );
buf ( n6394 , R_b09_15884f98 );
buf ( n6395 , R_d73_1580b4f8 );
buf ( n6396 , R_754_15811d58 );
buf ( n6397 , R_1128_10084d78 );
buf ( n6398 , R_1392_14a15db8 );
buf ( n6399 , R_1747_17018588 );
buf ( n6400 , R_19b1_13dd9f98 );
buf ( n6401 , R_d35_14a11858 );
buf ( n6402 , R_716_156b9c38 );
buf ( n6403 , R_b47_140af4b8 );
buf ( n6404 , R_1166_13ccdcf8 );
buf ( n6405 , R_1354_13d41738 );
buf ( n6406 , R_1785_1162d218 );
buf ( n6407 , R_1973_14a18338 );
buf ( n6408 , R_a2b_13c1e6d8 );
buf ( n6409 , R_832_13df5c58 );
buf ( n6410 , R_e51_156ab278 );
buf ( n6411 , R_104a_14a108b8 );
buf ( n6412 , R_1470_15887bf8 );
buf ( n6413 , R_1669_158828d8 );
buf ( n6414 , R_e81_1007dc58 );
buf ( n6415 , R_9fb_1486fb58 );
buf ( n6416 , R_862_156ab138 );
buf ( n6417 , R_101a_13d5a798 );
buf ( n6418 , R_14a0_13d38818 );
buf ( n6419 , R_1639_1162abf8 );
buf ( n6420 , R_ba5_140b4af8 );
buf ( n6421 , R_6b8_1580d898 );
buf ( n6422 , R_586_15ff8488 );
buf ( n6423 , R_cd7_156b7e38 );
buf ( n6424 , R_11c4_117ecad8 );
buf ( n6425 , R_12f6_17015ba8 );
buf ( n6426 , R_17e3_13c1dd78 );
buf ( n6427 , R_1915_14a17f78 );
buf ( n6428 , R_aff_140aba98 );
buf ( n6429 , R_d7d_148714f8 );
buf ( n6430 , R_75e_10084418 );
buf ( n6431 , R_111e_11635918 );
buf ( n6432 , R_139c_1580e0b8 );
buf ( n6433 , R_173d_13deffd8 );
buf ( n6434 , R_19bb_13df9df8 );
buf ( n6435 , R_7dd_13d28898 );
buf ( n6436 , R_dfc_156b9ff8 );
buf ( n6437 , R_a80_13ddc8d8 );
buf ( n6438 , R_109f_13cd2cf8 );
buf ( n6439 , R_141b_12fc10f8 );
buf ( n6440 , R_16be_13bf0098 );
buf ( n6441 , R_1a3a_156b79d8 );
buf ( n6442 , R_9d5_15ff1908 );
buf ( n6443 , R_ea7_14a124d8 );
buf ( n6444 , R_888_13deebd8 );
buf ( n6445 , R_ff4_13cd7b18 );
buf ( n6446 , R_14c6_13cd5d18 );
buf ( n6447 , R_1613_123bc198 );
buf ( n6448 , R_677_13c0c758 );
buf ( n6449 , R_c96_13c0d838 );
buf ( n6450 , R_be6_1162cf98 );
buf ( n6451 , R_5c7_1162f1f8 );
buf ( n6452 , R_1205_156b94b8 );
buf ( n6453 , R_12b5_158816b8 );
buf ( n6454 , R_1824_13c04f58 );
buf ( n6455 , R_18d4_13beb958 );
buf ( n6456 , R_f1a_124c4f38 );
buf ( n6457 , R_8fb_13c1e9f8 );
buf ( n6458 , R_962_14a15ef8 );
buf ( n6459 , R_f81_1580d438 );
buf ( n6460 , R_1539_14b267b8 );
buf ( n6461 , R_15a0_15ff32a8 );
buf ( n6462 , R_d28_156b3fb8 );
buf ( n6463 , R_709_117ea4b8 );
buf ( n6464 , R_b54_13c04c38 );
buf ( n6465 , R_1173_15810778 );
buf ( n6466 , R_1347_13dd5f38 );
buf ( n6467 , R_1792_13d39858 );
buf ( n6468 , R_1966_12fc2098 );
buf ( n6469 , R_a1b_123c17d8 );
buf ( n6470 , R_842_13bf4738 );
buf ( n6471 , R_e61_13cd0958 );
buf ( n6472 , R_103a_13ccdbb8 );
buf ( n6473 , R_1480_117f1e98 );
buf ( n6474 , R_1659_13c1fcb8 );
buf ( n6475 , R_820_17013088 );
buf ( n6476 , R_a3d_11c6bc78 );
buf ( n6477 , R_e3f_123c0e78 );
buf ( n6478 , R_105c_13dd87d8 );
buf ( n6479 , R_145e_13d5a3d8 );
buf ( n6480 , R_167b_14a19878 );
buf ( n6481 , R_ebb_13def998 );
buf ( n6482 , R_89c_1486e898 );
buf ( n6483 , R_9c1_13cd04f8 );
buf ( n6484 , R_fe0_15fee7a8 );
buf ( n6485 , R_14da_13b95818 );
buf ( n6486 , R_15ff_117f1538 );
buf ( n6487 , R_8d0_13ccd078 );
buf ( n6488 , R_98d_13cceab8 );
buf ( n6489 , R_eef_15ff2308 );
buf ( n6490 , R_fac_13df65b8 );
buf ( n6491 , R_150e_13bed398 );
buf ( n6492 , R_15cb_1580a558 );
buf ( n6493 , R_663_13c24218 );
buf ( n6494 , R_c82_11633bb8 );
buf ( n6495 , R_bfa_117f1d58 );
buf ( n6496 , R_5db_13c0d798 );
buf ( n6497 , R_1219_156b0f98 );
buf ( n6498 , R_12a1_15811e98 );
buf ( n6499 , R_1838_123c2098 );
buf ( n6500 , R_18c0_13ddb258 );
buf ( n6501 , R_bbb_13c08dd8 );
buf ( n6502 , R_6a2_14870cd8 );
buf ( n6503 , R_59c_1700ffc8 );
buf ( n6504 , R_cc1_13d5b0f8 );
buf ( n6505 , R_11da_14b1dcf8 );
buf ( n6506 , R_12e0_14b29c38 );
buf ( n6507 , R_17f9_13ddb438 );
buf ( n6508 , R_18ff_1162d538 );
buf ( n6509 , R_ecc_123bde58 );
buf ( n6510 , R_9b0_1587f458 );
buf ( n6511 , R_8ad_10082e38 );
buf ( n6512 , R_fcf_14a0e798 );
buf ( n6513 , R_14eb_140ad258 );
buf ( n6514 , R_15ee_117f3158 );
buf ( n6515 , R_d13_13c25e38 );
buf ( n6516 , R_6f4_156b4918 );
buf ( n6517 , R_b69_11c6e8d8 );
buf ( n6518 , R_1188_13cd35b8 );
buf ( n6519 , R_1332_11637d58 );
buf ( n6520 , R_17a7_117f6a38 );
buf ( n6521 , R_1951_156b6b78 );
buf ( n6522 , R_acf_13d503d8 );
buf ( n6523 , R_dad_13cd3838 );
buf ( n6524 , R_78e_13b929d8 );
buf ( n6525 , R_10ee_1587c438 );
buf ( n6526 , R_13cc_1587b3f8 );
buf ( n6527 , R_170d_12fbf9d8 );
buf ( n6528 , R_19eb_15ff53c8 );
buf ( n6529 , R_8c8_12fbe038 );
buf ( n6530 , R_ee7_13c03dd8 );
buf ( n6531 , R_995_13d50518 );
buf ( n6532 , R_fb4_156b0e58 );
buf ( n6533 , R_1506_156b9e18 );
buf ( n6534 , R_15d3_123b5ed8 );
buf ( n6535 , R_b9b_13dfa118 );
buf ( n6536 , R_6c2_14b1d618 );
buf ( n6537 , R_57c_13d464b8 );
buf ( n6538 , R_ce1_13d27358 );
buf ( n6539 , R_11ba_13cda458 );
buf ( n6540 , R_1300_13dec478 );
buf ( n6541 , R_17d9_156af918 );
buf ( n6542 , R_191f_14a0d578 );
buf ( n6543 , R_7e4_117f6c18 );
buf ( n6544 , R_e03_13b8c718 );
buf ( n6545 , R_a79_13d52db8 );
buf ( n6546 , R_1098_13cd2438 );
buf ( n6547 , R_1422_13cd7f78 );
buf ( n6548 , R_16b7_14b28518 );
buf ( n6549 , R_1a41_150e4d78 );
buf ( n6550 , R_ae5_17012048 );
buf ( n6551 , R_d97_1162ab58 );
buf ( n6552 , R_778_13d52098 );
buf ( n6553 , R_1104_13dd7a18 );
buf ( n6554 , R_13b6_14a17118 );
buf ( n6555 , R_1723_13d50018 );
buf ( n6556 , R_19d5_117edc58 );
buf ( n6557 , R_d53_13c0ae58 );
buf ( n6558 , R_b29_13b95c78 );
buf ( n6559 , R_734_14a0f558 );
buf ( n6560 , R_1148_117f6218 );
buf ( n6561 , R_1372_11c6cd58 );
buf ( n6562 , R_1767_11c691f8 );
buf ( n6563 , R_1991_13cd58b8 );
buf ( n6564 , R_f2c_15814d78 );
buf ( n6565 , R_90d_158848b8 );
buf ( n6566 , R_950_140b3798 );
buf ( n6567 , R_f6f_14a1a318 );
buf ( n6568 , R_154b_11632218 );
buf ( n6569 , R_158e_14a0b1d8 );
buf ( n6570 , R_ec6_13d37b98 );
buf ( n6571 , R_8a7_1580e6f8 );
buf ( n6572 , R_9b6_14a0cc18 );
buf ( n6573 , R_fd5_1580cc18 );
buf ( n6574 , R_14e5_13b8fd78 );
buf ( n6575 , R_15f4_170165a8 );
buf ( n6576 , R_7c0_100854f8 );
buf ( n6577 , R_ddf_13b92898 );
buf ( n6578 , R_a9d_1162c318 );
buf ( n6579 , R_10bc_140b7d98 );
buf ( n6580 , R_13fe_13cd60d8 );
buf ( n6581 , R_16db_156aaf58 );
buf ( n6582 , R_1a1d_13cd9ff8 );
buf ( n6583 , R_7f5_13b9a1d8 );
buf ( n6584 , R_e14_123bf078 );
buf ( n6585 , R_a68_150dbbd8 );
buf ( n6586 , R_1087_1587ad18 );
buf ( n6587 , R_1433_13dd7978 );
buf ( n6588 , R_16a6_13df8458 );
buf ( n6589 , R_1a52_11c70778 );
buf ( n6590 , R_646_156ad618 );
buf ( n6591 , R_c65_10086538 );
buf ( n6592 , R_c17_13ccb3b8 );
buf ( n6593 , R_5f8_1580f418 );
buf ( n6594 , R_1236_1587e558 );
buf ( n6595 , R_1284_14a1a458 );
buf ( n6596 , R_1855_10084a58 );
buf ( n6597 , R_18a3_1700b1a8 );
buf ( n6598 , R_69c_156b9058 );
buf ( n6599 , R_bc1_13bee298 );
buf ( n6600 , R_cbb_13ccbbd8 );
buf ( n6601 , R_5a2_15813658 );
buf ( n6602 , R_11e0_1587e878 );
buf ( n6603 , R_12da_14b29d78 );
buf ( n6604 , R_17ff_14a10b38 );
buf ( n6605 , R_18f9_14a16718 );
buf ( n6606 , R_adc_156ae6f8 );
buf ( n6607 , R_da0_13bf5db8 );
buf ( n6608 , R_781_13d42f98 );
buf ( n6609 , R_10fb_10085778 );
buf ( n6610 , R_13bf_123bf6b8 );
buf ( n6611 , R_171a_150deb58 );
buf ( n6612 , R_19de_117ef918 );
buf ( n6613 , R_9e7_13d54578 );
buf ( n6614 , R_e95_13d26ef8 );
buf ( n6615 , R_876_13d41698 );
buf ( n6616 , R_1006_13c08f18 );
buf ( n6617 , R_14b4_1700e268 );
buf ( n6618 , R_1625_13b96d58 );
buf ( n6619 , R_807_13cd8478 );
buf ( n6620 , R_e26_1700df48 );
buf ( n6621 , R_a56_124c4ad8 );
buf ( n6622 , R_1075_15883b98 );
buf ( n6623 , R_1445_15880218 );
buf ( n6624 , R_1694_13d218b8 );
buf ( n6625 , R_1a64_13ccac38 );
buf ( n6626 , R_a28_13cd9918 );
buf ( n6627 , R_835_140b35b8 );
buf ( n6628 , R_e54_14a179d8 );
buf ( n6629 , R_1047_14b26df8 );
buf ( n6630 , R_1473_156b60d8 );
buf ( n6631 , R_1666_14a165d8 );
buf ( n6632 , R_b0e_14a15818 );
buf ( n6633 , R_d6e_14a0c998 );
buf ( n6634 , R_74f_13c24678 );
buf ( n6635 , R_112d_1162be18 );
buf ( n6636 , R_138d_13b92258 );
buf ( n6637 , R_174c_116339d8 );
buf ( n6638 , R_19ac_14b1b4f8 );
buf ( n6639 , R_bb5_13cd29d8 );
buf ( n6640 , R_6a8_1162e618 );
buf ( n6641 , R_596_13dd6398 );
buf ( n6642 , R_cc7_123b4b78 );
buf ( n6643 , R_11d4_15ff30c8 );
buf ( n6644 , R_12e6_14a0ff58 );
buf ( n6645 , R_17f3_13ddb578 );
buf ( n6646 , R_1905_1486dfd8 );
buf ( n6647 , R_baa_14a15278 );
buf ( n6648 , R_6b3_17011288 );
buf ( n6649 , R_58b_140b1c18 );
buf ( n6650 , R_cd2_13d24dd8 );
buf ( n6651 , R_11c9_14b25278 );
buf ( n6652 , R_12f1_1587da18 );
buf ( n6653 , R_17e8_1587c078 );
buf ( n6654 , R_1910_12fc0978 );
buf ( n6655 , R_66e_17014348 );
buf ( n6656 , R_c8d_123b7ff8 );
buf ( n6657 , R_bef_14a167b8 );
buf ( n6658 , R_5d0_13c1db98 );
buf ( n6659 , R_120e_13c0d518 );
buf ( n6660 , R_12ac_13ccaf58 );
buf ( n6661 , R_182d_140b0098 );
buf ( n6662 , R_18cb_123b9e98 );
buf ( n6663 , R_8b3_13c0d298 );
buf ( n6664 , R_ed2_1580c538 );
buf ( n6665 , R_9aa_124c51b8 );
buf ( n6666 , R_fc9_13b8d118 );
buf ( n6667 , R_14f1_150e8978 );
buf ( n6668 , R_15e8_15884db8 );
buf ( n6669 , R_8e2_13bf6858 );
buf ( n6670 , R_97b_150e7a78 );
buf ( n6671 , R_f01_14a13e78 );
buf ( n6672 , R_f9a_116364f8 );
buf ( n6673 , R_1520_1162d678 );
buf ( n6674 , R_15b9_13d21a98 );
buf ( n6675 , R_7fa_123bbbf8 );
buf ( n6676 , R_e19_13d59ed8 );
buf ( n6677 , R_a63_14a16678 );
buf ( n6678 , R_1082_13c09d78 );
buf ( n6679 , R_1438_13bf2398 );
buf ( n6680 , R_16a1_14a16cb8 );
buf ( n6681 , R_1a57_13c28a98 );
buf ( n6682 , R_81d_1580d078 );
buf ( n6683 , R_a40_123bcd78 );
buf ( n6684 , R_e3c_117f2c58 );
buf ( n6685 , R_105f_13de2558 );
buf ( n6686 , R_145b_11633e38 );
buf ( n6687 , R_167e_1486d858 );
buf ( n6688 , R_7f0_13b90458 );
buf ( n6689 , R_e0f_140ab138 );
buf ( n6690 , R_a6d_117ee838 );
buf ( n6691 , R_108c_13bf90f8 );
buf ( n6692 , R_142e_11632538 );
buf ( n6693 , R_16ab_140b8d38 );
buf ( n6694 , R_1a4d_11c70bd8 );
buf ( n6695 , R_7d6_14b1e3d8 );
buf ( n6696 , R_df5_1580eab8 );
buf ( n6697 , R_a87_14a10138 );
buf ( n6698 , R_10a6_117efa58 );
buf ( n6699 , R_1414_1162b9b8 );
buf ( n6700 , R_16c5_14a10db8 );
buf ( n6701 , R_1a33_1486ebb8 );
buf ( n6702 , R_f0c_140b21b8 );
buf ( n6703 , R_8ed_11636d18 );
buf ( n6704 , R_970_13c0f818 );
buf ( n6705 , R_f8f_11632fd8 );
buf ( n6706 , R_152b_13beb778 );
buf ( n6707 , R_15ae_123b2eb8 );
buf ( n6708 , R_e6b_13b8ded8 );
buf ( n6709 , R_a11_158133d8 );
buf ( n6710 , R_84c_13bef918 );
buf ( n6711 , R_1030_140b72f8 );
buf ( n6712 , R_148a_140b0598 );
buf ( n6713 , R_164f_13d52778 );
buf ( n6714 , R_afa_123c0c98 );
buf ( n6715 , R_d82_13cd1858 );
buf ( n6716 , R_763_1580e298 );
buf ( n6717 , R_1119_1587c118 );
buf ( n6718 , R_13a1_158898b8 );
buf ( n6719 , R_1738_11c6f878 );
buf ( n6720 , R_19c0_1007ded8 );
buf ( n6721 , R_e7d_15811538 );
buf ( n6722 , R_9ff_13d245b8 );
buf ( n6723 , R_85e_13cd3018 );
buf ( n6724 , R_101e_13d5d8f8 );
buf ( n6725 , R_149c_13d5a978 );
buf ( n6726 , R_163d_13ccd438 );
buf ( n6727 , R_b8d_156aae18 );
buf ( n6728 , R_6d0_1162bb98 );
buf ( n6729 , R_56e_10086e98 );
buf ( n6730 , R_cef_14870eb8 );
buf ( n6731 , R_11ac_13c24498 );
buf ( n6732 , R_130e_14a17758 );
buf ( n6733 , R_17cb_14a0e478 );
buf ( n6734 , R_192d_123becb8 );
buf ( n6735 , R_d32_13d20558 );
buf ( n6736 , R_713_15882978 );
buf ( n6737 , R_b4a_13d22cb8 );
buf ( n6738 , R_1169_123b7c38 );
buf ( n6739 , R_1351_14a14558 );
buf ( n6740 , R_1788_13ccae18 );
buf ( n6741 , R_1970_124c43f8 );
buf ( n6742 , R_7cd_13d58df8 );
buf ( n6743 , R_dec_156ae518 );
buf ( n6744 , R_a90_13dd8058 );
buf ( n6745 , R_10af_117f0818 );
buf ( n6746 , R_140b_1580d1b8 );
buf ( n6747 , R_16ce_117ebe58 );
buf ( n6748 , R_1a2a_15810e58 );
buf ( n6749 , R_e72_13c1e8b8 );
buf ( n6750 , R_a0a_13d54438 );
buf ( n6751 , R_853_123bd778 );
buf ( n6752 , R_1029_13cd2898 );
buf ( n6753 , R_1491_117f33d8 );
buf ( n6754 , R_1648_15ff12c8 );
buf ( n6755 , R_80f_13d449d8 );
buf ( n6756 , R_a4e_13b8e798 );
buf ( n6757 , R_e2e_13dd57b8 );
buf ( n6758 , R_106d_13b8b598 );
buf ( n6759 , R_144d_13cd65d8 );
buf ( n6760 , R_168c_15ff1c28 );
buf ( R_187c_13cca558 , n30988 );
buf ( R_125d_156aaaf8 , n31654 );
buf ( R_c3e_13d2c178 , C0 );
buf ( R_61f_117eb278 , n31656 );
buf ( R_187d_117f5b38 , n32505 );
buf ( R_125e_13b8fe18 , C0 );
buf ( R_c3f_123b4358 , n32506 );
buf ( R_187b_13ccb278 , n32507 );
buf ( R_620_13dfb518 , n32508 );
buf ( R_125c_15816b78 , n32509 );
buf ( R_c3d_13c22918 , n33386 );
buf ( R_61e_14a0c538 , C0 );
buf ( R_5e7_10080958 , n33387 );
buf ( R_c06_170189e8 , C0 );
buf ( R_18b4_1162f978 , n33388 );
buf ( R_1225_13c08298 , n33982 );
buf ( R_1844_117ef378 , n33983 );
buf ( R_1295_123bcf58 , n34146 );
buf ( R_c76_15ff42e8 , C0 );
buf ( R_657_13bf5c78 , n34147 );
buf ( R_187e_140ac0d8 , C0 );
buf ( R_125f_13c0f638 , n34148 );
buf ( R_c40_1580a9b8 , n34149 );
buf ( R_621_11c70318 , n35066 );
buf ( R_187a_13ddd2d8 , C0 );
buf ( R_61d_123b84f8 , n35124 );
buf ( R_125b_1162bf58 , n35125 );
buf ( R_c3c_15ff9928 , n35126 );
buf ( R_12be_13ccf378 , C0 );
buf ( R_5be_11c6a738 , C0 );
buf ( R_bdd_17016508 , n35177 );
buf ( R_c9f_11636598 , n35178 );
buf ( R_11fc_13ddf7b8 , n35179 );
buf ( R_680_10085638 , n35180 );
buf ( R_181b_13d430d8 , n35181 );
buf ( R_18dd_13c062b8 , n35371 );
buf ( R_180c_156b4eb8 , n35372 );
buf ( R_12cd_13d535d8 , n35528 );
buf ( R_5af_1700c3c8 , n35550 );
buf ( R_cae_14a14ff8 , C0 );
buf ( R_bce_15ff4608 , C0 );
buf ( R_68f_13befcd8 , n35551 );
buf ( R_18ec_13d204b8 , n35552 );
buf ( R_11ed_116361d8 , n35587 );
buf ( R_187f_15811038 , n35588 );
buf ( R_1260_13d3b6f8 , n35589 );
buf ( R_c41_14a0bef8 , n35643 );
buf ( R_622_123b3bd8 , C0 );
buf ( R_61c_13d56378 , n35644 );
buf ( R_c3b_150e7c58 , n35645 );
buf ( R_1879_15ff5c88 , n35682 );
buf ( R_125a_13bf58b8 , C0 );
buf ( R_f82_13c1cd38 , C0 );
buf ( R_963_13c209d8 , n35683 );
buf ( R_8fa_117ec678 , C0 );
buf ( R_f19_15ff0648 , n37510 );
buf ( R_1538_13d29bf8 , n37511 );
buf ( R_15a1_150e22f8 , n39363 );
buf ( R_158f_13cd9058 , n39364 );
buf ( R_f70_17015608 , n39365 );
buf ( R_951_156b2578 , n39809 );
buf ( R_90c_13c0e0f8 , n39810 );
buf ( R_f2b_140b8838 , n39811 );
buf ( R_154a_1587f278 , C0 );
buf ( R_1880_13c22738 , n39812 );
buf ( R_1261_13ccc0d8 , n39867 );
buf ( R_c42_117eb818 , C0 );
buf ( R_623_140b3158 , n39868 );
buf ( R_61b_11c70458 , n39869 );
buf ( R_c3a_13b96218 , C0 );
buf ( R_1259_13d23578 , n39921 );
buf ( R_1878_1162da38 , n39922 );
buf ( R_ce6_14875d78 , C0 );
buf ( R_1924_13d1df38 , n39923 );
buf ( R_11b5_13d56f58 , n40158 );
buf ( R_577_1162c818 , n40160 );
buf ( R_6c7_10082438 , n40161 );
buf ( R_17d4_13cda278 , n40162 );
buf ( R_1305_10081fd8 , n41282 );
buf ( R_b96_15812b18 , C0 );
buf ( R_1881_156b0638 , n41328 );
buf ( R_1262_12fc1698 , C0 );
buf ( R_c43_140b0138 , n41329 );
buf ( R_624_13d421d8 , n41330 );
buf ( R_61a_14b2a318 , C0 );
buf ( R_c39_117eaeb8 , n41380 );
buf ( R_1258_117e8618 , n41381 );
buf ( R_1877_1162cdb8 , n41382 );
buf ( R_119b_15ffa3c8 , n41383 );
buf ( R_55d_13b8e5b8 , n41385 );
buf ( R_131f_158106d8 , n41386 );
buf ( R_6e1_13c0fb38 , n41442 );
buf ( R_17ba_15fed6c8 , C0 );
buf ( R_b7c_13b96e98 , n41443 );
buf ( R_193e_123b6018 , C0 );
buf ( R_d00_117ec358 , n41444 );
buf ( R_1323_13d5b878 , n41445 );
buf ( R_6e5_15ff5328 , n41509 );
buf ( R_559_13c024d8 , n41511 );
buf ( R_1197_13bf4918 , n41512 );
buf ( R_1942_11c6dd98 , C0 );
buf ( R_d04_14a16df8 , n41513 );
buf ( R_17b6_13dec158 , C0 );
buf ( R_b78_13c10c18 , n41514 );
buf ( R_13ca_13d2c718 , C0 );
buf ( R_19e9_13bf62b8 , n41539 );
buf ( R_170f_150defb8 , n41540 );
buf ( R_10f0_140b1ad8 , n41541 );
buf ( R_ad1_11c6ac38 , n41599 );
buf ( R_78c_13d5d3f8 , n41600 );
buf ( R_dab_140b3dd8 , n41601 );
buf ( R_883_13b936f8 , n41602 );
buf ( R_ff9_11631958 , n42165 );
buf ( R_ea2_150dd758 , C0 );
buf ( R_9da_13cd8018 , C0 );
buf ( R_1618_117f3658 , n42166 );
buf ( R_14c1_123ba4d8 , n42233 );
buf ( R_b5e_14a0f918 , C0 );
buf ( R_179c_123bb018 , n42234 );
buf ( R_133d_13cd4e18 , n42300 );
buf ( R_6ff_14a0a918 , n42301 );
buf ( R_195c_150ddf78 , n42302 );
buf ( R_117d_123b8c78 , n42372 );
buf ( R_d1e_124c2cd8 , C0 );
buf ( R_5f7_12fbf758 , n42373 );
buf ( R_c16_13df9858 , C0 );
buf ( R_1235_15880cb8 , n42449 );
buf ( R_1854_1580fd78 , n42450 );
buf ( R_18a4_13bf2d98 , n42451 );
buf ( R_1285_100890f8 , n42502 );
buf ( R_c66_13bed2f8 , C0 );
buf ( R_647_13d51af8 , n42503 );
buf ( R_1882_13d1fbf8 , C0 );
buf ( R_1263_123be498 , n42504 );
buf ( R_c44_13c229b8 , n42505 );
buf ( R_625_13c1e638 , n42548 );
buf ( R_619_156b6718 , n42606 );
buf ( R_c38_117efd78 , n42607 );
buf ( R_1257_14a0f0f8 , n42608 );
buf ( R_1876_15ffcb28 , C0 );
buf ( R_985_1587c4d8 , n42688 );
buf ( R_1516_12fc1eb8 , C0 );
buf ( R_15c3_13c02078 , n42689 );
buf ( R_8d8_13d22fd8 , n42690 );
buf ( R_fa4_13d1e898 , n42691 );
buf ( R_ef7_1162bd78 , n42692 );
buf ( R_1663_124c2698 , n42693 );
buf ( R_838_1580b8b8 , n42694 );
buf ( R_a25_13bf4ff8 , n42846 );
buf ( R_1476_1486bd78 , C0 );
buf ( R_1044_13d57818 , n42847 );
buf ( R_e57_13b8f738 , n42848 );
buf ( R_15fa_13c0bb78 , C0 );
buf ( R_ec0_13c1bf78 , n42849 );
buf ( R_fdb_15ff7308 , n42850 );
buf ( R_14df_14a0cdf8 , n42851 );
buf ( R_9bc_15812758 , n42852 );
buf ( R_8a1_13d21818 , n44699 );
buf ( R_1883_13d41058 , n44700 );
buf ( R_1264_13c02758 , n44701 );
buf ( R_c45_13d24c98 , n44724 );
buf ( R_626_123b86d8 , C0 );
buf ( R_618_1587ea58 , n44725 );
buf ( R_c37_13c0bfd8 , n44726 );
buf ( R_1256_13d54258 , C0 );
buf ( R_1875_158179d8 , n44762 );
buf ( R_1145_13b98658 , n45155 );
buf ( R_737_116313b8 , n45156 );
buf ( R_b26_1486a518 , C0 );
buf ( R_d56_117e9d38 , C0 );
buf ( R_1764_13ccf7d8 , n45157 );
buf ( R_1375_13c275f8 , n45223 );
buf ( R_1994_123bac58 , n45224 );
buf ( R_143d_13bf2258 , n45271 );
buf ( R_a5e_1587ed78 , C0 );
buf ( R_e1e_13c1bbb8 , C0 );
buf ( R_107d_15888418 , n45812 );
buf ( R_7ff_13cd45f8 , n45813 );
buf ( R_169c_15885fd8 , n45814 );
buf ( R_1a5c_13de04d8 , n45815 );
buf ( R_1a48_13c1ff38 , n45816 );
buf ( R_a72_1486d358 , C0 );
buf ( R_1429_13d23438 , n45874 );
buf ( R_1091_14a11d58 , n45907 );
buf ( R_e0a_13bfa3b8 , C0 );
buf ( R_16b0_140aae18 , n45908 );
buf ( R_7eb_123b8278 , n45909 );
buf ( R_12c6_13cd49b8 , C0 );
buf ( R_5b6_117f1f38 , C0 );
buf ( R_ca7_140b4418 , n45910 );
buf ( R_bd5_13d51698 , n45967 );
buf ( R_688_13b99af8 , n45968 );
buf ( R_11f4_13d1e6b8 , n45969 );
buf ( R_18e5_13d45658 , n46079 );
buf ( R_1813_13d29c98 , n46080 );
buf ( R_16d9_14a17cf8 , n46353 );
buf ( R_1a1f_11c70958 , n46354 );
buf ( R_1400_14b29b98 , n46355 );
buf ( R_de1_13cd0638 , n47281 );
buf ( R_7c2_15ffa508 , C0 );
buf ( R_a9b_100865d8 , n47282 );
buf ( R_10ba_15881938 , C0 );
buf ( R_1805_14b271b8 , n47413 );
buf ( R_5a8_123b8318 , n47420 );
buf ( R_cb5_170107e8 , n47512 );
buf ( R_bc7_13c2a758 , n47513 );
buf ( R_696_10082ed8 , C0 );
buf ( R_18f3_15ffc628 , n47514 );
buf ( R_11e6_14b222f8 , C0 );
buf ( R_12d4_11634d38 , n47515 );
buf ( R_119f_156b4738 , n47516 );
buf ( R_561_1162a658 , n47518 );
buf ( R_6dd_117f36f8 , n47561 );
buf ( R_131b_15ff76c8 , n47562 );
buf ( R_17be_15816538 , C0 );
buf ( R_b80_13cd8338 , n47563 );
buf ( R_cfc_1700d2c8 , n47564 );
buf ( R_193a_15885718 , C0 );
buf ( R_5da_13df70f8 , C0 );
buf ( R_18c1_11c6f738 , n47773 );
buf ( R_bf9_13d28ed8 , n47824 );
buf ( R_12a2_13bf2578 , C0 );
buf ( R_1218_13d28078 , n47825 );
buf ( R_c83_13d59f78 , n47826 );
buf ( R_1837_13deb9d8 , n47827 );
buf ( R_664_123b47b8 , n47828 );
buf ( R_e39_156b3518 , n47896 );
buf ( R_a43_14b1feb8 , n47897 );
buf ( R_81a_13cceb58 , C0 );
buf ( R_1062_117eedd8 , C0 );
buf ( R_1458_13df07f8 , n47898 );
buf ( R_1681_140b99b8 , n48140 );
buf ( R_1327_124c2b98 , n48141 );
buf ( R_6e9_156b3158 , n48205 );
buf ( R_555_13d59b18 , n48206 );
buf ( R_1193_13b97438 , n48207 );
buf ( R_1946_14a16858 , C0 );
buf ( R_d08_13d59938 , n48208 );
buf ( R_b74_123c0478 , n48209 );
buf ( R_17b2_13cd6498 , C0 );
buf ( R_113a_117eb458 , C0 );
buf ( R_742_14a129d8 , C0 );
buf ( R_b1b_11629758 , n48210 );
buf ( R_d61_11633618 , n48261 );
buf ( R_1380_15887338 , n48262 );
buf ( R_1759_14874518 , n48343 );
buf ( R_199f_13d3c9b8 , n48344 );
buf ( R_1884_13cd1c18 , n48345 );
buf ( R_1265_156b0818 , n48399 );
buf ( R_c46_1580b598 , C0 );
buf ( R_627_117efb98 , n48400 );
buf ( R_617_158807b8 , n48401 );
buf ( R_c36_156b63f8 , C0 );
buf ( R_1255_1580dbb8 , n48453 );
buf ( R_1874_13df9c18 , n48454 );
buf ( R_87a_13c286d8 , C0 );
buf ( R_1002_14a17938 , C0 );
buf ( R_e99_123ba258 , n48528 );
buf ( R_9e3_170110a8 , n48529 );
buf ( R_1621_117eacd8 , n48537 );
buf ( R_14b8_123b31d8 , n48538 );
buf ( R_edf_117f5bd8 , n48539 );
buf ( R_14fe_13d55518 , C0 );
buf ( R_15db_117f7258 , n48540 );
buf ( R_fbc_13beb9f8 , n48541 );
buf ( R_8c0_11631ef8 , n48542 );
buf ( R_99d_13cd4d78 , n48581 );
buf ( R_845_15888918 , n49290 );
buf ( R_1656_117f4af8 , C0 );
buf ( R_1483_13d53d58 , n49291 );
buf ( R_a18_12fbdef8 , n49292 );
buf ( R_e64_14875058 , n49293 );
buf ( R_1037_15815098 , n49294 );
buf ( R_d8e_11630878 , C0 );
buf ( R_172c_13d39d58 , n49295 );
buf ( R_13ad_14a12618 , n49357 );
buf ( R_19cc_13cda1d8 , n49358 );
buf ( R_110d_13dd5cb8 , n49423 );
buf ( R_aee_117e9478 , C0 );
buf ( R_76f_117f4378 , n49424 );
buf ( R_ccd_13b8c8f8 , n49486 );
buf ( R_590_13dd64d8 , n49487 );
buf ( R_17ed_156b36f8 , n49502 );
buf ( R_190b_14872038 , n49503 );
buf ( R_6ae_156ab958 , C0 );
buf ( R_baf_1700cd28 , n49504 );
buf ( R_12ec_124c3778 , n49505 );
buf ( R_11ce_11c6cad8 , C0 );
buf ( R_17a3_150e7398 , n49506 );
buf ( R_1336_148754b8 , C0 );
buf ( R_6f8_13c1c018 , n49507 );
buf ( R_1184_150e6498 , n49508 );
buf ( R_1955_14b235b8 , n49741 );
buf ( R_d17_14b27398 , n49742 );
buf ( R_b65_13dde318 , n49798 );
buf ( R_1885_1486cdb8 , n49830 );
buf ( R_1266_14a12438 , C0 );
buf ( R_c47_100803b8 , n49831 );
buf ( R_628_117eb098 , n49832 );
buf ( R_616_170152e8 , C0 );
buf ( R_c35_123b88b8 , n49882 );
buf ( R_1254_150e59f8 , n49883 );
buf ( R_1873_12fc2278 , n49884 );
buf ( R_74a_1008cb18 , C0 );
buf ( R_1132_15880e98 , C0 );
buf ( R_d69_14b23158 , n49942 );
buf ( R_b13_140b3d38 , n49943 );
buf ( R_1388_140aaf58 , n49944 );
buf ( R_19a7_140b9b98 , n49945 );
buf ( R_1751_1007feb8 , n49984 );
buf ( R_b57_13ccd6b8 , n49985 );
buf ( R_1344_117f3018 , n49986 );
buf ( R_1795_1008b678 , n50105 );
buf ( R_706_1580bd18 , C0 );
buf ( R_1963_13d1f478 , n50106 );
buf ( R_1176_17015b08 , C0 );
buf ( R_d25_15882298 , n50168 );
buf ( R_1590_150e4b98 , n50169 );
buf ( R_f71_124c4998 , n50273 );
buf ( R_952_14b26e98 , C0 );
buf ( R_90b_13d41af8 , n50274 );
buf ( R_f2a_1162a158 , C0 );
buf ( R_1549_1587ff98 , n50349 );
buf ( R_5c6_15816218 , C0 );
buf ( R_12b6_1587db58 , C0 );
buf ( R_be5_140b5818 , n50400 );
buf ( R_c97_156b09f8 , n50401 );
buf ( R_1204_13c23b38 , n50402 );
buf ( R_678_15884ef8 , n50403 );
buf ( R_1823_13d53df8 , n50404 );
buf ( R_18d5_11636098 , n50491 );
buf ( R_ed8_117e9c98 , n50492 );
buf ( R_15e2_14a140f8 , C0 );
buf ( R_14f7_13b965d8 , n50493 );
buf ( R_fc3_14b27e38 , n50494 );
buf ( R_8b9_14875e18 , n50535 );
buf ( R_9a4_117ee018 , n50536 );
buf ( R_1a04_13c22b98 , n50537 );
buf ( R_13e5_13de07f8 , n50584 );
buf ( R_16f4_123b9fd8 , n50585 );
buf ( R_dc6_14873f78 , C0 );
buf ( R_10d5_13b94a58 , n50619 );
buf ( R_7a7_116355f8 , n50620 );
buf ( R_ab6_15814e18 , C0 );
buf ( R_1886_11638c58 , C0 );
buf ( R_1267_14b23f18 , n50621 );
buf ( R_c48_13bf5e58 , n50622 );
buf ( R_629_150e7e38 , n50665 );
buf ( R_615_13c1d7d8 , n50723 );
buf ( R_c34_15ff1228 , n50724 );
buf ( R_1253_13d222b8 , n50725 );
buf ( R_1872_13ccb4f8 , C0 );
buf ( R_16f6_116389d8 , C0 );
buf ( R_10d7_156b5778 , n50726 );
buf ( R_ab8_156ac8f8 , n50727 );
buf ( R_1a02_13cd8298 , C0 );
buf ( R_13e3_14a0a7d8 , n50728 );
buf ( R_7a5_13d456f8 , n50775 );
buf ( R_dc4_11634b58 , n50776 );
buf ( R_b4d_1700f208 , n50811 );
buf ( R_710_156ac718 , n50812 );
buf ( R_178b_1580ca38 , n50813 );
buf ( R_196d_117eb8b8 , n50845 );
buf ( R_d2f_13dedf58 , n50846 );
buf ( R_116c_140b8338 , n50847 );
buf ( R_134e_13d282f8 , C0 );
buf ( R_1a06_1486e1b8 , C0 );
buf ( R_13e7_116377b8 , n50848 );
buf ( R_dc8_1162b058 , n50849 );
buf ( R_7a9_123bd458 , n50892 );
buf ( R_16f2_158857b8 , C0 );
buf ( R_ab4_12fbed58 , n50893 );
buf ( R_10d3_158899f8 , n50894 );
buf ( R_85a_156b1a38 , C0 );
buf ( R_1498_15811c18 , n50895 );
buf ( R_1641_150db8b8 , n51622 );
buf ( R_a03_123bd818 , n51623 );
buf ( R_e79_13cd8658 , n51672 );
buf ( R_1022_11c6cf38 , C0 );
buf ( R_150d_14b21678 , n51721 );
buf ( R_15cc_14a0ba98 , n51722 );
buf ( R_8cf_13ded9b8 , n51723 );
buf ( R_fad_140ac038 , n51751 );
buf ( R_eee_11632e98 , C0 );
buf ( R_98e_12fbecb8 , C0 );
buf ( R_13bd_13df6c98 , n51794 );
buf ( R_19dc_156b6858 , n51795 );
buf ( R_171c_117ecb78 , n51796 );
buf ( R_10fd_117eef18 , n51830 );
buf ( R_ade_13dd7658 , C0 );
buf ( R_77f_117f4558 , n51831 );
buf ( R_d9e_13ddc3d8 , C0 );
buf ( R_16f8_14a0e018 , n51832 );
buf ( R_10d9_123b9538 , n51866 );
buf ( R_aba_13c29678 , C0 );
buf ( R_7a3_13ccb138 , n51867 );
buf ( R_dc2_158108b8 , C0 );
buf ( R_13e1_156b8478 , n51910 );
buf ( R_1a00_123b7f58 , n51911 );
buf ( R_971_13df5618 , n51939 );
buf ( R_8ec_123bbd38 , n51940 );
buf ( R_15af_14866eb8 , n51941 );
buf ( R_f0b_13cd72f8 , n51942 );
buf ( R_f90_15812438 , n51943 );
buf ( R_152a_13df8818 , C0 );
buf ( R_c15_15fee528 , n51993 );
buf ( R_1234_15ff9e28 , n51994 );
buf ( R_1853_13dd8738 , n51995 );
buf ( R_18a5_170177c8 , n52027 );
buf ( R_1286_124c4858 , C0 );
buf ( R_c67_13ccba98 , n52028 );
buf ( R_648_15814058 , n52029 );
buf ( R_5f6_13cce018 , C0 );
buf ( R_c05_14866d78 , n52080 );
buf ( R_18b5_10087cf8 , n52112 );
buf ( R_1224_13ccff58 , n52113 );
buf ( R_1296_13dda7b8 , C0 );
buf ( R_1843_1580a878 , n52114 );
buf ( R_c77_13d523b8 , n52115 );
buf ( R_658_140ae1f8 , n52116 );
buf ( R_5e6_13d46698 , C0 );
buf ( R_1a08_14b1b958 , n52117 );
buf ( R_13e9_13d22358 , n52164 );
buf ( R_dca_14b297d8 , C0 );
buf ( R_7ab_15887ab8 , n52165 );
buf ( R_ab2_13df75f8 , C0 );
buf ( R_10d1_13d55d38 , n52199 );
buf ( R_16f0_14b1e978 , n52200 );
buf ( R_d87_123bae38 , n52201 );
buf ( R_1733_15ff79e8 , n52202 );
buf ( R_13a6_156b1718 , C0 );
buf ( R_1114_13d46ff8 , n52203 );
buf ( R_19c5_13bf6ad8 , n52215 );
buf ( R_af5_13c1b6b8 , n52294 );
buf ( R_768_158896d8 , n52295 );
buf ( R_964_123c1f58 , n52296 );
buf ( R_8f9_117ee658 , n52377 );
buf ( R_f18_14a19d78 , n52378 );
buf ( R_1537_117e9b58 , n52379 );
buf ( R_15a2_13ccce98 , C0 );
buf ( R_f83_14a0e978 , n52380 );
buf ( R_1887_17018da8 , n52381 );
buf ( R_1268_13d38278 , n52382 );
buf ( R_c49_123b36d8 , n52630 );
buf ( R_62a_13d42278 , C0 );
buf ( R_614_13c2a258 , n52631 );
buf ( R_c33_150e7bb8 , n52632 );
buf ( R_1252_116378f8 , C0 );
buf ( R_1871_13defad8 , n52667 );
buf ( R_11a3_13c1be38 , n52668 );
buf ( R_565_13ddbb18 , n52670 );
buf ( R_6d9_11636818 , n52713 );
buf ( R_1317_1580c5d8 , n52714 );
buf ( R_17c2_13c03518 , C0 );
buf ( R_b84_156b5278 , n52715 );
buf ( R_cf8_15881a78 , n52716 );
buf ( R_1936_13d2a558 , C0 );
buf ( R_13b4_156abb38 , n52717 );
buf ( R_19d3_13bf92d8 , n52718 );
buf ( R_1725_13cd9a58 , n52730 );
buf ( R_1106_14b1c718 , C0 );
buf ( R_ae7_13cd22f8 , n52731 );
buf ( R_776_14873bb8 , C0 );
buf ( R_d95_15815778 , n52778 );
buf ( R_feb_1486c818 , n52779 );
buf ( R_eb0_13d53498 , n52780 );
buf ( R_14cf_14b1bd18 , n52781 );
buf ( R_9cc_158172f8 , n52782 );
buf ( R_160a_17010ce8 , C0 );
buf ( R_891_13b8ab98 , n52799 );
buf ( R_132b_1007f7d8 , n52800 );
buf ( R_6ed_140b6538 , n52864 );
buf ( R_118f_14b1ee78 , n52865 );
buf ( R_194a_13d2ae18 , C0 );
buf ( R_d0c_13dee8b8 , n52866 );
buf ( R_b70_13d20f58 , n52867 );
buf ( R_17ae_13d29a18 , C0 );
buf ( R_1a3c_13b95278 , n52868 );
buf ( R_109d_10084878 , n52900 );
buf ( R_141d_13d441b8 , n52947 );
buf ( R_16bc_14a0bdb8 , n52948 );
buf ( R_dfe_15ff38e8 , C0 );
buf ( R_7df_1587d338 , n52949 );
buf ( R_a7e_14a0bb38 , C0 );
buf ( R_151f_12fbe998 , n52950 );
buf ( R_97c_13d528b8 , n52951 );
buf ( R_15ba_1008b0d8 , C0 );
buf ( R_8e1_15889818 , n52968 );
buf ( R_f00_17017ae8 , n52969 );
buf ( R_f9b_13b974d8 , n52970 );
buf ( R_16fa_14b299b8 , C0 );
buf ( R_10db_13cd6cb8 , n52971 );
buf ( R_abc_15882b58 , n52972 );
buf ( R_7a1_15ffcd08 , n53015 );
buf ( R_dc0_117f53b8 , n53016 );
buf ( R_13df_156b9238 , n53017 );
buf ( R_19fe_13c01fd8 , C0 );
buf ( R_5cf_124c4678 , n53018 );
buf ( R_12ad_13cca878 , n53068 );
buf ( R_bee_156ac498 , C0 );
buf ( R_c8e_156b6cb8 , C0 );
buf ( R_120d_123be218 , n53093 );
buf ( R_66f_13df8d18 , n53094 );
buf ( R_182c_13b90598 , n53095 );
buf ( R_18cc_170190c8 , n53096 );
buf ( R_1505_13d27858 , n53145 );
buf ( R_15d4_13d3a078 , n53146 );
buf ( R_fb5_13c265b8 , n53174 );
buf ( R_8c7_13ccf738 , n53175 );
buf ( R_996_13cd1498 , C0 );
buf ( R_ee6_156ae158 , C0 );
buf ( R_1a0a_140b9238 , C0 );
buf ( R_13eb_150e7438 , n53176 );
buf ( R_dcc_15815c78 , n53177 );
buf ( R_7ad_1008c078 , n53220 );
buf ( R_ab0_11629618 , n53221 );
buf ( R_10cf_1580df78 , n53222 );
buf ( R_16ee_123bf758 , C0 );
buf ( R_1660_13dd6258 , n53223 );
buf ( R_83b_117f03b8 , n53224 );
buf ( R_a22_156b92d8 , C0 );
buf ( R_1479_13ddc518 , n53286 );
buf ( R_1041_14a0db18 , n53315 );
buf ( R_e5a_11633118 , C0 );
buf ( R_1711_11c69d38 , n53349 );
buf ( R_10f2_1486ad38 , C0 );
buf ( R_ad3_13d5a5b8 , n53350 );
buf ( R_78a_13dfa2f8 , C0 );
buf ( R_da9_123bc9b8 , n53397 );
buf ( R_13c8_11628e98 , n53398 );
buf ( R_19e7_14a10098 , n53399 );
buf ( R_eb5_13cd9cd8 , n53455 );
buf ( R_fe6_13df1d38 , C0 );
buf ( R_14d4_13c27a58 , n53456 );
buf ( R_9c7_140af5f8 , n53457 );
buf ( R_896_123b6658 , C0 );
buf ( R_1605_156b1b78 , n53573 );
buf ( R_1888_1580c858 , n53574 );
buf ( R_1269_13b99c38 , n53625 );
buf ( R_c4a_14a0cb78 , C0 );
buf ( R_62b_1162a1f8 , n53626 );
buf ( R_613_124c47b8 , n53627 );
buf ( R_c32_14b23518 , C0 );
buf ( R_1251_13d3fed8 , n53670 );
buf ( R_1870_13b92bb8 , n53671 );
buf ( R_16cc_156ba318 , n53672 );
buf ( R_1a2c_156b08b8 , n53673 );
buf ( R_140d_11638258 , n53716 );
buf ( R_dee_13c0e058 , C0 );
buf ( R_7cf_123bbe78 , n53717 );
buf ( R_a8e_170160a8 , C0 );
buf ( R_10ad_10082618 , n53868 );
buf ( R_11b0_13b99f58 , n53869 );
buf ( R_572_140ab458 , n53871 );
buf ( R_6cc_117e8a78 , n53872 );
buf ( R_130a_13dda498 , C0 );
buf ( R_17cf_13d389f8 , n53873 );
buf ( R_b91_14b1f418 , n53916 );
buf ( R_ceb_13d56d78 , n53917 );
buf ( R_1929_13cd4af8 , n53968 );
buf ( R_f72_13c2a1b8 , C0 );
buf ( R_953_14b20a98 , n53969 );
buf ( R_90a_156ae658 , C0 );
buf ( R_f29_11630698 , n53985 );
buf ( R_1548_140ac538 , n53986 );
buf ( R_1591_13c25618 , n53992 );
buf ( R_16fc_156b9a58 , n53993 );
buf ( R_10dd_13d551f8 , n54027 );
buf ( R_abe_14a15958 , C0 );
buf ( R_79f_140af7d8 , n54028 );
buf ( R_dbe_13cd4c38 , C0 );
buf ( R_13dd_15884b38 , n54071 );
buf ( R_19fc_13b96fd8 , n54072 );
buf ( R_ff0_123b3b38 , n54073 );
buf ( R_eab_11634518 , n54074 );
buf ( R_9d1_13d4ed58 , n54599 );
buf ( R_14ca_11631e58 , C0 );
buf ( R_160f_170102e8 , n54600 );
buf ( R_88c_116319f8 , n54601 );
buf ( R_e36_13c05b38 , C0 );
buf ( R_a46_11637e98 , C0 );
buf ( R_817_116294d8 , n54602 );
buf ( R_1065_13c0b218 , n54626 );
buf ( R_1455_117ef238 , n54673 );
buf ( R_1684_13dd5ad8 , n54674 );
buf ( R_e2b_13d28578 , n54675 );
buf ( R_a51_11630ff8 , n54720 );
buf ( R_80c_13d2acd8 , n54721 );
buf ( R_1070_150e2d98 , n54722 );
buf ( R_1a69_11c6fe18 , n54745 );
buf ( R_168f_13d295b8 , n54746 );
buf ( R_144a_1580c678 , C0 );
buf ( R_1a0c_13ccacd8 , n54747 );
buf ( R_13ed_13cd4ff8 , n54790 );
buf ( R_dce_14871f98 , C0 );
buf ( R_7af_11633578 , n54791 );
buf ( R_aae_15814238 , C0 );
buf ( R_10cd_13d20878 , n54870 );
buf ( R_16ec_13df6a18 , n54871 );
buf ( R_1889_13bf9c38 , n54903 );
buf ( R_126a_15886a78 , C0 );
buf ( R_c4b_13cd76b8 , n54904 );
buf ( R_62c_10086038 , n54905 );
buf ( R_612_10088dd8 , C0 );
buf ( R_c31_13b90778 , n54955 );
buf ( R_1250_13d58c18 , n54956 );
buf ( R_186f_1162dcb8 , n54957 );
buf ( R_1a21_150e5598 , n54964 );
buf ( R_1402_140b1cb8 , C0 );
buf ( R_de3_140b0778 , n54965 );
buf ( R_7c4_13cd5138 , n54966 );
buf ( R_a99_13cd0a98 , n55257 );
buf ( R_10b8_13bea7d8 , n55258 );
buf ( R_16d7_15888a58 , n55259 );
buf ( R_b23_1587bc18 , n55260 );
buf ( R_d59_14868cb8 , n55307 );
buf ( R_1378_14b28158 , n55308 );
buf ( R_1761_11631f98 , n55342 );
buf ( R_1997_13d45158 , n55343 );
buf ( R_1142_117f06d8 , C0 );
buf ( R_73a_13de1158 , C0 );
buf ( R_1a35_1486d7b8 , n55350 );
buf ( R_16c3_13c01498 , n55351 );
buf ( R_1416_1162ee38 , C0 );
buf ( R_df7_117f35b8 , n55352 );
buf ( R_7d8_156abc78 , n55353 );
buf ( R_a85_17014168 , n55399 );
buf ( R_10a4_1486b0f8 , n55400 );
buf ( R_a59_14a1a1d8 , n55434 );
buf ( R_e23_13df5f78 , n55435 );
buf ( R_1078_1580f558 , n55436 );
buf ( R_804_156b6f38 , n55437 );
buf ( R_1697_13d59d98 , n55438 );
buf ( R_1a61_14a195f8 , n55445 );
buf ( R_1442_14a18c98 , C0 );
buf ( R_1096_13dd6f78 , C0 );
buf ( R_1424_13b906d8 , n55446 );
buf ( R_16b5_13c045f8 , n55470 );
buf ( R_e05_140ad938 , n55517 );
buf ( R_7e6_1486dd58 , C0 );
buf ( R_a77_100895f8 , n55518 );
buf ( R_1a43_170104c8 , n55519 );
buf ( R_15ef_15889318 , n55520 );
buf ( R_ecb_13df7198 , n55521 );
buf ( R_14ea_13cd2078 , C0 );
buf ( R_fd0_13cd59f8 , n55522 );
buf ( R_8ac_15889278 , n55523 );
buf ( R_9b1_1008a3b8 , n55542 );
buf ( R_cc2_14a11218 , C0 );
buf ( R_17f8_13c28d18 , n55543 );
buf ( R_59b_15812bb8 , n55550 );
buf ( R_1900_1486c318 , n55551 );
buf ( R_6a3_11c69658 , n55552 );
buf ( R_bba_13deb7f8 , C0 );
buf ( R_12e1_123bbf18 , n55804 );
buf ( R_11d9_14a18518 , n55839 );
buf ( R_1125_124c3e58 , n55885 );
buf ( R_d76_156b6218 , C0 );
buf ( R_b06_14b24af8 , C0 );
buf ( R_1395_13c0d978 , n55932 );
buf ( R_19b4_14a10598 , n55933 );
buf ( R_1744_11c6e3d8 , n55934 );
buf ( R_757_13d3ceb8 , n55935 );
buf ( R_16fe_123b51b8 , C0 );
buf ( R_10df_156b31f8 , n55936 );
buf ( R_ac0_123c19b8 , n55937 );
buf ( R_79d_13ddd698 , n55980 );
buf ( R_dbc_13d207d8 , n55981 );
buf ( R_13db_13d412d8 , n55982 );
buf ( R_19fa_140afeb8 , C0 );
buf ( R_188a_14a0dd98 , C0 );
buf ( R_126b_170193e8 , n55983 );
buf ( R_c4c_14874a18 , n55984 );
buf ( R_62d_123c23b8 , n56027 );
buf ( R_611_156aa558 , n56085 );
buf ( R_c30_13cd8158 , n56086 );
buf ( R_124f_13cd9418 , n56087 );
buf ( R_186e_1162cb38 , C0 );
buf ( R_1233_13d5c318 , n56088 );
buf ( R_1852_11635698 , C0 );
buf ( R_18a6_15885218 , C0 );
buf ( R_1287_13c29e98 , n56089 );
buf ( R_c68_12fc1cd8 , n56090 );
buf ( R_649_150e1f38 , n56137 );
buf ( R_5f5_13bf7398 , n56184 );
buf ( R_c14_13defe98 , n56185 );
buf ( R_18c2_13d5d998 , C0 );
buf ( R_bf8_13bf77f8 , n56186 );
buf ( R_12a3_14b20278 , n56187 );
buf ( R_1217_123bdd18 , n56188 );
buf ( R_c84_123bee98 , n56189 );
buf ( R_1836_14a16038 , C0 );
buf ( R_665_117eefb8 , n56236 );
buf ( R_5d9_15fed588 , n56283 );
buf ( R_84f_1587bdf8 , n56284 );
buf ( R_148d_156b2d98 , n56331 );
buf ( R_164c_156b65d8 , n56332 );
buf ( R_a0e_13cd5098 , C0 );
buf ( R_e6e_13c1e818 , C0 );
buf ( R_102d_14a14878 , n56357 );
buf ( R_d7b_1007dbb8 , n56358 );
buf ( R_1120_13cd3158 , n56359 );
buf ( R_139a_12fbf398 , C0 );
buf ( R_b01_1587af98 , n56393 );
buf ( R_19b9_116327b8 , n56405 );
buf ( R_75c_13d54b18 , n56406 );
buf ( R_173f_14a0d1b8 , n56407 );
buf ( R_ca0_117f3978 , n56408 );
buf ( R_bdc_14867a98 , n56409 );
buf ( R_11fb_13d26638 , n56410 );
buf ( R_681_13c02c58 , n56457 );
buf ( R_18de_1162c638 , C0 );
buf ( R_181a_15887fb8 , C0 );
buf ( R_12bf_12fbe3f8 , n56458 );
buf ( R_5bd_123b9678 , n56703 );
buf ( R_1a0e_1486b698 , C0 );
buf ( R_13ef_156ba1d8 , n56704 );
buf ( R_dd0_12fc0798 , n56705 );
buf ( R_7b1_14a13478 , n56752 );
buf ( R_aac_116311d8 , n56753 );
buf ( R_10cb_150dccb8 , n56754 );
buf ( R_16ea_140b6cb8 , C0 );
buf ( R_ffe_13ccf198 , C0 );
buf ( R_e9d_13d27038 , n56810 );
buf ( R_9df_14a17398 , n56811 );
buf ( R_161d_13b962b8 , n56823 );
buf ( R_14bc_117f0598 , n56824 );
buf ( R_87e_140b08b8 , C0 );
buf ( R_5a1_13d446b8 , n56831 );
buf ( R_cbc_12fc1b98 , n56832 );
buf ( R_bc0_13dfb338 , n56833 );
buf ( R_69d_11c69798 , n56880 );
buf ( R_18fa_140b5098 , C0 );
buf ( R_11df_15880998 , n56881 );
buf ( R_12db_156b4af8 , n56882 );
buf ( R_17fe_1580f5f8 , C0 );
buf ( R_191b_13c25f78 , n56883 );
buf ( R_580_1162b4b8 , n56884 );
buf ( R_6be_158101d8 , C0 );
buf ( R_17dd_14872358 , n56899 );
buf ( R_12fc_15813dd8 , n56900 );
buf ( R_b9f_140b49b8 , n56901 );
buf ( R_cdd_13bf42d8 , n56963 );
buf ( R_11be_150e4378 , C0 );
buf ( R_eba_13d29158 , C0 );
buf ( R_fe1_13d2bef8 , n56985 );
buf ( R_14d9_13c21338 , n57032 );
buf ( R_9c2_116297f8 , C0 );
buf ( R_89b_117ed118 , n57033 );
buf ( R_1600_117e96f8 , n57034 );
buf ( R_585_14a19b98 , n57035 );
buf ( R_1916_150e99b8 , C0 );
buf ( R_17e2_123c1d78 , C0 );
buf ( R_6b9_150dc998 , n57082 );
buf ( R_ba4_13c04d78 , n57083 );
buf ( R_12f7_117f4ff8 , n57084 );
buf ( R_11c3_117ee158 , n57085 );
buf ( R_cd8_150deab8 , n57086 );
buf ( R_15c4_13d46e18 , n57087 );
buf ( R_8d7_13de10b8 , n57088 );
buf ( R_fa5_13df4858 , n57116 );
buf ( R_ef6_13c1f358 , C0 );
buf ( R_986_11631278 , C0 );
buf ( R_1515_13ccb8b8 , n57165 );
buf ( R_11a7_123b9b78 , n57166 );
buf ( R_569_12fbfd98 , n57168 );
buf ( R_6d5_14b25958 , n57211 );
buf ( R_1313_1587dab8 , n57212 );
buf ( R_17c6_13d290b8 , C0 );
buf ( R_b88_14a0d9d8 , n57213 );
buf ( R_cf4_13bea558 , n57214 );
buf ( R_1932_13cd1538 , C0 );
buf ( R_1778_11631598 , n57215 );
buf ( R_d42_1580f918 , C0 );
buf ( R_1159_148722b8 , n57230 );
buf ( R_1361_14a18658 , n57277 );
buf ( R_b3a_11637678 , C0 );
buf ( R_1980_15883a58 , n57278 );
buf ( R_723_14a0aeb8 , n57279 );
buf ( R_ec5_123c1eb8 , n57344 );
buf ( R_fd6_15ff7448 , C0 );
buf ( R_14e4_14a121b8 , n57345 );
buf ( R_9b7_117eaaf8 , n57346 );
buf ( R_8a6_156b3018 , C0 );
buf ( R_15f5_140ade38 , n57362 );
buf ( R_d45_117f4418 , n57405 );
buf ( R_1775_140b5d18 , n57439 );
buf ( R_1364_13c1d918 , n57440 );
buf ( R_1156_15ff6fe8 , C0 );
buf ( R_1983_100863f8 , n57441 );
buf ( R_726_13d39498 , C0 );
buf ( R_b37_10089b98 , n57442 );
buf ( R_15e9_11636db8 , n57458 );
buf ( R_14f0_13b92398 , n57459 );
buf ( R_fca_156b44b8 , C0 );
buf ( R_8b2_11629078 , C0 );
buf ( R_9ab_14866698 , n57460 );
buf ( R_ed1_158870b8 , n57543 );
buf ( R_1632_117f1178 , C0 );
buf ( R_9f4_1486d2b8 , n57544 );
buf ( R_e88_124c4498 , n57545 );
buf ( R_1013_14a135b8 , n57546 );
buf ( R_14a7_15814af8 , n57547 );
buf ( R_869_14a19e18 , n57868 );
buf ( R_132f_13c0b8f8 , n57869 );
buf ( R_6f1_150df878 , n57916 );
buf ( R_118b_14b27618 , n57917 );
buf ( R_194e_14b236f8 , C0 );
buf ( R_d10_123b2d78 , n57918 );
buf ( R_b6c_123b8138 , n57919 );
buf ( R_17aa_13dfac58 , C0 );
buf ( R_188b_117e9978 , n57920 );
buf ( R_126c_1580edd8 , n57921 );
buf ( R_c4d_13d24b58 , n57947 );
buf ( R_62e_13bf7438 , C0 );
buf ( R_610_14a186f8 , n57948 );
buf ( R_c2f_14a0c038 , n57949 );
buf ( R_124e_117ee338 , C0 );
buf ( R_186d_15fee348 , n57984 );
buf ( R_e8c_1587e738 , n57985 );
buf ( R_162e_123b25f8 , C0 );
buf ( R_9f0_140abe58 , n57986 );
buf ( R_14ab_13dd50d8 , n57987 );
buf ( R_86d_14a18dd8 , n58011 );
buf ( R_100f_13d5dad8 , n58012 );
buf ( R_8f8_15ff8668 , n58013 );
buf ( R_f17_14a18e78 , n58014 );
buf ( R_1536_14a0dc58 , C0 );
buf ( R_15a3_12fc08d8 , n58015 );
buf ( R_f84_117e8d98 , n58016 );
buf ( R_965_140b2578 , n58044 );
buf ( R_d71_14b23018 , n58102 );
buf ( R_b0b_13c21e78 , n58103 );
buf ( R_1390_17016a08 , n58104 );
buf ( R_19af_11636458 , n58105 );
buf ( R_1749_117ec178 , n58114 );
buf ( R_752_15ff64a8 , C0 );
buf ( R_112a_1587e0f8 , C0 );
buf ( R_18b6_13bf3018 , C0 );
buf ( R_1223_13dd8418 , n58115 );
buf ( R_1297_13b99738 , n58116 );
buf ( R_1842_123b43f8 , C0 );
buf ( R_c78_15887018 , n58117 );
buf ( R_659_123b34f8 , n58160 );
buf ( R_5e5_13df0578 , n58203 );
buf ( R_c04_13cd6f38 , n58204 );
buf ( R_954_17014988 , n58205 );
buf ( R_909_13d3efd8 , n58212 );
buf ( R_f28_13bf6fd8 , n58213 );
buf ( R_1547_13df7b98 , n58214 );
buf ( R_1592_156b9918 , C0 );
buf ( R_f73_13d22a38 , n58215 );
buf ( R_70d_13beb098 , n58258 );
buf ( R_178e_13c1cb58 , C0 );
buf ( R_196a_156b6d58 , C0 );
buf ( R_d2c_14a0ec98 , n58259 );
buf ( R_116f_13d3e7b8 , n58260 );
buf ( R_134b_15ff6cc8 , n58261 );
buf ( R_b50_15815598 , n58262 );
buf ( R_caf_156adc58 , n58263 );
buf ( R_bcd_1162baf8 , n58315 );
buf ( R_690_13c1e098 , n58316 );
buf ( R_18ed_124c3278 , n58371 );
buf ( R_11ec_1008d0b8 , n58372 );
buf ( R_12ce_13c071b8 , C0 );
buf ( R_180b_1008abd8 , n58373 );
buf ( R_5ae_13cd7ed8 , n58379 );
buf ( R_177b_1007d6b8 , n58380 );
buf ( R_d3f_13cd10d8 , n58381 );
buf ( R_115c_150e8f18 , n58382 );
buf ( R_135e_11c696f8 , C0 );
buf ( R_b3d_13dddeb8 , n58609 );
buf ( R_720_13d395d8 , n58610 );
buf ( R_197d_14a15458 , n58622 );
buf ( R_1700_140ae8d8 , n58623 );
buf ( R_10e1_13c07758 , n58657 );
buf ( R_ac2_156ad2f8 , C0 );
buf ( R_79b_15886398 , n58658 );
buf ( R_dba_116373f8 , C0 );
buf ( R_13d9_14a14378 , n58701 );
buf ( R_19f8_117ef558 , n58702 );
buf ( R_595_13def178 , n58709 );
buf ( R_17f2_1580c998 , C0 );
buf ( R_1906_13ccad78 , C0 );
buf ( R_6a9_15ff4ba8 , n58752 );
buf ( R_bb4_117f4d78 , n58753 );
buf ( R_12e7_13cd42d8 , n58754 );
buf ( R_11d3_1162b0f8 , n58755 );
buf ( R_cc8_123b7738 , n58756 );
buf ( R_d48_13c21c98 , n58757 );
buf ( R_1772_14a16998 , C0 );
buf ( R_1367_15880858 , n58758 );
buf ( R_1153_117f1678 , n58759 );
buf ( R_1986_11c6c038 , C0 );
buf ( R_729_117f72f8 , n58806 );
buf ( R_b34_158825b8 , n58807 );
buf ( R_ff5_13c2a618 , n58835 );
buf ( R_ea6_150dd7f8 , C0 );
buf ( R_9d6_13c01f38 , C0 );
buf ( R_14c5_14a0e518 , n58878 );
buf ( R_1614_156b2b18 , n58879 );
buf ( R_887_14a18298 , n58880 );
buf ( R_848_13ddf218 , n58881 );
buf ( R_1653_14869438 , n58882 );
buf ( R_1486_156afe18 , C0 );
buf ( R_a15_1700ed08 , n58914 );
buf ( R_e67_117f4e18 , n58915 );
buf ( R_1034_156ac5d8 , n58916 );
buf ( R_8eb_150db1d8 , n58917 );
buf ( R_15b0_1580bdb8 , n58918 );
buf ( R_f0a_14a0ce98 , C0 );
buf ( R_f91_117f6f38 , n58931 );
buf ( R_1529_123bca58 , n58987 );
buf ( R_972_13ccc038 , C0 );
buf ( R_1a10_123b4718 , n58988 );
buf ( R_13f1_13d24298 , n59046 );
buf ( R_dd2_14a19198 , C0 );
buf ( R_7b3_13c07938 , n59047 );
buf ( R_aaa_13b8cfd8 , C0 );
buf ( R_10c9_15812a78 , n59097 );
buf ( R_16e8_13cd8d38 , n59098 );
buf ( R_d64_15ff5968 , n59099 );
buf ( R_b18_117f40f8 , n59100 );
buf ( R_1383_13c2a438 , n59101 );
buf ( R_19a2_117f01d8 , C0 );
buf ( R_1756_123c0f18 , C0 );
buf ( R_1137_13d20ff8 , n59102 );
buf ( R_745_13c1d5f8 , n59149 );
buf ( R_1636_14b22618 , C0 );
buf ( R_9f8_13decdd8 , n59150 );
buf ( R_e84_14875b98 , n59151 );
buf ( R_1017_13d3bbf8 , n59152 );
buf ( R_865_13d4e7b8 , n59157 );
buf ( R_14a3_11c6d078 , n59158 );
buf ( R_83e_13d43ad8 , C0 );
buf ( R_a1f_13d22d58 , n59159 );
buf ( R_147c_1580d398 , n59160 );
buf ( R_103e_13d57958 , C0 );
buf ( R_e5d_1486ddf8 , n59204 );
buf ( R_165d_13bec038 , n59250 );
buf ( R_1494_117f6718 , n59251 );
buf ( R_1645_11c6c178 , n59279 );
buf ( R_a07_14b251d8 , n59280 );
buf ( R_e75_1580a5f8 , n59339 );
buf ( R_1026_158103b8 , C0 );
buf ( R_856_13cd2a78 , C0 );
buf ( R_188c_13d39ad8 , n59340 );
buf ( R_126d_11636638 , n59391 );
buf ( R_c4e_13c0fe58 , C0 );
buf ( R_62f_116305f8 , n59392 );
buf ( R_60f_13bf44b8 , n59393 );
buf ( R_c2e_156b6c18 , C0 );
buf ( R_124d_123b5438 , n59449 );
buf ( R_186c_15817758 , n59450 );
buf ( R_57b_12fc1f58 , n59451 );
buf ( R_6c3_14a11718 , n59452 );
buf ( R_17d8_13bf24d8 , n59453 );
buf ( R_1301_13ccee78 , n59496 );
buf ( R_b9a_140b40f8 , C0 );
buf ( R_ce2_156b49b8 , C0 );
buf ( R_11b9_13d5d5d8 , n59513 );
buf ( R_1920_117ea198 , n59514 );
buf ( R_1713_14a0f878 , n59515 );
buf ( R_10f4_13de4c18 , n59516 );
buf ( R_ad5_117ed1b8 , n59531 );
buf ( R_788_117e8ed8 , n59532 );
buf ( R_da7_11635ff8 , n59533 );
buf ( R_13c6_123c10f8 , C0 );
buf ( R_19e5_1580eb58 , n59540 );
buf ( R_e90_11637038 , n59541 );
buf ( R_9ec_117eb958 , n59542 );
buf ( R_162a_117ec0d8 , C0 );
buf ( R_14af_156abdb8 , n59543 );
buf ( R_871_1587f138 , n59567 );
buf ( R_100b_11631d18 , n59568 );
buf ( R_111b_1580faf8 , n59569 );
buf ( R_139f_150df058 , n59570 );
buf ( R_afc_117f8158 , n59571 );
buf ( R_19be_13ccfff8 , C0 );
buf ( R_761_12fbf078 , n59618 );
buf ( R_173a_156b5a98 , C0 );
buf ( R_d80_13c1d418 , n59619 );
buf ( R_58a_13ddaf38 , n59620 );
buf ( R_1911_124c4038 , n59671 );
buf ( R_17e7_15883198 , n59672 );
buf ( R_6b4_15881bb8 , n59673 );
buf ( R_ba9_13d5c958 , n59711 );
buf ( R_12f2_17013c68 , C0 );
buf ( R_11c8_11634fb8 , n59712 );
buf ( R_cd3_13c06178 , n59713 );
buf ( R_6fc_13de34f8 , n59714 );
buf ( R_1180_13ddc298 , n59715 );
buf ( R_1959_14a14698 , n59768 );
buf ( R_d1b_13cd9558 , n59769 );
buf ( R_b61_13d22538 , n59804 );
buf ( R_179f_150e5818 , n59805 );
buf ( R_133a_13d57138 , C0 );
buf ( R_be4_15817bb8 , n59806 );
buf ( R_c98_13dec298 , n59807 );
buf ( R_1203_1587d978 , n59808 );
buf ( R_679_123b7918 , n59851 );
buf ( R_1822_117e9018 , C0 );
buf ( R_18d6_13c2ad98 , C0 );
buf ( R_5c5_1162b5f8 , n59878 );
buf ( R_12b7_117f83d8 , n59879 );
buf ( R_ca8_14a11038 , n59880 );
buf ( R_bd4_11637ad8 , n59881 );
buf ( R_689_158869d8 , n59924 );
buf ( R_11f3_116300f8 , n59925 );
buf ( R_18e6_156b1678 , C0 );
buf ( R_1812_11c6f558 , C0 );
buf ( R_12c7_13b97c58 , n59926 );
buf ( R_5b5_11637fd8 , n59927 );
buf ( R_177e_14b1a738 , C0 );
buf ( R_d3c_13b8b278 , n59928 );
buf ( R_115f_156ac7b8 , n59929 );
buf ( R_135b_13d38b38 , n59930 );
buf ( R_b40_158142d8 , n59931 );
buf ( R_71d_13c1ea98 , n59974 );
buf ( R_197a_13c0a318 , C0 );
buf ( R_e16_17018088 , C0 );
buf ( R_1085_13c03e78 , n59998 );
buf ( R_7f7_15888b98 , n59999 );
buf ( R_16a4_158821f8 , n60000 );
buf ( R_1a54_13de0438 , n60001 );
buf ( R_1435_10082258 , n60044 );
buf ( R_a66_15882838 , C0 );
buf ( R_703_14867bd8 , n60045 );
buf ( R_1960_1162c958 , n60046 );
buf ( R_1179_13d3c7d8 , n60077 );
buf ( R_d22_13d599d8 , C0 );
buf ( R_b5a_13bf68f8 , C0 );
buf ( R_1341_13d458d8 , n60120 );
buf ( R_1798_1700e9e8 , n60121 );
buf ( R_171e_13df60b8 , C0 );
buf ( R_10ff_13ddcab8 , n60122 );
buf ( R_ae0_14a11f38 , n60123 );
buf ( R_77d_13d27df8 , n60170 );
buf ( R_d9c_13ccd4d8 , n60171 );
buf ( R_13bb_1587d478 , n60172 );
buf ( R_19da_13dd5a38 , C0 );
buf ( R_108a_1486e938 , C0 );
buf ( R_e11_13cd8c98 , n60215 );
buf ( R_16a9_14a130b8 , n60239 );
buf ( R_7f2_156b2938 , C0 );
buf ( R_1a4f_13d3a618 , n60240 );
buf ( R_a6b_13b8e1f8 , n60241 );
buf ( R_1430_13dd84b8 , n60242 );
buf ( R_d4b_117f6178 , n60243 );
buf ( R_176f_13d447f8 , n60244 );
buf ( R_136a_13c26838 , C0 );
buf ( R_1150_15ff71c8 , n60245 );
buf ( R_1989_13ccbc78 , n60257 );
buf ( R_72c_10083c98 , n60258 );
buf ( R_b31_13d44c58 , n60273 );
buf ( R_814_13d51eb8 , n60274 );
buf ( R_1068_1580ea18 , n60275 );
buf ( R_1687_123b81d8 , n60276 );
buf ( R_1452_13df0938 , C0 );
buf ( R_e33_14a0c3f8 , n60277 );
buf ( R_a49_14a0eb58 , n60305 );
buf ( R_1851_13d5b058 , n60559 );
buf ( R_18a7_13b96858 , n60560 );
buf ( R_1288_13c1daf8 , n60561 );
buf ( R_c69_156af738 , n60608 );
buf ( R_64a_11629438 , C0 );
buf ( R_5f4_140b13f8 , n60609 );
buf ( R_c13_1162db78 , n60610 );
buf ( R_1232_156aaa58 , C0 );
buf ( R_15bb_117f3338 , n60611 );
buf ( R_8e0_14a0f698 , n60612 );
buf ( R_f9c_14a104f8 , n60613 );
buf ( R_eff_13d381d8 , n60614 );
buf ( R_151e_15883af8 , C0 );
buf ( R_97d_14a16178 , n60642 );
buf ( R_1702_13cd9198 , C0 );
buf ( R_10e3_117f2f78 , n60643 );
buf ( R_ac4_1700f028 , n60644 );
buf ( R_799_13d5a018 , n60687 );
buf ( R_db8_150e6998 , n60688 );
buf ( R_13d7_14b1d1b8 , n60689 );
buf ( R_19f6_1580aa58 , C0 );
buf ( R_14fd_156b56d8 , n60738 );
buf ( R_15dc_123bfd98 , n60739 );
buf ( R_fbd_14a0b098 , n60767 );
buf ( R_8bf_14875f58 , n60768 );
buf ( R_99e_15ff9388 , C0 );
buf ( R_ede_11634338 , C0 );
buf ( R_188d_17018e48 , n60800 );
buf ( R_126e_150e04f8 , C0 );
buf ( R_c4f_15814918 , n60801 );
buf ( R_630_13d25558 , n60802 );
buf ( R_60e_13cd3d38 , C0 );
buf ( R_c2d_1580aaf8 , n60852 );
buf ( R_124c_13d40018 , n60853 );
buf ( R_186b_13d42bd8 , n60854 );
buf ( R_1a23_13d52458 , n60855 );
buf ( R_1404_1486a8d8 , n60856 );
buf ( R_de5_11633a78 , n60899 );
buf ( R_7c6_156b9738 , C0 );
buf ( R_a97_13c05e58 , n60900 );
buf ( R_10b6_124c3638 , C0 );
buf ( R_16d5_123bc4b8 , n60925 );
buf ( R_bed_13b90db8 , n60976 );
buf ( R_c8f_117ef4b8 , n60977 );
buf ( R_120c_13ddcd38 , n60978 );
buf ( R_670_13ccfaf8 , n60979 );
buf ( R_182b_13cd80b8 , n60980 );
buf ( R_18cd_13c1ca18 , n61012 );
buf ( R_5ce_14b1ded8 , C0 );
buf ( R_12ae_13c1f178 , C0 );
buf ( R_bc6_13cd7bb8 , C0 );
buf ( R_697_13bf83d8 , n61013 );
buf ( R_18f4_15881cf8 , n61014 );
buf ( R_11e5_1162add8 , n61049 );
buf ( R_12d5_17015928 , n61069 );
buf ( R_1804_150e44b8 , n61070 );
buf ( R_5a7_12fbe178 , n61077 );
buf ( R_cb6_1162e398 , C0 );
buf ( R_110f_15887518 , n61078 );
buf ( R_19ca_156b8a18 , C0 );
buf ( R_af0_17012a48 , n61079 );
buf ( R_76d_156b1df8 , n61122 );
buf ( R_d8c_15814b98 , n61123 );
buf ( R_172e_117ed438 , C0 );
buf ( R_13ab_13b99878 , n61124 );
buf ( R_1a12_13d52ef8 , C0 );
buf ( R_13f3_156b74d8 , n61125 );
buf ( R_dd4_140ac5d8 , n61126 );
buf ( R_7b5_13c1f718 , n61169 );
buf ( R_aa8_14a0ea18 , n61170 );
buf ( R_10c7_13df2c38 , n61171 );
buf ( R_16e6_156b9eb8 , C0 );
buf ( R_15cd_13cd86f8 , n61187 );
buf ( R_8ce_13d1e2f8 , C0 );
buf ( R_fae_13bf6df8 , C0 );
buf ( R_eed_15812578 , n61224 );
buf ( R_98f_117f62b8 , n61225 );
buf ( R_150c_15ff3848 , n61226 );
buf ( R_908_123c0658 , n61227 );
buf ( R_f27_13cd08b8 , n61228 );
buf ( R_1546_14a18f18 , C0 );
buf ( R_1593_13d58e98 , n61229 );
buf ( R_f74_158805d8 , n61230 );
buf ( R_955_1580f0f8 , n61258 );
buf ( R_d5c_1580ed38 , n61259 );
buf ( R_137b_13d5cc78 , n61260 );
buf ( R_175e_15813478 , C0 );
buf ( R_199a_117e8b18 , C0 );
buf ( R_113f_123b3098 , n61261 );
buf ( R_73d_13c220f8 , n61304 );
buf ( R_b20_13c06c18 , n61305 );
buf ( R_163a_13d3ddb8 , C0 );
buf ( R_9fc_14a0b818 , n61306 );
buf ( R_e80_11633ed8 , n61307 );
buf ( R_101b_123b6518 , n61308 );
buf ( R_861_124c3bd8 , n61315 );
buf ( R_149f_123b5e38 , n61316 );
buf ( R_1080_14a149b8 , n61317 );
buf ( R_7fc_13d3f258 , n61318 );
buf ( R_169f_124c2d78 , n61319 );
buf ( R_1a59_117eded8 , n61325 );
buf ( R_143a_14a0edd8 , C0 );
buf ( R_a61_1700dd68 , n61359 );
buf ( R_e1b_13cd1178 , n61360 );
buf ( R_140f_117f1cb8 , n61361 );
buf ( R_df0_13c09cd8 , n61362 );
buf ( R_7d1_14b28978 , n61406 );
buf ( R_a8c_123c0338 , n61407 );
buf ( R_10ab_13df0398 , n61408 );
buf ( R_16ca_13d52f98 , C0 );
buf ( R_1a2e_13c22698 , C0 );
buf ( R_b10_14b21fd8 , n61409 );
buf ( R_138b_156b0318 , n61410 );
buf ( R_19aa_14a194b8 , C0 );
buf ( R_174e_15811a38 , C0 );
buf ( R_74d_117f0e58 , n61453 );
buf ( R_112f_156aac38 , n61454 );
buf ( R_d6c_156b62b8 , n61455 );
buf ( R_1781_1162d5d8 , n61506 );
buf ( R_d39_15811b78 , n61549 );
buf ( R_1162_124c2558 , C0 );
buf ( R_1358_156b8e78 , n61550 );
buf ( R_b43_13c06858 , n61551 );
buf ( R_71a_117ee798 , C0 );
buf ( R_1977_15880b78 , n61552 );
buf ( R_1108_13ccfb98 , n61553 );
buf ( R_ae9_1580cd58 , n61584 );
buf ( R_774_1700a7a8 , n61585 );
buf ( R_d93_13cce0b8 , n61586 );
buf ( R_13b2_15886898 , C0 );
buf ( R_1727_14870e18 , n61587 );
buf ( R_19d1_123b5b18 , n61599 );
buf ( R_188e_11c6a698 , C0 );
buf ( R_126f_14b23c98 , n61600 );
buf ( R_c50_13d471d8 , n61601 );
buf ( R_631_13ddd7d8 , n61644 );
buf ( R_60d_117f3a18 , n61687 );
buf ( R_c2c_13d2c498 , n61688 );
buf ( R_124b_156b97d8 , n61689 );
buf ( R_186a_13ddb118 , C0 );
buf ( R_fdc_1162ca98 , n61690 );
buf ( R_14de_13c202f8 , C0 );
buf ( R_9bd_11632cb8 , n61709 );
buf ( R_8a0_13bf81f8 , n61710 );
buf ( R_15fb_123ba078 , n61711 );
buf ( R_ebf_13b91678 , n61712 );
buf ( R_e94_148719f8 , n61713 );
buf ( R_9e8_15ff97e8 , n61714 );
buf ( R_1626_13de2918 , C0 );
buf ( R_14b3_13dde9f8 , n61715 );
buf ( R_875_156aea18 , n61730 );
buf ( R_1007_15881578 , n61731 );
buf ( R_14f6_11638938 , C0 );
buf ( R_fc4_1580d578 , n61732 );
buf ( R_8b8_123ba2f8 , n61733 );
buf ( R_9a5_117ecc18 , n61752 );
buf ( R_ed7_14a0da78 , n61753 );
buf ( R_15e3_123c0158 , n61754 );
buf ( R_e0c_1700d0e8 , n61755 );
buf ( R_16ae_123b38b8 , C0 );
buf ( R_7ed_117ef738 , n61804 );
buf ( R_1a4a_12fc1c38 , C0 );
buf ( R_a70_150dbc78 , n61805 );
buf ( R_142b_15889bd8 , n61806 );
buf ( R_108f_13de36d8 , n61807 );
buf ( R_d4e_11c6b6d8 , C0 );
buf ( R_176c_13ddfcb8 , n61808 );
buf ( R_136d_11634dd8 , n61851 );
buf ( R_114d_158861b8 , n61875 );
buf ( R_198c_13d53a38 , n61876 );
buf ( R_72f_11637498 , n61877 );
buf ( R_b2e_170098a8 , C0 );
buf ( R_8f7_13b8e298 , n61878 );
buf ( R_f16_1587d838 , C0 );
buf ( R_1535_13ded2d8 , n61934 );
buf ( R_15a4_1162bcd8 , n61935 );
buf ( R_f85_170174a8 , n61971 );
buf ( R_966_156acd58 , C0 );
buf ( R_12a4_13cd0db8 , n61972 );
buf ( R_1216_13c26518 , C0 );
buf ( R_c85_13d505b8 , n62019 );
buf ( R_1835_13b8eb58 , n62050 );
buf ( R_666_13cd8798 , C0 );
buf ( R_5d8_14a11fd8 , n62051 );
buf ( R_18c3_156b8c98 , n62052 );
buf ( R_bf7_156b4418 , n62053 );
buf ( R_15d5_117ed898 , n62069 );
buf ( R_fb6_14b24558 , C0 );
buf ( R_8c6_13d442f8 , C0 );
buf ( R_997_123bb478 , n62070 );
buf ( R_ee5_14a14af8 , n62119 );
buf ( R_1504_13d553d8 , n62120 );
buf ( R_6d1_158167b8 , n62163 );
buf ( R_130f_156ab4f8 , n62164 );
buf ( R_17ca_150df9b8 , C0 );
buf ( R_b8c_124c3ef8 , n62165 );
buf ( R_cf0_11c6a878 , n62166 );
buf ( R_192e_150e8a18 , C0 );
buf ( R_11ab_13d29d38 , n62167 );
buf ( R_56d_156b76b8 , n62169 );
buf ( R_1704_13bf4238 , n62170 );
buf ( R_10e5_14871778 , n62203 );
buf ( R_ac6_1587bcb8 , C0 );
buf ( R_797_14b1c178 , n62204 );
buf ( R_db6_13ddd058 , C0 );
buf ( R_13d5_1587c618 , n62247 );
buf ( R_19f4_150e3ab8 , n62248 );
buf ( R_1298_156b1d58 , n62249 );
buf ( R_1841_13d2c538 , n62264 );
buf ( R_c79_156b5598 , n62307 );
buf ( R_65a_14874ab8 , C0 );
buf ( R_5e4_13bf0278 , n62308 );
buf ( R_c03_14a0d2f8 , n62309 );
buf ( R_18b7_13ccd1b8 , n62310 );
buf ( R_1222_14b1acd8 , C0 );
buf ( R_1073_14b20f98 , n62311 );
buf ( R_809_13d3e678 , n62367 );
buf ( R_1a66_123b6158 , C0 );
buf ( R_1692_117f31f8 , C0 );
buf ( R_1447_13b93338 , n62368 );
buf ( R_e28_156abbd8 , n62369 );
buf ( R_a54_13cce838 , n62370 );
buf ( R_1054_13bf8ab8 , n62371 );
buf ( R_1466_13d5abf8 , C0 );
buf ( R_1673_1580e798 , n62372 );
buf ( R_e47_1587b178 , n62373 );
buf ( R_a35_117f5db8 , n62380 );
buf ( R_828_10081f38 , n62381 );
buf ( R_1469_1587ee18 , n62424 );
buf ( R_1051_11635c38 , n62457 );
buf ( R_e4a_11629118 , C0 );
buf ( R_1670_1007f238 , n62458 );
buf ( R_82b_13cd7258 , n62459 );
buf ( R_a32_1486afb8 , C0 );
buf ( R_1187_117f4198 , n62460 );
buf ( R_1952_14a0c0d8 , C0 );
buf ( R_d14_13dee778 , n62461 );
buf ( R_b68_10089d78 , n62462 );
buf ( R_17a6_15811f38 , C0 );
buf ( R_1333_117f21b8 , n62463 );
buf ( R_6f5_13d43678 , n62506 );
buf ( R_6c8_1580d758 , n62507 );
buf ( R_1306_1580d938 , C0 );
buf ( R_17d3_13d3a578 , n62508 );
buf ( R_b95_117f7618 , n62540 );
buf ( R_ce7_13d27218 , n62541 );
buf ( R_1925_15ff0328 , n62592 );
buf ( R_11b4_13b8ec98 , n62593 );
buf ( R_576_13d2bf98 , n62594 );
buf ( R_e00_13cd8bf8 , n62595 );
buf ( R_7e1_150e4058 , n62654 );
buf ( R_a7c_156b7118 , n62655 );
buf ( R_1a3e_14a0b278 , C0 );
buf ( R_109b_123bd4f8 , n62656 );
buf ( R_141f_1008c578 , n62657 );
buf ( R_16ba_156b6e98 , C0 );
buf ( R_188f_156b5458 , n62658 );
buf ( R_1270_14a103b8 , n62659 );
buf ( R_c51_11630af8 , n62686 );
buf ( R_632_13ccde38 , C0 );
buf ( R_60c_13dd9c78 , n62687 );
buf ( R_c2b_14b23478 , n62688 );
buf ( R_124a_140b7898 , C0 );
buf ( R_1869_14b29cd8 , n62723 );
buf ( R_1a14_117ebbd8 , n62724 );
buf ( R_13f5_13cd8a18 , n62767 );
buf ( R_dd6_13de0d98 , C0 );
buf ( R_7b7_15816a38 , n62768 );
buf ( R_aa6_13d28c58 , C0 );
buf ( R_10c5_11632998 , n62807 );
buf ( R_16e4_10087078 , n62808 );
buf ( R_190c_13d1d998 , n62809 );
buf ( R_6af_124c33b8 , n62810 );
buf ( R_bae_1587b5d8 , C0 );
buf ( R_12ed_14a176b8 , n62853 );
buf ( R_11cd_13cd27f8 , n62871 );
buf ( R_cce_116331b8 , C0 );
buf ( R_58f_156b9558 , n62872 );
buf ( R_17ec_13dd7fb8 , n62873 );
buf ( R_1057_123bd278 , n62874 );
buf ( R_1463_124c4b78 , n62875 );
buf ( R_1676_140ae6f8 , C0 );
buf ( R_e44_148741f8 , n62876 );
buf ( R_a38_150dc3f8 , n62877 );
buf ( R_825_123b3278 , n62933 );
buf ( R_18a8_1580c8f8 , n62934 );
buf ( R_1289_13c09738 , n62985 );
buf ( R_c6a_15811fd8 , C0 );
buf ( R_64b_1007d938 , n62986 );
buf ( R_5f3_116307d8 , n62987 );
buf ( R_c12_1162cc78 , C0 );
buf ( R_1231_13dee9f8 , n63019 );
buf ( R_1850_1587f778 , n63020 );
buf ( R_146c_14872f38 , n63021 );
buf ( R_104e_1580f7d8 , C0 );
buf ( R_e4d_14b20d18 , n63068 );
buf ( R_166d_13d20058 , n63096 );
buf ( R_82e_1580f2d8 , C0 );
buf ( R_a2f_123b3db8 , n63097 );
buf ( R_19c3_116340b8 , n63098 );
buf ( R_af7_13cd2d98 , n63099 );
buf ( R_766_13c07618 , C0 );
buf ( R_1735_13bf9f58 , n63126 );
buf ( R_d85_13dd7518 , n63169 );
buf ( R_13a4_150ea138 , n63170 );
buf ( R_1116_13c02438 , C0 );
buf ( R_df9_13dd9458 , n63213 );
buf ( R_7da_14a16fd8 , C0 );
buf ( R_a83_13b9a278 , n63214 );
buf ( R_10a2_123b3d18 , C0 );
buf ( R_1a37_1587f958 , n63215 );
buf ( R_16c1_13d3d458 , n63234 );
buf ( R_1418_13d2b1d8 , n63235 );
buf ( R_ea1_156b5c78 , n63291 );
buf ( R_9db_13c05bd8 , n63292 );
buf ( R_1619_15888d78 , n63299 );
buf ( R_14c0_17012fe8 , n63300 );
buf ( R_882_13dee458 , C0 );
buf ( R_ffa_11c68f78 , C0 );
buf ( R_1967_15ff9608 , n63301 );
buf ( R_1172_170122c8 , C0 );
buf ( R_d29_13bed898 , n63344 );
buf ( R_1348_156b1178 , n63345 );
buf ( R_b53_1162fe78 , n63346 );
buf ( R_1791_15ff73a8 , n63396 );
buf ( R_70a_13dee818 , C0 );
buf ( R_8ea_13b91c18 , C0 );
buf ( R_15b1_140b0d18 , n63412 );
buf ( R_f09_13d4f9d8 , n63418 );
buf ( R_f92_13b99238 , C0 );
buf ( R_1528_13cca918 , n63419 );
buf ( R_973_12fc1738 , n63420 );
buf ( R_907_13d1cef8 , n63421 );
buf ( R_f26_13d51378 , C0 );
buf ( R_1545_13ddab78 , n63477 );
buf ( R_1594_123b52f8 , n63478 );
buf ( R_f75_1587ec38 , n63494 );
buf ( R_956_117f3bf8 , C0 );
buf ( R_a1c_13d42098 , n63495 );
buf ( R_147f_15ffd208 , n63496 );
buf ( R_103b_12fbfbb8 , n63497 );
buf ( R_e60_13b98dd8 , n63498 );
buf ( R_165a_156b9418 , C0 );
buf ( R_841_13de1e78 , n63554 );
buf ( R_1715_13c03ab8 , n63578 );
buf ( R_10f6_1587fc78 , C0 );
buf ( R_ad7_11c6aaf8 , n63579 );
buf ( R_786_13bf7938 , C0 );
buf ( R_da5_13c24c18 , n63622 );
buf ( R_13c4_156adbb8 , n63623 );
buf ( R_19e3_13b8b4f8 , n63624 );
buf ( R_15c5_13cce478 , n63640 );
buf ( R_8d6_14a156d8 , C0 );
buf ( R_fa6_13ccd7f8 , C0 );
buf ( R_ef5_13c0f8b8 , n63874 );
buf ( R_987_148737f8 , n63875 );
buf ( R_1514_13d4ea38 , n63876 );
buf ( R_d36_13cd2938 , C0 );
buf ( R_1165_1700dae8 , n63891 );
buf ( R_1355_13c0e2d8 , n63934 );
buf ( R_b46_12fbedf8 , C0 );
buf ( R_717_13c1ebd8 , n63935 );
buf ( R_1974_13b938d8 , n63936 );
buf ( R_1784_14b1b3b8 , n63937 );
buf ( R_156d_13b91d58 , n63987 );
buf ( R_f4e_13d2bb38 , C0 );
buf ( R_156c_1486f8d8 , n63988 );
buf ( R_92f_1587e418 , n63989 );
buf ( R_f4d_158174d8 , n64005 );
buf ( R_92e_15880df8 , C0 );
buf ( R_156e_13bee0b8 , C0 );
buf ( R_f4f_13d1f298 , n64006 );
buf ( R_930_117f5818 , n64007 );
buf ( R_156b_13cd6a38 , n64008 );
buf ( R_f4c_13d4edf8 , n64009 );
buf ( R_92d_13b93838 , n64053 );
buf ( R_156f_1700c828 , n64054 );
buf ( R_f50_13d5d038 , n64055 );
buf ( R_931_1007f198 , n64087 );
buf ( R_92c_13bef238 , n64088 );
buf ( R_156a_14a0d7f8 , C0 );
buf ( R_f4b_1162df38 , n64089 );
buf ( R_682_13dd6a78 , C0 );
buf ( R_11fa_12fbfe38 , C0 );
buf ( R_18df_1162e1b8 , n64090 );
buf ( R_1819_117f44b8 , n64121 );
buf ( R_12c0_156b3478 , n64122 );
buf ( R_5bc_150db098 , n64123 );
buf ( R_ca1_15888af8 , n64166 );
buf ( R_bdb_123b9178 , n64167 );
buf ( R_1890_13c0a4f8 , n64168 );
buf ( R_1271_13cd3e78 , n64219 );
buf ( R_c52_11629cf8 , C0 );
buf ( R_633_1587c6b8 , n64220 );
buf ( R_60b_17014c08 , n64221 );
buf ( R_c2a_13c01d58 , C0 );
buf ( R_1249_150de798 , n64253 );
buf ( R_1868_13cd62b8 , n64254 );
buf ( R_105a_14a112b8 , C0 );
buf ( R_1460_158862f8 , n64255 );
buf ( R_1679_13cd44b8 , n64283 );
buf ( R_e41_14a14e18 , n64326 );
buf ( R_a3b_13cd1998 , n64327 );
buf ( R_822_117e9158 , C0 );
buf ( R_1570_13d44118 , n64328 );
buf ( R_f51_13ccb778 , n64344 );
buf ( R_932_15810d18 , C0 );
buf ( R_92b_14a180b8 , n64345 );
buf ( R_f4a_1162c8b8 , C0 );
buf ( R_1569_13bede38 , n64380 );
buf ( R_163e_12fc0338 , C0 );
buf ( R_a00_13df4df8 , n64381 );
buf ( R_e7c_13c08798 , n64382 );
buf ( R_101f_117ed9d8 , n64383 );
buf ( R_85d_117f4738 , n64392 );
buf ( R_149b_13cd1038 , n64393 );
buf ( R_146f_117f47d8 , n64394 );
buf ( R_104b_158885f8 , n64395 );
buf ( R_e50_12fbe858 , n64396 );
buf ( R_166a_1587c938 , C0 );
buf ( R_831_156b2398 , n64452 );
buf ( R_a2c_11c701d8 , n64453 );
buf ( R_801_150e6e98 , n64509 );
buf ( R_169a_13b94878 , C0 );
buf ( R_1a5e_1162d3f8 , C0 );
buf ( R_143f_13b8c218 , n64510 );
buf ( R_a5c_13b8c178 , n64511 );
buf ( R_e20_13ddd0f8 , n64512 );
buf ( R_107b_156b2118 , n64513 );
buf ( R_d51_13df3b38 , n64556 );
buf ( R_1769_14b21038 , n64590 );
buf ( R_1370_13cd2618 , n64591 );
buf ( R_114a_13c218d8 , C0 );
buf ( R_198f_13d28bb8 , n64592 );
buf ( R_732_13d55fb8 , C0 );
buf ( R_b2b_13ccd2f8 , n64593 );
buf ( R_1571_1580af58 , n64642 );
buf ( R_f52_12fc1ff8 , C0 );
buf ( R_933_14868718 , n64643 );
buf ( R_92a_13c01a38 , C0 );
buf ( R_f49_13d4f4d8 , n64659 );
buf ( R_1568_1580c218 , n64660 );
buf ( R_1706_15814eb8 , C0 );
buf ( R_10e7_14a160d8 , n64661 );
buf ( R_ac8_156afa58 , n64662 );
buf ( R_795_14a12b18 , n64705 );
buf ( R_db4_117edd98 , n64706 );
buf ( R_13d3_13b90f98 , n64707 );
buf ( R_19f2_12fbf258 , C0 );
buf ( R_17b9_156b0b38 , n64741 );
buf ( R_193f_13d3aa78 , n64742 );
buf ( R_b7b_13befeb8 , n64743 );
buf ( R_d01_140ab318 , n64790 );
buf ( R_119a_13b8a5f8 , C0 );
buf ( R_1320_14b27f78 , n64791 );
buf ( R_55c_11630e18 , n64793 );
buf ( R_6e2_158149b8 , C0 );
buf ( R_106b_117f3518 , n64794 );
buf ( R_168a_117eb598 , C0 );
buf ( R_144f_14b26718 , n64795 );
buf ( R_e30_123b3e58 , n64796 );
buf ( R_a4c_170172c8 , n64797 );
buf ( R_811_15882478 , n64853 );
buf ( R_1406_148665f8 , C0 );
buf ( R_de7_1007fcd8 , n64854 );
buf ( R_7c8_156b7f78 , n64855 );
buf ( R_a95_117f6cb8 , n64901 );
buf ( R_10b4_13d3d598 , n64902 );
buf ( R_16d3_1700be28 , n64903 );
buf ( R_1a25_13b9a318 , n64910 );
buf ( R_1572_156b67b8 , C0 );
buf ( R_f53_123c01f8 , n64911 );
buf ( R_934_156b0958 , n64912 );
buf ( R_929_13d5bf58 , n64940 );
buf ( R_f48_13c256b8 , n64941 );
buf ( R_1567_13b91e98 , n64942 );
buf ( R_1943_11c70598 , n64943 );
buf ( R_d05_13c0cd98 , n64986 );
buf ( R_b77_13d415f8 , n64987 );
buf ( R_17b5_14a12118 , n65011 );
buf ( R_1324_15887298 , n65012 );
buf ( R_6e6_13becb78 , C0 );
buf ( R_558_116299d8 , n65014 );
buf ( R_1196_13d4f398 , C0 );
buf ( R_e98_13d433f8 , n65015 );
buf ( R_9e4_13cccdf8 , n65016 );
buf ( R_1622_13c044b8 , C0 );
buf ( R_14b7_13d21318 , n65017 );
buf ( R_879_15884c78 , n65023 );
buf ( R_1003_124c39f8 , n65024 );
buf ( R_1a16_1486b418 , C0 );
buf ( R_13f7_13d24338 , n65025 );
buf ( R_dd8_1587fd18 , n65026 );
buf ( R_7b9_13c0f458 , n65069 );
buf ( R_aa4_13c1d0f8 , n65070 );
buf ( R_10c3_13ccbef8 , n65071 );
buf ( R_16e2_140b6df8 , C0 );
buf ( R_1573_14a0c498 , n65072 );
buf ( R_f54_11632858 , n65073 );
buf ( R_935_150e5318 , n65105 );
buf ( R_928_156aab98 , n65106 );
buf ( R_f47_13cd9238 , n65107 );
buf ( R_1566_123b2a58 , C0 );
buf ( R_a0b_11637858 , n65108 );
buf ( R_e71_14b21a38 , n65157 );
buf ( R_102a_11c6ccb8 , C0 );
buf ( R_852_14b1d938 , C0 );
buf ( R_1490_13bf8158 , n65158 );
buf ( R_1649_13dd4f98 , n65186 );
buf ( R_a12_1008b358 , C0 );
buf ( R_e6a_156b7a78 , C0 );
buf ( R_1031_14b25778 , n65211 );
buf ( R_84b_156ad1b8 , n65212 );
buf ( R_1650_13dd4e58 , n65213 );
buf ( R_1489_13c21978 , n65256 );
buf ( R_7e8_1486a0b8 , n65257 );
buf ( R_1a45_1162e2f8 , n65263 );
buf ( R_a75_156b0778 , n65291 );
buf ( R_1426_11637718 , C0 );
buf ( R_1094_13d28398 , n65292 );
buf ( R_16b3_117efeb8 , n65293 );
buf ( R_e07_13d453d8 , n65294 );
buf ( R_17bd_1162b918 , n65321 );
buf ( R_b7f_14a0be58 , n65322 );
buf ( R_cfd_13d1d038 , n65365 );
buf ( R_193b_13d39f38 , n65366 );
buf ( R_119e_13c1bcf8 , C0 );
buf ( R_560_12fbf118 , n65368 );
buf ( R_6de_13cd4058 , C0 );
buf ( R_131c_13c245d8 , n65369 );
buf ( R_1891_123b9858 , n65401 );
buf ( R_1272_13dd9ef8 , C0 );
buf ( R_c53_15ff5148 , n65402 );
buf ( R_634_11631818 , n65403 );
buf ( R_60a_156b2758 , C0 );
buf ( R_c29_13cd0598 , n65453 );
buf ( R_1248_12fbfcf8 , n65454 );
buf ( R_1867_14a0ded8 , n65455 );
buf ( R_9cd_13d1f518 , n65486 );
buf ( R_14ce_1008b5d8 , C0 );
buf ( R_160b_14b24cd8 , n65487 );
buf ( R_890_11628df8 , n65488 );
buf ( R_fec_13ccc5d8 , n65489 );
buf ( R_eaf_13d5baf8 , n65490 );
buf ( R_15bc_15889138 , n65491 );
buf ( R_8df_11637358 , n65492 );
buf ( R_f9d_158889b8 , n65520 );
buf ( R_efe_11632b78 , C0 );
buf ( R_97e_13c29718 , C0 );
buf ( R_151d_1700bc48 , n65569 );
buf ( R_ae2_123bdef8 , C0 );
buf ( R_77b_17011828 , n65570 );
buf ( R_d9a_13c047d8 , C0 );
buf ( R_13b9_15ffc948 , n65613 );
buf ( R_19d8_14870b98 , n65614 );
buf ( R_1720_156b9198 , n65615 );
buf ( R_1101_140b7398 , n65666 );
buf ( R_1202_15881898 , C0 );
buf ( R_67a_13de2878 , C0 );
buf ( R_1821_117f1c18 , n65697 );
buf ( R_18d7_1580f378 , n65698 );
buf ( R_5c4_14868fd8 , n65699 );
buf ( R_12b8_11631b38 , n65700 );
buf ( R_be3_13de2198 , n65701 );
buf ( R_c99_13c029d8 , n65744 );
buf ( R_fd1_13c1d058 , n65767 );
buf ( R_14e9_14868538 , n65811 );
buf ( R_9b2_1580b6d8 , C0 );
buf ( R_8ab_14a0fc38 , n65812 );
buf ( R_15f0_140ae3d8 , n65813 );
buf ( R_eca_14a11df8 , C0 );
buf ( R_1574_13cd7cf8 , n65814 );
buf ( R_f55_14b1ac38 , n65830 );
buf ( R_936_140acf38 , C0 );
buf ( R_927_124c4178 , n65831 );
buf ( R_f46_14a0af58 , C0 );
buf ( R_1565_1700e808 , n65896 );
buf ( R_14d3_1580e5b8 , n65897 );
buf ( R_9c8_15fef248 , n65898 );
buf ( R_895_13d532b8 , n65915 );
buf ( R_1606_1007ef18 , C0 );
buf ( R_eb4_117eda78 , n65916 );
buf ( R_fe7_1162ba58 , n65917 );
buf ( R_8f6_156b7b18 , C0 );
buf ( R_f15_158819d8 , n65933 );
buf ( R_15a5_158168f8 , n65949 );
buf ( R_1534_123b9c18 , n65950 );
buf ( R_f86_13c1ce78 , C0 );
buf ( R_967_11c68938 , n65951 );
buf ( R_1901_15817ed8 , n66002 );
buf ( R_6a4_1162c1d8 , n66003 );
buf ( R_bb9_156ab1d8 , n66032 );
buf ( R_12e2_11636a98 , C0 );
buf ( R_11d8_156aa738 , n66033 );
buf ( R_cc3_15887c98 , n66034 );
buf ( R_59a_117f76b8 , n66040 );
buf ( R_17f7_117e9838 , n66041 );
buf ( R_105d_123b4998 , n66064 );
buf ( R_145d_123bec18 , n66107 );
buf ( R_167c_140b6178 , n66108 );
buf ( R_e3e_150da7d8 , C0 );
buf ( R_a3e_11635cd8 , C0 );
buf ( R_81f_156b45f8 , n66109 );
buf ( R_120b_13def358 , n66110 );
buf ( R_671_140b4058 , n66153 );
buf ( R_182a_117ef698 , C0 );
buf ( R_18ce_156b4e18 , C0 );
buf ( R_5cd_14a185b8 , n66168 );
buf ( R_12af_15ff69a8 , n66169 );
buf ( R_bec_124c2878 , n66170 );
buf ( R_c90_117eb778 , n66171 );
buf ( R_1386_14a0c7b8 , C0 );
buf ( R_19a5_1008a598 , n66182 );
buf ( R_1753_13cd1218 , n66183 );
buf ( R_748_13d3b518 , n66184 );
buf ( R_1134_1580ad78 , n66185 );
buf ( R_d67_13d3caf8 , n66186 );
buf ( R_b15_156b2078 , n66200 );
buf ( R_128a_15880718 , C0 );
buf ( R_c6b_14a13518 , n66201 );
buf ( R_64c_148739d8 , n66202 );
buf ( R_5f2_13dd5538 , C0 );
buf ( R_c11_15ff5aa8 , n66253 );
buf ( R_1230_124c42b8 , n66254 );
buf ( R_184f_1587fa98 , n66255 );
buf ( R_18a9_11c6f918 , n66280 );
buf ( R_bbf_1587ddd8 , n66281 );
buf ( R_69e_123b5bb8 , C0 );
buf ( R_18fb_13df16f8 , n66282 );
buf ( R_11de_10089058 , C0 );
buf ( R_12dc_13c0bc18 , n66283 );
buf ( R_17fd_13d408d8 , n66314 );
buf ( R_5a0_11631db8 , n66321 );
buf ( R_cbd_14872df8 , n66364 );
buf ( R_691_15883378 , n66407 );
buf ( R_18ee_14a171b8 , C0 );
buf ( R_11eb_13d4f078 , n66408 );
buf ( R_12cf_158850d8 , n66409 );
buf ( R_180a_13d3fc58 , C0 );
buf ( R_5ad_14a0c2b8 , n66415 );
buf ( R_cb0_13de1658 , n66416 );
buf ( R_bcc_13df1f18 , n66417 );
buf ( R_1472_13d3c698 , C0 );
buf ( R_1048_13df8bd8 , n66418 );
buf ( R_e53_10087b18 , n66419 );
buf ( R_1667_13beaf58 , n66420 );
buf ( R_834_15888698 , n66421 );
buf ( R_a29_13de0618 , n66437 );
buf ( R_1575_13d42598 , n66486 );
buf ( R_f56_13c0c578 , C0 );
buf ( R_937_15886c58 , n66487 );
buf ( R_926_158846d8 , C0 );
buf ( R_f45_13d4f438 , n66503 );
buf ( R_1564_1587b038 , n66504 );
buf ( R_906_14a145f8 , C0 );
buf ( R_f25_13d24e78 , n66520 );
buf ( R_1544_124c4fd8 , n66521 );
buf ( R_1595_14b1f698 , n66527 );
buf ( R_f76_117f6fd8 , C0 );
buf ( R_957_15888878 , n66528 );
buf ( R_c7a_140ac998 , C0 );
buf ( R_65b_1580b778 , n66529 );
buf ( R_5e3_117eba98 , n66530 );
buf ( R_c02_123b2f58 , C0 );
buf ( R_18b8_12fc05b8 , n66531 );
buf ( R_1221_15812cf8 , n66563 );
buf ( R_1299_14b1fc38 , n66614 );
buf ( R_1840_13d549d8 , n66615 );
buf ( R_1947_156ac3f8 , n66616 );
buf ( R_d09_150dd438 , n66659 );
buf ( R_b73_117f7938 , n66660 );
buf ( R_17b1_14a0dcf8 , n66706 );
buf ( R_1328_13d2aeb8 , n66707 );
buf ( R_6ea_123bbb58 , C0 );
buf ( R_1192_1587dbf8 , C0 );
buf ( R_137e_13c27738 , C0 );
buf ( R_175b_15883ff8 , n66708 );
buf ( R_199d_1008a6d8 , n66720 );
buf ( R_113c_13d20eb8 , n66721 );
buf ( R_740_13bf6b78 , n66722 );
buf ( R_b1d_123c1918 , n66753 );
buf ( R_d5f_15888c38 , n66754 );
buf ( R_fcb_13def8f8 , n66755 );
buf ( R_8b1_170124a8 , n66772 );
buf ( R_9ac_14a190f8 , n66773 );
buf ( R_ed0_13d23d98 , n66774 );
buf ( R_15ea_1580e658 , C0 );
buf ( R_14ef_123bead8 , n66775 );
buf ( R_d33_123bd8b8 , n66776 );
buf ( R_1168_156b6fd8 , n66777 );
buf ( R_1352_13c10b78 , C0 );
buf ( R_b49_14a158b8 , n66811 );
buf ( R_714_1587c898 , n66812 );
buf ( R_1971_13ddfe98 , n66823 );
buf ( R_1787_1486e2f8 , n66824 );
buf ( R_68a_14a15b38 , C0 );
buf ( R_11f2_1162a6f8 , C0 );
buf ( R_18e7_13c08c98 , n66825 );
buf ( R_1811_117e9a18 , n66839 );
buf ( R_12c8_140aa878 , n66840 );
buf ( R_5b4_140b2a78 , n66841 );
buf ( R_ca9_15887e78 , n66884 );
buf ( R_bd3_13c0e9b8 , n66885 );
buf ( R_195d_15884818 , n66897 );
buf ( R_117c_14874838 , n66898 );
buf ( R_d1f_1007f698 , n66899 );
buf ( R_b5d_123bb8d8 , n66934 );
buf ( R_133e_13d55dd8 , C0 );
buf ( R_179b_12fbde58 , n66935 );
buf ( R_700_13cd9878 , n66936 );
buf ( R_1576_1700c6e8 , C0 );
buf ( R_f57_14a14198 , n66937 );
buf ( R_938_13bedc58 , n66938 );
buf ( R_925_13df1338 , n66961 );
buf ( R_f44_156b99b8 , n66962 );
buf ( R_1563_158841d8 , n66963 );
buf ( R_c86_14a12e38 , C0 );
buf ( R_1834_13cd3f18 , n66964 );
buf ( R_667_1486b558 , n66965 );
buf ( R_5d7_156b0c78 , n66966 );
buf ( R_18c4_11c709f8 , n66967 );
buf ( R_bf6_11c6f378 , C0 );
buf ( R_12a5_1162d718 , n67017 );
buf ( R_1215_117f51d8 , n67042 );
buf ( R_1892_13d3b1f8 , C0 );
buf ( R_1273_13dd5c18 , n67043 );
buf ( R_c54_13becd58 , n67044 );
buf ( R_635_13d2c678 , n67087 );
buf ( R_609_1580ef18 , n67130 );
buf ( R_c28_140ba098 , n67131 );
buf ( R_1247_13ccda78 , n67132 );
buf ( R_1866_13bf9eb8 , C0 );
buf ( R_9d2_13ccb958 , C0 );
buf ( R_14c9_117f80b8 , n67175 );
buf ( R_1610_1700a988 , n67176 );
buf ( R_88b_1587e5f8 , n67177 );
buf ( R_ff1_13b8bd18 , n67199 );
buf ( R_eaa_13dd6618 , C0 );
buf ( R_1708_11630558 , n67200 );
buf ( R_10e9_123c2138 , n67228 );
buf ( R_aca_14a131f8 , C0 );
buf ( R_793_12fc2138 , n67229 );
buf ( R_db2_123b68d8 , C0 );
buf ( R_13d1_156ac998 , n67272 );
buf ( R_19f0_13d47138 , n67273 );
buf ( R_7d3_13dd99f8 , n67274 );
buf ( R_a8a_150e0ef8 , C0 );
buf ( R_10a9_1486ae78 , n67293 );
buf ( R_16c8_13dfaed8 , n67294 );
buf ( R_1a30_14a19698 , n67295 );
buf ( R_1411_13dfa438 , n67338 );
buf ( R_df2_150e09f8 , C0 );
buf ( R_14e3_11634838 , n67339 );
buf ( R_9b8_13d43b78 , n67340 );
buf ( R_8a5_13bee798 , n67357 );
buf ( R_15f6_117f0458 , C0 );
buf ( R_ec4_11c68a78 , n67358 );
buf ( R_fd7_116387f8 , n67359 );
buf ( R_17c1_13d57d18 , n67391 );
buf ( R_b83_13bedd98 , n67392 );
buf ( R_cf9_1587d798 , n67435 );
buf ( R_1937_150e3c98 , n67436 );
buf ( R_11a2_13c05138 , C0 );
buf ( R_564_15815278 , n67437 );
buf ( R_6da_13c00f98 , C0 );
buf ( R_1318_1008a9f8 , n67438 );
buf ( R_faf_158866b8 , n67439 );
buf ( R_8cd_15ff2ee8 , n67456 );
buf ( R_eec_117f7078 , n67457 );
buf ( R_990_11633c58 , n67458 );
buf ( R_150b_13cd8dd8 , n67459 );
buf ( R_15ce_13df0898 , C0 );
buf ( R_1766_116318b8 , C0 );
buf ( R_1373_15810598 , n67460 );
buf ( R_1147_13b8d438 , n67461 );
buf ( R_1992_13b8d1b8 , C0 );
buf ( R_735_13cd4cd8 , n67504 );
buf ( R_b28_1162fab8 , n67505 );
buf ( R_d54_150e15d8 , n67506 );
buf ( R_1577_13d44ed8 , n67507 );
buf ( R_f58_13d3e178 , n67508 );
buf ( R_939_123b2878 , n67540 );
buf ( R_924_140b7118 , n67541 );
buf ( R_f43_140aeab8 , n67542 );
buf ( R_1562_100874d8 , C0 );
buf ( R_17ce_13d50b58 , C0 );
buf ( R_b90_14a17e38 , n67543 );
buf ( R_cec_156b8fb8 , n67544 );
buf ( R_192a_13df93f8 , C0 );
buf ( R_11af_156b2a78 , n67545 );
buf ( R_571_13b96ad8 , n67547 );
buf ( R_6cd_150dc5d8 , n67590 );
buf ( R_130b_14b1eab8 , n67591 );
buf ( R_19b7_117f7758 , n67592 );
buf ( R_75a_150de5b8 , C0 );
buf ( R_1741_100824d8 , n67741 );
buf ( R_d79_1008a638 , n67784 );
buf ( R_1122_150e9a58 , C0 );
buf ( R_1398_10083978 , n67785 );
buf ( R_b03_158129d8 , n67786 );
buf ( R_14d8_13cd4698 , n67787 );
buf ( R_9c3_13befa58 , n67788 );
buf ( R_89a_117edb18 , C0 );
buf ( R_1601_13d272b8 , n67804 );
buf ( R_eb9_11638438 , n67860 );
buf ( R_fe2_13defdf8 , C0 );
buf ( R_13f9_1580cb78 , n67903 );
buf ( R_dda_117f7118 , C0 );
buf ( R_7bb_13bf54f8 , n67904 );
buf ( R_aa2_12fc1a58 , C0 );
buf ( R_10c1_13b901d8 , n67911 );
buf ( R_16e0_158811b8 , n67912 );
buf ( R_1a18_156b8bf8 , n67913 );
buf ( R_fbe_13cd90f8 , C0 );
buf ( R_8be_13df3278 , C0 );
buf ( R_99f_123b6b58 , n67914 );
buf ( R_edd_13b99cd8 , n67923 );
buf ( R_15dd_156aef18 , n67939 );
buf ( R_14fc_140b09f8 , n67940 );
buf ( R_19b2_150e0318 , C0 );
buf ( R_1746_123b75f8 , C0 );
buf ( R_755_14a13338 , n67983 );
buf ( R_1127_13de3318 , n67984 );
buf ( R_d74_17011d28 , n67985 );
buf ( R_b08_150dce98 , n67986 );
buf ( R_1393_11c68c58 , n67987 );
buf ( R_1956_15813158 , C0 );
buf ( R_d18_156b9698 , n67988 );
buf ( R_b64_156b3a18 , n67989 );
buf ( R_17a2_117e8758 , C0 );
buf ( R_1337_13d20af8 , n67990 );
buf ( R_6f9_17012b88 , n68033 );
buf ( R_1183_1580f698 , n68034 );
buf ( R_bb3_17013d08 , n68035 );
buf ( R_12e8_14b1e158 , n68036 );
buf ( R_11d2_124c3318 , C0 );
buf ( R_cc9_11c6e018 , n68079 );
buf ( R_594_13cd9698 , n68085 );
buf ( R_17f1_13c0bdf8 , n68100 );
buf ( R_1907_13ccaa58 , n68101 );
buf ( R_6aa_13de4038 , C0 );
buf ( R_ba3_13cd5bd8 , n68102 );
buf ( R_12f8_13cd2758 , n68103 );
buf ( R_11c2_13c1fc18 , C0 );
buf ( R_cd9_14b1f878 , n68146 );
buf ( R_584_12fc0bf8 , n68147 );
buf ( R_1917_13d21f98 , n68148 );
buf ( R_17e1_13d37878 , n68163 );
buf ( R_6ba_11637b78 , C0 );
buf ( R_8e9_13cd6b78 , n68180 );
buf ( R_15b2_117f08b8 , C0 );
buf ( R_f08_156b5db8 , n68181 );
buf ( R_f93_13b92758 , n68182 );
buf ( R_1527_13ccaeb8 , n68183 );
buf ( R_974_13c0c2f8 , n68184 );
buf ( R_ad9_150e2a78 , n68199 );
buf ( R_784_13dfa4d8 , n68200 );
buf ( R_da3_14a0cd58 , n68201 );
buf ( R_13c2_13d2a4b8 , C0 );
buf ( R_19e1_1700c5a8 , n68208 );
buf ( R_1717_13df61f8 , n68209 );
buf ( R_10f8_156b7258 , n68210 );
buf ( R_1578_123bab18 , n68211 );
buf ( R_f59_13c10358 , n68227 );
buf ( R_93a_1486f978 , C0 );
buf ( R_923_11632178 , n68228 );
buf ( R_f42_14b1f9b8 , C0 );
buf ( R_1561_13bf4a58 , n68277 );
buf ( R_1060_13c0b358 , n68278 );
buf ( R_145a_14a12bb8 , C0 );
buf ( R_167f_14a19378 , n68279 );
buf ( R_e3b_13dd7f18 , n68280 );
buf ( R_a41_14a10d18 , n68359 );
buf ( R_81c_13bf79d8 , n68360 );
buf ( R_12fd_1007d9d8 , n68403 );
buf ( R_b9e_123ba618 , C0 );
buf ( R_cde_13d39218 , C0 );
buf ( R_11bd_11c6dcf8 , n68419 );
buf ( R_191c_1580c038 , n68420 );
buf ( R_57f_158160d8 , n68421 );
buf ( R_6bf_13df4e98 , n68422 );
buf ( R_17dc_15ff5508 , n68423 );
buf ( R_1893_117f0d18 , n68424 );
buf ( R_1274_156b1218 , n68425 );
buf ( R_c55_13cce338 , n68452 );
buf ( R_636_123c1238 , C0 );
buf ( R_608_13d58678 , n68453 );
buf ( R_c27_13bf2a78 , n68454 );
buf ( R_1246_14b229d8 , C0 );
buf ( R_1865_156b4d78 , n68489 );
buf ( R_772_11634a18 , C0 );
buf ( R_d91_13c0fdb8 , n68532 );
buf ( R_13b0_1486d0d8 , n68533 );
buf ( R_1729_123b6338 , n68579 );
buf ( R_19cf_11c70c78 , n68580 );
buf ( R_110a_156b12b8 , C0 );
buf ( R_aeb_11638758 , n68581 );
buf ( R_e78_117ef0f8 , n68582 );
buf ( R_1023_15ff3ac8 , n68583 );
buf ( R_859_13c0f098 , n68592 );
buf ( R_1497_116337f8 , n68593 );
buf ( R_1642_1162e578 , C0 );
buf ( R_a04_13c22e18 , n68594 );
buf ( R_76b_13ddaad8 , n68595 );
buf ( R_d8a_10085458 , C0 );
buf ( R_1730_11c6fd78 , n68596 );
buf ( R_13a9_15887978 , n68639 );
buf ( R_1111_11629c58 , n68680 );
buf ( R_19c8_123b61f8 , n68681 );
buf ( R_af2_11635558 , C0 );
buf ( R_1045_13c2abb8 , n68704 );
buf ( R_e56_13c1f0d8 , C0 );
buf ( R_1664_1700d9a8 , n68705 );
buf ( R_837_13d43c18 , n68706 );
buf ( R_a26_13c28c78 , C0 );
buf ( R_1475_123b8bd8 , n68749 );
buf ( R_e63_156b1358 , n68750 );
buf ( R_1038_10085f98 , n68751 );
buf ( R_1657_13cd2c58 , n68752 );
buf ( R_844_117f3ab8 , n68753 );
buf ( R_1482_140b29d8 , C0 );
buf ( R_a19_156ad4d8 , n68777 );
buf ( R_18f5_1587d518 , n68828 );
buf ( R_11e4_158159f8 , n68829 );
buf ( R_12d6_11c6c5d8 , C0 );
buf ( R_1803_123b54d8 , n68830 );
buf ( R_5a6_13ccf5f8 , n68836 );
buf ( R_cb7_1162c458 , n68837 );
buf ( R_bc5_14a0c5d8 , n68880 );
buf ( R_698_14a0feb8 , n68881 );
buf ( R_194b_15882658 , n68882 );
buf ( R_d0d_1580bef8 , n68925 );
buf ( R_b6f_117eb638 , n68926 );
buf ( R_17ad_156b4f58 , n68972 );
buf ( R_132c_158823d8 , n68973 );
buf ( R_6ee_14a0faf8 , C0 );
buf ( R_118e_156ab3b8 , C0 );
buf ( R_75f_14870918 , n68974 );
buf ( R_173c_123b9218 , n68975 );
buf ( R_d7e_11634018 , C0 );
buf ( R_111d_13beeb58 , n69021 );
buf ( R_139d_100868f8 , n69064 );
buf ( R_afe_15ff7ee8 , C0 );
buf ( R_19bc_17010248 , n69065 );
buf ( R_1175_11634c98 , n69096 );
buf ( R_d26_1587cf78 , C0 );
buf ( R_b56_13c236d8 , C0 );
buf ( R_1345_13cd4738 , n69139 );
buf ( R_1794_15813338 , n69140 );
buf ( R_707_13d580d8 , n69141 );
buf ( R_1964_13d42b38 , n69142 );
buf ( R_f24_13b92938 , n69143 );
buf ( R_1543_15ff0828 , n69144 );
buf ( R_1596_15ff8a28 , C0 );
buf ( R_f77_158124d8 , n69145 );
buf ( R_958_13df5bb8 , n69146 );
buf ( R_905_13d4f758 , n69158 );
buf ( R_1579_13b8d078 , n69193 );
buf ( R_f5a_15884d18 , C0 );
buf ( R_93b_1580c3f8 , n69194 );
buf ( R_922_140af198 , C0 );
buf ( R_f41_156b7cf8 , n69210 );
buf ( R_1560_14a14cd8 , n69211 );
buf ( R_c6c_14b20318 , n69212 );
buf ( R_64d_13ccebf8 , n69255 );
buf ( R_5f1_15814c38 , n69298 );
buf ( R_c10_15817898 , n69299 );
buf ( R_122f_13d22038 , n69300 );
buf ( R_184e_14b1b8b8 , C0 );
buf ( R_18aa_11638b18 , C0 );
buf ( R_128b_1587eaf8 , n69301 );
buf ( R_1695_14a12ed8 , n69323 );
buf ( R_1a63_1486ec58 , n69324 );
buf ( R_1444_15ff0788 , n69325 );
buf ( R_a57_13d5aa18 , n69326 );
buf ( R_e25_14a17078 , n69369 );
buf ( R_1076_1587b678 , C0 );
buf ( R_806_14a0bd18 , C0 );
buf ( R_fb7_15887158 , n69370 );
buf ( R_8c5_1008b2b8 , n69386 );
buf ( R_998_13d573b8 , n69387 );
buf ( R_ee4_15ff7da8 , n69388 );
buf ( R_1503_150daf58 , n69389 );
buf ( R_15d6_117ed398 , C0 );
buf ( R_7ca_150de978 , C0 );
buf ( R_a93_156af4b8 , n69390 );
buf ( R_10b2_100826b8 , C0 );
buf ( R_16d1_156b27f8 , n69414 );
buf ( R_1a27_13cd2118 , n69415 );
buf ( R_1408_1587fbd8 , n69416 );
buf ( R_de9_13cd12b8 , n69459 );
buf ( R_9e0_15ffc9e8 , n69460 );
buf ( R_161e_123b8a98 , C0 );
buf ( R_14bb_10081cb8 , n69461 );
buf ( R_87d_123b9498 , n69467 );
buf ( R_fff_12fbe5d8 , n69468 );
buf ( R_e9c_13df34f8 , n69469 );
buf ( R_ba8_123c12d8 , n69470 );
buf ( R_12f3_11634f18 , n69471 );
buf ( R_11c7_17013b28 , n69472 );
buf ( R_cd4_13c2b018 , n69473 );
buf ( R_589_14a19058 , n69474 );
buf ( R_1912_156aacd8 , C0 );
buf ( R_17e6_140b2758 , C0 );
buf ( R_6b5_1587d658 , n69517 );
buf ( R_f14_13d26458 , n69518 );
buf ( R_15a6_1162eb18 , C0 );
buf ( R_1533_14b268f8 , n69519 );
buf ( R_f87_11637998 , n69520 );
buf ( R_968_13d2b958 , n69521 );
buf ( R_8f5_13bebe58 , n69537 );
buf ( R_8d5_150e1c18 , n69554 );
buf ( R_fa7_12fbff78 , n69555 );
buf ( R_ef4_1162ea78 , n69556 );
buf ( R_988_15814198 , n69557 );
buf ( R_1513_13c06498 , n69558 );
buf ( R_15c6_12fbf2f8 , C0 );
buf ( R_8b7_15ffa468 , n69559 );
buf ( R_9a6_13d46058 , C0 );
buf ( R_ed6_13d57598 , C0 );
buf ( R_15e4_156aeb58 , n69560 );
buf ( R_14f5_13c29178 , n69609 );
buf ( R_fc5_13b8d258 , n69637 );
buf ( R_acc_13df8638 , n69638 );
buf ( R_791_13d42818 , n69681 );
buf ( R_db0_13bf9418 , n69682 );
buf ( R_13cf_123c2318 , n69683 );
buf ( R_19ee_11630cd8 , C0 );
buf ( R_170a_13d25698 , C0 );
buf ( R_10eb_13debbb8 , n69684 );
buf ( R_19ad_1587f9f8 , n69696 );
buf ( R_174b_15ff3528 , n69697 );
buf ( R_750_1008c9d8 , n69698 );
buf ( R_112c_13c015d8 , n69699 );
buf ( R_d6f_117eae18 , n69700 );
buf ( R_b0d_13d41c38 , n69731 );
buf ( R_138e_158113f8 , C0 );
buf ( R_168d_156b2f78 , n69759 );
buf ( R_144c_14a0dbb8 , n69760 );
buf ( R_e2d_1587d3d8 , n69803 );
buf ( R_a4f_15814418 , n69804 );
buf ( R_80e_156ac218 , C0 );
buf ( R_106e_14a15318 , C0 );
buf ( R_157a_156b4198 , C0 );
buf ( R_f5b_1162d7b8 , n69805 );
buf ( R_93c_13b933d8 , n69806 );
buf ( R_921_15813298 , n69829 );
buf ( R_f40_13cd1fd8 , n69830 );
buf ( R_155f_148745b8 , n69831 );
buf ( R_1275_13d26bd8 , n69882 );
buf ( R_c56_12fbf438 , C0 );
buf ( R_637_14b20db8 , n69883 );
buf ( R_607_15886258 , n69884 );
buf ( R_c26_13d3ac58 , C0 );
buf ( R_1245_13d261d8 , n69909 );
buf ( R_1864_13ddb2f8 , n69910 );
buf ( R_1894_13cd6998 , n69911 );
buf ( R_9d7_1580ac38 , n69912 );
buf ( R_1615_150e0598 , n69944 );
buf ( R_14c4_15ffa148 , n69945 );
buf ( R_886_156aa9b8 , C0 );
buf ( R_ff6_13d424f8 , C0 );
buf ( R_ea5_13d23b18 , n70001 );
buf ( R_1a51_13cda098 , n70007 );
buf ( R_a69_123b4f38 , n70035 );
buf ( R_1432_14b1d258 , C0 );
buf ( R_1088_13bec3f8 , n70036 );
buf ( R_e13_140ab1d8 , n70037 );
buf ( R_16a7_156afb98 , n70038 );
buf ( R_7f4_14b238d8 , n70039 );
buf ( R_17c5_12fc1058 , n70071 );
buf ( R_b87_140b0db8 , n70072 );
buf ( R_cf5_156ab818 , n70115 );
buf ( R_1933_11633258 , n70116 );
buf ( R_11a6_13c243f8 , C0 );
buf ( R_568_13ccd9d8 , n70117 );
buf ( R_6d6_13ccc498 , C0 );
buf ( R_1314_13b93158 , n70118 );
buf ( R_a81_11c6b098 , n70154 );
buf ( R_10a0_148694d8 , n70155 );
buf ( R_1a39_150e4cd8 , n70161 );
buf ( R_16bf_13d3e8f8 , n70162 );
buf ( R_141a_13ccc678 , C0 );
buf ( R_dfb_123b4c18 , n70163 );
buf ( R_7dc_14b22578 , n70164 );
buf ( R_116b_13ddcb58 , n70165 );
buf ( R_134f_14b1c7b8 , n70166 );
buf ( R_b4c_13d41eb8 , n70167 );
buf ( R_711_140b8798 , n70210 );
buf ( R_178a_13b96538 , C0 );
buf ( R_196e_150e3658 , C0 );
buf ( R_d30_13df5118 , n70211 );
buf ( R_b99_13df2ff8 , n70236 );
buf ( R_ce3_10088b58 , n70237 );
buf ( R_11b8_156b8798 , n70238 );
buf ( R_1921_13b91df8 , n70289 );
buf ( R_57a_13ccb818 , n70290 );
buf ( R_6c4_15887798 , n70291 );
buf ( R_17d7_11c6faf8 , n70292 );
buf ( R_1302_12fbe8f8 , C0 );
buf ( R_65c_117f0278 , n70293 );
buf ( R_5e2_117ef198 , C0 );
buf ( R_c01_13df0118 , n70344 );
buf ( R_18b9_13ded058 , n70369 );
buf ( R_1220_117f77f8 , n70370 );
buf ( R_129a_14a10ef8 , C0 );
buf ( R_183f_140b7f78 , n70371 );
buf ( R_c7b_1580c178 , n70372 );
buf ( R_7bd_12fc1558 , n70415 );
buf ( R_aa0_11c6be58 , n70416 );
buf ( R_10bf_13df54d8 , n70417 );
buf ( R_16de_13de3138 , C0 );
buf ( R_1a1a_156b8ab8 , C0 );
buf ( R_13fb_156b4b98 , n70418 );
buf ( R_ddc_11632df8 , n70419 );
buf ( R_a7a_11c6b1d8 , C0 );
buf ( R_1a40_140b6d58 , n70420 );
buf ( R_1099_116354b8 , n70465 );
buf ( R_1421_117ef7d8 , n70508 );
buf ( R_16b8_13d3ea38 , n70509 );
buf ( R_e02_15ff37a8 , C0 );
buf ( R_7e3_15812118 , n70510 );
buf ( R_1a56_13bf0818 , C0 );
buf ( R_1437_123bad98 , n70511 );
buf ( R_a64_13beb318 , n70512 );
buf ( R_e18_156afc38 , n70513 );
buf ( R_1083_123c0a18 , n70514 );
buf ( R_7f9_156b30b8 , n70570 );
buf ( R_16a2_150e9418 , C0 );
buf ( R_18e0_13c201b8 , n70571 );
buf ( R_1818_140b47d8 , n70572 );
buf ( R_12c1_123bb838 , n70622 );
buf ( R_5bb_156b5638 , n70623 );
buf ( R_ca2_13dd9d18 , C0 );
buf ( R_bda_13b985b8 , C0 );
buf ( R_683_11634478 , n70624 );
buf ( R_11f9_13ccd938 , n70656 );
buf ( R_157b_1486f0b8 , n70657 );
buf ( R_f5c_13de2378 , n70658 );
buf ( R_93d_117f0ef8 , n70690 );
buf ( R_920_13df90d8 , n70691 );
buf ( R_f3f_13bf1a38 , n70692 );
buf ( R_155e_123c0d38 , C0 );
buf ( R_8de_13d4e0d8 , C0 );
buf ( R_f9e_13b8a738 , C0 );
buf ( R_efd_123bfed8 , n70716 );
buf ( R_97f_123c21d8 , n70717 );
buf ( R_151c_13d5c4f8 , n70718 );
buf ( R_15bd_13df43f8 , n70734 );
buf ( R_1763_13d44618 , n70735 );
buf ( R_1995_17017548 , n70746 );
buf ( R_1144_17018948 , n70747 );
buf ( R_738_1700bce8 , n70748 );
buf ( R_b25_1162ad38 , n70763 );
buf ( R_d57_13c242b8 , n70764 );
buf ( R_1376_117f5098 , C0 );
buf ( R_9be_140aaaf8 , C0 );
buf ( R_89f_156b2ed8 , n70765 );
buf ( R_15fc_13c28db8 , n70766 );
buf ( R_ebe_13cd5c78 , C0 );
buf ( R_fdd_1162dd58 , n70788 );
buf ( R_14dd_123b8db8 , n70831 );
buf ( R_14aa_13c0f9f8 , C0 );
buf ( R_86c_13df77d8 , n70832 );
buf ( R_1010_15884278 , n70833 );
buf ( R_e8b_15880ad8 , n70834 );
buf ( R_162f_15ff7808 , n70835 );
buf ( R_9f1_123be718 , n70853 );
buf ( R_1457_13d54758 , n70854 );
buf ( R_1682_1587fb38 , C0 );
buf ( R_e38_150debf8 , n70855 );
buf ( R_a44_1580d618 , n70856 );
buf ( R_819_14873898 , n70912 );
buf ( R_1063_13cd8978 , n70913 );
buf ( R_1a4c_156b8b58 , n70914 );
buf ( R_a6e_117ec3f8 , C0 );
buf ( R_142d_14b1c998 , n70957 );
buf ( R_108d_14a0a878 , n70974 );
buf ( R_e0e_156b9f58 , C0 );
buf ( R_16ac_13bf1218 , n70975 );
buf ( R_7ef_1700c788 , n70976 );
buf ( R_1014_13c079d8 , n70977 );
buf ( R_868_1587de78 , n70978 );
buf ( R_14a6_10081998 , C0 );
buf ( R_1633_117e9ab8 , n70979 );
buf ( R_9f5_13d25c38 , n70997 );
buf ( R_e87_15ff9ce8 , n70998 );
buf ( R_1829_123b40d8 , n71029 );
buf ( R_18cf_13ded238 , n71030 );
buf ( R_5cc_156aa698 , n71031 );
buf ( R_12b0_14a177f8 , n71032 );
buf ( R_beb_13cca738 , n71033 );
buf ( R_c91_15ff1cc8 , n71076 );
buf ( R_120a_13cd9738 , C0 );
buf ( R_672_13c06fd8 , C0 );
buf ( R_779_13cd2258 , n71119 );
buf ( R_d98_13b958b8 , n71120 );
buf ( R_13b7_1700e308 , n71121 );
buf ( R_19d6_117ecfd8 , C0 );
buf ( R_1722_123b5a78 , C0 );
buf ( R_1103_117f7bb8 , n71122 );
buf ( R_ae4_11634ab8 , n71123 );
buf ( R_c57_15814f58 , n71124 );
buf ( R_638_14a151d8 , n71125 );
buf ( R_606_13d50838 , C0 );
buf ( R_c25_10083bf8 , n71175 );
buf ( R_1244_13ddb898 , n71176 );
buf ( R_1863_123b9f38 , n71177 );
buf ( R_1895_13df3a98 , n71209 );
buf ( R_1276_123bda98 , C0 );
buf ( R_1042_13cd6718 , C0 );
buf ( R_e59_1587dd38 , n71252 );
buf ( R_1661_13de0758 , n71284 );
buf ( R_83a_13d21598 , C0 );
buf ( R_a23_14869cf8 , n71285 );
buf ( R_1478_13cd7618 , n71286 );
buf ( R_668_11c6aff8 , n71287 );
buf ( R_5d6_13d24158 , C0 );
buf ( R_18c5_123b5f78 , n71319 );
buf ( R_bf5_123ba7f8 , n71370 );
buf ( R_12a6_148674f8 , C0 );
buf ( R_1214_15886cf8 , n71371 );
buf ( R_c87_13c21bf8 , n71372 );
buf ( R_1833_117f3838 , n71373 );
buf ( R_1820_14872a38 , n71374 );
buf ( R_18d8_13b8ef18 , n71375 );
buf ( R_5c3_10080778 , n71376 );
buf ( R_12b9_140abb38 , n71426 );
buf ( R_be2_13b98338 , C0 );
buf ( R_c9a_13cd1f38 , C0 );
buf ( R_1201_15ff65e8 , n71458 );
buf ( R_67b_13c02bb8 , n71459 );
buf ( R_1542_14a19cd8 , C0 );
buf ( R_1597_117ee478 , n71460 );
buf ( R_f78_156af198 , n71461 );
buf ( R_959_11631bd8 , n71483 );
buf ( R_904_13bebbd8 , n71484 );
buf ( R_f23_13c2b338 , n71485 );
buf ( R_157c_14a0eab8 , n71486 );
buf ( R_f5d_15817c58 , n71502 );
buf ( R_93e_13cd6858 , C0 );
buf ( R_91f_117f7d98 , n71503 );
buf ( R_f3e_1700a708 , C0 );
buf ( R_155d_1700fa28 , n71559 );
buf ( R_764_150dee78 , n71560 );
buf ( R_1737_13cd6538 , n71561 );
buf ( R_d83_150dc678 , n71562 );
buf ( R_1118_13cce3d8 , n71563 );
buf ( R_13a2_13df95d8 , C0 );
buf ( R_af9_14b1bc78 , n71594 );
buf ( R_19c1_15811358 , n71605 );
buf ( R_14ae_14b22438 , C0 );
buf ( R_870_158800d8 , n71606 );
buf ( R_100c_14b1bef8 , n71607 );
buf ( R_e8f_13c27cd8 , n71608 );
buf ( R_9ed_150e3a18 , n71625 );
buf ( R_162b_13d24478 , n71626 );
buf ( R_64e_12fbeb78 , C0 );
buf ( R_5f0_13d25738 , n71627 );
buf ( R_c0f_1587ef58 , n71628 );
buf ( R_122e_14a181f8 , C0 );
buf ( R_184d_1486ac98 , n71643 );
buf ( R_18ab_13bf9d78 , n71644 );
buf ( R_128c_11c6a378 , n71645 );
buf ( R_c6d_13d3be78 , n71688 );
buf ( R_d11_117f09f8 , n71731 );
buf ( R_b6b_13c0e878 , n71732 );
buf ( R_17a9_15ff62c8 , n71761 );
buf ( R_1330_1580d6b8 , n71762 );
buf ( R_6f2_123ba398 , C0 );
buf ( R_118a_13c1eef8 , C0 );
buf ( R_194f_13c0e738 , n71763 );
buf ( R_1758_14a14eb8 , n71764 );
buf ( R_19a0_13c204d8 , n71765 );
buf ( R_1139_117ef878 , n71790 );
buf ( R_743_13d5a478 , n71791 );
buf ( R_b1a_13c01038 , C0 );
buf ( R_d62_15811df8 , C0 );
buf ( R_1381_123b3a98 , n71834 );
buf ( R_e6d_123b7238 , n71893 );
buf ( R_102e_150ddd98 , C0 );
buf ( R_84e_15883418 , C0 );
buf ( R_164d_14a0c678 , n71916 );
buf ( R_148c_1580e8d8 , n71917 );
buf ( R_a0f_15ffbae8 , n71918 );
buf ( R_12ee_13d3d958 , C0 );
buf ( R_11cc_14a11a38 , n71919 );
buf ( R_ccf_15812258 , n71920 );
buf ( R_58e_150e4558 , n71921 );
buf ( R_17eb_150e6538 , n71922 );
buf ( R_190d_14b294b8 , n71973 );
buf ( R_6b0_14a172f8 , n71974 );
buf ( R_bad_15883c38 , n72006 );
buf ( R_1018_13d2a878 , n72007 );
buf ( R_864_13c09238 , n72008 );
buf ( R_14a2_13cd9e18 , C0 );
buf ( R_1637_1162fbf8 , n72009 );
buf ( R_9f9_156b7438 , n72026 );
buf ( R_e83_15886438 , n72027 );
buf ( R_1a5b_13df6158 , n72028 );
buf ( R_143c_15ff2a88 , n72029 );
buf ( R_a5f_13df1518 , n72030 );
buf ( R_e1d_13c288b8 , n72073 );
buf ( R_107e_13c1c298 , C0 );
buf ( R_7fe_117f30b8 , C0 );
buf ( R_169d_156abf98 , n72097 );
buf ( R_15b3_13cd6e98 , n72098 );
buf ( R_f07_13b953b8 , n72099 );
buf ( R_f94_13d25198 , n72100 );
buf ( R_1526_1486bf58 , C0 );
buf ( R_975_13d529f8 , n72128 );
buf ( R_8e8_117f0bd8 , n72129 );
buf ( R_78f_1162c9f8 , n72130 );
buf ( R_dae_11c6d578 , C0 );
buf ( R_13cd_14a162b8 , n72173 );
buf ( R_19ec_15814738 , n72174 );
buf ( R_170c_13ccdd98 , n72175 );
buf ( R_10ed_15882dd8 , n72203 );
buf ( R_ace_15885cb8 , C0 );
buf ( R_157d_13cd56d8 , n72242 );
buf ( R_f5e_140b53b8 , C0 );
buf ( R_93f_13d57778 , n72243 );
buf ( R_91e_15886f78 , C0 );
buf ( R_f3d_11634798 , n72259 );
buf ( R_155c_156adf78 , n72260 );
buf ( R_782_15ffd168 , C0 );
buf ( R_da1_14b290f8 , n72303 );
buf ( R_13c0_117f6b78 , n72304 );
buf ( R_19df_117eb318 , n72305 );
buf ( R_1719_13c1f8f8 , n72322 );
buf ( R_10fa_13decd38 , C0 );
buf ( R_adb_17014708 , n72323 );
buf ( R_a88_13cd40f8 , n72324 );
buf ( R_10a7_117eb1d8 , n72325 );
buf ( R_16c6_158880f8 , C0 );
buf ( R_1a32_15818018 , C0 );
buf ( R_1413_13d57ef8 , n72326 );
buf ( R_df4_17013f88 , n72327 );
buf ( R_7d5_15889098 , n72376 );
buf ( R_639_13df0cf8 , n72419 );
buf ( R_605_14b1c3f8 , n72462 );
buf ( R_c24_11632d58 , n72463 );
buf ( R_1243_158151d8 , n72464 );
buf ( R_1862_140b94b8 , C0 );
buf ( R_1896_13c0a598 , C0 );
buf ( R_1277_13c27378 , n72465 );
buf ( R_c58_13dddc38 , n72466 );
buf ( R_15a7_17013448 , n72467 );
buf ( R_1532_156b4ff8 , C0 );
buf ( R_f88_13d225d8 , n72468 );
buf ( R_969_13cce298 , n72490 );
buf ( R_8f4_156b9af8 , n72491 );
buf ( R_f13_13c2b478 , n72492 );
buf ( R_1750_14a13018 , n72493 );
buf ( R_74b_123b9998 , n72494 );
buf ( R_1131_13d21c78 , n72519 );
buf ( R_d6a_13c0c118 , C0 );
buf ( R_b12_1587bb78 , C0 );
buf ( R_1389_13c2a4d8 , n72562 );
buf ( R_19a8_124c5578 , n72563 );
buf ( R_a9e_13de43f8 , C0 );
buf ( R_10bd_1162e6b8 , n72572 );
buf ( R_16dc_14b1f058 , n72573 );
buf ( R_1a1c_13cda138 , n72574 );
buf ( R_13fd_14a0e0b8 , n72617 );
buf ( R_dde_15ffc448 , C0 );
buf ( R_7bf_123bb0b8 , n72618 );
buf ( R_1027_13c277d8 , n72619 );
buf ( R_855_14a117b8 , n72628 );
buf ( R_1493_13bee3d8 , n72629 );
buf ( R_1646_13ccbdb8 , C0 );
buf ( R_a08_15ffa5a8 , n72630 );
buf ( R_e74_123b4678 , n72631 );
buf ( R_12d0_14a11cb8 , n72632 );
buf ( R_1809_13d4f7f8 , n72663 );
buf ( R_5ac_11c6e838 , n72670 );
buf ( R_cb1_13d2c998 , n72713 );
buf ( R_bcb_1007e3d8 , n72714 );
buf ( R_692_1587be98 , C0 );
buf ( R_18ef_13d28758 , n72715 );
buf ( R_11ea_1580f238 , C0 );
buf ( R_991_1007ff58 , n72734 );
buf ( R_eeb_12fbe0d8 , n72735 );
buf ( R_150a_14a0b3b8 , C0 );
buf ( R_15cf_10085958 , n72736 );
buf ( R_fb0_117f5318 , n72737 );
buf ( R_8cc_13bf3338 , n72738 );
buf ( R_ce8_11c6a7d8 , n72739 );
buf ( R_1926_116372b8 , C0 );
buf ( R_11b3_13cd3fb8 , n72740 );
buf ( R_575_15817438 , n72741 );
buf ( R_6c9_13dee318 , n72784 );
buf ( R_1307_15ff2da8 , n72785 );
buf ( R_17d2_156b8978 , C0 );
buf ( R_b94_1587e198 , n72786 );
buf ( R_1810_117f12b8 , n72787 );
buf ( R_12c9_17017868 , n72837 );
buf ( R_5b3_123baa78 , n72838 );
buf ( R_caa_15fedbc8 , C0 );
buf ( R_bd2_1580d9d8 , C0 );
buf ( R_68b_13ddf038 , n72839 );
buf ( R_11f1_13c2a938 , n72871 );
buf ( R_18e8_123bd638 , n72872 );
buf ( R_157e_13dee278 , C0 );
buf ( R_f5f_1162d038 , n72873 );
buf ( R_940_1486f838 , n72874 );
buf ( R_91d_14b1cdf8 , n72902 );
buf ( R_f3c_148682b8 , n72903 );
buf ( R_155b_12fc0158 , n72904 );
buf ( R_14b2_15ff2628 , C0 );
buf ( R_874_123c0298 , n72905 );
buf ( R_1008_1587dc98 , n72906 );
buf ( R_e93_13cd4878 , n72907 );
buf ( R_9e9_123b4498 , n72924 );
buf ( R_1627_156b7578 , n72925 );
buf ( R_cf1_124c34f8 , n72968 );
buf ( R_192f_14a12cf8 , n72969 );
buf ( R_11aa_117e9bf8 , C0 );
buf ( R_56c_140ab598 , n72971 );
buf ( R_6d2_1162ec58 , C0 );
buf ( R_1310_13ddf538 , n72972 );
buf ( R_17c9_11638578 , n73004 );
buf ( R_b8b_13df36d8 , n73005 );
buf ( R_a91_13ccfeb8 , n73046 );
buf ( R_10b0_117ea418 , n73047 );
buf ( R_16cf_11c6b138 , n73048 );
buf ( R_1a29_13d384f8 , n73054 );
buf ( R_140a_140aa5f8 , C0 );
buf ( R_deb_140b71b8 , n73055 );
buf ( R_7cc_13cd94b8 , n73056 );
buf ( R_1a47_100862b8 , n73057 );
buf ( R_a73_123be538 , n73058 );
buf ( R_1428_13dde3b8 , n73059 );
buf ( R_1092_15ff41a8 , C0 );
buf ( R_e09_15887a18 , n73102 );
buf ( R_16b1_13c0c258 , n73126 );
buf ( R_7ea_11c6e518 , C0 );
buf ( R_e66_170138a8 , C0 );
buf ( R_1035_1162a478 , n73145 );
buf ( R_847_14a15a98 , n73146 );
buf ( R_1654_1580fff8 , n73147 );
buf ( R_1485_117f6358 , n73190 );
buf ( R_a16_14b25638 , C0 );
buf ( R_b60_13b97b18 , n73191 );
buf ( R_179e_156b3c98 , C0 );
buf ( R_133b_13ddde18 , n73192 );
buf ( R_6fd_156b8338 , n73235 );
buf ( R_117f_13cd7578 , n73236 );
buf ( R_195a_150e1218 , C0 );
buf ( R_d1c_13d3fd98 , n73237 );
buf ( R_134c_14a11ad8 , n73238 );
buf ( R_b4f_12fbee98 , n73239 );
buf ( R_70e_124c25f8 , C0 );
buf ( R_178d_11638a78 , n73284 );
buf ( R_196b_1580a918 , n73285 );
buf ( R_d2d_13cd54f8 , n73328 );
buf ( R_116e_117ebb38 , C0 );
buf ( R_5e1_14b286f8 , n73371 );
buf ( R_c00_150df558 , n73372 );
buf ( R_18ba_11638bb8 , C0 );
buf ( R_121f_13dfa1b8 , n73373 );
buf ( R_129b_13cd3298 , n73374 );
buf ( R_183e_1587c398 , C0 );
buf ( R_c7c_11c6a558 , n73375 );
buf ( R_65d_13cd74d8 , n73418 );
buf ( R_9b3_13df8138 , n73419 );
buf ( R_8aa_13dd9a98 , C0 );
buf ( R_15f1_156b5d18 , n73435 );
buf ( R_ec9_1587c1b8 , n73491 );
buf ( R_fd2_13c05098 , C0 );
buf ( R_14e8_1700a528 , n73492 );
buf ( R_11dd_14875918 , n73527 );
buf ( R_12dd_14a0e158 , n73553 );
buf ( R_17fc_11635eb8 , n73554 );
buf ( R_59f_14a14c38 , n73560 );
buf ( R_cbe_116357d8 , C0 );
buf ( R_bbe_15881438 , C0 );
buf ( R_18fc_17009bc8 , n73561 );
buf ( R_69f_13d56b98 , n73562 );
buf ( R_1598_13cd92d8 , n73563 );
buf ( R_f79_13bf2e38 , n73579 );
buf ( R_95a_13d37698 , C0 );
buf ( R_903_117ec7b8 , n73580 );
buf ( R_f22_14a13978 , C0 );
buf ( R_1541_15886758 , n73629 );
buf ( R_12e3_17014028 , n73630 );
buf ( R_11d7_1587d5b8 , n73631 );
buf ( R_cc4_13bead78 , n73632 );
buf ( R_599_150dcf38 , n73639 );
buf ( R_17f6_117f1498 , C0 );
buf ( R_1902_14b1af58 , C0 );
buf ( R_6a5_13df56b8 , n73682 );
buf ( R_bb8_124c3b38 , n73683 );
buf ( R_14bf_150dd938 , n73684 );
buf ( R_881_150db278 , n73690 );
buf ( R_ffb_15813ab8 , n73691 );
buf ( R_ea0_13b95778 , n73692 );
buf ( R_9dc_15ff19a8 , n73693 );
buf ( R_161a_14b23bf8 , C0 );
buf ( R_1454_123b4538 , n73694 );
buf ( R_e35_11c70098 , n73737 );
buf ( R_a47_1486f3d8 , n73738 );
buf ( R_816_13c06cb8 , C0 );
buf ( R_1066_13bee838 , C0 );
buf ( R_1685_15ff1d68 , n73766 );
buf ( R_8b0_15813c98 , n73767 );
buf ( R_9ad_13de0bb8 , n73791 );
buf ( R_ecf_13c26798 , n73792 );
buf ( R_15eb_140b6498 , n73793 );
buf ( R_14ee_13d5a298 , C0 );
buf ( R_fcc_150e33d8 , n73794 );
buf ( R_101c_11c6ce98 , n73795 );
buf ( R_860_14a17b18 , n73796 );
buf ( R_149e_11c6edd8 , C0 );
buf ( R_163b_13c04b98 , n73797 );
buf ( R_9fd_117ebf98 , n73822 );
buf ( R_e7f_117f6038 , n73823 );
buf ( R_604_15811718 , n73824 );
buf ( R_c23_123bfc58 , n73825 );
buf ( R_1242_10080c78 , C0 );
buf ( R_1861_12fbf7f8 , n73859 );
buf ( R_1897_13d3d1d8 , n73860 );
buf ( R_1278_117f4f58 , n73861 );
buf ( R_c59_116304b8 , n73876 );
buf ( R_63a_13c0a278 , C0 );
buf ( R_b59_15feff68 , n73911 );
buf ( R_1342_148716d8 , C0 );
buf ( R_1797_117f7e38 , n73912 );
buf ( R_704_123b2ff8 , n73913 );
buf ( R_1961_1162de98 , n73923 );
buf ( R_1178_13cd24d8 , n73924 );
buf ( R_d23_11c68618 , n73925 );
buf ( R_157f_13b8ce98 , n73926 );
buf ( R_f60_140af9b8 , n73927 );
buf ( R_941_13df8b38 , n73951 );
buf ( R_91c_13df6d38 , n73952 );
buf ( R_f3b_15810c78 , n73953 );
buf ( R_155a_15882338 , C0 );
buf ( R_e5c_117f6df8 , n73954 );
buf ( R_165e_117edf78 , C0 );
buf ( R_83d_13c24ad8 , n74010 );
buf ( R_a20_15883738 , n74011 );
buf ( R_147b_1700f5c8 , n74012 );
buf ( R_103f_123b9ad8 , n74013 );
buf ( R_5ef_1162a018 , n74014 );
buf ( R_c0e_158802b8 , C0 );
buf ( R_122d_150e4eb8 , n74039 );
buf ( R_184c_14a19418 , n74040 );
buf ( R_18ac_117f13f8 , n74041 );
buf ( R_128d_123b2af8 , n74092 );
buf ( R_c6e_15ff6408 , C0 );
buf ( R_64f_13bf1ad8 , n74093 );
buf ( R_9a0_13dd6078 , n74094 );
buf ( R_edc_123be678 , n74095 );
buf ( R_15de_15ff2268 , C0 );
buf ( R_14fb_13c29038 , n74096 );
buf ( R_fbf_150e4f58 , n74097 );
buf ( R_8bd_13cd5ef8 , n74114 );
buf ( R_1998_14b279d8 , n74115 );
buf ( R_1141_1580bbd8 , n74145 );
buf ( R_73b_14a15638 , n74146 );
buf ( R_b22_13cce8d8 , C0 );
buf ( R_d5a_13bf6178 , C0 );
buf ( R_1379_123bdbd8 , n74189 );
buf ( R_1760_117f7f78 , n74190 );
buf ( R_1981_1587b7b8 , n74202 );
buf ( R_b39_15ffae68 , n74217 );
buf ( R_724_117ec8f8 , n74218 );
buf ( R_1777_1587ccf8 , n74219 );
buf ( R_d43_13beedd8 , n74220 );
buf ( R_1362_150dfcd8 , C0 );
buf ( R_1158_13bf0f98 , n74221 );
buf ( R_770_15888058 , n74222 );
buf ( R_d8f_11629f78 , n74223 );
buf ( R_13ae_13bf3478 , C0 );
buf ( R_172b_156b88d8 , n74224 );
buf ( R_19cd_117ed578 , n74235 );
buf ( R_110c_15810458 , n74236 );
buf ( R_aed_14a0e298 , n74267 );
buf ( R_1449_14b26678 , n74310 );
buf ( R_e2a_13c29858 , C0 );
buf ( R_a52_140af378 , C0 );
buf ( R_80b_158154f8 , n74311 );
buf ( R_1071_123c1378 , n74328 );
buf ( R_1a68_117ed618 , n74329 );
buf ( R_1690_13c216f8 , n74330 );
buf ( R_ef3_13cd06d8 , n74331 );
buf ( R_989_13c068f8 , n74353 );
buf ( R_1512_1162e078 , C0 );
buf ( R_15c7_13d3c4b8 , n74354 );
buf ( R_8d4_123c1738 , n74355 );
buf ( R_fa8_123be858 , n74356 );
buf ( R_1984_1162e438 , n74357 );
buf ( R_727_1700aca8 , n74358 );
buf ( R_b36_123bb338 , C0 );
buf ( R_d46_13cd3338 , C0 );
buf ( R_1774_13c26c98 , n74359 );
buf ( R_1365_150db818 , n74402 );
buf ( R_1155_17012868 , n74417 );
buf ( R_b3c_13cd4eb8 , n74418 );
buf ( R_721_156b7d98 , n74461 );
buf ( R_197e_13d5c8b8 , C0 );
buf ( R_177a_123c1418 , C0 );
buf ( R_d40_11635af8 , n74462 );
buf ( R_115b_123bf2f8 , n74463 );
buf ( R_135f_11c6da78 , n74464 );
buf ( R_894_1587b2b8 , n74465 );
buf ( R_1607_123bd138 , n74466 );
buf ( R_eb3_123b5cf8 , n74467 );
buf ( R_fe8_15816678 , n74468 );
buf ( R_14d2_11636e58 , C0 );
buf ( R_9c9_13cce798 , n74486 );
buf ( R_160c_117f74d8 , n74487 );
buf ( R_88f_13c0d338 , n74488 );
buf ( R_fed_12fc1198 , n74505 );
buf ( R_eae_13cd1d58 , C0 );
buf ( R_9ce_1162c6d8 , C0 );
buf ( R_14cd_10081178 , n74548 );
buf ( R_dac_14a109f8 , n74549 );
buf ( R_13cb_13ccf0f8 , n74550 );
buf ( R_19ea_11629b18 , C0 );
buf ( R_170e_1580e338 , C0 );
buf ( R_10ef_14a199b8 , n74551 );
buf ( R_ad0_123b65b8 , n74552 );
buf ( R_78d_15817618 , n74595 );
buf ( R_999_1008a138 , n74613 );
buf ( R_ee3_158135b8 , n74614 );
buf ( R_1502_117ea238 , C0 );
buf ( R_15d7_11c6ab98 , n74615 );
buf ( R_fb8_156b7bb8 , n74616 );
buf ( R_8c4_117f8018 , n74617 );
buf ( R_efc_12fc14b8 , n74618 );
buf ( R_980_13d2b9f8 , n74619 );
buf ( R_151b_14a153b8 , n74620 );
buf ( R_15be_11629bb8 , C0 );
buf ( R_8dd_13d1dcb8 , n74636 );
buf ( R_f9f_13bf1858 , n74637 );
buf ( R_8a4_13cd4418 , n74638 );
buf ( R_15f7_117ea878 , n74639 );
buf ( R_ec3_14a15e58 , n74640 );
buf ( R_fd8_117f1718 , n74641 );
buf ( R_14e2_13ddc478 , C0 );
buf ( R_9b9_1008a458 , n74665 );
buf ( R_1580_123b3958 , n74666 );
buf ( R_f61_14867318 , n74682 );
buf ( R_942_140b3a18 , C0 );
buf ( R_91b_156b0d18 , n74683 );
buf ( R_f3a_1007f4b8 , C0 );
buf ( R_1559_13c234f8 , n74732 );
buf ( R_1441_13ded378 , n74775 );
buf ( R_a5a_13c097d8 , C0 );
buf ( R_e22_117eccb8 , C0 );
buf ( R_1079_13beb6d8 , n74793 );
buf ( R_803_140b8158 , n74794 );
buf ( R_1698_15811998 , n74795 );
buf ( R_1a60_14b1b778 , n74796 );
buf ( R_1987_140b7cf8 , n74797 );
buf ( R_72a_158127f8 , C0 );
buf ( R_b33_13d2aaf8 , n74798 );
buf ( R_d49_15811678 , n74841 );
buf ( R_1771_17009c68 , n74869 );
buf ( R_1368_1587e9b8 , n74870 );
buf ( R_1152_13c0bd58 , C0 );
buf ( R_5d5_123be038 , n74913 );
buf ( R_18c6_13d3a1b8 , C0 );
buf ( R_bf4_1587cb18 , n74914 );
buf ( R_12a7_15817cf8 , n74915 );
buf ( R_1213_140ad078 , n74916 );
buf ( R_c88_17017cc8 , n74917 );
buf ( R_1832_123bc2d8 , C0 );
buf ( R_669_116322b8 , n74960 );
buf ( R_769_150da558 , n75003 );
buf ( R_d88_117f22f8 , n75004 );
buf ( R_1732_123b2558 , C0 );
buf ( R_13a7_13c08ab8 , n75005 );
buf ( R_1113_123c1e18 , n75006 );
buf ( R_19c6_13cd18f8 , C0 );
buf ( R_af4_1580feb8 , n75007 );
buf ( R_b3f_13c22198 , n75008 );
buf ( R_71e_140aec98 , C0 );
buf ( R_197b_123c14b8 , n75009 );
buf ( R_177d_17012728 , n75037 );
buf ( R_d3d_13c053b8 , n75080 );
buf ( R_115e_15885c18 , C0 );
buf ( R_135c_13cda3b8 , n75081 );
buf ( R_12d7_13cd2578 , n75082 );
buf ( R_1802_13d3fbb8 , C0 );
buf ( R_5a5_13d375f8 , n75089 );
buf ( R_cb8_11c6c218 , n75090 );
buf ( R_bc4_14b2a138 , n75091 );
buf ( R_699_15888ff8 , n75134 );
buf ( R_18f6_124c27d8 , C0 );
buf ( R_11e3_1162fa18 , n75135 );
buf ( R_b67_13cd4f58 , n75136 );
buf ( R_17a5_116334d8 , n75182 );
buf ( R_1334_13cd5598 , n75183 );
buf ( R_6f6_117f1858 , C0 );
buf ( R_1186_11635d78 , C0 );
buf ( R_1953_117eb6d8 , n75184 );
buf ( R_d15_123b5578 , n75227 );
buf ( R_603_13ddbe38 , n75228 );
buf ( R_c22_117f71b8 , C0 );
buf ( R_1241_1162a5b8 , n75260 );
buf ( R_1860_13ccdf78 , n75261 );
buf ( R_1898_11c6bb38 , n75262 );
buf ( R_1279_15887478 , n75313 );
buf ( R_c5a_14a16538 , C0 );
buf ( R_63b_15883cd8 , n75314 );
buf ( R_10bb_1587d8d8 , n75315 );
buf ( R_16da_124c3db8 , C0 );
buf ( R_1a1e_11c6ed38 , C0 );
buf ( R_13ff_17012c28 , n75316 );
buf ( R_de0_13d3abb8 , n75317 );
buf ( R_7c1_156b3bf8 , n75360 );
buf ( R_a9c_1162e4d8 , n75361 );
buf ( R_18d0_117f1358 , n75362 );
buf ( R_5cb_12fc0d38 , n75363 );
buf ( R_12b1_124c38b8 , n75413 );
buf ( R_bea_13ccb098 , C0 );
buf ( R_c92_150e3838 , C0 );
buf ( R_1209_14a0aa58 , n75445 );
buf ( R_673_14a13fb8 , n75446 );
buf ( R_1828_1580ab98 , n75447 );
buf ( R_14b6_1587d1f8 , C0 );
buf ( R_878_13c100d8 , n75448 );
buf ( R_1004_156ab318 , n75449 );
buf ( R_e97_14866918 , n75450 );
buf ( R_9e5_1587d6f8 , n75468 );
buf ( R_1623_13b96178 , n75469 );
buf ( R_11d1_1162f6f8 , n75490 );
buf ( R_cca_117eebf8 , C0 );
buf ( R_593_117ee0b8 , n75497 );
buf ( R_17f0_100833d8 , n75498 );
buf ( R_1908_1162f5b8 , n75499 );
buf ( R_6ab_13ccbe58 , n75500 );
buf ( R_bb2_15810278 , C0 );
buf ( R_12e9_13d26818 , n75543 );
buf ( R_f89_13d51738 , n75563 );
buf ( R_96a_1587c258 , C0 );
buf ( R_8f3_10082b18 , n75564 );
buf ( R_f12_1162b2d8 , C0 );
buf ( R_15a8_14b25db8 , n75565 );
buf ( R_1531_13c0ac78 , n75614 );
buf ( R_12c2_13d4e2b8 , C0 );
buf ( R_5ba_13b94d78 , C0 );
buf ( R_ca3_13ddaa38 , n75615 );
buf ( R_bd9_13d54398 , n75669 );
buf ( R_684_117f5a98 , n75670 );
buf ( R_11f8_13bf1538 , n75671 );
buf ( R_18e1_17010388 , n75723 );
buf ( R_1817_1580f9b8 , n75724 );
buf ( R_a7f_117ebc78 , n75725 );
buf ( R_1a3b_13d275d8 , n75726 );
buf ( R_109e_14a11538 , C0 );
buf ( R_16bd_117eb9f8 , n75750 );
buf ( R_141c_123b3f98 , n75751 );
buf ( R_dfd_1700cf08 , n75794 );
buf ( R_7de_15881ed8 , C0 );
buf ( R_f95_13d51058 , n75800 );
buf ( R_1525_140b5598 , n75856 );
buf ( R_976_140b2f78 , C0 );
buf ( R_8e7_13dd8ff8 , n75857 );
buf ( R_15b4_13dee598 , n75858 );
buf ( R_f06_14b29238 , C0 );
buf ( R_899_13d5a8d8 , n75874 );
buf ( R_1602_13c28ef8 , C0 );
buf ( R_eb8_13c1c0b8 , n75875 );
buf ( R_fe3_13ccb598 , n75876 );
buf ( R_14d7_14a0fb98 , n75877 );
buf ( R_9c4_123c1a58 , n75878 );
buf ( R_1599_13bf40f8 , n75884 );
buf ( R_f7a_13d510f8 , C0 );
buf ( R_95b_15813838 , n75885 );
buf ( R_902_14a0aff8 , C0 );
buf ( R_f21_15812398 , n75901 );
buf ( R_1540_14871458 , n75902 );
buf ( R_1321_156b1038 , n75949 );
buf ( R_1199_13cd3bf8 , n75980 );
buf ( R_6e3_140b27f8 , n75981 );
buf ( R_55b_13d54f78 , n75982 );
buf ( R_1940_117ed758 , n75983 );
buf ( R_17b8_14b1ca38 , n75984 );
buf ( R_d02_14b21998 , C0 );
buf ( R_b7a_140b8298 , C0 );
buf ( R_ed5_123b27d8 , n76033 );
buf ( R_15e5_13d3e0d8 , n76049 );
buf ( R_14f4_1580cad8 , n76050 );
buf ( R_fc6_117f2078 , C0 );
buf ( R_8b6_12fbe7b8 , C0 );
buf ( R_9a7_13dd6118 , n76051 );
buf ( R_d96_13c23778 , C0 );
buf ( R_13b5_124c31d8 , n76094 );
buf ( R_19d4_123b6798 , n76095 );
buf ( R_1724_117edcf8 , n76096 );
buf ( R_1105_158130b8 , n76147 );
buf ( R_ae6_14873e38 , C0 );
buf ( R_777_17012228 , n76148 );
buf ( R_1581_10080458 , n76260 );
buf ( R_f62_13ccaff8 , C0 );
buf ( R_943_156b21b8 , n76261 );
buf ( R_91a_13d23e38 , C0 );
buf ( R_f39_117f5778 , n76277 );
buf ( R_1558_15ffb2c8 , n76278 );
buf ( R_88a_15880c18 , C0 );
buf ( R_ff2_13d42638 , C0 );
buf ( R_ea9_15810ef8 , n76334 );
buf ( R_9d3_12fc1e18 , n76335 );
buf ( R_14c8_13d50d38 , n76336 );
buf ( R_1611_13df2b98 , n76352 );
buf ( R_5c2_150db138 , C0 );
buf ( R_12ba_158138d8 , C0 );
buf ( R_be1_10082898 , n76403 );
buf ( R_c9b_13b977f8 , n76404 );
buf ( R_1200_13d3d778 , n76405 );
buf ( R_67c_13dec978 , n76406 );
buf ( R_181f_156b4558 , n76407 );
buf ( R_18d9_117f3e78 , n76433 );
buf ( R_1743_15ff3488 , n76434 );
buf ( R_758_13cd0ef8 , n76435 );
buf ( R_1124_14a17d98 , n76436 );
buf ( R_d77_14a0ca38 , n76437 );
buf ( R_1396_156ace98 , C0 );
buf ( R_b05_13d37d78 , n76451 );
buf ( R_19b5_13cd3c98 , n76462 );
buf ( R_d9f_1580b818 , n76463 );
buf ( R_13be_156af5f8 , C0 );
buf ( R_19dd_13d56238 , n76469 );
buf ( R_171b_14a0ac38 , n76470 );
buf ( R_10fc_13d52c78 , n76471 );
buf ( R_add_17015ce8 , n76486 );
buf ( R_780_13cd31f8 , n76487 );
buf ( R_198a_12fc1af8 , C0 );
buf ( R_72d_13d467d8 , n76530 );
buf ( R_b30_156ac358 , n76531 );
buf ( R_d4c_11633d98 , n76532 );
buf ( R_176e_12fbe678 , C0 );
buf ( R_136b_15810638 , n76533 );
buf ( R_114f_123ba1b8 , n76534 );
buf ( R_119d_123ba578 , n76548 );
buf ( R_55f_13cce658 , n76550 );
buf ( R_6df_13bf5ef8 , n76551 );
buf ( R_131d_14a11c18 , n76594 );
buf ( R_17bc_15886d98 , n76595 );
buf ( R_b7e_123b7eb8 , C0 );
buf ( R_cfe_123b7418 , C0 );
buf ( R_193c_123b6298 , n76596 );
buf ( R_b42_116296b8 , C0 );
buf ( R_71b_13cd8fb8 , n76597 );
buf ( R_1978_1587e698 , n76598 );
buf ( R_1780_1587b718 , n76599 );
buf ( R_d3a_117f6678 , C0 );
buf ( R_1161_13beb3b8 , n76614 );
buf ( R_1359_11c6d9d8 , n76657 );
buf ( R_1325_156ac178 , n76700 );
buf ( R_6e7_15882fb8 , n76701 );
buf ( R_557_15885f38 , n76703 );
buf ( R_1195_116363b8 , n76734 );
buf ( R_1944_124c2918 , n76735 );
buf ( R_d06_13dde818 , C0 );
buf ( R_b76_13d41b98 , C0 );
buf ( R_17b4_13d29ab8 , n76736 );
buf ( R_1020_117ed258 , n76737 );
buf ( R_85c_1580fc38 , n76738 );
buf ( R_149a_13bf0ef8 , C0 );
buf ( R_163f_13de4218 , n76739 );
buf ( R_a01_156b1498 , n76764 );
buf ( R_e7b_1486b738 , n76765 );
buf ( R_11c1_123b5618 , n76781 );
buf ( R_cda_156b9878 , C0 );
buf ( R_1918_15880f38 , n76782 );
buf ( R_583_13cccb78 , n76783 );
buf ( R_17e0_14a15d18 , n76784 );
buf ( R_6bb_117f2398 , n76785 );
buf ( R_ba2_14a0e5b8 , C0 );
buf ( R_12f9_13d5c9f8 , n76828 );
buf ( R_5ee_12fc0c98 , C0 );
buf ( R_c0d_13b93fb8 , n76879 );
buf ( R_122c_14b217b8 , n76880 );
buf ( R_18ad_13cd6358 , n76912 );
buf ( R_184b_1486d3f8 , n76913 );
buf ( R_128e_13b91a38 , C0 );
buf ( R_c6f_150e83d8 , n76914 );
buf ( R_650_116346f8 , n76915 );
buf ( R_5e0_13df04d8 , n76916 );
buf ( R_bff_123b92b8 , n76917 );
buf ( R_18bb_11c6f698 , n76918 );
buf ( R_121e_14b1d438 , C0 );
buf ( R_129c_1007ebf8 , n76919 );
buf ( R_183d_15882e78 , n76934 );
buf ( R_c7d_13c108f8 , n76977 );
buf ( R_65e_13d43998 , C0 );
buf ( R_75d_156ad118 , n77020 );
buf ( R_173e_148678b8 , C0 );
buf ( R_d7c_123be998 , n77021 );
buf ( R_111f_14a110d8 , n77022 );
buf ( R_139b_156b35b8 , n77023 );
buf ( R_b00_13ccf558 , n77024 );
buf ( R_19ba_17014d48 , C0 );
buf ( R_a78_13cd1cb8 , n77025 );
buf ( R_1a42_15817118 , C0 );
buf ( R_1097_13d240b8 , n77026 );
buf ( R_1423_13c05a98 , n77027 );
buf ( R_16b6_140aab98 , C0 );
buf ( R_e04_156b17b8 , n77028 );
buf ( R_7e5_14b1e798 , n77077 );
buf ( R_746_170166e8 , C0 );
buf ( R_1136_13d56558 , C0 );
buf ( R_d65_1008bb78 , n77120 );
buf ( R_b17_123bcc38 , n77121 );
buf ( R_1384_140b3298 , n77122 );
buf ( R_19a3_117eaa58 , n77123 );
buf ( R_1755_10087258 , n77172 );
buf ( R_c21_1700d4a8 , n77222 );
buf ( R_1240_11630238 , n77223 );
buf ( R_185f_13bf7118 , n77224 );
buf ( R_1899_156b1fd8 , n77249 );
buf ( R_127a_14b28298 , C0 );
buf ( R_c5b_13d26278 , n77250 );
buf ( R_63c_1587b538 , n77251 );
buf ( R_602_156afff8 , C0 );
buf ( R_753_116336b8 , n77252 );
buf ( R_1129_13ccc3f8 , n77293 );
buf ( R_d72_13b95e58 , C0 );
buf ( R_b0a_156ad438 , C0 );
buf ( R_1391_15886578 , n77336 );
buf ( R_19b0_17014a28 , n77337 );
buf ( R_1748_117eeab8 , n77338 );
buf ( R_e32_13c05c78 , C0 );
buf ( R_a4a_117e8bb8 , C0 );
buf ( R_813_11631318 , n77339 );
buf ( R_1069_116369f8 , n77356 );
buf ( R_1688_156b6a38 , n77357 );
buf ( R_1451_150e6b78 , n77400 );
buf ( R_cdf_150dfa58 , n77401 );
buf ( R_11bc_11c6a9b8 , n77402 );
buf ( R_191d_13c10678 , n77453 );
buf ( R_57e_1162f338 , n77454 );
buf ( R_6c0_13b98c98 , n77455 );
buf ( R_17db_117f6858 , n77456 );
buf ( R_12fe_116291b8 , C0 );
buf ( R_b9d_14872678 , n77488 );
buf ( R_1349_13d26db8 , n77531 );
buf ( R_b52_1162a978 , C0 );
buf ( R_1790_117e9798 , n77532 );
buf ( R_70b_17018808 , n77533 );
buf ( R_1968_13bf0318 , n77534 );
buf ( R_d2a_15fef568 , C0 );
buf ( R_1171_117f5278 , n77565 );
buf ( R_192b_11633cf8 , n77566 );
buf ( R_11ae_123bc238 , C0 );
buf ( R_570_117ec218 , n77567 );
buf ( R_6ce_13dee1d8 , C0 );
buf ( R_130c_15ff67c8 , n77568 );
buf ( R_17cd_13b91858 , n77600 );
buf ( R_b8f_14b25b38 , n77601 );
buf ( R_ced_14a0a558 , n77644 );
buf ( R_1582_150e7ed8 , C0 );
buf ( R_f63_13cca7d8 , n77645 );
buf ( R_944_13d1fab8 , n77646 );
buf ( R_919_123bdf98 , n77674 );
buf ( R_f38_13d26958 , n77675 );
buf ( R_1557_14a16c18 , n77676 );
buf ( R_10ae_123b9358 , C0 );
buf ( R_16cd_117eee78 , n77695 );
buf ( R_1a2b_140accb8 , n77696 );
buf ( R_140c_11c6f058 , n77697 );
buf ( R_ded_14a14738 , n77740 );
buf ( R_7ce_13d45d38 , C0 );
buf ( R_a8f_17014de8 , n77741 );
buf ( R_10a5_13d564b8 , n77768 );
buf ( R_16c4_1580f878 , n77769 );
buf ( R_1a34_14a19558 , n77770 );
buf ( R_1415_158165d8 , n77813 );
buf ( R_df6_156b2bb8 , C0 );
buf ( R_7d7_13c29998 , n77814 );
buf ( R_a86_123bc0f8 , C0 );
buf ( R_165b_13de0898 , n77815 );
buf ( R_840_156b26b8 , n77816 );
buf ( R_a1d_14a15778 , n77843 );
buf ( R_147e_11638078 , C0 );
buf ( R_103c_140b0ef8 , n77844 );
buf ( R_e5f_150e3d38 , n77845 );
buf ( R_11c6_13def038 , C0 );
buf ( R_cd5_13cd09f8 , n77888 );
buf ( R_588_13de09d8 , n77889 );
buf ( R_1913_13beef18 , n77890 );
buf ( R_17e5_150de518 , n77905 );
buf ( R_6b6_13d519b8 , C0 );
buf ( R_ba7_13d2ca38 , n77906 );
buf ( R_12f4_11c6ca38 , n77907 );
buf ( R_19e8_15888e18 , n77908 );
buf ( R_1710_13bf6718 , n77909 );
buf ( R_10f1_124c52f8 , n77937 );
buf ( R_ad2_156b8658 , C0 );
buf ( R_78b_1162ddf8 , n77938 );
buf ( R_daa_1008ced8 , C0 );
buf ( R_13c9_13de18d8 , n77981 );
buf ( R_11a1_117e91f8 , n78012 );
buf ( R_563_13d1ea78 , n78013 );
buf ( R_6db_13dd91d8 , n78014 );
buf ( R_1319_117f10d8 , n78057 );
buf ( R_17c0_15ff4888 , n78058 );
buf ( R_b82_13beff58 , C0 );
buf ( R_cfa_14b21ad8 , C0 );
buf ( R_1938_13df6ab8 , n78059 );
buf ( R_82a_14a0cfd8 , C0 );
buf ( R_a33_11c70278 , n78060 );
buf ( R_1468_158803f8 , n78061 );
buf ( R_1052_117f42d8 , C0 );
buf ( R_1671_13dd6898 , n78078 );
buf ( R_e49_15ff8f28 , n78121 );
buf ( R_1329_14a16ad8 , n78164 );
buf ( R_6eb_13d45b58 , n78165 );
buf ( R_1191_15881618 , n78179 );
buf ( R_1948_13c26a18 , n78180 );
buf ( R_d0a_158820b8 , C0 );
buf ( R_b72_13c103f8 , C0 );
buf ( R_17b0_13decf18 , n78181 );
buf ( R_a36_13b92438 , C0 );
buf ( R_827_123b8f98 , n78182 );
buf ( R_1055_11635738 , n78208 );
buf ( R_1465_14a18ab8 , n78251 );
buf ( R_1674_11636c78 , n78252 );
buf ( R_e46_15884098 , C0 );
buf ( R_851_11635238 , n78261 );
buf ( R_148f_13df4358 , n78262 );
buf ( R_164a_13c1e318 , C0 );
buf ( R_a0c_100899b8 , n78263 );
buf ( R_e70_117ec538 , n78264 );
buf ( R_102b_13d38d18 , n78265 );
buf ( R_198d_156b4378 , n78276 );
buf ( R_730_123bb518 , n78277 );
buf ( R_b2d_124c29b8 , n78292 );
buf ( R_d4f_13cd15d8 , n78293 );
buf ( R_176b_150e5bd8 , n78294 );
buf ( R_136e_15ff6b88 , C0 );
buf ( R_114c_140b06d8 , n78295 );
buf ( R_16f5_13d39b78 , n78318 );
buf ( R_1a03_14b23338 , n78319 );
buf ( R_10d6_150df4b8 , C0 );
buf ( R_13e4_13cd99b8 , n78320 );
buf ( R_ab7_1700b748 , n78321 );
buf ( R_dc5_15ff3f28 , n78368 );
buf ( R_7a6_150dad78 , C0 );
buf ( R_1a05_1162d498 , n78374 );
buf ( R_13e6_1486e578 , C0 );
buf ( R_dc7_13cd2398 , n78375 );
buf ( R_16f3_10088bf8 , n78376 );
buf ( R_7a8_13beac38 , n78377 );
buf ( R_10d4_13d1de98 , n78378 );
buf ( R_ab5_13df25f8 , n78415 );
buf ( R_82d_13c24b78 , n78471 );
buf ( R_a30_117ef9b8 , n78472 );
buf ( R_146b_150da9b8 , n78473 );
buf ( R_104f_170118c8 , n78474 );
buf ( R_e4c_13ddfd58 , n78475 );
buf ( R_166e_123be3f8 , C0 );
buf ( R_73e_15883878 , C0 );
buf ( R_b1f_11631098 , n78476 );
buf ( R_d5d_11636778 , n78519 );
buf ( R_137c_11634e78 , n78520 );
buf ( R_175d_13df13d8 , n78554 );
buf ( R_199b_150dc8f8 , n78555 );
buf ( R_113e_10081ad8 , C0 );
buf ( R_b45_13cce978 , n78576 );
buf ( R_718_123b4fd8 , n78577 );
buf ( R_1975_13deedb8 , n78587 );
buf ( R_1783_15817e38 , n78588 );
buf ( R_d37_13d26d18 , n78589 );
buf ( R_1164_13df29b8 , n78590 );
buf ( R_1356_15884958 , C0 );
buf ( R_16f7_140b9558 , n78591 );
buf ( R_10d8_13d55158 , n78592 );
buf ( R_ab9_14a16358 , n78626 );
buf ( R_1a01_14a0bf98 , n78632 );
buf ( R_7a4_13cca698 , n78633 );
buf ( R_13e2_13d50338 , C0 );
buf ( R_dc3_13d5b918 , n78634 );
buf ( R_1509_13c080b8 , n78683 );
buf ( R_15d0_13d5d7b8 , n78684 );
buf ( R_fb1_17011fa8 , n78707 );
buf ( R_8cb_1162afb8 , n78708 );
buf ( R_992_158117b8 , C0 );
buf ( R_eea_158843b8 , C0 );
buf ( R_1a07_15817f78 , n78709 );
buf ( R_13e8_13d57458 , n78710 );
buf ( R_dc9_13dedb98 , n78753 );
buf ( R_7aa_14a113f8 , C0 );
buf ( R_ab3_13ccea18 , n78754 );
buf ( R_16f1_13c2b298 , n78778 );
buf ( R_10d2_14a0f4b8 , C0 );
buf ( R_84a_1700eee8 , C0 );
buf ( R_1651_100849b8 , n78801 );
buf ( R_1488_15811858 , n78802 );
buf ( R_a13_117f7ed8 , n78803 );
buf ( R_e69_14b24ff8 , n78852 );
buf ( R_1032_15884638 , C0 );
buf ( R_1434_15884a98 , n78853 );
buf ( R_a67_1587c9d8 , n78854 );
buf ( R_e15_117f6538 , n78897 );
buf ( R_1086_158844f8 , C0 );
buf ( R_16a5_1587d018 , n78920 );
buf ( R_7f6_14a10318 , C0 );
buf ( R_1a53_11c70b38 , n78921 );
buf ( R_f7b_13c24f38 , n78922 );
buf ( R_95c_13b8ad78 , n78923 );
buf ( R_901_15ff0dc8 , n78929 );
buf ( R_f20_11633078 , n78930 );
buf ( R_153f_140abef8 , n78931 );
buf ( R_159a_13d58d58 , C0 );
buf ( R_1a20_117f5638 , n78932 );
buf ( R_1401_14a19918 , n78975 );
buf ( R_de2_123bef38 , C0 );
buf ( R_7c3_14a0f058 , n78976 );
buf ( R_a9a_15816f38 , C0 );
buf ( R_10b9_15ff6908 , n78982 );
buf ( R_16d8_14b209f8 , n78983 );
buf ( R_1583_13b8ba98 , n78984 );
buf ( R_f64_123b9718 , n78985 );
buf ( R_945_123bcaf8 , n79002 );
buf ( R_918_13c20ed8 , n79003 );
buf ( R_f37_158875b8 , n79004 );
buf ( R_1556_140b5db8 , C0 );
buf ( R_a39_17016d28 , n79043 );
buf ( R_824_140b4b98 , n79044 );
buf ( R_1058_13b8c7b8 , n79045 );
buf ( R_1462_13d228f8 , C0 );
buf ( R_1677_1008aef8 , n79046 );
buf ( R_e43_140ab8b8 , n79047 );
buf ( R_123f_12fc2458 , n79048 );
buf ( R_185e_100815d8 , C0 );
buf ( R_189a_15ff14a8 , C0 );
buf ( R_127b_13de1a18 , n79049 );
buf ( R_c5c_140b8518 , n79050 );
buf ( R_63d_13df0438 , n79093 );
buf ( R_601_14a12c58 , n79136 );
buf ( R_c20_1486b7d8 , n79137 );
buf ( R_15fd_156b4c38 , n79153 );
buf ( R_ebd_117f1ad8 , n79202 );
buf ( R_fde_13d429f8 , C0 );
buf ( R_14dc_13ddc5b8 , n79203 );
buf ( R_9bf_15ff2128 , n79204 );
buf ( R_89e_123bbdd8 , C0 );
buf ( R_16f9_13cd6218 , n79228 );
buf ( R_10da_14a0d4d8 , C0 );
buf ( R_abb_14b262b8 , n79229 );
buf ( R_7a2_13de1fb8 , C0 );
buf ( R_dc1_13c211f8 , n79272 );
buf ( R_13e0_1486e4d8 , n79273 );
buf ( R_19ff_123b42b8 , n79274 );
buf ( R_1739_15ff78a8 , n79293 );
buf ( R_d81_140ad4d8 , n79336 );
buf ( R_111a_13d42ef8 , C0 );
buf ( R_13a0_117f2bb8 , n79337 );
buf ( R_afb_13bf4af8 , n79338 );
buf ( R_19bf_117f5e58 , n79339 );
buf ( R_762_156b33d8 , C0 );
buf ( R_1a09_1162d358 , n79345 );
buf ( R_13ea_1580dc58 , C0 );
buf ( R_dcb_1162f798 , n79346 );
buf ( R_7ac_13c08838 , n79347 );
buf ( R_ab1_150e1b78 , n79372 );
buf ( R_10d0_150e7938 , n79373 );
buf ( R_16ef_14a136f8 , n79374 );
buf ( R_a6c_123b7378 , n79375 );
buf ( R_142f_117f79d8 , n79376 );
buf ( R_108b_156b83d8 , n79377 );
buf ( R_e10_14a0b4f8 , n79378 );
buf ( R_16aa_150e47d8 , C0 );
buf ( R_7f1_123bc378 , n79427 );
buf ( R_1a4e_123b60b8 , C0 );
buf ( R_5b2_1486f018 , n79428 );
buf ( R_cab_15fee028 , n79429 );
buf ( R_bd1_1587dfb8 , n79481 );
buf ( R_68c_123c1b98 , n79482 );
buf ( R_11f0_13cd3a18 , n79483 );
buf ( R_18e9_13b98a18 , n79535 );
buf ( R_180f_13c1cbf8 , n79536 );
buf ( R_12ca_14a13dd8 , C0 );
buf ( R_1000_13d4e858 , n79537 );
buf ( R_e9b_13cd5f98 , n79538 );
buf ( R_9e1_13bea878 , n79555 );
buf ( R_161f_10080098 , n79556 );
buf ( R_14ba_1580ba98 , C0 );
buf ( R_87c_13dee6d8 , n79557 );
buf ( R_830_1008cc58 , n79558 );
buf ( R_a2d_13d43f38 , n79570 );
buf ( R_146e_17010ba8 , C0 );
buf ( R_104c_13d1f658 , n79571 );
buf ( R_e4f_13ccef18 , n79572 );
buf ( R_166b_116345b8 , n79573 );
buf ( R_ff7_13c0cf78 , n79574 );
buf ( R_ea4_117ea738 , n79575 );
buf ( R_9d8_156b6ad8 , n79576 );
buf ( R_1616_17009da8 , C0 );
buf ( R_14c3_116384d8 , n79577 );
buf ( R_885_13de02f8 , n79583 );
buf ( R_11b7_11c6de38 , n79584 );
buf ( R_1922_13c26018 , C0 );
buf ( R_579_13d5d358 , n79585 );
buf ( R_6c5_13d59398 , n79628 );
buf ( R_17d6_11c6d258 , C0 );
buf ( R_1303_156b3d38 , n79629 );
buf ( R_b98_14b1aeb8 , n79630 );
buf ( R_ce4_117f17b8 , n79631 );
buf ( R_96b_15816c18 , n79632 );
buf ( R_8f2_158891d8 , C0 );
buf ( R_f11_124c3598 , n79638 );
buf ( R_15a9_1007e0b8 , n79654 );
buf ( R_1530_13c1c5b8 , n79655 );
buf ( R_f8a_1580da78 , C0 );
buf ( R_5ab_13d20b98 , n79662 );
buf ( R_cb2_15883eb8 , C0 );
buf ( R_bca_1162ecf8 , C0 );
buf ( R_693_1580e978 , n79663 );
buf ( R_18f0_14868178 , n79664 );
buf ( R_11e9_12fc0518 , n79689 );
buf ( R_12d1_15ff4388 , n79694 );
buf ( R_1808_117ec998 , n79695 );
buf ( R_112e_124c40d8 , C0 );
buf ( R_d6d_10080278 , n79738 );
buf ( R_b0f_150e1e98 , n79739 );
buf ( R_138c_14a12938 , n79740 );
buf ( R_19ab_1486d5d8 , n79741 );
buf ( R_174d_13c05318 , n79744 );
buf ( R_74e_117e9dd8 , C0 );
buf ( R_5d4_1587e918 , n79745 );
buf ( R_18c7_117ed7f8 , n79746 );
buf ( R_bf3_158826f8 , n79747 );
buf ( R_12a8_140b92d8 , n79748 );
buf ( R_1212_13debed8 , C0 );
buf ( R_c89_15886078 , n79791 );
buf ( R_1831_13b99eb8 , n79805 );
buf ( R_66a_117f7c58 , C0 );
buf ( R_16fb_13d39a38 , n79806 );
buf ( R_10dc_140acad8 , n79807 );
buf ( R_abd_12fbf938 , n79841 );
buf ( R_7a0_1162cef8 , n79842 );
buf ( R_dbf_13d1dd58 , n79843 );
buf ( R_13de_13bf51d8 , C0 );
buf ( R_19fd_13c22cd8 , n79849 );
buf ( R_a62_11630378 , C0 );
buf ( R_e1a_13d29f18 , C0 );
buf ( R_1081_156ae298 , n79866 );
buf ( R_7fb_13c27c38 , n79867 );
buf ( R_16a0_1007f9b8 , n79868 );
buf ( R_1a58_123b6a18 , n79869 );
buf ( R_1439_11637c18 , n79912 );
buf ( R_1511_1162c778 , n79961 );
buf ( R_15c8_10085a98 , n79962 );
buf ( R_8d3_15fefba8 , n79963 );
buf ( R_fa9_150dc218 , n79980 );
buf ( R_ef2_13d3af78 , C0 );
buf ( R_98a_11629578 , C0 );
buf ( R_151a_15ff8d48 , C0 );
buf ( R_15bf_15ff4f68 , n79981 );
buf ( R_8dc_13dd7b58 , n79982 );
buf ( R_fa0_1162a838 , n79983 );
buf ( R_efb_13ccc2b8 , n79984 );
buf ( R_981_156acad8 , n80012 );
buf ( R_133f_11636ef8 , n80013 );
buf ( R_179a_13ccf918 , C0 );
buf ( R_701_13dd6438 , n80056 );
buf ( R_195e_15817578 , C0 );
buf ( R_117b_156b5f98 , n80057 );
buf ( R_d20_1162aa18 , n80058 );
buf ( R_b5c_116370d8 , n80059 );
buf ( R_c0c_13d3f7f8 , n80060 );
buf ( R_122b_117ec498 , n80061 );
buf ( R_18ae_13d39998 , C0 );
buf ( R_184a_124c54d8 , C0 );
buf ( R_128f_123b97b8 , n80062 );
buf ( R_c70_15885998 , n80063 );
buf ( R_651_14a122f8 , n80106 );
buf ( R_5ed_13cccad8 , n80149 );
buf ( R_1a0b_1486ee38 , n80150 );
buf ( R_13ec_117f2758 , n80151 );
buf ( R_dcd_13d1e438 , n80194 );
buf ( R_7ae_13d3c058 , C0 );
buf ( R_aaf_140af698 , n80195 );
buf ( R_10ce_11637538 , C0 );
buf ( R_16ed_156af558 , n80218 );
buf ( R_a55_12fbef38 , n80251 );
buf ( R_e27_13d405b8 , n80252 );
buf ( R_1074_14b1a878 , n80253 );
buf ( R_808_13c22c38 , n80254 );
buf ( R_1693_13cd4558 , n80255 );
buf ( R_1a65_1587f8b8 , n80258 );
buf ( R_1446_1587eff8 , C0 );
buf ( R_a3c_150e6038 , n80259 );
buf ( R_821_117f1b78 , n80308 );
buf ( R_105b_13cd2f78 , n80309 );
buf ( R_145f_13b8d398 , n80310 );
buf ( R_167a_13df45d8 , C0 );
buf ( R_e40_13c26f18 , n80311 );
buf ( R_1584_1580b318 , n80312 );
buf ( R_f65_13d3b5b8 , n80328 );
buf ( R_946_14a10a98 , C0 );
buf ( R_917_117f5458 , n80329 );
buf ( R_f36_14a118f8 , C0 );
buf ( R_1555_15815638 , n80385 );
buf ( R_cd0_117f6d58 , n80386 );
buf ( R_58d_1587f3b8 , n80387 );
buf ( R_17ea_15ffadc8 , C0 );
buf ( R_190e_13bf3d38 , C0 );
buf ( R_6b1_15ffc808 , n80430 );
buf ( R_bac_13c0a098 , n80431 );
buf ( R_12ef_14b277f8 , n80432 );
buf ( R_11cb_15ff6f48 , n80433 );
buf ( R_977_1580b1d8 , n80434 );
buf ( R_8e6_1580c0d8 , C0 );
buf ( R_15b5_14866f58 , n80450 );
buf ( R_f05_123b8ef8 , n80456 );
buf ( R_f96_15885538 , C0 );
buf ( R_1524_1162d178 , n80457 );
buf ( R_11a5_156b5138 , n80471 );
buf ( R_567_13bf17b8 , n80473 );
buf ( R_6d7_12fc12d8 , n80474 );
buf ( R_1315_123b2698 , n80517 );
buf ( R_17c4_13ccc718 , n80518 );
buf ( R_b86_123b9a38 , C0 );
buf ( R_cf6_14b29738 , C0 );
buf ( R_1934_123bf7f8 , n80519 );
buf ( R_1338_116375d8 , n80520 );
buf ( R_6fa_13bec218 , C0 );
buf ( R_1182_13c1c658 , C0 );
buf ( R_1957_13d3ec18 , n80521 );
buf ( R_d19_13def3f8 , n80564 );
buf ( R_b63_15ffbb88 , n80565 );
buf ( R_17a1_117f24d8 , n80594 );
buf ( R_132d_1587ce38 , n80637 );
buf ( R_6ef_158893b8 , n80638 );
buf ( R_118d_124c3958 , n80652 );
buf ( R_194c_1587cbb8 , n80653 );
buf ( R_d0e_13c10998 , C0 );
buf ( R_b6e_117ef5f8 , C0 );
buf ( R_17ac_1486cb38 , n80654 );
buf ( R_12b2_156ab458 , C0 );
buf ( R_be9_14867638 , n80705 );
buf ( R_c93_14a12258 , n80706 );
buf ( R_1208_13bec358 , n80707 );
buf ( R_674_123c0018 , n80708 );
buf ( R_1827_13c01b78 , n80709 );
buf ( R_18d1_117e98d8 , n80734 );
buf ( R_5ca_13ccca38 , C0 );
buf ( R_16fd_13bf4378 , n80751 );
buf ( R_10de_140b68f8 , C0 );
buf ( R_abf_13befd78 , n80752 );
buf ( R_79e_15817b18 , C0 );
buf ( R_dbd_117f2b18 , n80795 );
buf ( R_13dc_13d1ce58 , n80796 );
buf ( R_19fb_150e3978 , n80797 );
buf ( R_858_150dae18 , n80798 );
buf ( R_1496_13b8b098 , C0 );
buf ( R_1643_1162c278 , n80799 );
buf ( R_a05_117f4cd8 , n80824 );
buf ( R_e77_1486b878 , n80825 );
buf ( R_1024_11635058 , n80826 );
buf ( R_733_10086998 , n80827 );
buf ( R_b2a_150dd2f8 , C0 );
buf ( R_d52_1580c498 , C0 );
buf ( R_1768_15813b58 , n80828 );
buf ( R_1371_156b10d8 , n80871 );
buf ( R_1149_156aff58 , n80921 );
buf ( R_1990_117f1df8 , n80922 );
buf ( R_185d_1162a0b8 , n80943 );
buf ( R_189b_123bccd8 , n80944 );
buf ( R_127c_1580f198 , n80945 );
buf ( R_c5d_13bf88d8 , n80988 );
buf ( R_63e_170163c8 , C0 );
buf ( R_600_150e8798 , n80989 );
buf ( R_c1f_117ebdb8 , n80990 );
buf ( R_123e_13ccb318 , C0 );
buf ( R_bfe_17018b28 , C0 );
buf ( R_18bc_123b9df8 , n80991 );
buf ( R_121d_11632718 , n81016 );
buf ( R_129d_117f6998 , n81067 );
buf ( R_183c_14b21498 , n81068 );
buf ( R_c7e_14a0d6b8 , C0 );
buf ( R_65f_14874978 , n81069 );
buf ( R_5df_13c24178 , n81070 );
buf ( R_833_117f3dd8 , n81071 );
buf ( R_a2a_14869bb8 , C0 );
buf ( R_1471_140adbb8 , n81114 );
buf ( R_1049_11636138 , n81137 );
buf ( R_e52_13d4e498 , C0 );
buf ( R_1668_13b909f8 , n81138 );
buf ( R_15df_14b24c38 , n81139 );
buf ( R_14fa_15ff7128 , C0 );
buf ( R_fc0_13beba98 , n81140 );
buf ( R_8bc_14a0e338 , n81141 );
buf ( R_9a1_123b5758 , n81165 );
buf ( R_edb_17017048 , n81166 );
buf ( R_1a0d_13ccaaf8 , n81172 );
buf ( R_13ee_13d23398 , C0 );
buf ( R_dcf_13cccfd8 , n81173 );
buf ( R_7b0_123bf4d8 , n81174 );
buf ( R_aad_14873a78 , n81199 );
buf ( R_10cc_13cd01d8 , n81200 );
buf ( R_16eb_150e81f8 , n81201 );
buf ( R_172d_13cda318 , n81231 );
buf ( R_13ac_116343d8 , n81232 );
buf ( R_110e_14a11998 , C0 );
buf ( R_19cb_13d3a758 , n81233 );
buf ( R_aef_13d50dd8 , n81234 );
buf ( R_76e_13bf8d38 , C0 );
buf ( R_d8d_13dd52b8 , n81277 );
buf ( R_715_13b94ff8 , n81320 );
buf ( R_1972_156aa918 , C0 );
buf ( R_1786_140b5778 , C0 );
buf ( R_d34_15ff3b68 , n81321 );
buf ( R_1167_1587c7f8 , n81322 );
buf ( R_1353_123c05b8 , n81323 );
buf ( R_b48_15814378 , n81324 );
buf ( R_17fb_11c6bd18 , n81325 );
buf ( R_59e_13cd0098 , n81332 );
buf ( R_cbf_15fed948 , n81333 );
buf ( R_bbd_13b8f418 , n81375 );
buf ( R_18fd_15882798 , n81426 );
buf ( R_6a0_117edbb8 , n81427 );
buf ( R_11dc_150db458 , n81428 );
buf ( R_12de_117e9658 , C0 );
buf ( R_19db_123b8458 , n81429 );
buf ( R_171d_13d45e78 , n81446 );
buf ( R_10fe_117ebd18 , C0 );
buf ( R_adf_13ccfcd8 , n81447 );
buf ( R_77e_123bcff8 , C0 );
buf ( R_d9d_12fc0298 , n81490 );
buf ( R_13bc_13c07cf8 , n81491 );
buf ( R_142a_14a0f2d8 , C0 );
buf ( R_1090_1486e7f8 , n81492 );
buf ( R_e0b_156b7758 , n81493 );
buf ( R_16af_1486be18 , n81494 );
buf ( R_7ec_123b4038 , n81495 );
buf ( R_1a49_13ccbb38 , n81501 );
buf ( R_a71_117f59f8 , n81551 );
buf ( R_15f2_13d4fe38 , C0 );
buf ( R_ec8_15883058 , n81552 );
buf ( R_fd3_10088798 , n81553 );
buf ( R_14e7_14b1ce98 , n81554 );
buf ( R_9b4_13bf5b38 , n81555 );
buf ( R_8a9_13c21298 , n81571 );
buf ( R_ece_11634bf8 , C0 );
buf ( R_15ec_13d3f4d8 , n81572 );
buf ( R_14ed_117f5f98 , n81621 );
buf ( R_fcd_1580d258 , n81644 );
buf ( R_8af_13ddfb78 , n81645 );
buf ( R_9ae_140b18f8 , C0 );
buf ( R_1501_117f0a98 , n81694 );
buf ( R_15d8_11c6ea18 , n81695 );
buf ( R_fb9_15ff0be8 , n81723 );
buf ( R_8c3_10081498 , n81724 );
buf ( R_99a_15ffaaa8 , C0 );
buf ( R_ee2_13cd1b78 , C0 );
buf ( R_1712_11637178 , C0 );
buf ( R_10f3_14a19238 , n81725 );
buf ( R_ad4_14a0a5f8 , n81726 );
buf ( R_789_140b2cf8 , n81769 );
buf ( R_da8_140b3838 , n81770 );
buf ( R_13c7_13df0ed8 , n81771 );
buf ( R_19e6_11636958 , C0 );
buf ( R_95d_117f8338 , n81788 );
buf ( R_900_140b74d8 , n81789 );
buf ( R_f1f_1587f1d8 , n81790 );
buf ( R_153e_13d410f8 , C0 );
buf ( R_159b_1162f658 , n81791 );
buf ( R_f7c_15ffc268 , n81792 );
buf ( R_cc5_13b8c858 , n81835 );
buf ( R_598_17015108 , n81841 );
buf ( R_17f5_13c1c798 , n81856 );
buf ( R_1903_1162d2b8 , n81857 );
buf ( R_6a6_15816df8 , C0 );
buf ( R_bb7_14a17a78 , n81858 );
buf ( R_12e4_13df4678 , n81859 );
buf ( R_11d6_13cccf38 , C0 );
buf ( R_a4d_14a159f8 , n81887 );
buf ( R_810_1007f918 , n81888 );
buf ( R_106c_13cd4238 , n81889 );
buf ( R_168b_13d20d78 , n81890 );
buf ( R_144e_17019028 , C0 );
buf ( R_e2f_123b83b8 , n81891 );
buf ( R_f66_1700e448 , C0 );
buf ( R_947_13cd36f8 , n81892 );
buf ( R_916_12fbefd8 , C0 );
buf ( R_f35_13dd5fd8 , n81908 );
buf ( R_1554_13c04918 , n81909 );
buf ( R_1585_117efe18 , n81933 );
buf ( R_16ff_13b95318 , n81934 );
buf ( R_10e0_1580e478 , n81935 );
buf ( R_ac1_13d23078 , n81958 );
buf ( R_79c_1162d8f8 , n81959 );
buf ( R_dbb_1580e018 , n81960 );
buf ( R_13da_123c03d8 , C0 );
buf ( R_19f9_13cd81f8 , n81966 );
buf ( R_a3f_13c012b8 , n81967 );
buf ( R_81e_140b4cd8 , C0 );
buf ( R_105e_156ba278 , C0 );
buf ( R_145c_13ddc0b8 , n81968 );
buf ( R_167d_124c5438 , n81985 );
buf ( R_e3d_15889778 , n82028 );
buf ( R_be0_117ea5f8 , n82029 );
buf ( R_c9c_13b8ed38 , n82030 );
buf ( R_11ff_14a17618 , n82031 );
buf ( R_67d_156b7398 , n82074 );
buf ( R_181e_13c04e18 , C0 );
buf ( R_18da_13cd38d8 , C0 );
buf ( R_5c1_13c0a818 , n82100 );
buf ( R_12bb_13b8a918 , n82101 );
buf ( R_ca4_156b1c18 , n82102 );
buf ( R_bd8_117e87f8 , n82103 );
buf ( R_685_13bf38d8 , n82146 );
buf ( R_11f7_10080b38 , n82147 );
buf ( R_18e2_13becfd8 , C0 );
buf ( R_1816_14b1ff58 , C0 );
buf ( R_12c3_10083478 , n82148 );
buf ( R_5b9_140b2bb8 , n82153 );
buf ( R_1630_123b9cb8 , n82154 );
buf ( R_e8a_14b1db18 , C0 );
buf ( R_9f2_10089418 , C0 );
buf ( R_14a9_156acb78 , n82197 );
buf ( R_1011_12fbe218 , n82219 );
buf ( R_86b_124c4e98 , n82220 );
buf ( R_1726_14869a78 , C0 );
buf ( R_19d2_13d533f8 , C0 );
buf ( R_1107_13df9038 , n82221 );
buf ( R_ae8_13bef5f8 , n82222 );
buf ( R_775_158109f8 , n82265 );
buf ( R_d94_12fbf6b8 , n82266 );
buf ( R_13b3_13d40158 , n82267 );
buf ( R_1658_13bf9ff8 , n82268 );
buf ( R_843_150e0458 , n82269 );
buf ( R_1481_117e8e38 , n82312 );
buf ( R_a1a_15fefd88 , C0 );
buf ( R_1039_13ddba78 , n82330 );
buf ( R_e62_13c23098 , C0 );
buf ( R_1a0f_13c24038 , n82331 );
buf ( R_13f0_11c6e338 , n82332 );
buf ( R_dd1_13de4a38 , n82375 );
buf ( R_7b2_13bf2898 , C0 );
buf ( R_aab_13c1cfb8 , n82376 );
buf ( R_10ca_1700ac08 , C0 );
buf ( R_16e9_15ff3668 , n82400 );
buf ( R_1793_150de018 , n82401 );
buf ( R_708_14a0d258 , n82402 );
buf ( R_1965_13ccb6d8 , n82413 );
buf ( R_1174_11c6c358 , n82414 );
buf ( R_d27_13dee138 , n82415 );
buf ( R_b55_15ffb0e8 , n82440 );
buf ( R_1346_13d3f2f8 , C0 );
buf ( R_e1f_123b6ab8 , n82441 );
buf ( R_107c_117f4058 , n82442 );
buf ( R_800_13d219f8 , n82443 );
buf ( R_169b_150e49b8 , n82444 );
buf ( R_1a5d_1486e398 , n82447 );
buf ( R_143e_14a19f58 , C0 );
buf ( R_a5d_15880498 , n82475 );
buf ( R_1a22_15810b38 , C0 );
buf ( R_1403_124c5398 , n82476 );
buf ( R_de4_117f6498 , n82477 );
buf ( R_7c5_15ffbe08 , n82520 );
buf ( R_a98_1486db78 , n82521 );
buf ( R_10b7_14a17578 , n82522 );
buf ( R_16d6_14a10458 , C0 );
buf ( R_1a2d_13b8fcd8 , n82528 );
buf ( R_140e_13def718 , C0 );
buf ( R_def_13d3eb78 , n82529 );
buf ( R_7d0_156b2e38 , n82530 );
buf ( R_a8d_11632678 , n82554 );
buf ( R_10ac_156b5958 , n82555 );
buf ( R_16cb_156b72f8 , n82556 );
buf ( R_1634_17018c68 , n82557 );
buf ( R_9f6_158867f8 , C0 );
buf ( R_e86_14a183d8 , C0 );
buf ( R_1015_14b1e6f8 , n82574 );
buf ( R_867_15881398 , n82575 );
buf ( R_14a5_11629ed8 , n82618 );
buf ( R_e8e_150da878 , C0 );
buf ( R_9ee_13d54618 , C0 );
buf ( R_162c_13b96c18 , n82619 );
buf ( R_14ad_12fbf618 , n82662 );
buf ( R_86f_15ff83e8 , n82663 );
buf ( R_100d_158136f8 , n82685 );
buf ( R_189c_14a10c78 , n82686 );
buf ( R_127d_11636318 , n82737 );
buf ( R_c5e_15882a18 , C0 );
buf ( R_63f_156b5b38 , n82738 );
buf ( R_5ff_13d40ab8 , n82739 );
buf ( R_c1e_14a0b958 , C0 );
buf ( R_123d_13ddd5f8 , n82764 );
buf ( R_185c_11630738 , n82765 );
buf ( R_141e_13b90818 , C0 );
buf ( R_16bb_123b7d78 , n82766 );
buf ( R_dff_117eeb58 , n82767 );
buf ( R_7e0_13dfacf8 , n82768 );
buf ( R_a7d_123b7af8 , n82813 );
buf ( R_1a3d_156b9cd8 , n82819 );
buf ( R_109c_13b98d38 , n82820 );
buf ( R_cb9_150db638 , n82863 );
buf ( R_bc3_156b6678 , n82864 );
buf ( R_69a_13b8b6d8 , C0 );
buf ( R_18f7_13b90bd8 , n82865 );
buf ( R_11e2_13d1e4d8 , C0 );
buf ( R_12d8_13d43718 , n82866 );
buf ( R_1801_13c013f8 , n82880 );
buf ( R_5a4_15ff7d08 , n82886 );
buf ( R_13a5_13d45338 , n82929 );
buf ( R_1115_11630b98 , n82958 );
buf ( R_19c4_17016fa8 , n82959 );
buf ( R_af6_117f49b8 , C0 );
buf ( R_767_117f2d98 , n82960 );
buf ( R_d86_15fef7e8 , C0 );
buf ( R_1734_1580c718 , n82961 );
buf ( R_836_123b33b8 , C0 );
buf ( R_a27_117ede38 , n82962 );
buf ( R_1474_13c042d8 , n82963 );
buf ( R_1046_123bc918 , C0 );
buf ( R_e55_124c3a98 , n83006 );
buf ( R_1665_156ac678 , n83023 );
buf ( R_122a_14a0b318 , C0 );
buf ( R_18af_11c6f7d8 , n83024 );
buf ( R_1849_140b6358 , n83039 );
buf ( R_1290_13dd8b98 , n83040 );
buf ( R_c71_14a11e98 , n83083 );
buf ( R_652_13d386d8 , C0 );
buf ( R_5ec_14868df8 , n83084 );
buf ( R_c0b_13b8c038 , n83085 );
buf ( R_574_13d4ec18 , n83087 );
buf ( R_6ca_156b3f18 , C0 );
buf ( R_1308_117f2438 , n83088 );
buf ( R_17d1_11c6fa58 , n83115 );
buf ( R_b93_15881078 , n83116 );
buf ( R_ce9_156b86f8 , n83159 );
buf ( R_1927_123bb6f8 , n83160 );
buf ( R_11b2_14a101d8 , C0 );
buf ( R_8f1_14a0fcd8 , n83177 );
buf ( R_f10_156ab778 , n83178 );
buf ( R_15aa_13c1f498 , C0 );
buf ( R_152f_158884b8 , n83179 );
buf ( R_f8b_13dda218 , n83180 );
buf ( R_96c_15ff4e28 , n83181 );
buf ( R_948_15ff1728 , n83182 );
buf ( R_915_158834b8 , n83204 );
buf ( R_f34_123bd958 , n83205 );
buf ( R_1553_1162fdd8 , n83206 );
buf ( R_1586_13cd7938 , C0 );
buf ( R_f67_156b54f8 , n83207 );
buf ( R_1701_117ee5b8 , n83224 );
buf ( R_10e2_13b97cf8 , C0 );
buf ( R_ac3_13d41ff8 , n83225 );
buf ( R_79a_13b8d758 , C0 );
buf ( R_db9_13d4e358 , n83268 );
buf ( R_13d8_13c10178 , n83269 );
buf ( R_19f7_123b4218 , n83270 );
buf ( R_ec2_156acdf8 , C0 );
buf ( R_fd9_13cd6038 , n83292 );
buf ( R_14e1_13d4fbb8 , n83335 );
buf ( R_9ba_13d3b018 , C0 );
buf ( R_8a3_117f3298 , n83336 );
buf ( R_15f8_150dd618 , n83337 );
buf ( R_b1c_10084238 , n83338 );
buf ( R_d60_1700c1e8 , n83339 );
buf ( R_137f_13d27fd8 , n83340 );
buf ( R_175a_15fedda8 , C0 );
buf ( R_199e_123b8d18 , C0 );
buf ( R_113b_11c703b8 , n83341 );
buf ( R_741_156b0278 , n83384 );
buf ( R_15e6_140b4238 , C0 );
buf ( R_14f3_10088a18 , n83385 );
buf ( R_fc7_117e8c58 , n83386 );
buf ( R_8b5_13ccefb8 , n83402 );
buf ( R_9a8_14a19af8 , n83403 );
buf ( R_ed4_150e1998 , n83404 );
buf ( R_d68_15885b78 , n83405 );
buf ( R_b14_11c6b8b8 , n83406 );
buf ( R_1387_117eaf58 , n83407 );
buf ( R_19a6_14a19738 , C0 );
buf ( R_1752_150e4738 , C0 );
buf ( R_749_123b2918 , n83450 );
buf ( R_1133_1587e378 , n83451 );
buf ( R_1417_15ff4428 , n83452 );
buf ( R_df8_15888eb8 , n83453 );
buf ( R_7d9_124c3098 , n83502 );
buf ( R_a84_13b8b778 , n83503 );
buf ( R_10a3_13c1e4f8 , n83504 );
buf ( R_1a36_14b1b318 , C0 );
buf ( R_16c2_156b1e98 , C0 );
buf ( R_1a11_123b7b98 , n83511 );
buf ( R_13f2_13de2738 , C0 );
buf ( R_dd3_14a19a58 , n83512 );
buf ( R_7b4_15885a38 , n83513 );
buf ( R_aa9_13cd5818 , n83538 );
buf ( R_10c8_14a14058 , n83539 );
buf ( R_16e7_117eea18 , n83540 );
buf ( R_b27_10087e38 , n83541 );
buf ( R_d55_117f0f98 , n83584 );
buf ( R_1765_12fbdf98 , n83612 );
buf ( R_1374_17015888 , n83613 );
buf ( R_1146_123bed58 , C0 );
buf ( R_1993_13d53b78 , n83614 );
buf ( R_736_15ff9108 , C0 );
buf ( R_56b_123b7558 , n83615 );
buf ( R_6d3_1007e1f8 , n83616 );
buf ( R_1311_10087a78 , n83659 );
buf ( R_17c8_13d50a18 , n83660 );
buf ( R_b8a_14b26858 , C0 );
buf ( R_cf2_14a17438 , C0 );
buf ( R_1930_13c083d8 , n83661 );
buf ( R_11a9_117f1038 , n83675 );
buf ( R_1638_15815818 , n83676 );
buf ( R_9fa_123b77d8 , C0 );
buf ( R_e82_13df3ef8 , C0 );
buf ( R_1019_158858f8 , n83694 );
buf ( R_863_13d47318 , n83695 );
buf ( R_14a1_117ed938 , n83738 );
buf ( R_eb2_11c6d2f8 , C0 );
buf ( R_fe9_1162ed98 , n83760 );
buf ( R_14d1_1587ae58 , n83803 );
buf ( R_9ca_1587bd58 , C0 );
buf ( R_893_13ccf238 , n83804 );
buf ( R_1608_117f45f8 , n83805 );
buf ( R_6f3_17012cc8 , n83806 );
buf ( R_1189_13de2d78 , n83837 );
buf ( R_1950_123b8098 , n83838 );
buf ( R_d12_13cd6d58 , C0 );
buf ( R_b6a_140afff8 , C0 );
buf ( R_17a8_13d3cf58 , n83839 );
buf ( R_1331_148755f8 , n83882 );
buf ( R_e9f_17016288 , n83883 );
buf ( R_9dd_156ab8b8 , n83900 );
buf ( R_161b_13d3ca58 , n83901 );
buf ( R_14be_13b98478 , C0 );
buf ( R_880_117ea2d8 , n83902 );
buf ( R_ffc_13b8acd8 , n83903 );
buf ( R_1789_13cca9b8 , n83936 );
buf ( R_196f_13bf01d8 , n83937 );
buf ( R_d31_156b13f8 , n83980 );
buf ( R_116a_13c23e58 , C0 );
buf ( R_1350_11632498 , n83981 );
buf ( R_b4b_156ad398 , n83982 );
buf ( R_712_13b90d18 , C0 );
buf ( R_e92_117f2ed8 , C0 );
buf ( R_9ea_123b7e18 , C0 );
buf ( R_1628_123b7698 , n83983 );
buf ( R_14b1_14a16e98 , n84026 );
buf ( R_873_14a14238 , n84027 );
buf ( R_1009_13b980b8 , n84044 );
buf ( R_bf2_170099e8 , C0 );
buf ( R_12a9_1162d0d8 , n84094 );
buf ( R_1211_150e5278 , n84119 );
buf ( R_c8a_150e3798 , C0 );
buf ( R_1830_13bf6358 , n84120 );
buf ( R_66b_150e1498 , n84121 );
buf ( R_5d3_158808f8 , n84122 );
buf ( R_18c8_13cd9f58 , n84123 );
buf ( R_a42_15888198 , C0 );
buf ( R_81b_12fbec18 , n84124 );
buf ( R_1061_13d3c558 , n84141 );
buf ( R_1459_17016aa8 , n84184 );
buf ( R_1680_1486aab8 , n84185 );
buf ( R_e3a_123bb798 , C0 );
buf ( R_17ef_15889958 , n84186 );
buf ( R_1909_15815e58 , n84237 );
buf ( R_6ac_12fc1918 , n84238 );
buf ( R_bb1_14874d38 , n84263 );
buf ( R_12ea_13ddf358 , C0 );
buf ( R_11d0_170096c8 , n84264 );
buf ( R_ccb_117ec038 , n84265 );
buf ( R_592_13c23958 , n84266 );
buf ( R_fee_14b29f58 , C0 );
buf ( R_ead_13c22378 , n84315 );
buf ( R_9cf_1162e118 , n84316 );
buf ( R_14cc_123c0b58 , n84317 );
buf ( R_160d_123bff78 , n84333 );
buf ( R_88e_123c0fb8 , C0 );
buf ( R_8ff_156b7c58 , n84334 );
buf ( R_f1e_15880038 , C0 );
buf ( R_153d_15811218 , n84390 );
buf ( R_159c_15815db8 , n84391 );
buf ( R_f7d_13cd0778 , n84407 );
buf ( R_95e_13b98018 , C0 );
buf ( R_189d_13cd3518 , n84432 );
buf ( R_127e_13d4f118 , C0 );
buf ( R_c5f_12fbfa78 , n84433 );
buf ( R_640_140b2258 , n84434 );
buf ( R_5fe_15888558 , C0 );
buf ( R_c1d_13dfb1f8 , n84484 );
buf ( R_123c_15fee708 , n84485 );
buf ( R_185b_14b21538 , n84486 );
buf ( R_15d1_123b63d8 , n84502 );
buf ( R_fb2_15810818 , C0 );
buf ( R_8ca_15815bd8 , C0 );
buf ( R_993_11c6b598 , n84503 );
buf ( R_ee9_1700fca8 , n84512 );
buf ( R_1508_156b7898 , n84513 );
buf ( R_121c_158871f8 , n84514 );
buf ( R_129e_13d3cb98 , C0 );
buf ( R_183b_13c20bb8 , n84515 );
buf ( R_c7f_13cd6ad8 , n84516 );
buf ( R_660_156ba458 , n84517 );
buf ( R_5de_123b7cd8 , C0 );
buf ( R_18bd_140b9878 , n84542 );
buf ( R_bfd_11c6f238 , n84593 );
buf ( R_16b4_117ead78 , n84594 );
buf ( R_e06_1580ff58 , C0 );
buf ( R_7e7_15885858 , n84595 );
buf ( R_1a44_1162c4f8 , n84596 );
buf ( R_a76_13d38638 , C0 );
buf ( R_1095_156b0ef8 , n84611 );
buf ( R_1425_13d571d8 , n84654 );
buf ( R_8e5_150db318 , n84670 );
buf ( R_15b6_1580e838 , C0 );
buf ( R_f04_15885038 , n84671 );
buf ( R_f97_1700c288 , n84672 );
buf ( R_1523_140b8e78 , n84673 );
buf ( R_978_156b6498 , n84674 );
buf ( R_914_13d54c58 , n84675 );
buf ( R_f33_13d59258 , n84676 );
buf ( R_1552_13ccfa58 , C0 );
buf ( R_1587_140aacd8 , n84677 );
buf ( R_f68_140acb78 , n84678 );
buf ( R_949_14b26a38 , n84695 );
buf ( R_15c0_158147d8 , n84696 );
buf ( R_8db_1580e158 , n84697 );
buf ( R_fa1_1162ffb8 , n84714 );
buf ( R_efa_13bf5818 , C0 );
buf ( R_982_13debcf8 , C0 );
buf ( R_1519_15813e78 , n84763 );
buf ( R_164e_117eb138 , C0 );
buf ( R_148b_15886118 , n84764 );
buf ( R_a10_13df0f78 , n84765 );
buf ( R_e6c_15ff0d28 , n84766 );
buf ( R_102f_123c08d8 , n84767 );
buf ( R_84d_15feee88 , n84832 );
buf ( R_1703_13c254d8 , n84833 );
buf ( R_10e4_158894f8 , n84834 );
buf ( R_ac5_15883558 , n84849 );
buf ( R_798_123beb78 , n84850 );
buf ( R_db7_14869938 , n84851 );
buf ( R_13d6_156ae8d8 , C0 );
buf ( R_19f5_13d2c2b8 , n84857 );
buf ( R_eb7_11c6d1b8 , n84858 );
buf ( R_fe4_12fc21d8 , n84859 );
buf ( R_14d6_1008b178 , C0 );
buf ( R_9c5_14b21d58 , n84878 );
buf ( R_898_123b5c58 , n84879 );
buf ( R_1603_14872fd8 , n84880 );
buf ( R_1714_15889638 , n84881 );
buf ( R_10f5_140b5f98 , n84915 );
buf ( R_ad6_14873258 , C0 );
buf ( R_787_14a0e838 , n84916 );
buf ( R_da6_13ddc158 , C0 );
buf ( R_13c5_15fee208 , n84959 );
buf ( R_19e4_13de3a98 , n84960 );
buf ( R_98b_13b8dcf8 , n84961 );
buf ( R_ef1_13b924d8 , n84966 );
buf ( R_8d2_156ad578 , C0 );
buf ( R_faa_156b0458 , C0 );
buf ( R_1510_13d1f0b8 , n84967 );
buf ( R_15c9_13bf0b38 , n84983 );
buf ( R_aa7_13d451f8 , n84984 );
buf ( R_7b6_14a18018 , C0 );
buf ( R_dd5_124c5258 , n85027 );
buf ( R_10c6_1700ff28 , C0 );
buf ( R_13f4_14a0b778 , n85028 );
buf ( R_16e5_13c07ed8 , n85058 );
buf ( R_1a13_117ef058 , n85059 );
buf ( R_839_14b28f18 , n85108 );
buf ( R_e58_158814d8 , n85109 );
buf ( R_a24_123b5938 , n85110 );
buf ( R_1043_14b26538 , n85111 );
buf ( R_1477_117f0098 , n85112 );
buf ( R_1662_13df1978 , C0 );
buf ( R_854_15ff3e88 , n85113 );
buf ( R_e73_14b288d8 , n85114 );
buf ( R_a09_123bb158 , n85129 );
buf ( R_1028_117f4eb8 , n85130 );
buf ( R_1492_13cd4378 , C0 );
buf ( R_1647_12fc19b8 , n85131 );
buf ( R_be8_15ffcee8 , n85132 );
buf ( R_5c9_14b27438 , n85159 );
buf ( R_675_156aec98 , n85202 );
buf ( R_c94_13b8fb98 , n85203 );
buf ( R_1207_156b81f8 , n85204 );
buf ( R_12b3_13ddf718 , n85205 );
buf ( R_1826_140b01d8 , C0 );
buf ( R_18d2_13c290d8 , C0 );
buf ( R_cac_123c1058 , n85206 );
buf ( R_5b1_13d28e38 , n85207 );
buf ( R_68d_1700f2a8 , n85250 );
buf ( R_bd0_13ccc538 , n85251 );
buf ( R_11ef_117f3d38 , n85252 );
buf ( R_12cb_123bfe38 , n85253 );
buf ( R_180e_1580c7b8 , C0 );
buf ( R_18ea_14a115d8 , C0 );
buf ( R_d75_1486bc38 , n85296 );
buf ( R_756_13b8ae18 , C0 );
buf ( R_b07_140aaa58 , n85297 );
buf ( R_1126_156aaeb8 , C0 );
buf ( R_1394_15814878 , n85298 );
buf ( R_1745_123b4cb8 , n85310 );
buf ( R_19b3_123bc558 , n85311 );
buf ( R_d7a_13b95ef8 , C0 );
buf ( R_75b_15814558 , n85312 );
buf ( R_b02_14a13f18 , C0 );
buf ( R_1121_150e9c38 , n85336 );
buf ( R_1399_158830f8 , n85379 );
buf ( R_1740_13cd6fd8 , n85380 );
buf ( R_19b8_15812c58 , n85381 );
buf ( R_c0a_14a19ff8 , C0 );
buf ( R_5eb_15feeac8 , n85382 );
buf ( R_653_123be358 , n85383 );
buf ( R_c72_13df6fb8 , C0 );
buf ( R_1229_156b7938 , n85408 );
buf ( R_1291_14a0d758 , n85459 );
buf ( R_1848_14a197d8 , n85460 );
buf ( R_18b0_15815a98 , n85461 );
buf ( R_a96_150e8478 , C0 );
buf ( R_7c7_13d45c98 , n85462 );
buf ( R_de6_13c05778 , C0 );
buf ( R_10b5_156ab6d8 , n85474 );
buf ( R_1405_14a192d8 , n85517 );
buf ( R_16d4_14868c18 , n85518 );
buf ( R_1a24_116348d8 , n85519 );
buf ( R_85f_13dd89b8 , n85520 );
buf ( R_e7e_140ad6b8 , C0 );
buf ( R_9fe_13c02d98 , C0 );
buf ( R_101d_123b5d98 , n85538 );
buf ( R_149d_156b8dd8 , n85581 );
buf ( R_163c_1486a6f8 , n85582 );
buf ( R_d9b_13d3dbd8 , n85583 );
buf ( R_77c_116359b8 , n85584 );
buf ( R_ae1_15fed768 , n85599 );
buf ( R_1100_10085818 , n85600 );
buf ( R_13ba_15881d98 , C0 );
buf ( R_171f_13bf08b8 , n85601 );
buf ( R_19d9_1700c508 , n85611 );
buf ( R_889_15ff9b08 , n85628 );
buf ( R_9d4_11c6e6f8 , n85629 );
buf ( R_ea8_13d1fe78 , n85630 );
buf ( R_ff3_117efc38 , n85631 );
buf ( R_14c7_140b4918 , n85632 );
buf ( R_1612_13cd0278 , C0 );
buf ( R_582_14869118 , n85633 );
buf ( R_cdb_14a0ae18 , n85634 );
buf ( R_ba1_13d29338 , n85659 );
buf ( R_6bc_13cd53b8 , n85660 );
buf ( R_11c0_13deef98 , n85661 );
buf ( R_12fa_11631638 , C0 );
buf ( R_17df_13cd0e58 , n85662 );
buf ( R_1919_1587e2d8 , n85713 );
buf ( R_e24_13ddcfb8 , n85714 );
buf ( R_a58_14a18a18 , n85715 );
buf ( R_805_1580a7d8 , n85771 );
buf ( R_1077_11c6d898 , n85772 );
buf ( R_1443_13d3f9d8 , n85773 );
buf ( R_1696_156afd78 , C0 );
buf ( R_1a62_14b1b138 , C0 );
buf ( R_94a_156b24d8 , C0 );
buf ( R_f32_116350f8 , C0 );
buf ( R_913_100840f8 , n85774 );
buf ( R_f69_117f0c78 , n85790 );
buf ( R_1551_150dde38 , n85839 );
buf ( R_1588_150e7d98 , n85840 );
buf ( R_a50_13df7698 , n85841 );
buf ( R_e2c_15881e38 , n85842 );
buf ( R_80d_14a16a38 , n85898 );
buf ( R_106f_156ad938 , n85899 );
buf ( R_144b_1486ce58 , n85900 );
buf ( R_168e_123bbc98 , C0 );
buf ( R_6fe_13bf5318 , C0 );
buf ( R_b5f_13cd4918 , n85901 );
buf ( R_d1d_13def2b8 , n85944 );
buf ( R_117e_14a0ccb8 , C0 );
buf ( R_133c_117f2938 , n85945 );
buf ( R_179d_10085138 , n85991 );
buf ( R_195b_14b1c8f8 , n85992 );
buf ( R_cb3_1587b358 , n85993 );
buf ( R_5aa_13dd5678 , n85999 );
buf ( R_694_11636b38 , n86000 );
buf ( R_bc9_124c3d18 , n86052 );
buf ( R_11e8_13ccd258 , n86053 );
buf ( R_12d2_123bdc78 , C0 );
buf ( R_1807_117ee298 , n86054 );
buf ( R_18f1_156aba98 , n86108 );
buf ( R_c1c_156ba3b8 , n86109 );
buf ( R_5fd_14a10958 , n86152 );
buf ( R_641_123b90d8 , n86195 );
buf ( R_c60_158171b8 , n86196 );
buf ( R_123b_1162cd18 , n86197 );
buf ( R_127f_13b8a558 , n86198 );
buf ( R_185a_15814cd8 , C0 );
buf ( R_189e_13bf8e78 , C0 );
buf ( R_877_13d3e498 , n86199 );
buf ( R_9e6_14b28838 , C0 );
buf ( R_e96_156b4a58 , C0 );
buf ( R_1005_13c1edb8 , n86216 );
buf ( R_14b5_15882018 , n86259 );
buf ( R_1624_10086cb8 , n86260 );
buf ( R_db5_117ece98 , n86303 );
buf ( R_796_156b0138 , C0 );
buf ( R_ac7_148725d8 , n86304 );
buf ( R_10e6_11630918 , C0 );
buf ( R_13d4_15882bf8 , n86305 );
buf ( R_1705_10085db8 , n86323 );
buf ( R_19f3_1008c618 , n86324 );
buf ( R_96d_1162e7f8 , n86346 );
buf ( R_f0f_13d3d9f8 , n86347 );
buf ( R_8f0_13d29838 , n86348 );
buf ( R_f8c_117f2578 , n86349 );
buf ( R_152e_117f3f18 , C0 );
buf ( R_15ab_13ccc358 , n86350 );
buf ( R_587_124c5118 , n86351 );
buf ( R_cd6_13d39178 , C0 );
buf ( R_ba6_156ad9d8 , C0 );
buf ( R_6b7_13c0b718 , n86352 );
buf ( R_11c5_13d39538 , n86368 );
buf ( R_12f5_158104f8 , n86411 );
buf ( R_17e4_156acf38 , n86412 );
buf ( R_1914_10084f58 , n86413 );
buf ( R_846_100885b8 , C0 );
buf ( R_e65_15810318 , n86462 );
buf ( R_a17_13ccf878 , n86463 );
buf ( R_1036_140b5278 , C0 );
buf ( R_1484_11c6b778 , n86464 );
buf ( R_1655_1700cdc8 , n86481 );
buf ( R_a45_17017188 , n86515 );
buf ( R_e37_10083018 , n86516 );
buf ( R_818_13b8dbb8 , n86517 );
buf ( R_1064_1700d5e8 , n86518 );
buf ( R_1456_13cd8518 , C0 );
buf ( R_1683_1587f6d8 , n86519 );
buf ( R_57d_14b1ef18 , n86520 );
buf ( R_ce0_1580ccb8 , n86521 );
buf ( R_b9c_15884e58 , n86522 );
buf ( R_6c1_156b1538 , n86565 );
buf ( R_11bb_117ed2f8 , n86566 );
buf ( R_12ff_17012408 , n86567 );
buf ( R_17da_123bf398 , C0 );
buf ( R_191e_140b0c78 , C0 );
buf ( R_d58_13df39f8 , n86568 );
buf ( R_b24_15815958 , n86569 );
buf ( R_739_123c1698 , n86612 );
buf ( R_1143_13cd7078 , n86613 );
buf ( R_1377_158873d8 , n86614 );
buf ( R_1762_140aef18 , C0 );
buf ( R_1996_156b4058 , C0 );
buf ( R_95f_13bf9918 , n86615 );
buf ( R_f1d_15ff80c8 , n86631 );
buf ( R_8fe_13d4f898 , C0 );
buf ( R_f7e_156b42d8 , C0 );
buf ( R_153c_13c1d698 , n86632 );
buf ( R_159d_1162b198 , n86638 );
buf ( R_aa5_156b4238 , n86663 );
buf ( R_7b8_1162e9d8 , n86664 );
buf ( R_dd7_140b62b8 , n86665 );
buf ( R_10c4_12fc1878 , n86666 );
buf ( R_13f6_1700d728 , C0 );
buf ( R_16e3_123b4d58 , n86667 );
buf ( R_1a15_13d3e998 , n86673 );
buf ( R_b0c_123c1878 , n86674 );
buf ( R_d70_13b96038 , n86675 );
buf ( R_751_13bf12b8 , n86718 );
buf ( R_112b_13d5c3b8 , n86719 );
buf ( R_138f_13df66f8 , n86720 );
buf ( R_174a_13d24658 , C0 );
buf ( R_19ae_1587f818 , C0 );
buf ( R_a8b_117f7898 , n86721 );
buf ( R_7d2_10082a78 , C0 );
buf ( R_df1_15884778 , n86764 );
buf ( R_10aa_13c28458 , C0 );
buf ( R_1410_13cd5a98 , n86765 );
buf ( R_16c9_13c03018 , n86788 );
buf ( R_1a2f_15886b18 , n86789 );
buf ( R_d7f_117f5ef8 , n86790 );
buf ( R_760_13cce6f8 , n86791 );
buf ( R_afd_156ae018 , n86805 );
buf ( R_111c_13c0f138 , n86806 );
buf ( R_139e_15ff9428 , C0 );
buf ( R_173b_13d23758 , n86807 );
buf ( R_19bd_150e0c78 , n86817 );
buf ( R_70f_14b26038 , n86818 );
buf ( R_b4e_158835f8 , C0 );
buf ( R_d2e_15ff2d08 , C0 );
buf ( R_116d_14a0bc78 , n86833 );
buf ( R_134d_13cd26b8 , n86876 );
buf ( R_178c_13d39718 , n86877 );
buf ( R_196c_117ef418 , n86878 );
buf ( R_705_17018768 , n86921 );
buf ( R_b58_12fc00b8 , n86922 );
buf ( R_d24_13c0ca78 , n86923 );
buf ( R_1177_13d5b558 , n86924 );
buf ( R_1343_13d298d8 , n86925 );
buf ( R_1796_156ae338 , C0 );
buf ( R_1962_13d5d218 , C0 );
buf ( R_c9d_13c00ef8 , n86968 );
buf ( R_bdf_117f0638 , n86969 );
buf ( R_5c0_117ea0f8 , n86970 );
buf ( R_67e_14a0b8b8 , C0 );
buf ( R_11fe_124c36d8 , C0 );
buf ( R_12bc_13b981f8 , n86971 );
buf ( R_181d_123ba758 , n86985 );
buf ( R_18db_11c6d7f8 , n86986 );
buf ( R_ebc_1580cfd8 , n86987 );
buf ( R_89d_11c693d8 , n87003 );
buf ( R_9c0_13d46b98 , n87004 );
buf ( R_fdf_158176b8 , n87005 );
buf ( R_14db_156b5e58 , n87006 );
buf ( R_15fe_140b97d8 , C0 );
buf ( R_ee1_13d40c98 , n87015 );
buf ( R_99b_156b3838 , n87016 );
buf ( R_8c2_15813518 , C0 );
buf ( R_fba_140aebf8 , C0 );
buf ( R_1500_1700e8a8 , n87017 );
buf ( R_15d9_13d53538 , n87033 );
buf ( R_eda_13d57638 , C0 );
buf ( R_9a2_13c28bd8 , C0 );
buf ( R_8bb_13d43498 , n87034 );
buf ( R_fc1_156b40f8 , n87056 );
buf ( R_14f9_13cd6178 , n87105 );
buf ( R_15e0_13cd0458 , n87106 );
buf ( R_d8b_150dc7b8 , n87107 );
buf ( R_76c_150e63f8 , n87108 );
buf ( R_af1_13b8c3f8 , n87122 );
buf ( R_1110_13d5cdb8 , n87123 );
buf ( R_13aa_14b1d898 , C0 );
buf ( R_172f_11c6dbb8 , n87124 );
buf ( R_19c9_1509b4f8 , n87134 );
buf ( R_55a_158145f8 , n87135 );
buf ( R_6e4_11630a58 , n87136 );
buf ( R_b79_13ccfd78 , n87161 );
buf ( R_d03_124c2eb8 , n87162 );
buf ( R_1198_117f3b58 , n87163 );
buf ( R_1322_15ff6ea8 , C0 );
buf ( R_17b7_15810bd8 , n87164 );
buf ( R_1941_117ed4d8 , n87214 );
buf ( R_6cf_1486c6d8 , n87215 );
buf ( R_56f_14a0b598 , n87216 );
buf ( R_cee_13cd9c38 , C0 );
buf ( R_b8e_150e97d8 , C0 );
buf ( R_11ad_13d569b8 , n87231 );
buf ( R_130d_124c3818 , n87274 );
buf ( R_17cc_117e9298 , n87275 );
buf ( R_192c_13b94918 , n87276 );
buf ( R_94b_100881f8 , n87277 );
buf ( R_f31_13c231d8 , n87293 );
buf ( R_912_11630f58 , C0 );
buf ( R_f6a_117ea058 , C0 );
buf ( R_1550_17014668 , n87294 );
buf ( R_1589_123b7198 , n87318 );
buf ( R_bd7_14a0ef18 , n87319 );
buf ( R_ca5_1007eb58 , n87362 );
buf ( R_5b8_170170e8 , n87363 );
buf ( R_686_15810f98 , C0 );
buf ( R_11f6_14b22bb8 , C0 );
buf ( R_12c4_15ff0008 , n87364 );
buf ( R_1815_156b1cb8 , n87378 );
buf ( R_18e3_13ccb9f8 , n87379 );
buf ( R_6e0_14a15f98 , n87380 );
buf ( R_55e_148707d8 , n87381 );
buf ( R_cff_14a0b458 , n87382 );
buf ( R_b7d_156b6df8 , n87407 );
buf ( R_119c_14872ad8 , n87408 );
buf ( R_131e_13dd6e38 , C0 );
buf ( R_17bb_13bf1d58 , n87409 );
buf ( R_193d_11c70638 , n87459 );
buf ( R_d92_14b21358 , C0 );
buf ( R_773_117f54f8 , n87460 );
buf ( R_aea_17012908 , C0 );
buf ( R_1109_15ff3de8 , n87488 );
buf ( R_13b1_150dc358 , n87531 );
buf ( R_1728_13d5beb8 , n87532 );
buf ( R_19d0_14870af8 , n87533 );
buf ( R_e12_13b8cc18 , C0 );
buf ( R_a6a_13d1d218 , C0 );
buf ( R_7f3_148688f8 , n87534 );
buf ( R_1089_123b6838 , n87551 );
buf ( R_1431_15812ed8 , n87594 );
buf ( R_16a8_123bf118 , n87595 );
buf ( R_1a50_117ed6b8 , n87596 );
buf ( R_6f7_117e93d8 , n87597 );
buf ( R_b66_14a0f238 , C0 );
buf ( R_d16_13c1b7f8 , C0 );
buf ( R_1185_13d1ecf8 , n87611 );
buf ( R_1335_13bf1f38 , n87654 );
buf ( R_17a4_14b1ea18 , n87655 );
buf ( R_1954_15ff1ae8 , n87656 );
buf ( R_e17_13df86d8 , n87657 );
buf ( R_a65_14b22b18 , n87702 );
buf ( R_7f8_1700bec8 , n87703 );
buf ( R_1084_13d39038 , n87704 );
buf ( R_1436_15fef608 , C0 );
buf ( R_16a3_15ff2768 , n87705 );
buf ( R_1a55_123b5898 , n87711 );
buf ( R_a21_1587bad8 , n87729 );
buf ( R_83c_13cd7398 , n87730 );
buf ( R_e5b_123bf898 , n87731 );
buf ( R_1040_1008ac78 , n87732 );
buf ( R_147a_13c04378 , C0 );
buf ( R_165f_13cd97d8 , n87733 );
buf ( R_bfc_13d53cb8 , n87734 );
buf ( R_5dd_123b45d8 , n87777 );
buf ( R_661_13d3c2d8 , n87820 );
buf ( R_c80_1008ca78 , n87821 );
buf ( R_121b_14b24698 , n87822 );
buf ( R_129f_1008b7b8 , n87823 );
buf ( R_183a_156acc18 , C0 );
buf ( R_18be_14a0de38 , C0 );
buf ( R_c1b_123b48f8 , n87824 );
buf ( R_5fc_140b3518 , n87825 );
buf ( R_642_14a0d118 , C0 );
buf ( R_c61_13c06718 , n87868 );
buf ( R_123a_15ffcf88 , C0 );
buf ( R_1280_14a106d8 , n87869 );
buf ( R_1859_13d25378 , n87884 );
buf ( R_189f_14a13c98 , n87885 );
buf ( R_556_13d2a2d8 , n87886 );
buf ( R_6e8_12fbf4d8 , n87887 );
buf ( R_b75_156ae838 , n87912 );
buf ( R_d07_156abe58 , n87913 );
buf ( R_1194_1580f058 , n87914 );
buf ( R_1326_11c684d8 , C0 );
buf ( R_17b3_13ddb4d8 , n87915 );
buf ( R_1945_14b22898 , n87965 );
buf ( R_bf1_13df18d8 , n88016 );
buf ( R_5d2_10088f18 , C0 );
buf ( R_66c_123c06f8 , n88017 );
buf ( R_c8b_13c0e5f8 , n88018 );
buf ( R_1210_117f56d8 , n88019 );
buf ( R_12aa_140afb98 , C0 );
buf ( R_182f_13d58998 , n88020 );
buf ( R_18c9_11c6eb58 , n88045 );
buf ( R_cc0_1580fcd8 , n88046 );
buf ( R_59d_13df9d58 , n88052 );
buf ( R_6a1_13cd9b98 , n88095 );
buf ( R_bbc_13d4e678 , n88096 );
buf ( R_11db_124c45d8 , n88097 );
buf ( R_12df_13d27178 , n88098 );
buf ( R_17fa_13beb8b8 , C0 );
buf ( R_18fe_1587ca78 , C0 );
buf ( R_d63_117f68f8 , n88099 );
buf ( R_b19_158882d8 , n88113 );
buf ( R_744_123bea38 , n88114 );
buf ( R_1138_14869ed8 , n88115 );
buf ( R_1382_13b8b958 , C0 );
buf ( R_1757_13de1978 , n88116 );
buf ( R_19a1_123b3598 , n88126 );
buf ( R_db3_14869898 , n88127 );
buf ( R_794_17016788 , n88128 );
buf ( R_ac9_15811cb8 , n88143 );
buf ( R_10e8_140b1538 , n88144 );
buf ( R_13d2_13c292b8 , C0 );
buf ( R_1707_13ddd9b8 , n88145 );
buf ( R_19f1_13cce518 , n88151 );
buf ( R_ecd_13d5b5f8 , n88200 );
buf ( R_9af_1587fdb8 , n88201 );
buf ( R_8ae_11631778 , C0 );
buf ( R_fce_13c051d8 , C0 );
buf ( R_14ec_156b01d8 , n88202 );
buf ( R_15ed_1008af98 , n88218 );
buf ( R_da4_13cd7438 , n88219 );
buf ( R_785_116381b8 , n88262 );
buf ( R_ad8_117f7a78 , n88263 );
buf ( R_10f7_1587f598 , n88264 );
buf ( R_13c3_13cd0b38 , n88265 );
buf ( R_1716_123b6bf8 , C0 );
buf ( R_19e2_13d567d8 , C0 );
buf ( R_58c_1587fe58 , n88266 );
buf ( R_cd1_1486dc18 , n88309 );
buf ( R_bab_13df0e38 , n88310 );
buf ( R_6b2_14867ef8 , C0 );
buf ( R_11ca_123bd9f8 , C0 );
buf ( R_12f0_158817f8 , n88311 );
buf ( R_17e9_123bb5b8 , n88326 );
buf ( R_190f_15881b18 , n88327 );
buf ( R_979_117efcd8 , n88344 );
buf ( R_f03_13c06f38 , n88345 );
buf ( R_8e4_123b2b98 , n88346 );
buf ( R_f98_13d588f8 , n88347 );
buf ( R_1522_15817d98 , C0 );
buf ( R_15b7_11636bd8 , n88348 );
buf ( R_c09_14a18bf8 , n88399 );
buf ( R_5ea_1162b558 , C0 );
buf ( R_654_150e54f8 , n88400 );
buf ( R_c73_15810958 , n88401 );
buf ( R_1228_150e4ff8 , n88402 );
buf ( R_1292_117e9fb8 , C0 );
buf ( R_1847_13d54898 , n88403 );
buf ( R_18b1_1162ae78 , n88428 );
buf ( R_ec7_10083838 , n88429 );
buf ( R_8a8_140b6858 , n88430 );
buf ( R_9b5_156b6038 , n88449 );
buf ( R_fd4_13bef878 , n88450 );
buf ( R_14e6_123be178 , C0 );
buf ( R_15f3_1580b958 , n88451 );
buf ( R_6dc_13d56738 , n88452 );
buf ( R_562_11630198 , n88454 );
buf ( R_cfb_156b77f8 , n88455 );
buf ( R_b81_14b23658 , n88480 );
buf ( R_11a0_117f1a38 , n88481 );
buf ( R_131a_13cd6678 , C0 );
buf ( R_17bf_1162eed8 , n88482 );
buf ( R_1939_13b99198 , n88532 );
buf ( R_85b_150e9ff8 , n88533 );
buf ( R_e7a_13df06b8 , C0 );
buf ( R_a02_13d20378 , C0 );
buf ( R_1021_14873438 , n88551 );
buf ( R_1499_13c056d8 , n88594 );
buf ( R_1640_15816e98 , n88595 );
buf ( R_6c6_14b27a78 , C0 );
buf ( R_578_13c06678 , n88596 );
buf ( R_ce5_117e9518 , n88639 );
buf ( R_b97_116328f8 , n88640 );
buf ( R_11b6_123b6478 , C0 );
buf ( R_1304_150e5a98 , n88641 );
buf ( R_17d5_13cd9eb8 , n88685 );
buf ( R_1923_10086ad8 , n88686 );
buf ( R_aa3_123ba9d8 , n88687 );
buf ( R_7ba_17013308 , C0 );
buf ( R_dd9_1587f4f8 , n88730 );
buf ( R_10c2_13de4358 , C0 );
buf ( R_13f8_14866c38 , n88731 );
buf ( R_16e1_1587e058 , n88756 );
buf ( R_1a17_13d3a398 , n88757 );
buf ( R_ea3_117f04f8 , n88758 );
buf ( R_884_124c4358 , n88759 );
buf ( R_9d9_14a0c178 , n88776 );
buf ( R_ff8_14a15098 , n88777 );
buf ( R_14c2_13d50e78 , C0 );
buf ( R_1617_13de3e58 , n88778 );
buf ( R_e0d_13c081f8 , n88821 );
buf ( R_a6f_140ab4f8 , n88822 );
buf ( R_7ee_117eb4f8 , C0 );
buf ( R_108e_117ecf38 , C0 );
buf ( R_142c_13d55f18 , n88823 );
buf ( R_16ad_15885df8 , n88841 );
buf ( R_1a4b_13d3a118 , n88842 );
buf ( R_e01_13b8ca38 , n88885 );
buf ( R_a7b_150e6f38 , n88886 );
buf ( R_7e2_116332f8 , C0 );
buf ( R_109a_140adc58 , C0 );
buf ( R_1420_1580acd8 , n88887 );
buf ( R_16b9_13b972f8 , n88905 );
buf ( R_1a3f_13cd8f18 , n88906 );
buf ( R_597_156aeab8 , n88913 );
buf ( R_cc6_1486fd38 , C0 );
buf ( R_bb6_13d58fd8 , C0 );
buf ( R_6a7_140b7938 , n88914 );
buf ( R_11d5_14871bd8 , n88948 );
buf ( R_12e5_14b28bf8 , n88963 );
buf ( R_17f4_156b4cd8 , n88964 );
buf ( R_1904_140b9058 , n88965 );
buf ( R_dfa_1486ff18 , C0 );
buf ( R_a82_116368b8 , C0 );
buf ( R_7db_150dd1b8 , n88966 );
buf ( R_10a1_123b8598 , n88990 );
buf ( R_1419_13df1b58 , n89033 );
buf ( R_16c0_13b994b8 , n89034 );
buf ( R_1a38_13ccab98 , n89035 );
buf ( R_911_14b22078 , n89052 );
buf ( R_94c_123bc7d8 , n89053 );
buf ( R_f30_12fbf898 , n89054 );
buf ( R_f6b_13c0a6d8 , n89055 );
buf ( R_154f_1700ea88 , n89056 );
buf ( R_158a_13c25758 , C0 );
buf ( R_d44_13b99418 , n89057 );
buf ( R_b38_13d23618 , n89058 );
buf ( R_725_13d4f618 , n89101 );
buf ( R_1157_14a13298 , n89102 );
buf ( R_1363_124c4718 , n89103 );
buf ( R_1776_15882518 , C0 );
buf ( R_1982_15816fd8 , C0 );
buf ( R_983_1700b4c8 , n89104 );
buf ( R_ef9_1007e338 , n89128 );
buf ( R_8da_1587ba38 , C0 );
buf ( R_fa2_15ffaf08 , C0 );
buf ( R_1518_13c09ff8 , n89129 );
buf ( R_15c1_13c1e138 , n89145 );
buf ( R_d41_13bf8f18 , n89188 );
buf ( R_722_14b26fd8 , C0 );
buf ( R_b3b_14a0f378 , n89189 );
buf ( R_115a_156af9b8 , C0 );
buf ( R_1360_156aa5f8 , n89190 );
buf ( R_1779_13dec3d8 , n89218 );
buf ( R_197f_1700ba68 , n89219 );
buf ( R_7fd_13d29658 , n89275 );
buf ( R_e1c_156b8158 , n89276 );
buf ( R_a60_124c2738 , n89277 );
buf ( R_107f_13d55ab8 , n89278 );
buf ( R_143b_13cd5458 , n89279 );
buf ( R_169e_13d59618 , C0 );
buf ( R_1a5a_117ecd58 , C0 );
buf ( R_a94_158121b8 , n89280 );
buf ( R_7c9_13c1bb18 , n89323 );
buf ( R_de8_13df22d8 , n89324 );
buf ( R_10b3_17011328 , n89325 );
buf ( R_1407_140b9cd8 , n89326 );
buf ( R_16d2_150e0098 , C0 );
buf ( R_1a26_14868678 , C0 );
buf ( R_e9a_14a0e1f8 , C0 );
buf ( R_87b_123b2e18 , n89327 );
buf ( R_9e2_148680d8 , C0 );
buf ( R_1001_100877f8 , n89349 );
buf ( R_14b9_150dda78 , n89392 );
buf ( R_1620_117efff8 , n89393 );
buf ( R_bc2_1580b098 , C0 );
buf ( R_cba_13c20118 , C0 );
buf ( R_5a3_13b98298 , n89399 );
buf ( R_69b_13bf94b8 , n89400 );
buf ( R_11e1_1486a798 , n89425 );
buf ( R_12d9_123ba118 , n89451 );
buf ( R_1800_15888378 , n89452 );
buf ( R_18f8_156ac538 , n89453 );
buf ( R_960_13ccf418 , n89454 );
buf ( R_f1c_13df79b8 , n89455 );
buf ( R_8fd_123b6fb8 , n89475 );
buf ( R_f7f_140aa558 , n89476 );
buf ( R_153b_117f5d18 , n89477 );
buf ( R_159e_14871db8 , C0 );
buf ( R_d47_13d27998 , n89478 );
buf ( R_b35_1587cc58 , n89493 );
buf ( R_728_140ba318 , n89494 );
buf ( R_1154_117e95b8 , n89495 );
buf ( R_1366_17015568 , C0 );
buf ( R_1773_156ac2b8 , n89496 );
buf ( R_1985_1162c3b8 , n89506 );
buf ( R_b11_15883698 , n89520 );
buf ( R_d6b_123b8958 , n89521 );
buf ( R_74c_150e17b8 , n89522 );
buf ( R_1130_13bef0f8 , n89523 );
buf ( R_138a_13d25cd8 , C0 );
buf ( R_174f_13df2058 , n89524 );
buf ( R_19a9_1486eed8 , n89534 );
buf ( R_6ec_13c03b58 , n89535 );
buf ( R_b71_140afd78 , n89560 );
buf ( R_d0b_1587d158 , n89561 );
buf ( R_1190_13c09198 , n89562 );
buf ( R_132a_13d44bb8 , C0 );
buf ( R_17af_123b9d58 , n89563 );
buf ( R_1949_140b51d8 , n89613 );
buf ( R_815_158140f8 , n89669 );
buf ( R_a48_13bed6b8 , n89670 );
buf ( R_e34_13cd7e38 , n89671 );
buf ( R_1067_13b93ab8 , n89672 );
buf ( R_1453_15ff99c8 , n89673 );
buf ( R_1686_1008c258 , C0 );
buf ( R_af8_148696b8 , n89674 );
buf ( R_d84_156b3e78 , n89675 );
buf ( R_765_13df9678 , n89718 );
buf ( R_1117_140b2398 , n89719 );
buf ( R_13a3_123bd598 , n89720 );
buf ( R_1736_117f1218 , C0 );
buf ( R_19c2_14871098 , C0 );
buf ( R_d3e_14870198 , C0 );
buf ( R_71f_123b6e78 , n89721 );
buf ( R_b3e_11631138 , C0 );
buf ( R_115d_1008bd58 , n89736 );
buf ( R_135d_13cd9d78 , n89779 );
buf ( R_177c_11629258 , n89780 );
buf ( R_197c_13bec8f8 , n89781 );
buf ( R_96e_1162bff8 , C0 );
buf ( R_f0e_17010f68 , C0 );
buf ( R_8ef_13dd96d8 , n89782 );
buf ( R_f8d_13cd51d8 , n89788 );
buf ( R_152d_13d1f8d8 , n89844 );
buf ( R_15ac_12fc1418 , n89845 );
buf ( R_ee8_13d55658 , n89846 );
buf ( R_994_13c086f8 , n89847 );
buf ( R_8c9_1162f838 , n89863 );
buf ( R_fb3_11c6c7b8 , n89864 );
buf ( R_1507_14b218f8 , n89865 );
buf ( R_15d2_11c6e978 , C0 );
buf ( R_ed3_13b93018 , n89866 );
buf ( R_9a9_140ac3f8 , n89884 );
buf ( R_8b4_150e2e38 , n89885 );
buf ( R_fc8_14875238 , n89886 );
buf ( R_14f2_13cd1718 , C0 );
buf ( R_15e7_150e0e58 , n89887 );
buf ( R_c1a_13d3c198 , C0 );
buf ( R_5fb_156b22f8 , n89888 );
buf ( R_643_117ea698 , n89889 );
buf ( R_c62_1162c598 , C0 );
buf ( R_1239_15817938 , n89914 );
buf ( R_1281_158887d8 , n89965 );
buf ( R_1858_13bea9b8 , n89966 );
buf ( R_18a0_123bfcf8 , n89967 );
buf ( R_98c_13c21f18 , n89968 );
buf ( R_ef0_13d51418 , n89969 );
buf ( R_8d1_12fc06f8 , n89985 );
buf ( R_fab_14a127f8 , n89986 );
buf ( R_150f_15817398 , n89987 );
buf ( R_15ca_156b71b8 , C0 );
buf ( R_c95_123be2b8 , n90030 );
buf ( R_be7_1162d858 , n90031 );
buf ( R_5c8_15feeca8 , n90032 );
buf ( R_676_13d37e18 , C0 );
buf ( R_1206_13ddcc98 , C0 );
buf ( R_12b4_10087938 , n90033 );
buf ( R_1825_1486a298 , n90047 );
buf ( R_18d3_17018f88 , n90048 );
buf ( R_d5b_150e0958 , n90049 );
buf ( R_b21_14b21e98 , n90064 );
buf ( R_73c_13bec858 , n90065 );
buf ( R_1140_13b98798 , n90066 );
buf ( R_137a_13dd7018 , C0 );
buf ( R_175f_15ff7f88 , n90067 );
buf ( R_1999_117f2118 , n90077 );
buf ( R_d4a_13df40d8 , C0 );
buf ( R_b32_13c268d8 , C0 );
buf ( R_72b_11632c18 , n90078 );
buf ( R_1151_11638898 , n90093 );
buf ( R_1369_117f5138 , n90136 );
buf ( R_1770_124c2a58 , n90137 );
buf ( R_1988_150dfaf8 , n90138 );
buf ( R_db1_13bf06d8 , n90181 );
buf ( R_792_13ccb638 , C0 );
buf ( R_acb_13d2a378 , n90182 );
buf ( R_10ea_13d2b598 , C0 );
buf ( R_13d0_1700b388 , n90183 );
buf ( R_1709_1162a298 , n90200 );
buf ( R_19ef_150de1f8 , n90201 );
buf ( R_ae3_14b24738 , n90202 );
buf ( R_d99_156abef8 , n90245 );
buf ( R_77a_13c0f3b8 , C0 );
buf ( R_1102_11632358 , C0 );
buf ( R_13b8_13c29c18 , n90246 );
buf ( R_1721_14870f58 , n90261 );
buf ( R_19d7_13de38b8 , n90262 );
buf ( R_6d8_1580ebf8 , n90263 );
buf ( R_566_140b4f58 , n90264 );
buf ( R_cf7_13d26778 , n90265 );
buf ( R_b85_13df3958 , n90290 );
buf ( R_11a4_140b1178 , n90291 );
buf ( R_1316_13c24718 , C0 );
buf ( R_17c3_13df1e78 , n90292 );
buf ( R_1935_14a13798 , n90342 );
buf ( R_a0d_14a0f198 , n90349 );
buf ( R_850_1700cbe8 , n90350 );
buf ( R_e6f_117ee6f8 , n90351 );
buf ( R_102c_156ae3d8 , n90352 );
buf ( R_148e_17014208 , C0 );
buf ( R_164b_123b8638 , n90353 );
buf ( R_f2f_13ccded8 , n90354 );
buf ( R_910_158144b8 , n90355 );
buf ( R_94d_13de1dd8 , n90377 );
buf ( R_f6c_140aca38 , n90378 );
buf ( R_154e_158131f8 , C0 );
buf ( R_158b_123b5078 , n90379 );
buf ( R_70c_1162a338 , n90380 );
buf ( R_b51_13df4c18 , n90415 );
buf ( R_d2b_123bacf8 , n90416 );
buf ( R_1170_13ddca18 , n90417 );
buf ( R_134a_123bdb38 , C0 );
buf ( R_178f_14a0df78 , n90418 );
buf ( R_1969_13c0e918 , n90428 );
buf ( R_ec1_13c0ddd8 , n90477 );
buf ( R_8a2_13dd9638 , C0 );
buf ( R_9bb_14a13d38 , n90478 );
buf ( R_fda_14876098 , C0 );
buf ( R_14e0_117ea9b8 , n90479 );
buf ( R_15f9_13d4fcf8 , n90495 );
buf ( R_d3b_150e4a58 , n90496 );
buf ( R_71c_150dba98 , n90497 );
buf ( R_b41_100844b8 , n90511 );
buf ( R_1160_14a16498 , n90512 );
buf ( R_135a_156b8838 , C0 );
buf ( R_177f_13ccedd8 , n90513 );
buf ( R_1979_156ad7f8 , n90523 );
buf ( R_80a_11c686b8 , C0 );
buf ( R_a53_13d54ed8 , n90524 );
buf ( R_e29_124c3138 , n90567 );
buf ( R_1072_13d5c598 , C0 );
buf ( R_1448_156b5098 , n90568 );
buf ( R_1691_13bf8478 , n90585 );
buf ( R_1a67_13d3a898 , n90586 );
buf ( R_aa1_13ccbd18 , n90611 );
buf ( R_7bc_13ccc218 , n90612 );
buf ( R_ddb_15812618 , n90613 );
buf ( R_10c0_15816d58 , n90614 );
buf ( R_13fa_14b29a58 , C0 );
buf ( R_16df_10084eb8 , n90615 );
buf ( R_1a19_11c70a98 , n90621 );
buf ( R_a1e_13de1338 , C0 );
buf ( R_83f_123bc5f8 , n90622 );
buf ( R_e5e_13c25258 , C0 );
buf ( R_103d_123b2738 , n90645 );
buf ( R_147d_13d53e98 , n90688 );
buf ( R_165c_123b57f8 , n90689 );
buf ( R_c74_14b242d8 , n90690 );
buf ( R_c08_13ded7d8 , n90691 );
buf ( R_5e9_15816178 , n90734 );
buf ( R_655_13c026b8 , n90777 );
buf ( R_1227_123b72d8 , n90778 );
buf ( R_1293_1008c6b8 , n90779 );
buf ( R_1846_13c22af8 , C0 );
buf ( R_18b2_150dd4d8 , C0 );
buf ( R_a14_11632038 , n90780 );
buf ( R_849_123c1af8 , n90829 );
buf ( R_e68_15887658 , n90830 );
buf ( R_1033_13bf8518 , n90831 );
buf ( R_1487_1007fc38 , n90832 );
buf ( R_1652_11635418 , C0 );
buf ( R_68e_11630eb8 , C0 );
buf ( R_bcf_1486c4f8 , n90833 );
buf ( R_cad_150e5c78 , n90876 );
buf ( R_5b0_13d20c38 , n90882 );
buf ( R_11ee_13df5938 , C0 );
buf ( R_12cc_156aee78 , n90883 );
buf ( R_180d_13d29dd8 , n90897 );
buf ( R_18eb_13cd2bb8 , n90898 );
buf ( R_7e9_13b903b8 , n90947 );
buf ( R_e08_14a11498 , n90948 );
buf ( R_a74_13c02a78 , n90949 );
buf ( R_1093_123bddb8 , n90950 );
buf ( R_1427_1580dd98 , n90951 );
buf ( R_16b2_123b89f8 , C0 );
buf ( R_1a46_150dff58 , C0 );
buf ( R_c81_140ac718 , n90994 );
buf ( R_bfb_117e8f78 , n90995 );
buf ( R_5dc_13cd21b8 , n90996 );
buf ( R_662_11c6af58 , C0 );
buf ( R_121a_13dd6bb8 , C0 );
buf ( R_12a0_156af7d8 , n90997 );
buf ( R_1839_10083a18 , n91012 );
buf ( R_18bf_13cd63f8 , n91013 );
buf ( R_d4d_14b1c218 , n91056 );
buf ( R_b2f_14a168f8 , n91057 );
buf ( R_72e_15885178 , C0 );
buf ( R_114e_14866878 , C0 );
buf ( R_136c_13d5ce58 , n91058 );
buf ( R_176d_15883e18 , n91091 );
buf ( R_198b_123ba938 , n91092 );
buf ( R_bb0_11635198 , n91093 );
buf ( R_6ad_14b295f8 , n91136 );
buf ( R_591_123b56b8 , n91137 );
buf ( R_ccc_13c02f78 , n91138 );
buf ( R_11cf_13dedd78 , n91139 );
buf ( R_12eb_156ab598 , n91140 );
buf ( R_17ee_117f2a78 , C0 );
buf ( R_190a_1162b238 , C0 );
buf ( R_7d4_14a0fe18 , n91141 );
buf ( R_df3_14b1e478 , n91142 );
buf ( R_a89_13dd9278 , n91183 );
buf ( R_10a8_13d52958 , n91184 );
buf ( R_1412_11c6f198 , C0 );
buf ( R_16c7_13d27d58 , n91185 );
buf ( R_1a31_140b9d78 , n91192 );
buf ( R_c19_1700d408 , n91242 );
buf ( R_5fa_13df88b8 , C0 );
buf ( R_644_13d23938 , n91243 );
buf ( R_c63_1162e258 , n91244 );
buf ( R_1238_13df9a38 , n91245 );
buf ( R_1282_13c2acf8 , C0 );
buf ( R_1857_13cd2ed8 , n91246 );
buf ( R_18a1_156aefb8 , n91271 );
buf ( R_6f0_140ae658 , n91272 );
buf ( R_b6d_123b4178 , n91297 );
buf ( R_d0f_150df0f8 , n91298 );
buf ( R_118c_14a17898 , n91299 );
buf ( R_132e_13bed758 , C0 );
buf ( R_17ab_13cd0d18 , n91300 );
buf ( R_194d_1008c438 , n91350 );
buf ( R_802_13d3e5d8 , C0 );
buf ( R_e21_14a0aaf8 , n91393 );
buf ( R_a5b_13bf7e38 , n91394 );
buf ( R_107a_13d1ed98 , C0 );
buf ( R_1440_124c4d58 , n91395 );
buf ( R_1699_140b0318 , n91412 );
buf ( R_1a5f_124c5618 , n91413 );
buf ( R_8fc_13bebd18 , n91414 );
buf ( R_961_12fbe358 , n91431 );
buf ( R_f1b_13ddafd8 , n91432 );
buf ( R_f80_1486f478 , n91433 );
buf ( R_153a_116341f8 , C0 );
buf ( R_159f_1008d338 , n91434 );
buf ( R_ada_15812f78 , C0 );
buf ( R_da2_156b5ef8 , C0 );
buf ( R_783_123ba898 , n91435 );
buf ( R_10f9_123b7a58 , n91463 );
buf ( R_13c1_13d3bfb8 , n91506 );
buf ( R_1718_156b8018 , n91507 );
buf ( R_19e0_13dd4ef8 , n91508 );
buf ( R_6cb_117f2258 , n91509 );
buf ( R_573_1162dfd8 , n91510 );
buf ( R_cea_13d5be18 , C0 );
buf ( R_b92_13c01998 , C0 );
buf ( R_11b1_1700a208 , n91525 );
buf ( R_1309_117e8898 , n91568 );
buf ( R_17d0_156b8d38 , n91569 );
buf ( R_1928_14a0f738 , n91570 );
buf ( R_eb1_156b8f18 , n91619 );
buf ( R_892_11c69018 , C0 );
buf ( R_9cb_13bed1b8 , n91620 );
buf ( R_fea_13d2b3b8 , C0 );
buf ( R_14d0_13ccf698 , n91621 );
buf ( R_1609_13cd30b8 , n91637 );
buf ( R_67f_13cd88d8 , n91638 );
buf ( R_c9e_1580ee78 , C0 );
buf ( R_bde_123b3138 , C0 );
buf ( R_5bf_117f0b38 , n91639 );
buf ( R_11fd_1162f3d8 , n91671 );
buf ( R_12bd_13bf9698 , n91721 );
buf ( R_181c_13bf7758 , n91722 );
buf ( R_18dc_15817258 , n91723 );
buf ( R_c8c_13b97258 , n91724 );
buf ( R_bf0_13c26d38 , n91725 );
buf ( R_5d1_14875af8 , n91768 );
buf ( R_66d_1700eda8 , n91811 );
buf ( R_120f_156b0a98 , n91812 );
buf ( R_12ab_1486c278 , n91813 );
buf ( R_182e_116366d8 , C0 );
buf ( R_18ca_11c708b8 , C0 );
buf ( R_f2e_13dddb98 , C0 );
buf ( R_90f_13b8e3d8 , n91814 );
buf ( R_94e_117f3c98 , C0 );
buf ( R_f6d_13bf7a78 , n91830 );
buf ( R_154d_13df8c78 , n91879 );
buf ( R_158c_13d278f8 , n91880 );
buf ( R_702_13de3598 , C0 );
buf ( R_b5b_13d45bf8 , n91881 );
buf ( R_d21_156ac038 , n91924 );
buf ( R_117a_14b292d8 , C0 );
buf ( R_1340_123bbab8 , n91925 );
buf ( R_1799_13df1018 , n91960 );
buf ( R_195f_13b92e38 , n91961 );
buf ( R_d38_156afaf8 , n91962 );
buf ( R_719_13d1d498 , n92005 );
buf ( R_b44_13df7238 , n92006 );
buf ( R_1163_13b91358 , n92007 );
buf ( R_1357_13d5bcd8 , n92008 );
buf ( R_1782_1486c138 , C0 );
buf ( R_1976_14b1de38 , C0 );
buf ( R_695_13b93b58 , n92051 );
buf ( R_bc8_13dfb3d8 , n92052 );
buf ( R_cb4_15817078 , n92053 );
buf ( R_5a9_156b6998 , n92059 );
buf ( R_11e7_13bf3298 , n92060 );
buf ( R_12d3_14b28338 , n92061 );
buf ( R_1806_123b6dd8 , C0 );
buf ( R_18f2_13d40338 , C0 );
buf ( R_a06_158876f8 , C0 );
buf ( R_857_14874dd8 , n92062 );
buf ( R_e76_13bf0958 , C0 );
buf ( R_1025_13d59438 , n92085 );
buf ( R_1495_14870238 , n92128 );
buf ( R_1644_15ff4d88 , n92129 );
buf ( R_6fb_156b9378 , n92130 );
buf ( R_b62_123bb298 , C0 );
buf ( R_d1a_117ee1f8 , C0 );
buf ( R_1181_148748d8 , n92144 );
buf ( R_1339_1580de38 , n92187 );
buf ( R_17a0_13dd7478 , n92188 );
buf ( R_1958_156ae5b8 , n92189 );
buf ( R_97a_117eaff8 , C0 );
buf ( R_f02_13d538f8 , C0 );
buf ( R_8e3_13c107b8 , n92190 );
buf ( R_f99_1580efb8 , n92199 );
buf ( R_1521_148676d8 , n92248 );
buf ( R_15b8_13b93e78 , n92249 );
buf ( R_829_13b954f8 , n92298 );
buf ( R_a34_156b03b8 , n92299 );
buf ( R_e48_15813d38 , n92300 );
buf ( R_1053_13cd3478 , n92301 );
buf ( R_1467_13b8be58 , n92302 );
buf ( R_1672_13cd1df8 , C0 );
buf ( R_e89_13de0078 , n92351 );
buf ( R_9f3_156b0598 , n92352 );
buf ( R_86a_13b94378 , C0 );
buf ( R_1012_123bf618 , C0 );
buf ( R_14a8_13becdf8 , n92353 );
buf ( R_1631_1486c9f8 , n92370 );
buf ( R_acd_1008bfd8 , n92385 );
buf ( R_daf_123b59d8 , n92386 );
buf ( R_790_13d2bd18 , n92387 );
buf ( R_10ec_1700b6a8 , n92388 );
buf ( R_13ce_13df2a58 , C0 );
buf ( R_170b_14b26178 , n92389 );
buf ( R_19ed_148709b8 , n92395 );
buf ( R_a31_13cd7d98 , n92403 );
buf ( R_82c_140b1e98 , n92404 );
buf ( R_e4b_116316d8 , n92405 );
buf ( R_1050_13d3d138 , n92406 );
buf ( R_146a_123bd318 , C0 );
buf ( R_166f_140ad118 , n92407 );
buf ( R_eac_1007f418 , n92408 );
buf ( R_88d_13bf99b8 , n92424 );
buf ( R_9d0_17010748 , n92425 );
buf ( R_fef_1580b138 , n92426 );
buf ( R_14cb_13d44258 , n92427 );
buf ( R_160e_11632a38 , C0 );
buf ( R_826_13c24cb8 , C0 );
buf ( R_a37_158112b8 , n92428 );
buf ( R_e45_15fee168 , n92471 );
buf ( R_1056_15fedc68 , C0 );
buf ( R_1464_13d3fa78 , n92472 );
buf ( R_1675_14b28dd8 , n92489 );
buf ( R_eb6_11c69518 , C0 );
buf ( R_897_11c69338 , n92490 );
buf ( R_9c6_156ad258 , C0 );
buf ( R_fe5_14b1f4b8 , n92507 );
buf ( R_14d5_14871a98 , n92550 );
buf ( R_1604_13beed38 , n92551 );
buf ( R_9ef_14a126b8 , n92552 );
buf ( R_e8d_13c07578 , n92601 );
buf ( R_86e_13ded738 , C0 );
buf ( R_100e_100810d8 , C0 );
buf ( R_14ac_13cce158 , n92602 );
buf ( R_162d_13c0adb8 , n92619 );
buf ( R_7cb_14a0acd8 , n92620 );
buf ( R_dea_123c0798 , C0 );
buf ( R_a92_13d25238 , C0 );
buf ( R_10b1_13d55478 , n92635 );
buf ( R_1409_1587f638 , n92678 );
buf ( R_16d0_13c02ed8 , n92679 );
buf ( R_1a28_14a12398 , n92680 );
buf ( R_ee0_13d1ffb8 , n92681 );
buf ( R_99c_14a0f418 , n92682 );
buf ( R_8c1_14b25818 , n92699 );
buf ( R_fbb_123b70f8 , n92700 );
buf ( R_14ff_1580bf98 , n92701 );
buf ( R_15da_140ba138 , C0 );
buf ( R_687_14b23fb8 , n92702 );
buf ( R_bd6_13dd71f8 , C0 );
buf ( R_ca6_123bd098 , C0 );
buf ( R_5b7_117e8cf8 , n92703 );
buf ( R_11f5_15815318 , n92735 );
buf ( R_12c5_14a0f7d8 , n92785 );
buf ( R_1814_170116e8 , n92786 );
buf ( R_18e4_12fc1d78 , n92787 );
buf ( R_812_12fc0018 , C0 );
buf ( R_a4b_13bf22f8 , n92788 );
buf ( R_e31_13bee338 , n92831 );
buf ( R_106a_13d56a58 , C0 );
buf ( R_1450_1580a738 , n92832 );
buf ( R_1689_14a0c218 , n92849 );
buf ( R_e85_156aa878 , n92898 );
buf ( R_9f7_13d246f8 , n92899 );
buf ( R_866_15ffb868 , C0 );
buf ( R_1016_156af698 , C0 );
buf ( R_14a4_11c6ec98 , n92900 );
buf ( R_1635_15ff7588 , n92917 );
buf ( R_8ee_140ae338 , C0 );
buf ( R_96f_13d3b8d8 , n92918 );
buf ( R_f0d_13d4fa78 , n92924 );
buf ( R_f8e_13d541b8 , C0 );
buf ( R_152c_156b2258 , n92925 );
buf ( R_15ad_13d58218 , n92941 );
buf ( R_9de_124c3458 , C0 );
buf ( R_e9e_123b9038 , C0 );
buf ( R_87f_117f0958 , n92942 );
buf ( R_ffd_13c27f58 , n92959 );
buf ( R_14bd_13cd71b8 , n93002 );
buf ( R_161c_156b6178 , n93003 );
buf ( R_aec_14866b98 , n93004 );
buf ( R_d90_10081718 , n93005 );
buf ( R_771_1007ee78 , n93048 );
buf ( R_110b_14b24f58 , n93049 );
buf ( R_13af_158110d8 , n93050 );
buf ( R_172a_11c6feb8 , C0 );
buf ( R_19ce_11c6fc38 , C0 );
buf ( R_6d4_15ff47e8 , n93051 );
buf ( R_56a_17018268 , n93052 );
buf ( R_cf3_150e21b8 , n93053 );
buf ( R_b89_13cd67b8 , n93078 );
buf ( R_11a8_13c0ab38 , n93079 );
buf ( R_1312_15881758 , C0 );
buf ( R_17c7_1580cf38 , n93080 );
buf ( R_1931_11c6b4f8 , n93130 );
buf ( R_7be_13d51918 , C0 );
buf ( R_ddd_10083fb8 , n93173 );
buf ( R_a9f_140b7b18 , n93174 );
buf ( R_10be_1162c138 , C0 );
buf ( R_13fc_13b967b8 , n93175 );
buf ( R_16dd_15ffb728 , n93193 );
buf ( R_1a1b_13d3ab18 , n93194 );
buf ( R_a2e_1580aeb8 , C0 );
buf ( R_82f_14b26cb8 , n93195 );
buf ( R_e4e_13dec798 , C0 );
buf ( R_104d_13de2af8 , n93213 );
buf ( R_146d_156b1998 , n93256 );
buf ( R_166c_117f5958 , n93257 );
buf ( R_d50_156b51d8 , n93258 );
buf ( R_b2c_12fc0478 , n93259 );
buf ( R_731_15ffaa08 , n93302 );
buf ( R_114b_13ddbed8 , n93303 );
buf ( R_136f_11c6c718 , n93304 );
buf ( R_176a_11628f38 , C0 );
buf ( R_198e_150e3518 , C0 );
buf ( R_ed9_15ff7948 , n93353 );
buf ( R_9a3_13c1fad8 , n93354 );
buf ( R_8ba_116386b8 , C0 );
buf ( R_fc2_1700f7a8 , C0 );
buf ( R_14f8_117f15d8 , n93355 );
buf ( R_15e1_150dcd58 , n93371 );
buf ( R_b16_13c1c1f8 , C0 );
buf ( R_d66_13b8b1d8 , C0 );
buf ( R_747_158864d8 , n93372 );
buf ( R_1135_156b68f8 , n93397 );
buf ( R_1385_1580b278 , n93440 );
buf ( R_1754_156add98 , n93441 );
buf ( R_19a4_13d4fd98 , n93442 );
buf ( R_823_11c6f2d8 , n93443 );
buf ( R_a3a_14871318 , C0 );
buf ( R_e42_156ade38 , C0 );
buf ( R_1059_13c0f318 , n93465 );
buf ( R_1461_14a1a138 , n93508 );
buf ( R_1678_14a0fd78 , n93509 );
buf ( R_8d9_158837d8 , n93526 );
buf ( R_984_15882d38 , n93527 );
buf ( R_ef8_15816998 , n93528 );
buf ( R_fa3_15815458 , n93529 );
buf ( R_1517_156ad898 , n93530 );
buf ( R_15c2_11630c38 , C0 );
buf ( R_af3_13beae18 , n93531 );
buf ( R_d89_117e8938 , n93574 );
buf ( R_76a_123bceb8 , C0 );
buf ( R_1112_13c20c58 , C0 );
buf ( R_13a8_117f4a58 , n93575 );
buf ( R_1731_1008a818 , n93599 );
buf ( R_19c7_13d38bd8 , n93600 );
buf ( R_b04_156aed38 , n93601 );
buf ( R_d78_13cd7758 , n93602 );
buf ( R_759_11629938 , n93645 );
buf ( R_1123_15ffb908 , n93646 );
buf ( R_1397_13d37a58 , n93647 );
buf ( R_1742_13d237f8 , C0 );
buf ( R_19b6_14b20778 , C0 );
buf ( R_c64_13c1fdf8 , n93648 );
buf ( R_c18_12fc23b8 , n93649 );
buf ( R_5f9_13b8f238 , n93692 );
buf ( R_645_140b2118 , n93735 );
buf ( R_1237_1162dad8 , n93736 );
buf ( R_1283_14a18798 , n93737 );
buf ( R_1856_117f4878 , C0 );
buf ( R_18a2_13d53998 , C0 );
buf ( R_f2d_100818f8 , n93753 );
buf ( R_90e_11629898 , C0 );
buf ( R_94f_15888738 , n93754 );
buf ( R_f6e_14a188d8 , C0 );
buf ( R_154c_14a147d8 , n93755 );
buf ( R_158d_15ff0a08 , n93770 );
buf ( R_9eb_117ef2d8 , n93771 );
buf ( R_e91_1580e3d8 , n93827 );
buf ( R_872_13c0c7f8 , C0 );
buf ( R_100a_117f81f8 , C0 );
buf ( R_14b0_124c2f58 , n93828 );
buf ( R_1629_14a0b6d8 , n93845 );
buf ( R_656_15886bb8 , C0 );
buf ( R_c75_156b0db8 , n93888 );
buf ( R_c07_124c4cb8 , n93889 );
buf ( R_5e8_1162f298 , n93890 );
buf ( R_1226_13b8e018 , C0 );
buf ( R_1294_13b91ad8 , n93891 );
buf ( R_1845_13cd83d8 , n93906 );
buf ( R_18b3_13d1e118 , n93907 );
buf ( R_ba0_156b4698 , n93908 );
buf ( R_6bd_13c0ec38 , n93951 );
buf ( R_581_13d1d8f8 , n93952 );
buf ( R_cdc_13cd9378 , n93953 );
buf ( R_11bf_123b6c98 , n93954 );
buf ( R_12fb_150e3018 , n93955 );
buf ( R_17de_14b20458 , C0 );
buf ( R_191a_123b2cd8 , C0 );
buf ( R_d5e_14a10278 , C0 );
buf ( R_b1e_13df7418 , C0 );
buf ( R_73f_1587b998 , n93956 );
buf ( R_113d_13d58498 , n93986 );
buf ( R_137d_14a11b78 , n94029 );
buf ( R_175c_1587b218 , n94030 );
buf ( R_199c_17017408 , n94031 );
buf ( R_b09_15884f98 , n94045 );
buf ( R_d73_1580b4f8 , n94046 );
buf ( R_754_15811d58 , n94047 );
buf ( R_1128_10084d78 , n94048 );
buf ( R_1392_14a15db8 , C0 );
buf ( R_1747_17018588 , n94049 );
buf ( R_19b1_13dd9f98 , n94059 );
buf ( R_d35_14a11858 , n94102 );
buf ( R_716_156b9c38 , C0 );
buf ( R_b47_140af4b8 , n94103 );
buf ( R_1166_13ccdcf8 , C0 );
buf ( R_1354_13d41738 , n94104 );
buf ( R_1785_1162d218 , n94132 );
buf ( R_1973_14a18338 , n94133 );
buf ( R_a2b_13c1e6d8 , n94134 );
buf ( R_832_13df5c58 , C0 );
buf ( R_e51_156ab278 , n94177 );
buf ( R_104a_14a108b8 , C0 );
buf ( R_1470_15887bf8 , n94178 );
buf ( R_1669_158828d8 , n94195 );
buf ( R_e81_1007dc58 , n94244 );
buf ( R_9fb_1486fb58 , n94245 );
buf ( R_862_156ab138 , C0 );
buf ( R_101a_13d5a798 , C0 );
buf ( R_14a0_13d38818 , n94246 );
buf ( R_1639_1162abf8 , n94263 );
buf ( R_ba5_140b4af8 , n94288 );
buf ( R_6b8_1580d898 , n94289 );
buf ( R_586_15ff8488 , n94290 );
buf ( R_cd7_156b7e38 , n94291 );
buf ( R_11c4_117ecad8 , n94292 );
buf ( R_12f6_17015ba8 , C0 );
buf ( R_17e3_13c1dd78 , n94293 );
buf ( R_1915_14a17f78 , n94344 );
buf ( R_aff_140aba98 , n94345 );
buf ( R_d7d_148714f8 , n94388 );
buf ( R_75e_10084418 , C0 );
buf ( R_111e_11635918 , C0 );
buf ( R_139c_1580e0b8 , n94389 );
buf ( R_173d_13deffd8 , n94405 );
buf ( R_19bb_13df9df8 , n94406 );
buf ( R_7dd_13d28898 , n94455 );
buf ( R_dfc_156b9ff8 , n94456 );
buf ( R_a80_13ddc8d8 , n94457 );
buf ( R_109f_13cd2cf8 , n94458 );
buf ( R_141b_12fc10f8 , n94459 );
buf ( R_16be_13bf0098 , C0 );
buf ( R_1a3a_156b79d8 , C0 );
buf ( R_9d5_15ff1908 , n94476 );
buf ( R_ea7_14a124d8 , n94477 );
buf ( R_888_13deebd8 , n94478 );
buf ( R_ff4_13cd7b18 , n94479 );
buf ( R_14c6_13cd5d18 , C0 );
buf ( R_1613_123bc198 , n94480 );
buf ( R_677_13c0c758 , n94481 );
buf ( R_c96_13c0d838 , C0 );
buf ( R_be6_1162cf98 , C0 );
buf ( R_5c7_1162f1f8 , n94482 );
buf ( R_1205_156b94b8 , n94507 );
buf ( R_12b5_158816b8 , n94557 );
buf ( R_1824_13c04f58 , n94558 );
buf ( R_18d4_13beb958 , n94559 );
buf ( R_f1a_124c4f38 , C0 );
buf ( R_8fb_13c1e9f8 , n94560 );
buf ( R_962_14a15ef8 , C0 );
buf ( R_f81_1580d438 , n94576 );
buf ( R_1539_14b267b8 , n94625 );
buf ( R_15a0_15ff32a8 , n94626 );
buf ( R_d28_156b3fb8 , n94627 );
buf ( R_709_117ea4b8 , n94670 );
buf ( R_b54_13c04c38 , n94671 );
buf ( R_1173_15810778 , n94672 );
buf ( R_1347_13dd5f38 , n94673 );
buf ( R_1792_13d39858 , C0 );
buf ( R_1966_12fc2098 , C0 );
buf ( R_a1b_123c17d8 , n94674 );
buf ( R_842_13bf4738 , C0 );
buf ( R_e61_13cd0958 , n94723 );
buf ( R_103a_13ccdbb8 , C0 );
buf ( R_1480_117f1e98 , n94724 );
buf ( R_1659_13c1fcb8 , n94741 );
buf ( R_820_17013088 , n94742 );
buf ( R_a3d_11c6bc78 , n94791 );
buf ( R_e3f_123c0e78 , n94792 );
buf ( R_105c_13dd87d8 , n94793 );
buf ( R_145e_13d5a3d8 , C0 );
buf ( R_167b_14a19878 , n94794 );
buf ( R_ebb_13def998 , n94795 );
buf ( R_89c_1486e898 , n94796 );
buf ( R_9c1_13cd04f8 , n94814 );
buf ( R_fe0_15fee7a8 , n94815 );
buf ( R_14da_13b95818 , C0 );
buf ( R_15ff_117f1538 , n94816 );
buf ( R_8d0_13ccd078 , n94817 );
buf ( R_98d_13cceab8 , n94835 );
buf ( R_eef_15ff2308 , n94836 );
buf ( R_fac_13df65b8 , n94837 );
buf ( R_150e_13bed398 , C0 );
buf ( R_15cb_1580a558 , n94838 );
buf ( R_663_13c24218 , n94839 );
buf ( R_c82_11633bb8 , C0 );
buf ( R_bfa_117f1d58 , C0 );
buf ( R_5db_13c0d798 , n94840 );
buf ( R_1219_156b0f98 , n94865 );
buf ( R_12a1_15811e98 , n94915 );
buf ( R_1838_123c2098 , n94916 );
buf ( R_18c0_13ddb258 , n94917 );
buf ( R_bbb_13c08dd8 , n94918 );
buf ( R_6a2_14870cd8 , C0 );
buf ( R_59c_1700ffc8 , n94924 );
buf ( R_cc1_13d5b0f8 , n94967 );
buf ( R_11da_14b1dcf8 , C0 );
buf ( R_12e0_14b29c38 , n94968 );
buf ( R_17f9_13ddb438 , n94983 );
buf ( R_18ff_1162d538 , n94984 );
buf ( R_ecc_123bde58 , n94985 );
buf ( R_9b0_1587f458 , n94986 );
buf ( R_8ad_10082e38 , n95002 );
buf ( R_fcf_14a0e798 , n95003 );
buf ( R_14eb_140ad258 , n95004 );
buf ( R_15ee_117f3158 , C0 );
buf ( R_d13_13c25e38 , n95005 );
buf ( R_6f4_156b4918 , n95006 );
buf ( R_b69_11c6e8d8 , n95038 );
buf ( R_1188_13cd35b8 , n95039 );
buf ( R_1332_11637d58 , C0 );
buf ( R_17a7_117f6a38 , n95040 );
buf ( R_1951_156b6b78 , n95090 );
buf ( R_acf_13d503d8 , n95091 );
buf ( R_dad_13cd3838 , n95134 );
buf ( R_78e_13b929d8 , C0 );
buf ( R_10ee_1587c438 , C0 );
buf ( R_13cc_1587b3f8 , n95135 );
buf ( R_170d_12fbf9d8 , n95152 );
buf ( R_19eb_15ff53c8 , n95153 );
buf ( R_8c8_12fbe038 , n95154 );
buf ( R_ee7_13c03dd8 , n95155 );
buf ( R_995_13d50518 , n95173 );
buf ( R_fb4_156b0e58 , n95174 );
buf ( R_1506_156b9e18 , C0 );
buf ( R_15d3_123b5ed8 , n95175 );
buf ( R_b9b_13dfa118 , n95176 );
buf ( R_6c2_14b1d618 , C0 );
buf ( R_57c_13d464b8 , n95177 );
buf ( R_ce1_13d27358 , n95220 );
buf ( R_11ba_13cda458 , C0 );
buf ( R_1300_13dec478 , n95221 );
buf ( R_17d9_156af918 , n95244 );
buf ( R_191f_14a0d578 , n95245 );
buf ( R_7e4_117f6c18 , n95246 );
buf ( R_e03_13b8c718 , n95247 );
buf ( R_a79_13d52db8 , n95275 );
buf ( R_1098_13cd2438 , n95276 );
buf ( R_1422_13cd7f78 , C0 );
buf ( R_16b7_14b28518 , n95277 );
buf ( R_1a41_150e4d78 , n95283 );
buf ( R_ae5_17012048 , n95297 );
buf ( R_d97_1162ab58 , n95298 );
buf ( R_778_13d52098 , n95299 );
buf ( R_1104_13dd7a18 , n95300 );
buf ( R_13b6_14a17118 , C0 );
buf ( R_1723_13d50018 , n95301 );
buf ( R_19d5_117edc58 , n95311 );
buf ( R_d53_13c0ae58 , n95312 );
buf ( R_b29_13b95c78 , n95327 );
buf ( R_734_14a0f558 , n95328 );
buf ( R_1148_117f6218 , n95329 );
buf ( R_1372_11c6cd58 , C0 );
buf ( R_1767_11c691f8 , n95330 );
buf ( R_1991_13cd58b8 , n95340 );
buf ( R_f2c_15814d78 , n95341 );
buf ( R_90d_158848b8 , n95350 );
buf ( R_950_140b3798 , n95351 );
buf ( R_f6f_14a1a318 , n95352 );
buf ( R_154b_11632218 , n95353 );
buf ( R_158e_14a0b1d8 , C0 );
buf ( R_ec6_13d37b98 , C0 );
buf ( R_8a7_1580e6f8 , n95354 );
buf ( R_9b6_14a0cc18 , C0 );
buf ( R_fd5_1580cc18 , n95371 );
buf ( R_14e5_13b8fd78 , n95414 );
buf ( R_15f4_170165a8 , n95415 );
buf ( R_7c0_100854f8 , n95416 );
buf ( R_ddf_13b92898 , n95417 );
buf ( R_a9d_1162c318 , n95441 );
buf ( R_10bc_140b7d98 , n95442 );
buf ( R_13fe_13cd60d8 , C0 );
buf ( R_16db_156aaf58 , n95443 );
buf ( R_1a1d_13cd9ff8 , n95449 );
buf ( R_7f5_13b9a1d8 , n95498 );
buf ( R_e14_123bf078 , n95499 );
buf ( R_a68_150dbbd8 , n95500 );
buf ( R_1087_1587ad18 , n95501 );
buf ( R_1433_13dd7978 , n95502 );
buf ( R_16a6_13df8458 , C0 );
buf ( R_1a52_11c70778 , C0 );
buf ( R_646_156ad618 , C0 );
buf ( R_c65_10086538 , n95545 );
buf ( R_c17_13ccb3b8 , n95546 );
buf ( R_5f8_1580f418 , n95547 );
buf ( R_1236_1587e558 , C0 );
buf ( R_1284_14a1a458 , n95548 );
buf ( R_1855_10084a58 , n95564 );
buf ( R_18a3_1700b1a8 , n95565 );
buf ( R_69c_156b9058 , n95566 );
buf ( R_bc1_13bee298 , n95592 );
buf ( R_cbb_13ccbbd8 , n95593 );
buf ( R_5a2_15813658 , n95599 );
buf ( R_11e0_1587e878 , n95600 );
buf ( R_12da_14b29d78 , C0 );
buf ( R_17ff_14a10b38 , n95601 );
buf ( R_18f9_14a16718 , n95652 );
buf ( R_adc_156ae6f8 , n95653 );
buf ( R_da0_13bf5db8 , n95654 );
buf ( R_781_13d42f98 , n95697 );
buf ( R_10fb_10085778 , n95698 );
buf ( R_13bf_123bf6b8 , n95699 );
buf ( R_171a_150deb58 , C0 );
buf ( R_19de_117ef918 , C0 );
buf ( R_9e7_13d54578 , n95700 );
buf ( R_e95_13d26ef8 , n95749 );
buf ( R_876_13d41698 , C0 );
buf ( R_1006_13c08f18 , C0 );
buf ( R_14b4_1700e268 , n95750 );
buf ( R_1625_13b96d58 , n95759 );
buf ( R_807_13cd8478 , n95760 );
buf ( R_e26_1700df48 , C0 );
buf ( R_a56_124c4ad8 , C0 );
buf ( R_1075_15883b98 , n95777 );
buf ( R_1445_15880218 , n95820 );
buf ( R_1694_13d218b8 , n95821 );
buf ( R_1a64_13ccac38 , n95822 );
buf ( R_a28_13cd9918 , n95823 );
buf ( R_835_140b35b8 , n95872 );
buf ( R_e54_14a179d8 , n95873 );
buf ( R_1047_14b26df8 , n95874 );
buf ( R_1473_156b60d8 , n95875 );
buf ( R_1666_14a165d8 , C0 );
buf ( R_b0e_14a15818 , C0 );
buf ( R_d6e_14a0c998 , C0 );
buf ( R_74f_13c24678 , n95876 );
buf ( R_112d_1162be18 , n95901 );
buf ( R_138d_13b92258 , n95944 );
buf ( R_174c_116339d8 , n95945 );
buf ( R_19ac_14b1b4f8 , n95946 );
buf ( R_bb5_13cd29d8 , n95971 );
buf ( R_6a8_1162e618 , n95972 );
buf ( R_596_13dd6398 , n95978 );
buf ( R_cc7_123b4b78 , n95979 );
buf ( R_11d4_15ff30c8 , n95980 );
buf ( R_12e6_14a0ff58 , C0 );
buf ( R_17f3_13ddb578 , n95981 );
buf ( R_1905_1486dfd8 , n96032 );
buf ( R_baa_14a15278 , C0 );
buf ( R_6b3_17011288 , n96033 );
buf ( R_58b_140b1c18 , n96034 );
buf ( R_cd2_13d24dd8 , C0 );
buf ( R_11c9_14b25278 , n96050 );
buf ( R_12f1_1587da18 , n96093 );
buf ( R_17e8_1587c078 , n96094 );
buf ( R_1910_12fc0978 , n96095 );
buf ( R_66e_17014348 , C0 );
buf ( R_c8d_123b7ff8 , n96138 );
buf ( R_bef_14a167b8 , n96139 );
buf ( R_5d0_13c1db98 , n96140 );
buf ( R_120e_13c0d518 , C0 );
buf ( R_12ac_13ccaf58 , n96141 );
buf ( R_182d_140b0098 , n96155 );
buf ( R_18cb_123b9e98 , n96156 );
buf ( R_8b3_13c0d298 , n96157 );
buf ( R_ed2_1580c538 , C0 );
buf ( R_9aa_124c51b8 , C0 );
buf ( R_fc9_13b8d118 , n96174 );
buf ( R_14f1_150e8978 , n96223 );
buf ( R_15e8_15884db8 , n96224 );
buf ( R_8e2_13bf6858 , C0 );
buf ( R_97b_150e7a78 , n96225 );
buf ( R_f01_14a13e78 , n96240 );
buf ( R_f9a_116364f8 , C0 );
buf ( R_1520_1162d678 , n96241 );
buf ( R_15b9_13d21a98 , n96257 );
buf ( R_7fa_123bbbf8 , C0 );
buf ( R_e19_13d59ed8 , n96300 );
buf ( R_a63_14a16678 , n96301 );
buf ( R_1082_13c09d78 , C0 );
buf ( R_1438_13bf2398 , n96302 );
buf ( R_16a1_14a16cb8 , n96319 );
buf ( R_1a57_13c28a98 , n96320 );
buf ( R_81d_1580d078 , n96369 );
buf ( R_a40_123bcd78 , n96370 );
buf ( R_e3c_117f2c58 , n96371 );
buf ( R_105f_13de2558 , n96372 );
buf ( R_145b_11633e38 , n96373 );
buf ( R_167e_1486d858 , C0 );
buf ( R_7f0_13b90458 , n96374 );
buf ( R_e0f_140ab138 , n96375 );
buf ( R_a6d_117ee838 , n96403 );
buf ( R_108c_13bf90f8 , n96404 );
buf ( R_142e_11632538 , C0 );
buf ( R_16ab_140b8d38 , n96405 );
buf ( R_1a4d_11c70bd8 , n96411 );
buf ( R_7d6_14b1e3d8 , C0 );
buf ( R_df5_1580eab8 , n96454 );
buf ( R_a87_14a10138 , n96455 );
buf ( R_10a6_117efa58 , C0 );
buf ( R_1414_1162b9b8 , n96456 );
buf ( R_16c5_14a10db8 , n96474 );
buf ( R_1a33_1486ebb8 , n96475 );
buf ( R_f0c_140b21b8 , n96476 );
buf ( R_8ed_11636d18 , n96492 );
buf ( R_970_13c0f818 , n96493 );
buf ( R_f8f_11632fd8 , n96494 );
buf ( R_152b_13beb778 , n96495 );
buf ( R_15ae_123b2eb8 , C0 );
buf ( R_e6b_13b8ded8 , n96496 );
buf ( R_a11_158133d8 , n96541 );
buf ( R_84c_13bef918 , n96542 );
buf ( R_1030_140b72f8 , n96543 );
buf ( R_148a_140b0598 , C0 );
buf ( R_164f_13d52778 , n96544 );
buf ( R_afa_123c0c98 , C0 );
buf ( R_d82_13cd1858 , C0 );
buf ( R_763_1580e298 , n96545 );
buf ( R_1119_1587c118 , n96569 );
buf ( R_13a1_158898b8 , n96612 );
buf ( R_1738_11c6f878 , n96613 );
buf ( R_19c0_1007ded8 , n96614 );
buf ( R_e7d_15811538 , n96663 );
buf ( R_9ff_13d245b8 , n96664 );
buf ( R_85e_13cd3018 , C0 );
buf ( R_101e_13d5d8f8 , C0 );
buf ( R_149c_13d5a978 , n96665 );
buf ( R_163d_13ccd438 , n96682 );
buf ( R_b8d_156aae18 , n96707 );
buf ( R_6d0_1162bb98 , n96708 );
buf ( R_56e_10086e98 , n96709 );
buf ( R_cef_14870eb8 , n96710 );
buf ( R_11ac_13c24498 , n96711 );
buf ( R_130e_14a17758 , C0 );
buf ( R_17cb_14a0e478 , n96712 );
buf ( R_192d_123becb8 , n96762 );
buf ( R_d32_13d20558 , C0 );
buf ( R_713_15882978 , n96763 );
buf ( R_b4a_13d22cb8 , C0 );
buf ( R_1169_123b7c38 , n96778 );
buf ( R_1351_14a14558 , n96821 );
buf ( R_1788_13ccae18 , n96822 );
buf ( R_1970_124c43f8 , n96823 );
buf ( R_7cd_13d58df8 , n96866 );
buf ( R_dec_156ae518 , n96867 );
buf ( R_a90_13dd8058 , n96868 );
buf ( R_10af_117f0818 , n96869 );
buf ( R_140b_1580d1b8 , n96870 );
buf ( R_16ce_117ebe58 , C0 );
buf ( R_1a2a_15810e58 , C0 );
buf ( R_e72_13c1e8b8 , C0 );
buf ( R_a0a_13d54438 , C0 );
buf ( R_853_123bd778 , n96871 );
buf ( R_1029_13cd2898 , n96889 );
buf ( R_1491_117f33d8 , n96932 );
buf ( R_1648_15ff12c8 , n96933 );
buf ( R_80f_13d449d8 , n96934 );
buf ( R_a4e_13b8e798 , C0 );
buf ( R_e2e_13dd57b8 , C0 );
buf ( R_106d_13b8b598 , n96951 );
buf ( R_144d_13cd65d8 , n96994 );
buf ( R_168c_15ff1c28 , n96995 );
buf ( n30987 , RI15b3e9d0_1);
buf ( n30988 , n30987 );
buf ( n30989 , RI15b56850_817);
buf ( n30990 , RI15b51120_631);
not ( n30991 , n30990 );
buf ( n30992 , RI15b51288_634);
buf ( n30993 , RI15b51198_632);
buf ( n30994 , RI15b51210_633);
or ( n30995 , n30993 , n30994 );
nand ( n30996 , n30992 , n30995 );
not ( n30997 , n30996 );
and ( n30998 , n30997 , n30993 );
buf ( n30999 , n30998 );
not ( n31000 , n30996 );
and ( n31001 , n31000 , n30994 );
buf ( n31002 , n31001 );
not ( n31003 , n30996 );
and ( n31004 , n31003 , n30992 );
buf ( n31005 , n31004 );
not ( n31006 , n31005 );
nor ( n31007 , n30991 , n30999 , n31002 , n31006 );
and ( n31008 , n30989 , n31007 );
buf ( n31009 , RI15b4c2d8_464);
buf ( n31010 , RI15b51030_629);
not ( n31011 , n31010 );
and ( n31012 , n31009 , n31011 );
buf ( n31013 , RI15b4c260_463);
buf ( n31014 , RI15b50fb8_628);
not ( n31015 , n31014 );
and ( n31016 , n31013 , n31015 );
buf ( n31017 , RI15b4c1e8_462);
buf ( n31018 , RI15b50f40_627);
not ( n31019 , n31018 );
and ( n31020 , n31017 , n31019 );
buf ( n31021 , RI15b4c170_461);
buf ( n31022 , RI15b50ec8_626);
not ( n31023 , n31022 );
and ( n31024 , n31021 , n31023 );
buf ( n31025 , RI15b4c0f8_460);
buf ( n31026 , RI15b50e50_625);
not ( n31027 , n31026 );
or ( n31028 , n31025 , n31027 );
and ( n31029 , n31023 , n31028 );
and ( n31030 , n31021 , n31028 );
or ( n31031 , n31024 , n31029 , n31030 );
and ( n31032 , n31019 , n31031 );
and ( n31033 , n31017 , n31031 );
or ( n31034 , n31020 , n31032 , n31033 );
and ( n31035 , n31015 , n31034 );
and ( n31036 , n31013 , n31034 );
or ( n31037 , n31016 , n31035 , n31036 );
and ( n31038 , n31011 , n31037 );
and ( n31039 , n31009 , n31037 );
or ( n31040 , n31012 , n31038 , n31039 );
not ( n31041 , n31040 );
not ( n31042 , n31041 );
xor ( n31043 , n31017 , n31019 );
xor ( n31044 , n31043 , n31031 );
xor ( n31045 , n31013 , n31015 );
xor ( n31046 , n31045 , n31034 );
xor ( n31047 , n31009 , n31011 );
xor ( n31048 , n31047 , n31037 );
buf ( n31049 , n31041 );
buf ( n31050 , n31041 );
buf ( n31051 , n31041 );
buf ( n31052 , n31041 );
buf ( n31053 , n31041 );
buf ( n31054 , n31041 );
buf ( n31055 , n31041 );
buf ( n31056 , n31041 );
buf ( n31057 , n31041 );
buf ( n31058 , n31041 );
buf ( n31059 , n31041 );
buf ( n31060 , n31041 );
buf ( n31061 , n31041 );
buf ( n31062 , n31041 );
buf ( n31063 , n31041 );
buf ( n31064 , n31041 );
buf ( n31065 , n31041 );
buf ( n31066 , n31041 );
buf ( n31067 , n31041 );
buf ( n31068 , n31041 );
buf ( n31069 , n31041 );
buf ( n31070 , n31041 );
buf ( n31071 , n31041 );
buf ( n31072 , n31041 );
buf ( n31073 , n31041 );
xor ( n31074 , n31021 , n31023 );
xor ( n31075 , n31074 , n31028 );
or ( n31076 , n31044 , n31046 , n31048 , n31041 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31075 );
and ( n31077 , n31042 , n31076 );
not ( n31078 , n31077 );
buf ( n31079 , RI15b57750_849);
and ( n31080 , n31078 , n31079 );
and ( n31081 , n31022 , n31026 );
and ( n31082 , n31018 , n31081 );
xor ( n31083 , n31014 , n31082 );
and ( n31084 , n31083 , n31077 );
or ( n31085 , n31080 , n31084 );
buf ( n31086 , RI15b4fb90_585);
not ( n31087 , n31010 );
and ( n31088 , n31026 , n31022 , n31018 , n31014 , n31087 );
and ( n31089 , n31086 , n31088 );
buf ( n31090 , RI15b4f7d0_577);
not ( n31091 , n31026 );
and ( n31092 , n31091 , n31022 , n31018 , n31014 , n31087 );
and ( n31093 , n31090 , n31092 );
buf ( n31094 , RI15b4f410_569);
not ( n31095 , n31022 );
and ( n31096 , n31026 , n31095 , n31018 , n31014 , n31087 );
and ( n31097 , n31094 , n31096 );
buf ( n31098 , RI15b4f050_561);
and ( n31099 , n31091 , n31095 , n31018 , n31014 , n31087 );
and ( n31100 , n31098 , n31099 );
buf ( n31101 , RI15b4ec90_553);
not ( n31102 , n31018 );
and ( n31103 , n31026 , n31022 , n31102 , n31014 , n31087 );
and ( n31104 , n31101 , n31103 );
buf ( n31105 , RI15b4e8d0_545);
and ( n31106 , n31091 , n31022 , n31102 , n31014 , n31087 );
and ( n31107 , n31105 , n31106 );
buf ( n31108 , RI15b4e510_537);
and ( n31109 , n31026 , n31095 , n31102 , n31014 , n31087 );
and ( n31110 , n31108 , n31109 );
buf ( n31111 , RI15b4e150_529);
and ( n31112 , n31091 , n31095 , n31102 , n31014 , n31087 );
and ( n31113 , n31111 , n31112 );
buf ( n31114 , RI15b4dd90_521);
nor ( n31115 , n31091 , n31095 , n31102 , n31014 , n31010 );
and ( n31116 , n31114 , n31115 );
buf ( n31117 , RI15b4d9d0_513);
nor ( n31118 , n31026 , n31095 , n31102 , n31014 , n31010 );
and ( n31119 , n31117 , n31118 );
buf ( n31120 , RI15b4d610_505);
nor ( n31121 , n31091 , n31022 , n31102 , n31014 , n31010 );
and ( n31122 , n31120 , n31121 );
buf ( n31123 , RI15b4d250_497);
nor ( n31124 , n31026 , n31022 , n31102 , n31014 , n31010 );
and ( n31125 , n31123 , n31124 );
buf ( n31126 , RI15b4ce90_489);
nor ( n31127 , n31091 , n31095 , n31018 , n31014 , n31010 );
and ( n31128 , n31126 , n31127 );
buf ( n31129 , RI15b4cad0_481);
nor ( n31130 , n31026 , n31095 , n31018 , n31014 , n31010 );
and ( n31131 , n31129 , n31130 );
buf ( n31132 , RI15b4c710_473);
nor ( n31133 , n31091 , n31022 , n31018 , n31014 , n31010 );
and ( n31134 , n31132 , n31133 );
buf ( n31135 , RI15b4c350_465);
nor ( n31136 , n31026 , n31022 , n31018 , n31014 , n31010 );
and ( n31137 , n31135 , n31136 );
or ( n31138 , n31089 , n31093 , n31097 , n31100 , n31104 , n31107 , n31110 , n31113 , n31116 , n31119 , n31122 , n31125 , n31128 , n31131 , n31134 , n31137 );
not ( n31139 , n31138 );
buf ( n31140 , RI15b4fc08_586);
and ( n31141 , n31140 , n31088 );
buf ( n31142 , RI15b4f848_578);
and ( n31143 , n31142 , n31092 );
buf ( n31144 , RI15b4f488_570);
and ( n31145 , n31144 , n31096 );
buf ( n31146 , RI15b4f0c8_562);
and ( n31147 , n31146 , n31099 );
buf ( n31148 , RI15b4ed08_554);
and ( n31149 , n31148 , n31103 );
buf ( n31150 , RI15b4e948_546);
and ( n31151 , n31150 , n31106 );
buf ( n31152 , RI15b4e588_538);
and ( n31153 , n31152 , n31109 );
buf ( n31154 , RI15b4e1c8_530);
and ( n31155 , n31154 , n31112 );
buf ( n31156 , RI15b4de08_522);
and ( n31157 , n31156 , n31115 );
buf ( n31158 , RI15b4da48_514);
and ( n31159 , n31158 , n31118 );
buf ( n31160 , RI15b4d688_506);
and ( n31161 , n31160 , n31121 );
buf ( n31162 , RI15b4d2c8_498);
and ( n31163 , n31162 , n31124 );
buf ( n31164 , RI15b4cf08_490);
and ( n31165 , n31164 , n31127 );
buf ( n31166 , RI15b4cb48_482);
and ( n31167 , n31166 , n31130 );
buf ( n31168 , RI15b4c788_474);
and ( n31169 , n31168 , n31133 );
buf ( n31170 , RI15b4c3c8_466);
and ( n31171 , n31170 , n31136 );
or ( n31172 , n31141 , n31143 , n31145 , n31147 , n31149 , n31151 , n31153 , n31155 , n31157 , n31159 , n31161 , n31163 , n31165 , n31167 , n31169 , n31171 );
buf ( n31173 , RI15b4fc80_587);
and ( n31174 , n31173 , n31088 );
buf ( n31175 , RI15b4f8c0_579);
and ( n31176 , n31175 , n31092 );
buf ( n31177 , RI15b4f500_571);
and ( n31178 , n31177 , n31096 );
buf ( n31179 , RI15b4f140_563);
and ( n31180 , n31179 , n31099 );
buf ( n31181 , RI15b4ed80_555);
and ( n31182 , n31181 , n31103 );
buf ( n31183 , RI15b4e9c0_547);
and ( n31184 , n31183 , n31106 );
buf ( n31185 , RI15b4e600_539);
and ( n31186 , n31185 , n31109 );
buf ( n31187 , RI15b4e240_531);
and ( n31188 , n31187 , n31112 );
buf ( n31189 , RI15b4de80_523);
and ( n31190 , n31189 , n31115 );
buf ( n31191 , RI15b4dac0_515);
and ( n31192 , n31191 , n31118 );
buf ( n31193 , RI15b4d700_507);
and ( n31194 , n31193 , n31121 );
buf ( n31195 , RI15b4d340_499);
and ( n31196 , n31195 , n31124 );
buf ( n31197 , RI15b4cf80_491);
and ( n31198 , n31197 , n31127 );
buf ( n31199 , RI15b4cbc0_483);
and ( n31200 , n31199 , n31130 );
buf ( n31201 , RI15b4c800_475);
and ( n31202 , n31201 , n31133 );
buf ( n31203 , RI15b4c440_467);
and ( n31204 , n31203 , n31136 );
or ( n31205 , n31174 , n31176 , n31178 , n31180 , n31182 , n31184 , n31186 , n31188 , n31190 , n31192 , n31194 , n31196 , n31198 , n31200 , n31202 , n31204 );
buf ( n31206 , RI15b4fcf8_588);
and ( n31207 , n31206 , n31088 );
buf ( n31208 , RI15b4f938_580);
and ( n31209 , n31208 , n31092 );
buf ( n31210 , RI15b4f578_572);
and ( n31211 , n31210 , n31096 );
buf ( n31212 , RI15b4f1b8_564);
and ( n31213 , n31212 , n31099 );
buf ( n31214 , RI15b4edf8_556);
and ( n31215 , n31214 , n31103 );
buf ( n31216 , RI15b4ea38_548);
and ( n31217 , n31216 , n31106 );
buf ( n31218 , RI15b4e678_540);
and ( n31219 , n31218 , n31109 );
buf ( n31220 , RI15b4e2b8_532);
and ( n31221 , n31220 , n31112 );
buf ( n31222 , RI15b4def8_524);
and ( n31223 , n31222 , n31115 );
buf ( n31224 , RI15b4db38_516);
and ( n31225 , n31224 , n31118 );
buf ( n31226 , RI15b4d778_508);
and ( n31227 , n31226 , n31121 );
buf ( n31228 , RI15b4d3b8_500);
and ( n31229 , n31228 , n31124 );
buf ( n31230 , RI15b4cff8_492);
and ( n31231 , n31230 , n31127 );
buf ( n31232 , RI15b4cc38_484);
and ( n31233 , n31232 , n31130 );
buf ( n31234 , RI15b4c878_476);
and ( n31235 , n31234 , n31133 );
buf ( n31236 , RI15b4c4b8_468);
and ( n31237 , n31236 , n31136 );
or ( n31238 , n31207 , n31209 , n31211 , n31213 , n31215 , n31217 , n31219 , n31221 , n31223 , n31225 , n31227 , n31229 , n31231 , n31233 , n31235 , n31237 );
not ( n31239 , n31238 );
buf ( n31240 , RI15b4fd70_589);
and ( n31241 , n31240 , n31088 );
buf ( n31242 , RI15b4f9b0_581);
and ( n31243 , n31242 , n31092 );
buf ( n31244 , RI15b4f5f0_573);
and ( n31245 , n31244 , n31096 );
buf ( n31246 , RI15b4f230_565);
and ( n31247 , n31246 , n31099 );
buf ( n31248 , RI15b4ee70_557);
and ( n31249 , n31248 , n31103 );
buf ( n31250 , RI15b4eab0_549);
and ( n31251 , n31250 , n31106 );
buf ( n31252 , RI15b4e6f0_541);
and ( n31253 , n31252 , n31109 );
buf ( n31254 , RI15b4e330_533);
and ( n31255 , n31254 , n31112 );
buf ( n31256 , RI15b4df70_525);
and ( n31257 , n31256 , n31115 );
buf ( n31258 , RI15b4dbb0_517);
and ( n31259 , n31258 , n31118 );
buf ( n31260 , RI15b4d7f0_509);
and ( n31261 , n31260 , n31121 );
buf ( n31262 , RI15b4d430_501);
and ( n31263 , n31262 , n31124 );
buf ( n31264 , RI15b4d070_493);
and ( n31265 , n31264 , n31127 );
buf ( n31266 , RI15b4ccb0_485);
and ( n31267 , n31266 , n31130 );
buf ( n31268 , RI15b4c8f0_477);
and ( n31269 , n31268 , n31133 );
buf ( n31270 , RI15b4c530_469);
and ( n31271 , n31270 , n31136 );
or ( n31272 , n31241 , n31243 , n31245 , n31247 , n31249 , n31251 , n31253 , n31255 , n31257 , n31259 , n31261 , n31263 , n31265 , n31267 , n31269 , n31271 );
not ( n31273 , n31272 );
buf ( n31274 , RI15b4fde8_590);
and ( n31275 , n31274 , n31088 );
buf ( n31276 , RI15b4fa28_582);
and ( n31277 , n31276 , n31092 );
buf ( n31278 , RI15b4f668_574);
and ( n31279 , n31278 , n31096 );
buf ( n31280 , RI15b4f2a8_566);
and ( n31281 , n31280 , n31099 );
buf ( n31282 , RI15b4eee8_558);
and ( n31283 , n31282 , n31103 );
buf ( n31284 , RI15b4eb28_550);
and ( n31285 , n31284 , n31106 );
buf ( n31286 , RI15b4e768_542);
and ( n31287 , n31286 , n31109 );
buf ( n31288 , RI15b4e3a8_534);
and ( n31289 , n31288 , n31112 );
buf ( n31290 , RI15b4dfe8_526);
and ( n31291 , n31290 , n31115 );
buf ( n31292 , RI15b4dc28_518);
and ( n31293 , n31292 , n31118 );
buf ( n31294 , RI15b4d868_510);
and ( n31295 , n31294 , n31121 );
buf ( n31296 , RI15b4d4a8_502);
and ( n31297 , n31296 , n31124 );
buf ( n31298 , RI15b4d0e8_494);
and ( n31299 , n31298 , n31127 );
buf ( n31300 , RI15b4cd28_486);
and ( n31301 , n31300 , n31130 );
buf ( n31302 , RI15b4c968_478);
and ( n31303 , n31302 , n31133 );
buf ( n31304 , RI15b4c5a8_470);
and ( n31305 , n31304 , n31136 );
or ( n31306 , n31275 , n31277 , n31279 , n31281 , n31283 , n31285 , n31287 , n31289 , n31291 , n31293 , n31295 , n31297 , n31299 , n31301 , n31303 , n31305 );
buf ( n31307 , RI15b4fe60_591);
and ( n31308 , n31307 , n31088 );
buf ( n31309 , RI15b4faa0_583);
and ( n31310 , n31309 , n31092 );
buf ( n31311 , RI15b4f6e0_575);
and ( n31312 , n31311 , n31096 );
buf ( n31313 , RI15b4f320_567);
and ( n31314 , n31313 , n31099 );
buf ( n31315 , RI15b4ef60_559);
and ( n31316 , n31315 , n31103 );
buf ( n31317 , RI15b4eba0_551);
and ( n31318 , n31317 , n31106 );
buf ( n31319 , RI15b4e7e0_543);
and ( n31320 , n31319 , n31109 );
buf ( n31321 , RI15b4e420_535);
and ( n31322 , n31321 , n31112 );
buf ( n31323 , RI15b4e060_527);
and ( n31324 , n31323 , n31115 );
buf ( n31325 , RI15b4dca0_519);
and ( n31326 , n31325 , n31118 );
buf ( n31327 , RI15b4d8e0_511);
and ( n31328 , n31327 , n31121 );
buf ( n31329 , RI15b4d520_503);
and ( n31330 , n31329 , n31124 );
buf ( n31331 , RI15b4d160_495);
and ( n31332 , n31331 , n31127 );
buf ( n31333 , RI15b4cda0_487);
and ( n31334 , n31333 , n31130 );
buf ( n31335 , RI15b4c9e0_479);
and ( n31336 , n31335 , n31133 );
buf ( n31337 , RI15b4c620_471);
and ( n31338 , n31337 , n31136 );
or ( n31339 , n31308 , n31310 , n31312 , n31314 , n31316 , n31318 , n31320 , n31322 , n31324 , n31326 , n31328 , n31330 , n31332 , n31334 , n31336 , n31338 );
buf ( n31340 , RI15b4fed8_592);
and ( n31341 , n31340 , n31088 );
buf ( n31342 , RI15b4fb18_584);
and ( n31343 , n31342 , n31092 );
buf ( n31344 , RI15b4f758_576);
and ( n31345 , n31344 , n31096 );
buf ( n31346 , RI15b4f398_568);
and ( n31347 , n31346 , n31099 );
buf ( n31348 , RI15b4efd8_560);
and ( n31349 , n31348 , n31103 );
buf ( n31350 , RI15b4ec18_552);
and ( n31351 , n31350 , n31106 );
buf ( n31352 , RI15b4e858_544);
and ( n31353 , n31352 , n31109 );
buf ( n31354 , RI15b4e498_536);
and ( n31355 , n31354 , n31112 );
buf ( n31356 , RI15b4e0d8_528);
and ( n31357 , n31356 , n31115 );
buf ( n31358 , RI15b4dd18_520);
and ( n31359 , n31358 , n31118 );
buf ( n31360 , RI15b4d958_512);
and ( n31361 , n31360 , n31121 );
buf ( n31362 , RI15b4d598_504);
and ( n31363 , n31362 , n31124 );
buf ( n31364 , RI15b4d1d8_496);
and ( n31365 , n31364 , n31127 );
buf ( n31366 , RI15b4ce18_488);
and ( n31367 , n31366 , n31130 );
buf ( n31368 , RI15b4ca58_480);
and ( n31369 , n31368 , n31133 );
buf ( n31370 , RI15b4c698_472);
and ( n31371 , n31370 , n31136 );
or ( n31372 , n31341 , n31343 , n31345 , n31347 , n31349 , n31351 , n31353 , n31355 , n31357 , n31359 , n31361 , n31363 , n31365 , n31367 , n31369 , n31371 );
and ( n31373 , n31139 , n31172 , n31205 , n31239 , n31273 , n31306 , n31339 , n31372 );
and ( n31374 , n31085 , n31373 );
not ( n31375 , n31041 );
buf ( n31376 , n31041 );
buf ( n31377 , n31041 );
buf ( n31378 , n31041 );
buf ( n31379 , n31041 );
buf ( n31380 , n31041 );
buf ( n31381 , n31041 );
buf ( n31382 , n31041 );
buf ( n31383 , n31041 );
buf ( n31384 , n31041 );
buf ( n31385 , n31041 );
buf ( n31386 , n31041 );
buf ( n31387 , n31041 );
buf ( n31388 , n31041 );
buf ( n31389 , n31041 );
buf ( n31390 , n31041 );
buf ( n31391 , n31041 );
buf ( n31392 , n31041 );
buf ( n31393 , n31041 );
buf ( n31394 , n31041 );
buf ( n31395 , n31041 );
buf ( n31396 , n31041 );
buf ( n31397 , n31041 );
buf ( n31398 , n31041 );
buf ( n31399 , n31041 );
buf ( n31400 , n31041 );
or ( n31401 , n31044 , n31046 , n31048 , n31041 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31075 );
and ( n31402 , n31375 , n31401 );
not ( n31403 , n31402 );
and ( n31404 , n31403 , n31079 );
and ( n31405 , n31083 , n31402 );
or ( n31406 , n31404 , n31405 );
not ( n31407 , n31172 );
and ( n31408 , n31139 , n31407 , n31205 , n31239 , n31273 , n31306 , n31339 , n31372 );
and ( n31409 , n31406 , n31408 );
not ( n31410 , n31041 );
buf ( n31411 , n31041 );
buf ( n31412 , n31041 );
buf ( n31413 , n31041 );
buf ( n31414 , n31041 );
buf ( n31415 , n31041 );
buf ( n31416 , n31041 );
buf ( n31417 , n31041 );
buf ( n31418 , n31041 );
buf ( n31419 , n31041 );
buf ( n31420 , n31041 );
buf ( n31421 , n31041 );
buf ( n31422 , n31041 );
buf ( n31423 , n31041 );
buf ( n31424 , n31041 );
buf ( n31425 , n31041 );
buf ( n31426 , n31041 );
buf ( n31427 , n31041 );
buf ( n31428 , n31041 );
buf ( n31429 , n31041 );
buf ( n31430 , n31041 );
buf ( n31431 , n31041 );
buf ( n31432 , n31041 );
buf ( n31433 , n31041 );
buf ( n31434 , n31041 );
buf ( n31435 , n31041 );
or ( n31436 , n31044 , n31046 , n31048 , n31041 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31075 );
and ( n31437 , n31410 , n31436 );
not ( n31438 , n31437 );
and ( n31439 , n31438 , n31079 );
buf ( n31440 , RI15b54780_747);
buf ( n31441 , RI15b547f8_748);
not ( n31442 , n31441 );
buf ( n31443 , RI15b54870_749);
nor ( n31444 , n31440 , n31442 , n31443 );
not ( n31445 , n31440 );
and ( n31446 , n31445 , n31442 , n31443 );
or ( n31447 , n31444 , n31446 );
buf ( n31448 , RI15b667c8_1362);
buf ( n31449 , RI15b66840_1363);
and ( n31450 , n31448 , n31449 );
not ( n31451 , n31450 );
buf ( n31452 , RI15b54690_745);
not ( n31453 , n31452 );
and ( n31454 , n31451 , n31453 );
and ( n31455 , n31447 , n31454 );
not ( n31456 , n31455 );
buf ( n31457 , RI15b55950_785);
and ( n31458 , n31456 , n31457 );
buf ( n31459 , RI15b576d8_848);
buf ( n31460 , RI15b57660_847);
and ( n31461 , n31459 , n31460 );
xor ( n31462 , n31079 , n31461 );
and ( n31463 , n31462 , n31455 );
or ( n31464 , n31458 , n31463 );
and ( n31465 , n31464 , n31437 );
or ( n31466 , n31439 , n31465 );
not ( n31467 , n31372 );
nor ( n31468 , n31139 , n31172 , n31205 , n31239 , n31272 , n31306 , n31339 , n31467 );
and ( n31469 , n31466 , n31468 );
not ( n31470 , n31041 );
buf ( n31471 , n31041 );
buf ( n31472 , n31041 );
buf ( n31473 , n31041 );
buf ( n31474 , n31041 );
buf ( n31475 , n31041 );
buf ( n31476 , n31041 );
buf ( n31477 , n31041 );
buf ( n31478 , n31041 );
buf ( n31479 , n31041 );
buf ( n31480 , n31041 );
buf ( n31481 , n31041 );
buf ( n31482 , n31041 );
buf ( n31483 , n31041 );
buf ( n31484 , n31041 );
buf ( n31485 , n31041 );
buf ( n31486 , n31041 );
buf ( n31487 , n31041 );
buf ( n31488 , n31041 );
buf ( n31489 , n31041 );
buf ( n31490 , n31041 );
buf ( n31491 , n31041 );
buf ( n31492 , n31041 );
buf ( n31493 , n31041 );
buf ( n31494 , n31041 );
buf ( n31495 , n31041 );
or ( n31496 , n31044 , n31046 , n31048 , n31041 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31075 );
and ( n31497 , n31470 , n31496 );
not ( n31498 , n31497 );
and ( n31499 , n31498 , n31079 );
not ( n31500 , n31454 );
buf ( n31501 , RI15b56670_813);
not ( n31502 , n31501 );
and ( n31503 , n31502 , n31457 );
not ( n31504 , n31457 );
buf ( n31505 , RI15b558d8_784);
not ( n31506 , n31505 );
buf ( n31507 , RI15b55860_783);
not ( n31508 , n31507 );
buf ( n31509 , RI15b557e8_782);
not ( n31510 , n31509 );
and ( n31511 , n31508 , n31510 );
and ( n31512 , n31506 , n31511 );
xor ( n31513 , n31504 , n31512 );
and ( n31514 , n31513 , n31501 );
or ( n31515 , n31503 , n31514 );
and ( n31516 , n31500 , n31515 );
and ( n31517 , n31462 , n31454 );
or ( n31518 , n31516 , n31517 );
and ( n31519 , n31518 , n31497 );
or ( n31520 , n31499 , n31519 );
nor ( n31521 , n31139 , n31407 , n31205 , n31239 , n31272 , n31306 , n31339 , n31467 );
and ( n31522 , n31520 , n31521 );
and ( n31523 , n31139 , n31172 , n31205 , n31239 , n31273 , n31306 , n31339 , n31467 );
nor ( n31524 , n31138 , n31172 , n31205 , n31238 , n31273 , n31306 , n31339 , n31467 );
or ( n31525 , n31523 , n31524 );
not ( n31526 , n31205 );
and ( n31527 , n31138 , n31172 , n31526 , n31238 , n31273 , n31306 , n31339 , n31372 );
or ( n31528 , n31525 , n31527 );
and ( n31529 , n31138 , n31407 , n31526 , n31238 , n31273 , n31306 , n31339 , n31372 );
or ( n31530 , n31528 , n31529 );
and ( n31531 , n31139 , n31172 , n31526 , n31238 , n31273 , n31306 , n31339 , n31372 );
or ( n31532 , n31530 , n31531 );
not ( n31533 , n31339 );
and ( n31534 , n31139 , n31407 , n31526 , n31239 , n31272 , n31306 , n31533 , n31372 );
or ( n31535 , n31532 , n31534 );
and ( n31536 , n31139 , n31407 , n31526 , n31238 , n31272 , n31306 , n31533 , n31372 );
or ( n31537 , n31535 , n31536 );
and ( n31538 , n31138 , n31172 , n31526 , n31238 , n31272 , n31306 , n31533 , n31372 );
or ( n31539 , n31537 , n31538 );
nor ( n31540 , n31138 , n31172 , n31526 , n31238 , n31272 , n31306 , n31339 , n31372 );
or ( n31541 , n31539 , n31540 );
nor ( n31542 , n31139 , n31172 , n31526 , n31238 , n31272 , n31306 , n31339 , n31372 );
or ( n31543 , n31541 , n31542 );
nor ( n31544 , n31138 , n31172 , n31205 , n31238 , n31273 , n31306 , n31533 , n31467 );
or ( n31545 , n31543 , n31544 );
nor ( n31546 , n31138 , n31172 , n31205 , n31238 , n31272 , n31306 , n31533 , n31467 );
or ( n31547 , n31545 , n31546 );
nor ( n31548 , n31138 , n31172 , n31205 , n31238 , n31272 , n31306 , n31533 , n31372 );
or ( n31549 , n31547 , n31548 );
nor ( n31550 , n31139 , n31407 , n31205 , n31238 , n31272 , n31306 , n31533 , n31372 );
or ( n31551 , n31549 , n31550 );
nor ( n31552 , n31524 , n31523 , n31527 , n31529 , n31531 , n31534 , n31536 , n31538 , n31521 , n31468 , n31408 , n31373 , n31540 , n31542 , n31544 , n31546 , n31548 , n31550 );
or ( n31553 , n31551 , n31552 );
and ( n31554 , n31079 , n31553 );
or ( n31555 , n31374 , n31409 , n31469 , n31522 , n31554 );
not ( n31556 , n30999 );
and ( n31557 , n30990 , n31556 , n31002 , n31006 );
and ( n31558 , n31555 , n31557 );
not ( n31559 , n31452 );
buf ( n31560 , RI15b57570_845);
buf ( n31561 , RI15b574f8_844);
buf ( n31562 , RI15b57480_843);
buf ( n31563 , RI15b57408_842);
buf ( n31564 , RI15b57390_841);
buf ( n31565 , RI15b57318_840);
buf ( n31566 , RI15b572a0_839);
buf ( n31567 , RI15b57228_838);
buf ( n31568 , RI15b571b0_837);
buf ( n31569 , RI15b57138_836);
buf ( n31570 , RI15b570c0_835);
buf ( n31571 , RI15b57048_834);
buf ( n31572 , RI15b56fd0_833);
buf ( n31573 , RI15b56f58_832);
buf ( n31574 , RI15b56ee0_831);
buf ( n31575 , RI15b56e68_830);
buf ( n31576 , RI15b56df0_829);
buf ( n31577 , RI15b56d78_828);
buf ( n31578 , RI15b56d00_827);
buf ( n31579 , RI15b56c88_826);
buf ( n31580 , RI15b56c10_825);
buf ( n31581 , RI15b56b98_824);
buf ( n31582 , RI15b56b20_823);
buf ( n31583 , RI15b56aa8_822);
buf ( n31584 , RI15b56a30_821);
buf ( n31585 , RI15b569b8_820);
buf ( n31586 , RI15b56940_819);
buf ( n31587 , RI15b568c8_818);
buf ( n31588 , RI15b567d8_816);
buf ( n31589 , RI15b56760_815);
and ( n31590 , n31588 , n31589 );
and ( n31591 , n30989 , n31590 );
and ( n31592 , n31587 , n31591 );
and ( n31593 , n31586 , n31592 );
and ( n31594 , n31585 , n31593 );
and ( n31595 , n31584 , n31594 );
and ( n31596 , n31583 , n31595 );
and ( n31597 , n31582 , n31596 );
and ( n31598 , n31581 , n31597 );
and ( n31599 , n31580 , n31598 );
and ( n31600 , n31579 , n31599 );
and ( n31601 , n31578 , n31600 );
and ( n31602 , n31577 , n31601 );
and ( n31603 , n31576 , n31602 );
and ( n31604 , n31575 , n31603 );
and ( n31605 , n31574 , n31604 );
and ( n31606 , n31573 , n31605 );
and ( n31607 , n31572 , n31606 );
and ( n31608 , n31571 , n31607 );
and ( n31609 , n31570 , n31608 );
and ( n31610 , n31569 , n31609 );
and ( n31611 , n31568 , n31610 );
and ( n31612 , n31567 , n31611 );
and ( n31613 , n31566 , n31612 );
and ( n31614 , n31565 , n31613 );
and ( n31615 , n31564 , n31614 );
and ( n31616 , n31563 , n31615 );
and ( n31617 , n31562 , n31616 );
and ( n31618 , n31561 , n31617 );
xor ( n31619 , n31560 , n31618 );
not ( n31620 , n31619 );
xor ( n31621 , n30989 , n31590 );
and ( n31622 , n31620 , n31621 );
not ( n31623 , n31621 );
xor ( n31624 , n31588 , n31589 );
not ( n31625 , n31624 );
not ( n31626 , n31589 );
not ( n31627 , n31626 );
buf ( n31628 , RI15b566e8_814);
not ( n31629 , n31628 );
and ( n31630 , n31627 , n31629 );
and ( n31631 , n31625 , n31630 );
xor ( n31632 , n31623 , n31631 );
and ( n31633 , n31632 , n31619 );
or ( n31634 , n31622 , n31633 );
and ( n31635 , n31559 , n31634 );
and ( n31636 , n31079 , n31452 );
or ( n31637 , n31635 , n31636 );
nor ( n31638 , n30990 , n31556 , n31002 , n31005 );
and ( n31639 , n31637 , n31638 );
nor ( n31640 , n30991 , n30999 , n31002 , n31005 );
nor ( n31641 , n30991 , n31556 , n31002 , n31005 );
or ( n31642 , n31640 , n31641 );
and ( n31643 , n30991 , n31556 , n31002 , n31006 );
or ( n31644 , n31642 , n31643 );
and ( n31645 , n30991 , n30999 , n31002 , n31006 );
or ( n31646 , n31644 , n31645 );
and ( n31647 , n30990 , n30999 , n31002 , n31006 );
or ( n31648 , n31646 , n31647 );
nor ( n31649 , n30990 , n30999 , n31002 , n31006 );
or ( n31650 , n31648 , n31649 );
and ( n31651 , n31079 , n31650 );
or ( n31652 , C0 , n31008 , n31558 , n31639 , C0 , n31651 );
buf ( n31653 , n31652 );
buf ( n31654 , n31653 );
buf ( n31655 , RI15b3ea48_2);
buf ( n31656 , n31655 );
buf ( n31657 , RI15b58740_883);
buf ( n31658 , RI15b5d498_1048);
not ( n31659 , n31658 );
and ( n31660 , n31657 , n31659 );
buf ( n31661 , RI15b586c8_882);
buf ( n31662 , RI15b5d420_1047);
not ( n31663 , n31662 );
and ( n31664 , n31661 , n31663 );
buf ( n31665 , RI15b58650_881);
buf ( n31666 , RI15b5d3a8_1046);
not ( n31667 , n31666 );
and ( n31668 , n31665 , n31667 );
buf ( n31669 , RI15b585d8_880);
buf ( n31670 , RI15b5d330_1045);
not ( n31671 , n31670 );
and ( n31672 , n31669 , n31671 );
buf ( n31673 , RI15b58560_879);
buf ( n31674 , RI15b5d2b8_1044);
not ( n31675 , n31674 );
or ( n31676 , n31673 , n31675 );
and ( n31677 , n31671 , n31676 );
and ( n31678 , n31669 , n31676 );
or ( n31679 , n31672 , n31677 , n31678 );
and ( n31680 , n31667 , n31679 );
and ( n31681 , n31665 , n31679 );
or ( n31682 , n31668 , n31680 , n31681 );
and ( n31683 , n31663 , n31682 );
and ( n31684 , n31661 , n31682 );
or ( n31685 , n31664 , n31683 , n31684 );
and ( n31686 , n31659 , n31685 );
and ( n31687 , n31657 , n31685 );
or ( n31688 , n31660 , n31686 , n31687 );
not ( n31689 , n31688 );
not ( n31690 , n31689 );
xor ( n31691 , n31661 , n31663 );
xor ( n31692 , n31691 , n31682 );
xor ( n31693 , n31657 , n31659 );
xor ( n31694 , n31693 , n31685 );
buf ( n31695 , n31689 );
buf ( n31696 , n31689 );
buf ( n31697 , n31689 );
buf ( n31698 , n31689 );
buf ( n31699 , n31689 );
buf ( n31700 , n31689 );
buf ( n31701 , n31689 );
buf ( n31702 , n31689 );
buf ( n31703 , n31689 );
buf ( n31704 , n31689 );
buf ( n31705 , n31689 );
buf ( n31706 , n31689 );
buf ( n31707 , n31689 );
buf ( n31708 , n31689 );
buf ( n31709 , n31689 );
buf ( n31710 , n31689 );
buf ( n31711 , n31689 );
buf ( n31712 , n31689 );
buf ( n31713 , n31689 );
buf ( n31714 , n31689 );
buf ( n31715 , n31689 );
buf ( n31716 , n31689 );
buf ( n31717 , n31689 );
buf ( n31718 , n31689 );
buf ( n31719 , n31689 );
xor ( n31720 , n31665 , n31667 );
xor ( n31721 , n31720 , n31679 );
xor ( n31722 , n31669 , n31671 );
xor ( n31723 , n31722 , n31676 );
xor ( n31724 , n31673 , n31674 );
or ( n31725 , n31723 , n31724 );
and ( n31726 , n31721 , n31725 );
or ( n31727 , n31692 , n31694 , n31689 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31726 );
and ( n31728 , n31690 , n31727 );
not ( n31729 , n31728 );
buf ( n31730 , RI15b62f10_1241);
and ( n31731 , n31729 , n31730 );
buf ( n31732 , RI15b5c778_1020);
buf ( n31733 , RI15b5c700_1019);
buf ( n31734 , RI15b5c688_1018);
buf ( n31735 , RI15b5c610_1017);
buf ( n31736 , RI15b5c598_1016);
buf ( n31737 , RI15b5c520_1015);
buf ( n31738 , RI15b5c4a8_1014);
buf ( n31739 , RI15b5c430_1013);
buf ( n31740 , RI15b5c3b8_1012);
and ( n31741 , n31739 , n31740 );
or ( n31742 , n31738 , n31741 );
and ( n31743 , n31737 , n31742 );
and ( n31744 , n31736 , n31743 );
and ( n31745 , n31735 , n31744 );
and ( n31746 , n31734 , n31745 );
and ( n31747 , n31733 , n31746 );
xor ( n31748 , n31732 , n31747 );
xor ( n31749 , n31733 , n31746 );
buf ( n31750 , RI15b5c340_1011);
not ( n31751 , n31674 );
not ( n31752 , n31751 );
buf ( n31753 , n31752 );
not ( n31754 , n31753 );
not ( n31755 , n31754 );
xor ( n31756 , n31670 , n31674 );
not ( n31757 , n31756 );
buf ( n31758 , n31757 );
buf ( n31759 , n31758 );
not ( n31760 , n31759 );
not ( n31761 , n31760 );
and ( n31762 , n31670 , n31674 );
xor ( n31763 , n31666 , n31762 );
not ( n31764 , n31763 );
buf ( n31765 , n31764 );
buf ( n31766 , n31765 );
not ( n31767 , n31766 );
not ( n31768 , n31767 );
and ( n31769 , n31666 , n31762 );
xor ( n31770 , n31662 , n31769 );
not ( n31771 , n31770 );
buf ( n31772 , n31771 );
buf ( n31773 , n31772 );
not ( n31774 , n31773 );
not ( n31775 , n31774 );
nor ( n31776 , n31755 , n31761 , n31768 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31777 , n31750 , n31776 );
buf ( n31778 , RI15b5bf80_1003);
nor ( n31779 , n31754 , n31761 , n31768 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31780 , n31778 , n31779 );
buf ( n31781 , RI15b5bbc0_995);
nor ( n31782 , n31755 , n31760 , n31768 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31783 , n31781 , n31782 );
buf ( n31784 , RI15b5b800_987);
nor ( n31785 , n31754 , n31760 , n31768 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31786 , n31784 , n31785 );
buf ( n31787 , RI15b5b440_979);
nor ( n31788 , n31755 , n31761 , n31767 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31789 , n31787 , n31788 );
buf ( n31790 , RI15b5b080_971);
nor ( n31791 , n31754 , n31761 , n31767 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31792 , n31790 , n31791 );
buf ( n31793 , RI15b5acc0_963);
nor ( n31794 , n31755 , n31760 , n31767 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31795 , n31793 , n31794 );
buf ( n31796 , RI15b5a900_955);
nor ( n31797 , n31754 , n31760 , n31767 , n31775 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31798 , n31796 , n31797 );
buf ( n31799 , RI15b5a540_947);
nor ( n31800 , n31755 , n31761 , n31768 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31801 , n31799 , n31800 );
buf ( n31802 , RI15b5a180_939);
nor ( n31803 , n31754 , n31761 , n31768 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31804 , n31802 , n31803 );
buf ( n31805 , RI15b59dc0_931);
nor ( n31806 , n31755 , n31760 , n31768 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31807 , n31805 , n31806 );
buf ( n31808 , RI15b59a00_923);
nor ( n31809 , n31754 , n31760 , n31768 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31810 , n31808 , n31809 );
buf ( n31811 , RI15b59640_915);
nor ( n31812 , n31755 , n31761 , n31767 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31813 , n31811 , n31812 );
buf ( n31814 , RI15b59280_907);
nor ( n31815 , n31754 , n31761 , n31767 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31816 , n31814 , n31815 );
buf ( n31817 , RI15b58ec0_899);
nor ( n31818 , n31755 , n31760 , n31767 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31819 , n31817 , n31818 );
buf ( n31820 , RI15b58b00_891);
nor ( n31821 , n31754 , n31760 , n31767 , n31774 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n31822 , n31820 , n31821 );
or ( n31823 , n31777 , n31780 , n31783 , n31786 , n31789 , n31792 , n31795 , n31798 , n31801 , n31804 , n31807 , n31810 , n31813 , n31816 , n31819 , n31822 );
and ( n31824 , n31749 , n31823 );
xor ( n31825 , n31734 , n31745 );
buf ( n31826 , RI15b5c2c8_1010);
and ( n31827 , n31826 , n31776 );
buf ( n31828 , RI15b5bf08_1002);
and ( n31829 , n31828 , n31779 );
buf ( n31830 , RI15b5bb48_994);
and ( n31831 , n31830 , n31782 );
buf ( n31832 , RI15b5b788_986);
and ( n31833 , n31832 , n31785 );
buf ( n31834 , RI15b5b3c8_978);
and ( n31835 , n31834 , n31788 );
buf ( n31836 , RI15b5b008_970);
and ( n31837 , n31836 , n31791 );
buf ( n31838 , RI15b5ac48_962);
and ( n31839 , n31838 , n31794 );
buf ( n31840 , RI15b5a888_954);
and ( n31841 , n31840 , n31797 );
buf ( n31842 , RI15b5a4c8_946);
and ( n31843 , n31842 , n31800 );
buf ( n31844 , RI15b5a108_938);
and ( n31845 , n31844 , n31803 );
buf ( n31846 , RI15b59d48_930);
and ( n31847 , n31846 , n31806 );
buf ( n31848 , RI15b59988_922);
and ( n31849 , n31848 , n31809 );
buf ( n31850 , RI15b595c8_914);
and ( n31851 , n31850 , n31812 );
buf ( n31852 , RI15b59208_906);
and ( n31853 , n31852 , n31815 );
buf ( n31854 , RI15b58e48_898);
and ( n31855 , n31854 , n31818 );
buf ( n31856 , RI15b58a88_890);
and ( n31857 , n31856 , n31821 );
or ( n31858 , n31827 , n31829 , n31831 , n31833 , n31835 , n31837 , n31839 , n31841 , n31843 , n31845 , n31847 , n31849 , n31851 , n31853 , n31855 , n31857 );
and ( n31859 , n31825 , n31858 );
xor ( n31860 , n31735 , n31744 );
buf ( n31861 , RI15b5c250_1009);
and ( n31862 , n31861 , n31776 );
buf ( n31863 , RI15b5be90_1001);
and ( n31864 , n31863 , n31779 );
buf ( n31865 , RI15b5bad0_993);
and ( n31866 , n31865 , n31782 );
buf ( n31867 , RI15b5b710_985);
and ( n31868 , n31867 , n31785 );
buf ( n31869 , RI15b5b350_977);
and ( n31870 , n31869 , n31788 );
buf ( n31871 , RI15b5af90_969);
and ( n31872 , n31871 , n31791 );
buf ( n31873 , RI15b5abd0_961);
and ( n31874 , n31873 , n31794 );
buf ( n31875 , RI15b5a810_953);
and ( n31876 , n31875 , n31797 );
buf ( n31877 , RI15b5a450_945);
and ( n31878 , n31877 , n31800 );
buf ( n31879 , RI15b5a090_937);
and ( n31880 , n31879 , n31803 );
buf ( n31881 , RI15b59cd0_929);
and ( n31882 , n31881 , n31806 );
buf ( n31883 , RI15b59910_921);
and ( n31884 , n31883 , n31809 );
buf ( n31885 , RI15b59550_913);
and ( n31886 , n31885 , n31812 );
buf ( n31887 , RI15b59190_905);
and ( n31888 , n31887 , n31815 );
buf ( n31889 , RI15b58dd0_897);
and ( n31890 , n31889 , n31818 );
buf ( n31891 , RI15b58a10_889);
and ( n31892 , n31891 , n31821 );
or ( n31893 , n31862 , n31864 , n31866 , n31868 , n31870 , n31872 , n31874 , n31876 , n31878 , n31880 , n31882 , n31884 , n31886 , n31888 , n31890 , n31892 );
and ( n31894 , n31860 , n31893 );
xor ( n31895 , n31736 , n31743 );
buf ( n31896 , RI15b5c1d8_1008);
and ( n31897 , n31896 , n31776 );
buf ( n31898 , RI15b5be18_1000);
and ( n31899 , n31898 , n31779 );
buf ( n31900 , RI15b5ba58_992);
and ( n31901 , n31900 , n31782 );
buf ( n31902 , RI15b5b698_984);
and ( n31903 , n31902 , n31785 );
buf ( n31904 , RI15b5b2d8_976);
and ( n31905 , n31904 , n31788 );
buf ( n31906 , RI15b5af18_968);
and ( n31907 , n31906 , n31791 );
buf ( n31908 , RI15b5ab58_960);
and ( n31909 , n31908 , n31794 );
buf ( n31910 , RI15b5a798_952);
and ( n31911 , n31910 , n31797 );
buf ( n31912 , RI15b5a3d8_944);
and ( n31913 , n31912 , n31800 );
buf ( n31914 , RI15b5a018_936);
and ( n31915 , n31914 , n31803 );
buf ( n31916 , RI15b59c58_928);
and ( n31917 , n31916 , n31806 );
buf ( n31918 , RI15b59898_920);
and ( n31919 , n31918 , n31809 );
buf ( n31920 , RI15b594d8_912);
and ( n31921 , n31920 , n31812 );
buf ( n31922 , RI15b59118_904);
and ( n31923 , n31922 , n31815 );
buf ( n31924 , RI15b58d58_896);
and ( n31925 , n31924 , n31818 );
buf ( n31926 , RI15b58998_888);
and ( n31927 , n31926 , n31821 );
or ( n31928 , n31897 , n31899 , n31901 , n31903 , n31905 , n31907 , n31909 , n31911 , n31913 , n31915 , n31917 , n31919 , n31921 , n31923 , n31925 , n31927 );
and ( n31929 , n31895 , n31928 );
xor ( n31930 , n31737 , n31742 );
buf ( n31931 , RI15b5c160_1007);
and ( n31932 , n31931 , n31776 );
buf ( n31933 , RI15b5bda0_999);
and ( n31934 , n31933 , n31779 );
buf ( n31935 , RI15b5b9e0_991);
and ( n31936 , n31935 , n31782 );
buf ( n31937 , RI15b5b620_983);
and ( n31938 , n31937 , n31785 );
buf ( n31939 , RI15b5b260_975);
and ( n31940 , n31939 , n31788 );
buf ( n31941 , RI15b5aea0_967);
and ( n31942 , n31941 , n31791 );
buf ( n31943 , RI15b5aae0_959);
and ( n31944 , n31943 , n31794 );
buf ( n31945 , RI15b5a720_951);
and ( n31946 , n31945 , n31797 );
buf ( n31947 , RI15b5a360_943);
and ( n31948 , n31947 , n31800 );
buf ( n31949 , RI15b59fa0_935);
and ( n31950 , n31949 , n31803 );
buf ( n31951 , RI15b59be0_927);
and ( n31952 , n31951 , n31806 );
buf ( n31953 , RI15b59820_919);
and ( n31954 , n31953 , n31809 );
buf ( n31955 , RI15b59460_911);
and ( n31956 , n31955 , n31812 );
buf ( n31957 , RI15b590a0_903);
and ( n31958 , n31957 , n31815 );
buf ( n31959 , RI15b58ce0_895);
and ( n31960 , n31959 , n31818 );
buf ( n31961 , RI15b58920_887);
and ( n31962 , n31961 , n31821 );
or ( n31963 , n31932 , n31934 , n31936 , n31938 , n31940 , n31942 , n31944 , n31946 , n31948 , n31950 , n31952 , n31954 , n31956 , n31958 , n31960 , n31962 );
and ( n31964 , n31930 , n31963 );
xnor ( n31965 , n31738 , n31741 );
buf ( n31966 , RI15b5c0e8_1006);
and ( n31967 , n31966 , n31776 );
buf ( n31968 , RI15b5bd28_998);
and ( n31969 , n31968 , n31779 );
buf ( n31970 , RI15b5b968_990);
and ( n31971 , n31970 , n31782 );
buf ( n31972 , RI15b5b5a8_982);
and ( n31973 , n31972 , n31785 );
buf ( n31974 , RI15b5b1e8_974);
and ( n31975 , n31974 , n31788 );
buf ( n31976 , RI15b5ae28_966);
and ( n31977 , n31976 , n31791 );
buf ( n31978 , RI15b5aa68_958);
and ( n31979 , n31978 , n31794 );
buf ( n31980 , RI15b5a6a8_950);
and ( n31981 , n31980 , n31797 );
buf ( n31982 , RI15b5a2e8_942);
and ( n31983 , n31982 , n31800 );
buf ( n31984 , RI15b59f28_934);
and ( n31985 , n31984 , n31803 );
buf ( n31986 , RI15b59b68_926);
and ( n31987 , n31986 , n31806 );
buf ( n31988 , RI15b597a8_918);
and ( n31989 , n31988 , n31809 );
buf ( n31990 , RI15b593e8_910);
and ( n31991 , n31990 , n31812 );
buf ( n31992 , RI15b59028_902);
and ( n31993 , n31992 , n31815 );
buf ( n31994 , RI15b58c68_894);
and ( n31995 , n31994 , n31818 );
buf ( n31996 , RI15b588a8_886);
and ( n31997 , n31996 , n31821 );
or ( n31998 , n31967 , n31969 , n31971 , n31973 , n31975 , n31977 , n31979 , n31981 , n31983 , n31985 , n31987 , n31989 , n31991 , n31993 , n31995 , n31997 );
and ( n31999 , n31965 , n31998 );
xor ( n32000 , n31739 , n31740 );
buf ( n32001 , RI15b5c070_1005);
and ( n32002 , n32001 , n31776 );
buf ( n32003 , RI15b5bcb0_997);
and ( n32004 , n32003 , n31779 );
buf ( n32005 , RI15b5b8f0_989);
and ( n32006 , n32005 , n31782 );
buf ( n32007 , RI15b5b530_981);
and ( n32008 , n32007 , n31785 );
buf ( n32009 , RI15b5b170_973);
and ( n32010 , n32009 , n31788 );
buf ( n32011 , RI15b5adb0_965);
and ( n32012 , n32011 , n31791 );
buf ( n32013 , RI15b5a9f0_957);
and ( n32014 , n32013 , n31794 );
buf ( n32015 , RI15b5a630_949);
and ( n32016 , n32015 , n31797 );
buf ( n32017 , RI15b5a270_941);
and ( n32018 , n32017 , n31800 );
buf ( n32019 , RI15b59eb0_933);
and ( n32020 , n32019 , n31803 );
buf ( n32021 , RI15b59af0_925);
and ( n32022 , n32021 , n31806 );
buf ( n32023 , RI15b59730_917);
and ( n32024 , n32023 , n31809 );
buf ( n32025 , RI15b59370_909);
and ( n32026 , n32025 , n31812 );
buf ( n32027 , RI15b58fb0_901);
and ( n32028 , n32027 , n31815 );
buf ( n32029 , RI15b58bf0_893);
and ( n32030 , n32029 , n31818 );
buf ( n32031 , RI15b58830_885);
and ( n32032 , n32031 , n31821 );
or ( n32033 , n32002 , n32004 , n32006 , n32008 , n32010 , n32012 , n32014 , n32016 , n32018 , n32020 , n32022 , n32024 , n32026 , n32028 , n32030 , n32032 );
and ( n32034 , n32000 , n32033 );
not ( n32035 , n31740 );
buf ( n32036 , RI15b5bff8_1004);
and ( n32037 , n32036 , n31776 );
buf ( n32038 , RI15b5bc38_996);
and ( n32039 , n32038 , n31779 );
buf ( n32040 , RI15b5b878_988);
and ( n32041 , n32040 , n31782 );
buf ( n32042 , RI15b5b4b8_980);
and ( n32043 , n32042 , n31785 );
buf ( n32044 , RI15b5b0f8_972);
and ( n32045 , n32044 , n31788 );
buf ( n32046 , RI15b5ad38_964);
and ( n32047 , n32046 , n31791 );
buf ( n32048 , RI15b5a978_956);
and ( n32049 , n32048 , n31794 );
buf ( n32050 , RI15b5a5b8_948);
and ( n32051 , n32050 , n31797 );
buf ( n32052 , RI15b5a1f8_940);
and ( n32053 , n32052 , n31800 );
buf ( n32054 , RI15b59e38_932);
and ( n32055 , n32054 , n31803 );
buf ( n32056 , RI15b59a78_924);
and ( n32057 , n32056 , n31806 );
buf ( n32058 , RI15b596b8_916);
and ( n32059 , n32058 , n31809 );
buf ( n32060 , RI15b592f8_908);
and ( n32061 , n32060 , n31812 );
buf ( n32062 , RI15b58f38_900);
and ( n32063 , n32062 , n31815 );
buf ( n32064 , RI15b58b78_892);
and ( n32065 , n32064 , n31818 );
buf ( n32066 , RI15b587b8_884);
and ( n32067 , n32066 , n31821 );
or ( n32068 , n32037 , n32039 , n32041 , n32043 , n32045 , n32047 , n32049 , n32051 , n32053 , n32055 , n32057 , n32059 , n32061 , n32063 , n32065 , n32067 );
and ( n32069 , n32035 , n32068 );
and ( n32070 , n32033 , n32069 );
and ( n32071 , n32000 , n32069 );
or ( n32072 , n32034 , n32070 , n32071 );
and ( n32073 , n31998 , n32072 );
and ( n32074 , n31965 , n32072 );
or ( n32075 , n31999 , n32073 , n32074 );
and ( n32076 , n31963 , n32075 );
and ( n32077 , n31930 , n32075 );
or ( n32078 , n31964 , n32076 , n32077 );
and ( n32079 , n31928 , n32078 );
and ( n32080 , n31895 , n32078 );
or ( n32081 , n31929 , n32079 , n32080 );
and ( n32082 , n31893 , n32081 );
and ( n32083 , n31860 , n32081 );
or ( n32084 , n31894 , n32082 , n32083 );
and ( n32085 , n31858 , n32084 );
and ( n32086 , n31825 , n32084 );
or ( n32087 , n31859 , n32085 , n32086 );
and ( n32088 , n31823 , n32087 );
and ( n32089 , n31749 , n32087 );
or ( n32090 , n31824 , n32088 , n32089 );
xor ( n32091 , n31748 , n32090 );
and ( n32092 , n32091 , n31728 );
or ( n32093 , n31731 , n32092 );
not ( n32094 , n31658 );
and ( n32095 , n31674 , n31670 , n31666 , n31662 , n32094 );
and ( n32096 , n32036 , n32095 );
not ( n32097 , n31674 );
and ( n32098 , n32097 , n31670 , n31666 , n31662 , n32094 );
and ( n32099 , n32038 , n32098 );
not ( n32100 , n31670 );
and ( n32101 , n31674 , n32100 , n31666 , n31662 , n32094 );
and ( n32102 , n32040 , n32101 );
and ( n32103 , n32097 , n32100 , n31666 , n31662 , n32094 );
and ( n32104 , n32042 , n32103 );
not ( n32105 , n31666 );
and ( n32106 , n31674 , n31670 , n32105 , n31662 , n32094 );
and ( n32107 , n32044 , n32106 );
and ( n32108 , n32097 , n31670 , n32105 , n31662 , n32094 );
and ( n32109 , n32046 , n32108 );
and ( n32110 , n31674 , n32100 , n32105 , n31662 , n32094 );
and ( n32111 , n32048 , n32110 );
and ( n32112 , n32097 , n32100 , n32105 , n31662 , n32094 );
and ( n32113 , n32050 , n32112 );
nor ( n32114 , n32097 , n32100 , n32105 , n31662 , n31658 );
and ( n32115 , n32052 , n32114 );
nor ( n32116 , n31674 , n32100 , n32105 , n31662 , n31658 );
and ( n32117 , n32054 , n32116 );
nor ( n32118 , n32097 , n31670 , n32105 , n31662 , n31658 );
and ( n32119 , n32056 , n32118 );
nor ( n32120 , n31674 , n31670 , n32105 , n31662 , n31658 );
and ( n32121 , n32058 , n32120 );
nor ( n32122 , n32097 , n32100 , n31666 , n31662 , n31658 );
and ( n32123 , n32060 , n32122 );
nor ( n32124 , n31674 , n32100 , n31666 , n31662 , n31658 );
and ( n32125 , n32062 , n32124 );
nor ( n32126 , n32097 , n31670 , n31666 , n31662 , n31658 );
and ( n32127 , n32064 , n32126 );
nor ( n32128 , n31674 , n31670 , n31666 , n31662 , n31658 );
and ( n32129 , n32066 , n32128 );
or ( n32130 , n32096 , n32099 , n32102 , n32104 , n32107 , n32109 , n32111 , n32113 , n32115 , n32117 , n32119 , n32121 , n32123 , n32125 , n32127 , n32129 );
and ( n32131 , n32001 , n32095 );
and ( n32132 , n32003 , n32098 );
and ( n32133 , n32005 , n32101 );
and ( n32134 , n32007 , n32103 );
and ( n32135 , n32009 , n32106 );
and ( n32136 , n32011 , n32108 );
and ( n32137 , n32013 , n32110 );
and ( n32138 , n32015 , n32112 );
and ( n32139 , n32017 , n32114 );
and ( n32140 , n32019 , n32116 );
and ( n32141 , n32021 , n32118 );
and ( n32142 , n32023 , n32120 );
and ( n32143 , n32025 , n32122 );
and ( n32144 , n32027 , n32124 );
and ( n32145 , n32029 , n32126 );
and ( n32146 , n32031 , n32128 );
or ( n32147 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 );
not ( n32148 , n32147 );
and ( n32149 , n31966 , n32095 );
and ( n32150 , n31968 , n32098 );
and ( n32151 , n31970 , n32101 );
and ( n32152 , n31972 , n32103 );
and ( n32153 , n31974 , n32106 );
and ( n32154 , n31976 , n32108 );
and ( n32155 , n31978 , n32110 );
and ( n32156 , n31980 , n32112 );
and ( n32157 , n31982 , n32114 );
and ( n32158 , n31984 , n32116 );
and ( n32159 , n31986 , n32118 );
and ( n32160 , n31988 , n32120 );
and ( n32161 , n31990 , n32122 );
and ( n32162 , n31992 , n32124 );
and ( n32163 , n31994 , n32126 );
and ( n32164 , n31996 , n32128 );
or ( n32165 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 );
not ( n32166 , n32165 );
and ( n32167 , n31931 , n32095 );
and ( n32168 , n31933 , n32098 );
and ( n32169 , n31935 , n32101 );
and ( n32170 , n31937 , n32103 );
and ( n32171 , n31939 , n32106 );
and ( n32172 , n31941 , n32108 );
and ( n32173 , n31943 , n32110 );
and ( n32174 , n31945 , n32112 );
and ( n32175 , n31947 , n32114 );
and ( n32176 , n31949 , n32116 );
and ( n32177 , n31951 , n32118 );
and ( n32178 , n31953 , n32120 );
and ( n32179 , n31955 , n32122 );
and ( n32180 , n31957 , n32124 );
and ( n32181 , n31959 , n32126 );
and ( n32182 , n31961 , n32128 );
or ( n32183 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 );
and ( n32184 , n31896 , n32095 );
and ( n32185 , n31898 , n32098 );
and ( n32186 , n31900 , n32101 );
and ( n32187 , n31902 , n32103 );
and ( n32188 , n31904 , n32106 );
and ( n32189 , n31906 , n32108 );
and ( n32190 , n31908 , n32110 );
and ( n32191 , n31910 , n32112 );
and ( n32192 , n31912 , n32114 );
and ( n32193 , n31914 , n32116 );
and ( n32194 , n31916 , n32118 );
and ( n32195 , n31918 , n32120 );
and ( n32196 , n31920 , n32122 );
and ( n32197 , n31922 , n32124 );
and ( n32198 , n31924 , n32126 );
and ( n32199 , n31926 , n32128 );
or ( n32200 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 );
not ( n32201 , n32200 );
and ( n32202 , n31861 , n32095 );
and ( n32203 , n31863 , n32098 );
and ( n32204 , n31865 , n32101 );
and ( n32205 , n31867 , n32103 );
and ( n32206 , n31869 , n32106 );
and ( n32207 , n31871 , n32108 );
and ( n32208 , n31873 , n32110 );
and ( n32209 , n31875 , n32112 );
and ( n32210 , n31877 , n32114 );
and ( n32211 , n31879 , n32116 );
and ( n32212 , n31881 , n32118 );
and ( n32213 , n31883 , n32120 );
and ( n32214 , n31885 , n32122 );
and ( n32215 , n31887 , n32124 );
and ( n32216 , n31889 , n32126 );
and ( n32217 , n31891 , n32128 );
or ( n32218 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 );
and ( n32219 , n31826 , n32095 );
and ( n32220 , n31828 , n32098 );
and ( n32221 , n31830 , n32101 );
and ( n32222 , n31832 , n32103 );
and ( n32223 , n31834 , n32106 );
and ( n32224 , n31836 , n32108 );
and ( n32225 , n31838 , n32110 );
and ( n32226 , n31840 , n32112 );
and ( n32227 , n31842 , n32114 );
and ( n32228 , n31844 , n32116 );
and ( n32229 , n31846 , n32118 );
and ( n32230 , n31848 , n32120 );
and ( n32231 , n31850 , n32122 );
and ( n32232 , n31852 , n32124 );
and ( n32233 , n31854 , n32126 );
and ( n32234 , n31856 , n32128 );
or ( n32235 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 );
and ( n32236 , n31750 , n32095 );
and ( n32237 , n31778 , n32098 );
and ( n32238 , n31781 , n32101 );
and ( n32239 , n31784 , n32103 );
and ( n32240 , n31787 , n32106 );
and ( n32241 , n31790 , n32108 );
and ( n32242 , n31793 , n32110 );
and ( n32243 , n31796 , n32112 );
and ( n32244 , n31799 , n32114 );
and ( n32245 , n31802 , n32116 );
and ( n32246 , n31805 , n32118 );
and ( n32247 , n31808 , n32120 );
and ( n32248 , n31811 , n32122 );
and ( n32249 , n31814 , n32124 );
and ( n32250 , n31817 , n32126 );
and ( n32251 , n31820 , n32128 );
or ( n32252 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 );
and ( n32253 , n32130 , n32148 , n32166 , n32183 , n32201 , n32218 , n32235 , n32252 );
and ( n32254 , n32093 , n32253 );
not ( n32255 , n31689 );
buf ( n32256 , n31689 );
buf ( n32257 , n31689 );
buf ( n32258 , n31689 );
buf ( n32259 , n31689 );
buf ( n32260 , n31689 );
buf ( n32261 , n31689 );
buf ( n32262 , n31689 );
buf ( n32263 , n31689 );
buf ( n32264 , n31689 );
buf ( n32265 , n31689 );
buf ( n32266 , n31689 );
buf ( n32267 , n31689 );
buf ( n32268 , n31689 );
buf ( n32269 , n31689 );
buf ( n32270 , n31689 );
buf ( n32271 , n31689 );
buf ( n32272 , n31689 );
buf ( n32273 , n31689 );
buf ( n32274 , n31689 );
buf ( n32275 , n31689 );
buf ( n32276 , n31689 );
buf ( n32277 , n31689 );
buf ( n32278 , n31689 );
buf ( n32279 , n31689 );
buf ( n32280 , n31689 );
and ( n32281 , n31724 , n31723 );
or ( n32282 , n31721 , n31692 , n31694 , n31689 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 );
and ( n32283 , n32255 , n32282 );
not ( n32284 , n32283 );
and ( n32285 , n32284 , n31730 );
not ( n32286 , n31823 );
and ( n32287 , n31738 , n31739 );
and ( n32288 , n31737 , n32287 );
and ( n32289 , n31736 , n32288 );
and ( n32290 , n31735 , n32289 );
and ( n32291 , n31734 , n32290 );
and ( n32292 , n31733 , n32291 );
xor ( n32293 , n31732 , n32292 );
xor ( n32294 , n31733 , n32291 );
and ( n32295 , n32294 , n31823 );
xor ( n32296 , n31734 , n32290 );
and ( n32297 , n32296 , n31858 );
xor ( n32298 , n31735 , n32289 );
and ( n32299 , n32298 , n31893 );
xor ( n32300 , n31736 , n32288 );
and ( n32301 , n32300 , n31928 );
xor ( n32302 , n31737 , n32287 );
and ( n32303 , n32302 , n31963 );
xor ( n32304 , n31738 , n31739 );
and ( n32305 , n32304 , n31998 );
not ( n32306 , n31739 );
and ( n32307 , n32306 , n32033 );
and ( n32308 , n31740 , n32068 );
and ( n32309 , n32033 , n32308 );
and ( n32310 , n32306 , n32308 );
or ( n32311 , n32307 , n32309 , n32310 );
and ( n32312 , n31998 , n32311 );
and ( n32313 , n32304 , n32311 );
or ( n32314 , n32305 , n32312 , n32313 );
and ( n32315 , n31963 , n32314 );
and ( n32316 , n32302 , n32314 );
or ( n32317 , n32303 , n32315 , n32316 );
and ( n32318 , n31928 , n32317 );
and ( n32319 , n32300 , n32317 );
or ( n32320 , n32301 , n32318 , n32319 );
and ( n32321 , n31893 , n32320 );
and ( n32322 , n32298 , n32320 );
or ( n32323 , n32299 , n32321 , n32322 );
and ( n32324 , n31858 , n32323 );
and ( n32325 , n32296 , n32323 );
or ( n32326 , n32297 , n32324 , n32325 );
and ( n32327 , n31823 , n32326 );
and ( n32328 , n32294 , n32326 );
or ( n32329 , n32295 , n32327 , n32328 );
xor ( n32330 , n32293 , n32329 );
and ( n32331 , n32286 , n32330 );
and ( n32332 , n31739 , n31740 );
and ( n32333 , n31738 , n32332 );
and ( n32334 , n31737 , n32333 );
and ( n32335 , n31736 , n32334 );
and ( n32336 , n31735 , n32335 );
and ( n32337 , n31734 , n32336 );
and ( n32338 , n31733 , n32337 );
xor ( n32339 , n31732 , n32338 );
xor ( n32340 , n31733 , n32337 );
not ( n32341 , n31823 );
not ( n32342 , n32341 );
and ( n32343 , n32340 , n32342 );
xor ( n32344 , n31734 , n32336 );
not ( n32345 , n31858 );
not ( n32346 , n32345 );
and ( n32347 , n32344 , n32346 );
xor ( n32348 , n31735 , n32335 );
not ( n32349 , n31893 );
not ( n32350 , n32349 );
and ( n32351 , n32348 , n32350 );
xor ( n32352 , n31736 , n32334 );
not ( n32353 , n31928 );
not ( n32354 , n32353 );
and ( n32355 , n32352 , n32354 );
xor ( n32356 , n31737 , n32333 );
not ( n32357 , n31963 );
not ( n32358 , n32357 );
and ( n32359 , n32356 , n32358 );
xor ( n32360 , n31738 , n32332 );
not ( n32361 , n31998 );
not ( n32362 , n32361 );
and ( n32363 , n32360 , n32362 );
xor ( n32364 , n31739 , n31740 );
not ( n32365 , n32033 );
not ( n32366 , n32365 );
and ( n32367 , n32364 , n32366 );
not ( n32368 , n31740 );
not ( n32369 , n32068 );
not ( n32370 , n32369 );
or ( n32371 , n32368 , n32370 );
and ( n32372 , n32366 , n32371 );
and ( n32373 , n32364 , n32371 );
or ( n32374 , n32367 , n32372 , n32373 );
and ( n32375 , n32362 , n32374 );
and ( n32376 , n32360 , n32374 );
or ( n32377 , n32363 , n32375 , n32376 );
and ( n32378 , n32358 , n32377 );
and ( n32379 , n32356 , n32377 );
or ( n32380 , n32359 , n32378 , n32379 );
and ( n32381 , n32354 , n32380 );
and ( n32382 , n32352 , n32380 );
or ( n32383 , n32355 , n32381 , n32382 );
and ( n32384 , n32350 , n32383 );
and ( n32385 , n32348 , n32383 );
or ( n32386 , n32351 , n32384 , n32385 );
and ( n32387 , n32346 , n32386 );
and ( n32388 , n32344 , n32386 );
or ( n32389 , n32347 , n32387 , n32388 );
and ( n32390 , n32342 , n32389 );
and ( n32391 , n32340 , n32389 );
or ( n32392 , n32343 , n32390 , n32391 );
xnor ( n32393 , n32339 , n32392 );
and ( n32394 , n32393 , n31823 );
or ( n32395 , n32331 , n32394 );
and ( n32396 , n32395 , n32283 );
or ( n32397 , n32285 , n32396 );
and ( n32398 , n32130 , n32147 , n32166 , n32183 , n32201 , n32218 , n32235 , n32252 );
and ( n32399 , n32397 , n32398 );
not ( n32400 , n32130 );
not ( n32401 , n32183 );
not ( n32402 , n32252 );
and ( n32403 , n32400 , n32147 , n32165 , n32401 , n32201 , n32218 , n32235 , n32402 );
nor ( n32404 , n32130 , n32147 , n32165 , n32183 , n32201 , n32218 , n32235 , n32402 );
or ( n32405 , n32403 , n32404 );
and ( n32406 , n32400 , n32147 , n32166 , n32183 , n32201 , n32218 , n32235 , n32252 );
or ( n32407 , n32405 , n32406 );
not ( n32408 , n32235 );
and ( n32409 , n32400 , n32148 , n32166 , n32401 , n32200 , n32218 , n32408 , n32252 );
or ( n32410 , n32407 , n32409 );
and ( n32411 , n32400 , n32148 , n32166 , n32183 , n32200 , n32218 , n32408 , n32252 );
or ( n32412 , n32410 , n32411 );
and ( n32413 , n32130 , n32147 , n32166 , n32183 , n32200 , n32218 , n32408 , n32252 );
or ( n32414 , n32412 , n32413 );
nor ( n32415 , n32400 , n32148 , n32165 , n32401 , n32200 , n32218 , n32235 , n32402 );
or ( n32416 , n32414 , n32415 );
nor ( n32417 , n32400 , n32147 , n32165 , n32401 , n32200 , n32218 , n32235 , n32402 );
or ( n32418 , n32416 , n32417 );
and ( n32419 , n32400 , n32148 , n32165 , n32401 , n32201 , n32218 , n32235 , n32252 );
or ( n32420 , n32418 , n32419 );
and ( n32421 , n32400 , n32147 , n32165 , n32401 , n32201 , n32218 , n32235 , n32252 );
or ( n32422 , n32420 , n32421 );
nor ( n32423 , n32130 , n32147 , n32166 , n32183 , n32200 , n32218 , n32235 , n32252 );
or ( n32424 , n32422 , n32423 );
nor ( n32425 , n32400 , n32147 , n32166 , n32183 , n32200 , n32218 , n32235 , n32252 );
or ( n32426 , n32424 , n32425 );
nor ( n32427 , n32130 , n32147 , n32165 , n32183 , n32201 , n32218 , n32408 , n32402 );
or ( n32428 , n32426 , n32427 );
nor ( n32429 , n32130 , n32147 , n32165 , n32183 , n32200 , n32218 , n32408 , n32402 );
or ( n32430 , n32428 , n32429 );
nor ( n32431 , n32130 , n32147 , n32165 , n32183 , n32200 , n32218 , n32408 , n32252 );
or ( n32432 , n32430 , n32431 );
nor ( n32433 , n32400 , n32148 , n32165 , n32183 , n32200 , n32218 , n32408 , n32252 );
or ( n32434 , n32432 , n32433 );
nor ( n32435 , n32404 , n32403 , n32398 , n32253 , n32406 , n32409 , n32411 , n32413 , n32415 , n32417 , n32419 , n32421 , n32423 , n32425 , n32427 , n32429 , n32431 , n32433 );
or ( n32436 , n32434 , n32435 );
and ( n32437 , n31730 , n32436 );
or ( n32438 , n32254 , n32399 , n32437 );
buf ( n32439 , RI15b5d588_1050);
buf ( n32440 , RI15b5d6f0_1053);
buf ( n32441 , RI15b5d600_1051);
buf ( n32442 , RI15b5d678_1052);
or ( n32443 , n32441 , n32442 );
and ( n32444 , n32440 , n32443 );
not ( n32445 , n32444 );
and ( n32446 , n32445 , n32441 );
buf ( n32447 , n32446 );
not ( n32448 , n32447 );
not ( n32449 , n32444 );
and ( n32450 , n32449 , n32442 );
buf ( n32451 , n32450 );
not ( n32452 , n32444 );
and ( n32453 , n32452 , n32440 );
buf ( n32454 , n32453 );
not ( n32455 , n32454 );
and ( n32456 , n32439 , n32448 , n32451 , n32455 );
and ( n32457 , n32438 , n32456 );
buf ( n32458 , RI15b62e98_1240);
buf ( n32459 , RI15b62e20_1239);
buf ( n32460 , RI15b62da8_1238);
buf ( n32461 , RI15b62d30_1237);
buf ( n32462 , RI15b62cb8_1236);
buf ( n32463 , RI15b62c40_1235);
buf ( n32464 , RI15b62bc8_1234);
and ( n32465 , n32463 , n32464 );
and ( n32466 , n32462 , n32465 );
and ( n32467 , n32461 , n32466 );
and ( n32468 , n32460 , n32467 );
and ( n32469 , n32459 , n32468 );
and ( n32470 , n32458 , n32469 );
xor ( n32471 , n31730 , n32470 );
not ( n32472 , n32439 );
and ( n32473 , n32472 , n32448 , n32451 , n32455 );
and ( n32474 , n32471 , n32473 );
buf ( n32475 , RI15b606c0_1155);
not ( n32476 , n32475 );
and ( n32477 , n32476 , n32471 );
and ( n32478 , n32462 , n32463 );
and ( n32479 , n32461 , n32478 );
and ( n32480 , n32460 , n32479 );
and ( n32481 , n32459 , n32480 );
and ( n32482 , n32458 , n32481 );
xor ( n32483 , n31730 , n32482 );
and ( n32484 , n32483 , n32475 );
or ( n32485 , n32477 , n32484 );
nor ( n32486 , n32439 , n32448 , n32451 , n32454 );
and ( n32487 , n32485 , n32486 );
buf ( n32488 , RI15b63e10_1273);
nor ( n32489 , n32439 , n32447 , n32451 , n32454 );
and ( n32490 , n32488 , n32489 );
nor ( n32491 , n32472 , n32447 , n32451 , n32454 );
nor ( n32492 , n32472 , n32448 , n32451 , n32454 );
or ( n32493 , n32491 , n32492 );
and ( n32494 , n32472 , n32447 , n32451 , n32455 );
or ( n32495 , n32493 , n32494 );
and ( n32496 , n32439 , n32447 , n32451 , n32455 );
or ( n32497 , n32495 , n32496 );
nor ( n32498 , n32439 , n32447 , n32451 , n32455 );
or ( n32499 , n32497 , n32498 );
nor ( n32500 , n32472 , n32447 , n32451 , n32455 );
or ( n32501 , n32499 , n32500 );
and ( n32502 , n31730 , n32501 );
or ( n32503 , C0 , n32457 , n32474 , n32487 , n32490 , n32502 );
buf ( n32504 , n32503 );
buf ( n32505 , n32504 );
buf ( n32506 , n31655 );
buf ( n32507 , n31655 );
buf ( n32508 , n30987 );
buf ( n32509 , n30987 );
buf ( n32510 , RI15b4b090_425);
buf ( n32511 , RI15b44cb8_212);
not ( n32512 , n32511 );
buf ( n32513 , RI15b44e20_215);
buf ( n32514 , RI15b44d30_213);
buf ( n32515 , RI15b44da8_214);
or ( n32516 , n32514 , n32515 );
and ( n32517 , n32513 , n32516 );
not ( n32518 , n32517 );
and ( n32519 , n32518 , n32514 );
buf ( n32520 , n32519 );
not ( n32521 , n32517 );
and ( n32522 , n32521 , n32515 );
buf ( n32523 , n32522 );
not ( n32524 , n32517 );
and ( n32525 , n32524 , n32513 );
buf ( n32526 , n32525 );
not ( n32527 , n32526 );
nor ( n32528 , n32512 , n32520 , n32523 , n32527 );
and ( n32529 , n32510 , n32528 );
buf ( n32530 , RI15b3fe70_45);
buf ( n32531 , RI15b44bc8_210);
not ( n32532 , n32531 );
and ( n32533 , n32530 , n32532 );
buf ( n32534 , RI15b3fdf8_44);
buf ( n32535 , RI15b44b50_209);
not ( n32536 , n32535 );
and ( n32537 , n32534 , n32536 );
buf ( n32538 , RI15b3fd80_43);
buf ( n32539 , RI15b44ad8_208);
not ( n32540 , n32539 );
and ( n32541 , n32538 , n32540 );
buf ( n32542 , RI15b3fd08_42);
buf ( n32543 , RI15b44a60_207);
not ( n32544 , n32543 );
and ( n32545 , n32542 , n32544 );
buf ( n32546 , RI15b3fc90_41);
buf ( n32547 , RI15b449e8_206);
not ( n32548 , n32547 );
or ( n32549 , n32546 , n32548 );
and ( n32550 , n32544 , n32549 );
and ( n32551 , n32542 , n32549 );
or ( n32552 , n32545 , n32550 , n32551 );
and ( n32553 , n32540 , n32552 );
and ( n32554 , n32538 , n32552 );
or ( n32555 , n32541 , n32553 , n32554 );
and ( n32556 , n32536 , n32555 );
and ( n32557 , n32534 , n32555 );
or ( n32558 , n32537 , n32556 , n32557 );
and ( n32559 , n32532 , n32558 );
and ( n32560 , n32530 , n32558 );
or ( n32561 , n32533 , n32559 , n32560 );
not ( n32562 , n32561 );
not ( n32563 , n32562 );
xor ( n32564 , n32538 , n32540 );
xor ( n32565 , n32564 , n32552 );
xor ( n32566 , n32534 , n32536 );
xor ( n32567 , n32566 , n32555 );
xor ( n32568 , n32530 , n32532 );
xor ( n32569 , n32568 , n32558 );
buf ( n32570 , n32562 );
buf ( n32571 , n32562 );
buf ( n32572 , n32562 );
buf ( n32573 , n32562 );
buf ( n32574 , n32562 );
buf ( n32575 , n32562 );
buf ( n32576 , n32562 );
buf ( n32577 , n32562 );
buf ( n32578 , n32562 );
buf ( n32579 , n32562 );
buf ( n32580 , n32562 );
buf ( n32581 , n32562 );
buf ( n32582 , n32562 );
buf ( n32583 , n32562 );
buf ( n32584 , n32562 );
buf ( n32585 , n32562 );
buf ( n32586 , n32562 );
buf ( n32587 , n32562 );
buf ( n32588 , n32562 );
buf ( n32589 , n32562 );
buf ( n32590 , n32562 );
buf ( n32591 , n32562 );
buf ( n32592 , n32562 );
buf ( n32593 , n32562 );
buf ( n32594 , n32562 );
xor ( n32595 , n32542 , n32544 );
xor ( n32596 , n32595 , n32549 );
or ( n32597 , n32565 , n32567 , n32569 , n32562 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32596 );
and ( n32598 , n32563 , n32597 );
not ( n32599 , n32598 );
buf ( n32600 , RI15b4bf90_457);
and ( n32601 , n32599 , n32600 );
buf ( n32602 , n32601 );
buf ( n32603 , RI15b43728_166);
not ( n32604 , n32531 );
and ( n32605 , n32547 , n32543 , n32539 , n32535 , n32604 );
and ( n32606 , n32603 , n32605 );
buf ( n32607 , RI15b43368_158);
not ( n32608 , n32547 );
and ( n32609 , n32608 , n32543 , n32539 , n32535 , n32604 );
and ( n32610 , n32607 , n32609 );
buf ( n32611 , RI15b42fa8_150);
not ( n32612 , n32543 );
and ( n32613 , n32547 , n32612 , n32539 , n32535 , n32604 );
and ( n32614 , n32611 , n32613 );
buf ( n32615 , RI15b42be8_142);
and ( n32616 , n32608 , n32612 , n32539 , n32535 , n32604 );
and ( n32617 , n32615 , n32616 );
buf ( n32618 , RI15b42828_134);
not ( n32619 , n32539 );
and ( n32620 , n32547 , n32543 , n32619 , n32535 , n32604 );
and ( n32621 , n32618 , n32620 );
buf ( n32622 , RI15b42468_126);
and ( n32623 , n32608 , n32543 , n32619 , n32535 , n32604 );
and ( n32624 , n32622 , n32623 );
buf ( n32625 , RI15b420a8_118);
and ( n32626 , n32547 , n32612 , n32619 , n32535 , n32604 );
and ( n32627 , n32625 , n32626 );
buf ( n32628 , RI15b41ce8_110);
and ( n32629 , n32608 , n32612 , n32619 , n32535 , n32604 );
and ( n32630 , n32628 , n32629 );
buf ( n32631 , RI15b41928_102);
nor ( n32632 , n32608 , n32612 , n32619 , n32535 , n32531 );
and ( n32633 , n32631 , n32632 );
buf ( n32634 , RI15b41568_94);
nor ( n32635 , n32547 , n32612 , n32619 , n32535 , n32531 );
and ( n32636 , n32634 , n32635 );
buf ( n32637 , RI15b411a8_86);
nor ( n32638 , n32608 , n32543 , n32619 , n32535 , n32531 );
and ( n32639 , n32637 , n32638 );
buf ( n32640 , RI15b40de8_78);
nor ( n32641 , n32547 , n32543 , n32619 , n32535 , n32531 );
and ( n32642 , n32640 , n32641 );
buf ( n32643 , RI15b40a28_70);
nor ( n32644 , n32608 , n32612 , n32539 , n32535 , n32531 );
and ( n32645 , n32643 , n32644 );
buf ( n32646 , RI15b40668_62);
nor ( n32647 , n32547 , n32612 , n32539 , n32535 , n32531 );
and ( n32648 , n32646 , n32647 );
buf ( n32649 , RI15b402a8_54);
nor ( n32650 , n32608 , n32543 , n32539 , n32535 , n32531 );
and ( n32651 , n32649 , n32650 );
buf ( n32652 , RI15b3fee8_46);
nor ( n32653 , n32547 , n32543 , n32539 , n32535 , n32531 );
and ( n32654 , n32652 , n32653 );
or ( n32655 , n32606 , n32610 , n32614 , n32617 , n32621 , n32624 , n32627 , n32630 , n32633 , n32636 , n32639 , n32642 , n32645 , n32648 , n32651 , n32654 );
not ( n32656 , n32655 );
buf ( n32657 , RI15b437a0_167);
and ( n32658 , n32657 , n32605 );
buf ( n32659 , RI15b433e0_159);
and ( n32660 , n32659 , n32609 );
buf ( n32661 , RI15b43020_151);
and ( n32662 , n32661 , n32613 );
buf ( n32663 , RI15b42c60_143);
and ( n32664 , n32663 , n32616 );
buf ( n32665 , RI15b428a0_135);
and ( n32666 , n32665 , n32620 );
buf ( n32667 , RI15b424e0_127);
and ( n32668 , n32667 , n32623 );
buf ( n32669 , RI15b42120_119);
and ( n32670 , n32669 , n32626 );
buf ( n32671 , RI15b41d60_111);
and ( n32672 , n32671 , n32629 );
buf ( n32673 , RI15b419a0_103);
and ( n32674 , n32673 , n32632 );
buf ( n32675 , RI15b415e0_95);
and ( n32676 , n32675 , n32635 );
buf ( n32677 , RI15b41220_87);
and ( n32678 , n32677 , n32638 );
buf ( n32679 , RI15b40e60_79);
and ( n32680 , n32679 , n32641 );
buf ( n32681 , RI15b40aa0_71);
and ( n32682 , n32681 , n32644 );
buf ( n32683 , RI15b406e0_63);
and ( n32684 , n32683 , n32647 );
buf ( n32685 , RI15b40320_55);
and ( n32686 , n32685 , n32650 );
buf ( n32687 , RI15b3ff60_47);
and ( n32688 , n32687 , n32653 );
or ( n32689 , n32658 , n32660 , n32662 , n32664 , n32666 , n32668 , n32670 , n32672 , n32674 , n32676 , n32678 , n32680 , n32682 , n32684 , n32686 , n32688 );
buf ( n32690 , RI15b43818_168);
and ( n32691 , n32690 , n32605 );
buf ( n32692 , RI15b43458_160);
and ( n32693 , n32692 , n32609 );
buf ( n32694 , RI15b43098_152);
and ( n32695 , n32694 , n32613 );
buf ( n32696 , RI15b42cd8_144);
and ( n32697 , n32696 , n32616 );
buf ( n32698 , RI15b42918_136);
and ( n32699 , n32698 , n32620 );
buf ( n32700 , RI15b42558_128);
and ( n32701 , n32700 , n32623 );
buf ( n32702 , RI15b42198_120);
and ( n32703 , n32702 , n32626 );
buf ( n32704 , RI15b41dd8_112);
and ( n32705 , n32704 , n32629 );
buf ( n32706 , RI15b41a18_104);
and ( n32707 , n32706 , n32632 );
buf ( n32708 , RI15b41658_96);
and ( n32709 , n32708 , n32635 );
buf ( n32710 , RI15b41298_88);
and ( n32711 , n32710 , n32638 );
buf ( n32712 , RI15b40ed8_80);
and ( n32713 , n32712 , n32641 );
buf ( n32714 , RI15b40b18_72);
and ( n32715 , n32714 , n32644 );
buf ( n32716 , RI15b40758_64);
and ( n32717 , n32716 , n32647 );
buf ( n32718 , RI15b40398_56);
and ( n32719 , n32718 , n32650 );
buf ( n32720 , RI15b3ffd8_48);
and ( n32721 , n32720 , n32653 );
or ( n32722 , n32691 , n32693 , n32695 , n32697 , n32699 , n32701 , n32703 , n32705 , n32707 , n32709 , n32711 , n32713 , n32715 , n32717 , n32719 , n32721 );
buf ( n32723 , RI15b43890_169);
and ( n32724 , n32723 , n32605 );
buf ( n32725 , RI15b434d0_161);
and ( n32726 , n32725 , n32609 );
buf ( n32727 , RI15b43110_153);
and ( n32728 , n32727 , n32613 );
buf ( n32729 , RI15b42d50_145);
and ( n32730 , n32729 , n32616 );
buf ( n32731 , RI15b42990_137);
and ( n32732 , n32731 , n32620 );
buf ( n32733 , RI15b425d0_129);
and ( n32734 , n32733 , n32623 );
buf ( n32735 , RI15b42210_121);
and ( n32736 , n32735 , n32626 );
buf ( n32737 , RI15b41e50_113);
and ( n32738 , n32737 , n32629 );
buf ( n32739 , RI15b41a90_105);
and ( n32740 , n32739 , n32632 );
buf ( n32741 , RI15b416d0_97);
and ( n32742 , n32741 , n32635 );
buf ( n32743 , RI15b41310_89);
and ( n32744 , n32743 , n32638 );
buf ( n32745 , RI15b40f50_81);
and ( n32746 , n32745 , n32641 );
buf ( n32747 , RI15b40b90_73);
and ( n32748 , n32747 , n32644 );
buf ( n32749 , RI15b407d0_65);
and ( n32750 , n32749 , n32647 );
buf ( n32751 , RI15b40410_57);
and ( n32752 , n32751 , n32650 );
buf ( n32753 , RI15b40050_49);
and ( n32754 , n32753 , n32653 );
or ( n32755 , n32724 , n32726 , n32728 , n32730 , n32732 , n32734 , n32736 , n32738 , n32740 , n32742 , n32744 , n32746 , n32748 , n32750 , n32752 , n32754 );
not ( n32756 , n32755 );
buf ( n32757 , RI15b43908_170);
and ( n32758 , n32757 , n32605 );
buf ( n32759 , RI15b43548_162);
and ( n32760 , n32759 , n32609 );
buf ( n32761 , RI15b43188_154);
and ( n32762 , n32761 , n32613 );
buf ( n32763 , RI15b42dc8_146);
and ( n32764 , n32763 , n32616 );
buf ( n32765 , RI15b42a08_138);
and ( n32766 , n32765 , n32620 );
buf ( n32767 , RI15b42648_130);
and ( n32768 , n32767 , n32623 );
buf ( n32769 , RI15b42288_122);
and ( n32770 , n32769 , n32626 );
buf ( n32771 , RI15b41ec8_114);
and ( n32772 , n32771 , n32629 );
buf ( n32773 , RI15b41b08_106);
and ( n32774 , n32773 , n32632 );
buf ( n32775 , RI15b41748_98);
and ( n32776 , n32775 , n32635 );
buf ( n32777 , RI15b41388_90);
and ( n32778 , n32777 , n32638 );
buf ( n32779 , RI15b40fc8_82);
and ( n32780 , n32779 , n32641 );
buf ( n32781 , RI15b40c08_74);
and ( n32782 , n32781 , n32644 );
buf ( n32783 , RI15b40848_66);
and ( n32784 , n32783 , n32647 );
buf ( n32785 , RI15b40488_58);
and ( n32786 , n32785 , n32650 );
buf ( n32787 , RI15b400c8_50);
and ( n32788 , n32787 , n32653 );
or ( n32789 , n32758 , n32760 , n32762 , n32764 , n32766 , n32768 , n32770 , n32772 , n32774 , n32776 , n32778 , n32780 , n32782 , n32784 , n32786 , n32788 );
not ( n32790 , n32789 );
buf ( n32791 , RI15b43980_171);
and ( n32792 , n32791 , n32605 );
buf ( n32793 , RI15b435c0_163);
and ( n32794 , n32793 , n32609 );
buf ( n32795 , RI15b43200_155);
and ( n32796 , n32795 , n32613 );
buf ( n32797 , RI15b42e40_147);
and ( n32798 , n32797 , n32616 );
buf ( n32799 , RI15b42a80_139);
and ( n32800 , n32799 , n32620 );
buf ( n32801 , RI15b426c0_131);
and ( n32802 , n32801 , n32623 );
buf ( n32803 , RI15b42300_123);
and ( n32804 , n32803 , n32626 );
buf ( n32805 , RI15b41f40_115);
and ( n32806 , n32805 , n32629 );
buf ( n32807 , RI15b41b80_107);
and ( n32808 , n32807 , n32632 );
buf ( n32809 , RI15b417c0_99);
and ( n32810 , n32809 , n32635 );
buf ( n32811 , RI15b41400_91);
and ( n32812 , n32811 , n32638 );
buf ( n32813 , RI15b41040_83);
and ( n32814 , n32813 , n32641 );
buf ( n32815 , RI15b40c80_75);
and ( n32816 , n32815 , n32644 );
buf ( n32817 , RI15b408c0_67);
and ( n32818 , n32817 , n32647 );
buf ( n32819 , RI15b40500_59);
and ( n32820 , n32819 , n32650 );
buf ( n32821 , RI15b40140_51);
and ( n32822 , n32821 , n32653 );
or ( n32823 , n32792 , n32794 , n32796 , n32798 , n32800 , n32802 , n32804 , n32806 , n32808 , n32810 , n32812 , n32814 , n32816 , n32818 , n32820 , n32822 );
buf ( n32824 , RI15b439f8_172);
and ( n32825 , n32824 , n32605 );
buf ( n32826 , RI15b43638_164);
and ( n32827 , n32826 , n32609 );
buf ( n32828 , RI15b43278_156);
and ( n32829 , n32828 , n32613 );
buf ( n32830 , RI15b42eb8_148);
and ( n32831 , n32830 , n32616 );
buf ( n32832 , RI15b42af8_140);
and ( n32833 , n32832 , n32620 );
buf ( n32834 , RI15b42738_132);
and ( n32835 , n32834 , n32623 );
buf ( n32836 , RI15b42378_124);
and ( n32837 , n32836 , n32626 );
buf ( n32838 , RI15b41fb8_116);
and ( n32839 , n32838 , n32629 );
buf ( n32840 , RI15b41bf8_108);
and ( n32841 , n32840 , n32632 );
buf ( n32842 , RI15b41838_100);
and ( n32843 , n32842 , n32635 );
buf ( n32844 , RI15b41478_92);
and ( n32845 , n32844 , n32638 );
buf ( n32846 , RI15b410b8_84);
and ( n32847 , n32846 , n32641 );
buf ( n32848 , RI15b40cf8_76);
and ( n32849 , n32848 , n32644 );
buf ( n32850 , RI15b40938_68);
and ( n32851 , n32850 , n32647 );
buf ( n32852 , RI15b40578_60);
and ( n32853 , n32852 , n32650 );
buf ( n32854 , RI15b401b8_52);
and ( n32855 , n32854 , n32653 );
or ( n32856 , n32825 , n32827 , n32829 , n32831 , n32833 , n32835 , n32837 , n32839 , n32841 , n32843 , n32845 , n32847 , n32849 , n32851 , n32853 , n32855 );
buf ( n32857 , RI15b43a70_173);
and ( n32858 , n32857 , n32605 );
buf ( n32859 , RI15b436b0_165);
and ( n32860 , n32859 , n32609 );
buf ( n32861 , RI15b432f0_157);
and ( n32862 , n32861 , n32613 );
buf ( n32863 , RI15b42f30_149);
and ( n32864 , n32863 , n32616 );
buf ( n32865 , RI15b42b70_141);
and ( n32866 , n32865 , n32620 );
buf ( n32867 , RI15b427b0_133);
and ( n32868 , n32867 , n32623 );
buf ( n32869 , RI15b423f0_125);
and ( n32870 , n32869 , n32626 );
buf ( n32871 , RI15b42030_117);
and ( n32872 , n32871 , n32629 );
buf ( n32873 , RI15b41c70_109);
and ( n32874 , n32873 , n32632 );
buf ( n32875 , RI15b418b0_101);
and ( n32876 , n32875 , n32635 );
buf ( n32877 , RI15b414f0_93);
and ( n32878 , n32877 , n32638 );
buf ( n32879 , RI15b41130_85);
and ( n32880 , n32879 , n32641 );
buf ( n32881 , RI15b40d70_77);
and ( n32882 , n32881 , n32644 );
buf ( n32883 , RI15b409b0_69);
and ( n32884 , n32883 , n32647 );
buf ( n32885 , RI15b405f0_61);
and ( n32886 , n32885 , n32650 );
buf ( n32887 , RI15b40230_53);
and ( n32888 , n32887 , n32653 );
or ( n32889 , n32858 , n32860 , n32862 , n32864 , n32866 , n32868 , n32870 , n32872 , n32874 , n32876 , n32878 , n32880 , n32882 , n32884 , n32886 , n32888 );
and ( n32890 , n32656 , n32689 , n32722 , n32756 , n32790 , n32823 , n32856 , n32889 );
and ( n32891 , n32602 , n32890 );
not ( n32892 , n32562 );
buf ( n32893 , n32562 );
buf ( n32894 , n32562 );
buf ( n32895 , n32562 );
buf ( n32896 , n32562 );
buf ( n32897 , n32562 );
buf ( n32898 , n32562 );
buf ( n32899 , n32562 );
buf ( n32900 , n32562 );
buf ( n32901 , n32562 );
buf ( n32902 , n32562 );
buf ( n32903 , n32562 );
buf ( n32904 , n32562 );
buf ( n32905 , n32562 );
buf ( n32906 , n32562 );
buf ( n32907 , n32562 );
buf ( n32908 , n32562 );
buf ( n32909 , n32562 );
buf ( n32910 , n32562 );
buf ( n32911 , n32562 );
buf ( n32912 , n32562 );
buf ( n32913 , n32562 );
buf ( n32914 , n32562 );
buf ( n32915 , n32562 );
buf ( n32916 , n32562 );
buf ( n32917 , n32562 );
or ( n32918 , n32565 , n32567 , n32569 , n32562 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32596 );
and ( n32919 , n32892 , n32918 );
not ( n32920 , n32919 );
and ( n32921 , n32920 , n32600 );
buf ( n32922 , n32921 );
not ( n32923 , n32689 );
and ( n32924 , n32656 , n32923 , n32722 , n32756 , n32790 , n32823 , n32856 , n32889 );
and ( n32925 , n32922 , n32924 );
not ( n32926 , n32562 );
buf ( n32927 , n32562 );
buf ( n32928 , n32562 );
buf ( n32929 , n32562 );
buf ( n32930 , n32562 );
buf ( n32931 , n32562 );
buf ( n32932 , n32562 );
buf ( n32933 , n32562 );
buf ( n32934 , n32562 );
buf ( n32935 , n32562 );
buf ( n32936 , n32562 );
buf ( n32937 , n32562 );
buf ( n32938 , n32562 );
buf ( n32939 , n32562 );
buf ( n32940 , n32562 );
buf ( n32941 , n32562 );
buf ( n32942 , n32562 );
buf ( n32943 , n32562 );
buf ( n32944 , n32562 );
buf ( n32945 , n32562 );
buf ( n32946 , n32562 );
buf ( n32947 , n32562 );
buf ( n32948 , n32562 );
buf ( n32949 , n32562 );
buf ( n32950 , n32562 );
buf ( n32951 , n32562 );
or ( n32952 , n32565 , n32567 , n32569 , n32562 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32596 );
and ( n32953 , n32926 , n32952 );
not ( n32954 , n32953 );
and ( n32955 , n32954 , n32600 );
buf ( n32956 , RI15b48318_328);
buf ( n32957 , RI15b48390_329);
not ( n32958 , n32957 );
buf ( n32959 , RI15b48408_330);
nor ( n32960 , n32956 , n32958 , n32959 );
not ( n32961 , n32956 );
and ( n32962 , n32961 , n32958 , n32959 );
or ( n32963 , n32960 , n32962 );
buf ( n32964 , RI15b668b8_1364);
buf ( n32965 , RI15b3fba0_39);
and ( n32966 , n32964 , n32965 );
not ( n32967 , n32966 );
buf ( n32968 , RI15b47df0_317);
not ( n32969 , n32968 );
and ( n32970 , n32967 , n32969 );
and ( n32971 , n32963 , n32970 );
not ( n32972 , n32971 );
buf ( n32973 , RI15b4a190_393);
and ( n32974 , n32972 , n32973 );
buf ( n32975 , RI15b4bf18_456);
buf ( n32976 , RI15b4bea0_455);
buf ( n32977 , RI15b4be28_454);
buf ( n32978 , RI15b4bdb0_453);
buf ( n32979 , RI15b4bd38_452);
buf ( n32980 , RI15b4bcc0_451);
buf ( n32981 , RI15b4bc48_450);
buf ( n32982 , RI15b4bbd0_449);
buf ( n32983 , RI15b4bb58_448);
buf ( n32984 , RI15b4bae0_447);
buf ( n32985 , RI15b4ba68_446);
buf ( n32986 , RI15b4b9f0_445);
buf ( n32987 , RI15b4b978_444);
buf ( n32988 , RI15b4b900_443);
buf ( n32989 , RI15b4b888_442);
buf ( n32990 , RI15b4b810_441);
buf ( n32991 , RI15b4b798_440);
buf ( n32992 , RI15b4b720_439);
buf ( n32993 , RI15b4b6a8_438);
buf ( n32994 , RI15b4b630_437);
buf ( n32995 , RI15b4b5b8_436);
buf ( n32996 , RI15b4b540_435);
buf ( n32997 , RI15b4b4c8_434);
buf ( n32998 , RI15b4b450_433);
buf ( n32999 , RI15b4b3d8_432);
buf ( n33000 , RI15b4b360_431);
buf ( n33001 , RI15b4b2e8_430);
buf ( n33002 , RI15b4b270_429);
buf ( n33003 , RI15b4b1f8_428);
and ( n33004 , n33002 , n33003 );
and ( n33005 , n33001 , n33004 );
and ( n33006 , n33000 , n33005 );
and ( n33007 , n32999 , n33006 );
and ( n33008 , n32998 , n33007 );
and ( n33009 , n32997 , n33008 );
and ( n33010 , n32996 , n33009 );
and ( n33011 , n32995 , n33010 );
and ( n33012 , n32994 , n33011 );
and ( n33013 , n32993 , n33012 );
and ( n33014 , n32992 , n33013 );
and ( n33015 , n32991 , n33014 );
and ( n33016 , n32990 , n33015 );
and ( n33017 , n32989 , n33016 );
and ( n33018 , n32988 , n33017 );
and ( n33019 , n32987 , n33018 );
and ( n33020 , n32986 , n33019 );
and ( n33021 , n32985 , n33020 );
and ( n33022 , n32984 , n33021 );
and ( n33023 , n32983 , n33022 );
and ( n33024 , n32982 , n33023 );
and ( n33025 , n32981 , n33024 );
and ( n33026 , n32980 , n33025 );
and ( n33027 , n32979 , n33026 );
and ( n33028 , n32978 , n33027 );
and ( n33029 , n32977 , n33028 );
and ( n33030 , n32976 , n33029 );
and ( n33031 , n32975 , n33030 );
xor ( n33032 , n32600 , n33031 );
and ( n33033 , n33032 , n32971 );
or ( n33034 , n32974 , n33033 );
and ( n33035 , n33034 , n32953 );
or ( n33036 , n32955 , n33035 );
not ( n33037 , n32889 );
nor ( n33038 , n32656 , n32689 , n32722 , n32756 , n32789 , n32823 , n32856 , n33037 );
and ( n33039 , n33036 , n33038 );
not ( n33040 , n32562 );
buf ( n33041 , n32562 );
buf ( n33042 , n32562 );
buf ( n33043 , n32562 );
buf ( n33044 , n32562 );
buf ( n33045 , n32562 );
buf ( n33046 , n32562 );
buf ( n33047 , n32562 );
buf ( n33048 , n32562 );
buf ( n33049 , n32562 );
buf ( n33050 , n32562 );
buf ( n33051 , n32562 );
buf ( n33052 , n32562 );
buf ( n33053 , n32562 );
buf ( n33054 , n32562 );
buf ( n33055 , n32562 );
buf ( n33056 , n32562 );
buf ( n33057 , n32562 );
buf ( n33058 , n32562 );
buf ( n33059 , n32562 );
buf ( n33060 , n32562 );
buf ( n33061 , n32562 );
buf ( n33062 , n32562 );
buf ( n33063 , n32562 );
buf ( n33064 , n32562 );
buf ( n33065 , n32562 );
or ( n33066 , n32565 , n32567 , n32569 , n32562 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n32596 );
and ( n33067 , n33040 , n33066 );
not ( n33068 , n33067 );
and ( n33069 , n33068 , n32600 );
not ( n33070 , n32970 );
buf ( n33071 , RI15b4a208_394);
not ( n33072 , n33071 );
and ( n33073 , n33072 , n32973 );
not ( n33074 , n32973 );
buf ( n33075 , RI15b4a118_392);
not ( n33076 , n33075 );
buf ( n33077 , RI15b4a0a0_391);
not ( n33078 , n33077 );
buf ( n33079 , RI15b4a028_390);
not ( n33080 , n33079 );
buf ( n33081 , RI15b49fb0_389);
not ( n33082 , n33081 );
buf ( n33083 , RI15b49f38_388);
not ( n33084 , n33083 );
buf ( n33085 , RI15b49ec0_387);
not ( n33086 , n33085 );
buf ( n33087 , RI15b49e48_386);
not ( n33088 , n33087 );
buf ( n33089 , RI15b49dd0_385);
not ( n33090 , n33089 );
buf ( n33091 , RI15b49d58_384);
not ( n33092 , n33091 );
buf ( n33093 , RI15b49ce0_383);
not ( n33094 , n33093 );
buf ( n33095 , RI15b49c68_382);
not ( n33096 , n33095 );
buf ( n33097 , RI15b49bf0_381);
not ( n33098 , n33097 );
buf ( n33099 , RI15b49b78_380);
not ( n33100 , n33099 );
buf ( n33101 , RI15b49b00_379);
not ( n33102 , n33101 );
buf ( n33103 , RI15b49a88_378);
not ( n33104 , n33103 );
buf ( n33105 , RI15b49a10_377);
not ( n33106 , n33105 );
buf ( n33107 , RI15b49998_376);
not ( n33108 , n33107 );
buf ( n33109 , RI15b49920_375);
not ( n33110 , n33109 );
buf ( n33111 , RI15b498a8_374);
not ( n33112 , n33111 );
buf ( n33113 , RI15b49830_373);
not ( n33114 , n33113 );
buf ( n33115 , RI15b497b8_372);
not ( n33116 , n33115 );
buf ( n33117 , RI15b49740_371);
not ( n33118 , n33117 );
buf ( n33119 , RI15b496c8_370);
not ( n33120 , n33119 );
buf ( n33121 , RI15b49650_369);
not ( n33122 , n33121 );
buf ( n33123 , RI15b495d8_368);
not ( n33124 , n33123 );
buf ( n33125 , RI15b49560_367);
not ( n33126 , n33125 );
buf ( n33127 , RI15b494e8_366);
not ( n33128 , n33127 );
buf ( n33129 , RI15b49470_365);
not ( n33130 , n33129 );
buf ( n33131 , RI15b493f8_364);
not ( n33132 , n33131 );
buf ( n33133 , RI15b49380_363);
not ( n33134 , n33133 );
and ( n33135 , n33132 , n33134 );
and ( n33136 , n33130 , n33135 );
and ( n33137 , n33128 , n33136 );
and ( n33138 , n33126 , n33137 );
and ( n33139 , n33124 , n33138 );
and ( n33140 , n33122 , n33139 );
and ( n33141 , n33120 , n33140 );
and ( n33142 , n33118 , n33141 );
and ( n33143 , n33116 , n33142 );
and ( n33144 , n33114 , n33143 );
and ( n33145 , n33112 , n33144 );
and ( n33146 , n33110 , n33145 );
and ( n33147 , n33108 , n33146 );
and ( n33148 , n33106 , n33147 );
and ( n33149 , n33104 , n33148 );
and ( n33150 , n33102 , n33149 );
and ( n33151 , n33100 , n33150 );
and ( n33152 , n33098 , n33151 );
and ( n33153 , n33096 , n33152 );
and ( n33154 , n33094 , n33153 );
and ( n33155 , n33092 , n33154 );
and ( n33156 , n33090 , n33155 );
and ( n33157 , n33088 , n33156 );
and ( n33158 , n33086 , n33157 );
and ( n33159 , n33084 , n33158 );
and ( n33160 , n33082 , n33159 );
and ( n33161 , n33080 , n33160 );
and ( n33162 , n33078 , n33161 );
and ( n33163 , n33076 , n33162 );
xor ( n33164 , n33074 , n33163 );
and ( n33165 , n33164 , n33071 );
or ( n33166 , n33073 , n33165 );
and ( n33167 , n33070 , n33166 );
and ( n33168 , n33032 , n32970 );
or ( n33169 , n33167 , n33168 );
and ( n33170 , n33169 , n33067 );
or ( n33171 , n33069 , n33170 );
nor ( n33172 , n32656 , n32923 , n32722 , n32756 , n32789 , n32823 , n32856 , n33037 );
and ( n33173 , n33171 , n33172 );
and ( n33174 , n32656 , n32689 , n32722 , n32756 , n32790 , n32823 , n32856 , n33037 );
nor ( n33175 , n32655 , n32689 , n32722 , n32755 , n32790 , n32823 , n32856 , n33037 );
or ( n33176 , n33174 , n33175 );
not ( n33177 , n32722 );
and ( n33178 , n32655 , n32689 , n33177 , n32755 , n32790 , n32823 , n32856 , n32889 );
or ( n33179 , n33176 , n33178 );
and ( n33180 , n32655 , n32923 , n33177 , n32755 , n32790 , n32823 , n32856 , n32889 );
or ( n33181 , n33179 , n33180 );
and ( n33182 , n32656 , n32689 , n33177 , n32755 , n32790 , n32823 , n32856 , n32889 );
or ( n33183 , n33181 , n33182 );
not ( n33184 , n32856 );
and ( n33185 , n32656 , n32923 , n33177 , n32756 , n32789 , n32823 , n33184 , n32889 );
or ( n33186 , n33183 , n33185 );
and ( n33187 , n32656 , n32923 , n33177 , n32755 , n32789 , n32823 , n33184 , n32889 );
or ( n33188 , n33186 , n33187 );
and ( n33189 , n32655 , n32689 , n33177 , n32755 , n32789 , n32823 , n33184 , n32889 );
or ( n33190 , n33188 , n33189 );
nor ( n33191 , n32655 , n32689 , n33177 , n32755 , n32789 , n32823 , n32856 , n32889 );
or ( n33192 , n33190 , n33191 );
nor ( n33193 , n32656 , n32689 , n33177 , n32755 , n32789 , n32823 , n32856 , n32889 );
or ( n33194 , n33192 , n33193 );
nor ( n33195 , n32655 , n32689 , n32722 , n32755 , n32790 , n32823 , n33184 , n33037 );
or ( n33196 , n33194 , n33195 );
nor ( n33197 , n32655 , n32689 , n32722 , n32755 , n32789 , n32823 , n33184 , n33037 );
or ( n33198 , n33196 , n33197 );
nor ( n33199 , n32655 , n32689 , n32722 , n32755 , n32789 , n32823 , n33184 , n32889 );
or ( n33200 , n33198 , n33199 );
nor ( n33201 , n32656 , n32923 , n32722 , n32755 , n32789 , n32823 , n33184 , n32889 );
or ( n33202 , n33200 , n33201 );
nor ( n33203 , n33175 , n33174 , n33178 , n33180 , n33182 , n33185 , n33187 , n33189 , n33172 , n33038 , n32924 , n32890 , n33191 , n33193 , n33195 , n33197 , n33199 , n33201 );
or ( n33204 , n33202 , n33203 );
and ( n33205 , n32600 , n33204 );
or ( n33206 , n32891 , n32925 , n33039 , n33173 , n33205 );
not ( n33207 , n32520 );
and ( n33208 , n32511 , n33207 , n32523 , n32527 );
and ( n33209 , n33206 , n33208 );
not ( n33210 , n32968 );
buf ( n33211 , RI15b4b108_426);
buf ( n33212 , RI15b4b018_424);
buf ( n33213 , RI15b4afa0_423);
buf ( n33214 , RI15b4af28_422);
buf ( n33215 , RI15b4aeb0_421);
buf ( n33216 , RI15b4ae38_420);
buf ( n33217 , RI15b4adc0_419);
buf ( n33218 , RI15b4ad48_418);
buf ( n33219 , RI15b4acd0_417);
buf ( n33220 , RI15b4ac58_416);
buf ( n33221 , RI15b4abe0_415);
buf ( n33222 , RI15b4ab68_414);
buf ( n33223 , RI15b4aaf0_413);
buf ( n33224 , RI15b4aa78_412);
buf ( n33225 , RI15b4aa00_411);
buf ( n33226 , RI15b4a988_410);
buf ( n33227 , RI15b4a910_409);
buf ( n33228 , RI15b4a898_408);
buf ( n33229 , RI15b4a820_407);
buf ( n33230 , RI15b4a7a8_406);
buf ( n33231 , RI15b4a730_405);
buf ( n33232 , RI15b4a6b8_404);
buf ( n33233 , RI15b4a640_403);
buf ( n33234 , RI15b4a5c8_402);
buf ( n33235 , RI15b4a550_401);
buf ( n33236 , RI15b4a4d8_400);
buf ( n33237 , RI15b4a460_399);
buf ( n33238 , RI15b4a3e8_398);
buf ( n33239 , RI15b4a370_397);
buf ( n33240 , RI15b4a2f8_396);
and ( n33241 , n33239 , n33240 );
and ( n33242 , n33238 , n33241 );
and ( n33243 , n33237 , n33242 );
and ( n33244 , n33236 , n33243 );
and ( n33245 , n33235 , n33244 );
and ( n33246 , n33234 , n33245 );
and ( n33247 , n33233 , n33246 );
and ( n33248 , n33232 , n33247 );
and ( n33249 , n33231 , n33248 );
and ( n33250 , n33230 , n33249 );
and ( n33251 , n33229 , n33250 );
and ( n33252 , n33228 , n33251 );
and ( n33253 , n33227 , n33252 );
and ( n33254 , n33226 , n33253 );
and ( n33255 , n33225 , n33254 );
and ( n33256 , n33224 , n33255 );
and ( n33257 , n33223 , n33256 );
and ( n33258 , n33222 , n33257 );
and ( n33259 , n33221 , n33258 );
and ( n33260 , n33220 , n33259 );
and ( n33261 , n33219 , n33260 );
and ( n33262 , n33218 , n33261 );
and ( n33263 , n33217 , n33262 );
and ( n33264 , n33216 , n33263 );
and ( n33265 , n33215 , n33264 );
and ( n33266 , n33214 , n33265 );
and ( n33267 , n33213 , n33266 );
and ( n33268 , n33212 , n33267 );
and ( n33269 , n32510 , n33268 );
xor ( n33270 , n33211 , n33269 );
not ( n33271 , n33270 );
xor ( n33272 , n32510 , n33268 );
and ( n33273 , n33271 , n33272 );
not ( n33274 , n33272 );
xor ( n33275 , n33212 , n33267 );
not ( n33276 , n33275 );
xor ( n33277 , n33213 , n33266 );
not ( n33278 , n33277 );
xor ( n33279 , n33214 , n33265 );
not ( n33280 , n33279 );
xor ( n33281 , n33215 , n33264 );
not ( n33282 , n33281 );
xor ( n33283 , n33216 , n33263 );
not ( n33284 , n33283 );
xor ( n33285 , n33217 , n33262 );
not ( n33286 , n33285 );
xor ( n33287 , n33218 , n33261 );
not ( n33288 , n33287 );
xor ( n33289 , n33219 , n33260 );
not ( n33290 , n33289 );
xor ( n33291 , n33220 , n33259 );
not ( n33292 , n33291 );
xor ( n33293 , n33221 , n33258 );
not ( n33294 , n33293 );
xor ( n33295 , n33222 , n33257 );
not ( n33296 , n33295 );
xor ( n33297 , n33223 , n33256 );
not ( n33298 , n33297 );
xor ( n33299 , n33224 , n33255 );
not ( n33300 , n33299 );
xor ( n33301 , n33225 , n33254 );
not ( n33302 , n33301 );
xor ( n33303 , n33226 , n33253 );
not ( n33304 , n33303 );
xor ( n33305 , n33227 , n33252 );
not ( n33306 , n33305 );
xor ( n33307 , n33228 , n33251 );
not ( n33308 , n33307 );
xor ( n33309 , n33229 , n33250 );
not ( n33310 , n33309 );
xor ( n33311 , n33230 , n33249 );
not ( n33312 , n33311 );
xor ( n33313 , n33231 , n33248 );
not ( n33314 , n33313 );
xor ( n33315 , n33232 , n33247 );
not ( n33316 , n33315 );
xor ( n33317 , n33233 , n33246 );
not ( n33318 , n33317 );
xor ( n33319 , n33234 , n33245 );
not ( n33320 , n33319 );
xor ( n33321 , n33235 , n33244 );
not ( n33322 , n33321 );
xor ( n33323 , n33236 , n33243 );
not ( n33324 , n33323 );
xor ( n33325 , n33237 , n33242 );
not ( n33326 , n33325 );
xor ( n33327 , n33238 , n33241 );
not ( n33328 , n33327 );
xor ( n33329 , n33239 , n33240 );
not ( n33330 , n33329 );
not ( n33331 , n33240 );
not ( n33332 , n33331 );
buf ( n33333 , RI15b4a280_395);
not ( n33334 , n33333 );
and ( n33335 , n33332 , n33334 );
and ( n33336 , n33330 , n33335 );
and ( n33337 , n33328 , n33336 );
and ( n33338 , n33326 , n33337 );
and ( n33339 , n33324 , n33338 );
and ( n33340 , n33322 , n33339 );
and ( n33341 , n33320 , n33340 );
and ( n33342 , n33318 , n33341 );
and ( n33343 , n33316 , n33342 );
and ( n33344 , n33314 , n33343 );
and ( n33345 , n33312 , n33344 );
and ( n33346 , n33310 , n33345 );
and ( n33347 , n33308 , n33346 );
and ( n33348 , n33306 , n33347 );
and ( n33349 , n33304 , n33348 );
and ( n33350 , n33302 , n33349 );
and ( n33351 , n33300 , n33350 );
and ( n33352 , n33298 , n33351 );
and ( n33353 , n33296 , n33352 );
and ( n33354 , n33294 , n33353 );
and ( n33355 , n33292 , n33354 );
and ( n33356 , n33290 , n33355 );
and ( n33357 , n33288 , n33356 );
and ( n33358 , n33286 , n33357 );
and ( n33359 , n33284 , n33358 );
and ( n33360 , n33282 , n33359 );
and ( n33361 , n33280 , n33360 );
and ( n33362 , n33278 , n33361 );
and ( n33363 , n33276 , n33362 );
xor ( n33364 , n33274 , n33363 );
and ( n33365 , n33364 , n33270 );
or ( n33366 , n33273 , n33365 );
and ( n33367 , n33210 , n33366 );
and ( n33368 , n32600 , n32968 );
or ( n33369 , n33367 , n33368 );
nor ( n33370 , n32511 , n33207 , n32523 , n32526 );
and ( n33371 , n33369 , n33370 );
nor ( n33372 , n32512 , n32520 , n32523 , n32526 );
nor ( n33373 , n32512 , n33207 , n32523 , n32526 );
or ( n33374 , n33372 , n33373 );
and ( n33375 , n32512 , n33207 , n32523 , n32527 );
or ( n33376 , n33374 , n33375 );
and ( n33377 , n32512 , n32520 , n32523 , n32527 );
or ( n33378 , n33376 , n33377 );
and ( n33379 , n32511 , n32520 , n32523 , n32527 );
or ( n33380 , n33378 , n33379 );
nor ( n33381 , n32511 , n32520 , n32523 , n32527 );
or ( n33382 , n33380 , n33381 );
and ( n33383 , n32600 , n33382 );
or ( n33384 , C0 , n32529 , n33209 , n33371 , C0 , n33383 );
buf ( n33385 , n33384 );
buf ( n33386 , n33385 );
buf ( n33387 , n31655 );
buf ( n33388 , n30987 );
not ( n33389 , n31041 );
buf ( n33390 , n31041 );
buf ( n33391 , n31041 );
buf ( n33392 , n31041 );
buf ( n33393 , n31041 );
buf ( n33394 , n31041 );
buf ( n33395 , n31041 );
buf ( n33396 , n31041 );
buf ( n33397 , n31041 );
buf ( n33398 , n31041 );
buf ( n33399 , n31041 );
buf ( n33400 , n31041 );
buf ( n33401 , n31041 );
buf ( n33402 , n31041 );
buf ( n33403 , n31041 );
buf ( n33404 , n31041 );
buf ( n33405 , n31041 );
buf ( n33406 , n31041 );
buf ( n33407 , n31041 );
buf ( n33408 , n31041 );
buf ( n33409 , n31041 );
buf ( n33410 , n31041 );
buf ( n33411 , n31041 );
buf ( n33412 , n31041 );
buf ( n33413 , n31041 );
buf ( n33414 , n31041 );
xor ( n33415 , n31025 , n31026 );
or ( n33416 , n31075 , n33415 );
and ( n33417 , n31044 , n33416 );
or ( n33418 , n31046 , n31048 , n31041 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33417 );
and ( n33419 , n33389 , n33418 );
not ( n33420 , n33419 );
and ( n33421 , n33420 , n31570 );
buf ( n33422 , RI15b50928_614);
buf ( n33423 , RI15b508b0_613);
buf ( n33424 , RI15b50838_612);
buf ( n33425 , RI15b507c0_611);
buf ( n33426 , RI15b50748_610);
buf ( n33427 , RI15b506d0_609);
buf ( n33428 , RI15b50658_608);
buf ( n33429 , RI15b505e0_607);
buf ( n33430 , RI15b50568_606);
buf ( n33431 , RI15b504f0_605);
buf ( n33432 , RI15b50478_604);
buf ( n33433 , RI15b50400_603);
buf ( n33434 , RI15b50388_602);
buf ( n33435 , RI15b50310_601);
buf ( n33436 , RI15b50298_600);
buf ( n33437 , RI15b50220_599);
buf ( n33438 , RI15b501a8_598);
buf ( n33439 , RI15b50130_597);
buf ( n33440 , RI15b500b8_596);
buf ( n33441 , RI15b50040_595);
buf ( n33442 , RI15b4ffc8_594);
buf ( n33443 , RI15b4ff50_593);
and ( n33444 , n33442 , n33443 );
or ( n33445 , n33441 , n33444 );
and ( n33446 , n33440 , n33445 );
and ( n33447 , n33439 , n33446 );
and ( n33448 , n33438 , n33447 );
and ( n33449 , n33437 , n33448 );
and ( n33450 , n33436 , n33449 );
and ( n33451 , n33435 , n33450 );
and ( n33452 , n33434 , n33451 );
and ( n33453 , n33433 , n33452 );
and ( n33454 , n33432 , n33453 );
and ( n33455 , n33431 , n33454 );
and ( n33456 , n33430 , n33455 );
and ( n33457 , n33429 , n33456 );
and ( n33458 , n33428 , n33457 );
and ( n33459 , n33427 , n33458 );
and ( n33460 , n33426 , n33459 );
and ( n33461 , n33425 , n33460 );
and ( n33462 , n33424 , n33461 );
and ( n33463 , n33423 , n33462 );
xor ( n33464 , n33422 , n33463 );
xor ( n33465 , n33423 , n33462 );
xor ( n33466 , n33424 , n33461 );
xor ( n33467 , n33425 , n33460 );
xor ( n33468 , n33426 , n33459 );
xor ( n33469 , n33427 , n33458 );
xor ( n33470 , n33428 , n33457 );
xor ( n33471 , n33429 , n33456 );
xor ( n33472 , n33430 , n33455 );
xor ( n33473 , n33431 , n33454 );
xor ( n33474 , n33432 , n33453 );
xor ( n33475 , n33433 , n33452 );
xor ( n33476 , n33434 , n33451 );
xor ( n33477 , n33435 , n33450 );
xor ( n33478 , n33436 , n33449 );
not ( n33479 , n31026 );
not ( n33480 , n33479 );
buf ( n33481 , n33480 );
not ( n33482 , n33481 );
not ( n33483 , n33482 );
xor ( n33484 , n31022 , n31026 );
not ( n33485 , n33484 );
buf ( n33486 , n33485 );
buf ( n33487 , n33486 );
not ( n33488 , n33487 );
not ( n33489 , n33488 );
xor ( n33490 , n31018 , n31081 );
not ( n33491 , n33490 );
buf ( n33492 , n33491 );
buf ( n33493 , n33492 );
not ( n33494 , n33493 );
not ( n33495 , n33494 );
not ( n33496 , n31083 );
buf ( n33497 , n33496 );
buf ( n33498 , n33497 );
not ( n33499 , n33498 );
not ( n33500 , n33499 );
nor ( n33501 , n33483 , n33489 , n33495 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33502 , n31340 , n33501 );
nor ( n33503 , n33482 , n33489 , n33495 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33504 , n31342 , n33503 );
nor ( n33505 , n33483 , n33488 , n33495 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33506 , n31344 , n33505 );
nor ( n33507 , n33482 , n33488 , n33495 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33508 , n31346 , n33507 );
nor ( n33509 , n33483 , n33489 , n33494 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33510 , n31348 , n33509 );
nor ( n33511 , n33482 , n33489 , n33494 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33512 , n31350 , n33511 );
nor ( n33513 , n33483 , n33488 , n33494 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33514 , n31352 , n33513 );
nor ( n33515 , n33482 , n33488 , n33494 , n33500 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33516 , n31354 , n33515 );
nor ( n33517 , n33483 , n33489 , n33495 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33518 , n31356 , n33517 );
nor ( n33519 , n33482 , n33489 , n33495 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33520 , n31358 , n33519 );
nor ( n33521 , n33483 , n33488 , n33495 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33522 , n31360 , n33521 );
nor ( n33523 , n33482 , n33488 , n33495 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33524 , n31362 , n33523 );
nor ( n33525 , n33483 , n33489 , n33494 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33526 , n31364 , n33525 );
nor ( n33527 , n33482 , n33489 , n33494 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33528 , n31366 , n33527 );
nor ( n33529 , n33483 , n33488 , n33494 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33530 , n31368 , n33529 );
nor ( n33531 , n33482 , n33488 , n33494 , n33499 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n33532 , n31370 , n33531 );
or ( n33533 , n33502 , n33504 , n33506 , n33508 , n33510 , n33512 , n33514 , n33516 , n33518 , n33520 , n33522 , n33524 , n33526 , n33528 , n33530 , n33532 );
and ( n33534 , n33478 , n33533 );
xor ( n33535 , n33437 , n33448 );
and ( n33536 , n31307 , n33501 );
and ( n33537 , n31309 , n33503 );
and ( n33538 , n31311 , n33505 );
and ( n33539 , n31313 , n33507 );
and ( n33540 , n31315 , n33509 );
and ( n33541 , n31317 , n33511 );
and ( n33542 , n31319 , n33513 );
and ( n33543 , n31321 , n33515 );
and ( n33544 , n31323 , n33517 );
and ( n33545 , n31325 , n33519 );
and ( n33546 , n31327 , n33521 );
and ( n33547 , n31329 , n33523 );
and ( n33548 , n31331 , n33525 );
and ( n33549 , n31333 , n33527 );
and ( n33550 , n31335 , n33529 );
and ( n33551 , n31337 , n33531 );
or ( n33552 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 );
and ( n33553 , n33535 , n33552 );
xor ( n33554 , n33438 , n33447 );
and ( n33555 , n31274 , n33501 );
and ( n33556 , n31276 , n33503 );
and ( n33557 , n31278 , n33505 );
and ( n33558 , n31280 , n33507 );
and ( n33559 , n31282 , n33509 );
and ( n33560 , n31284 , n33511 );
and ( n33561 , n31286 , n33513 );
and ( n33562 , n31288 , n33515 );
and ( n33563 , n31290 , n33517 );
and ( n33564 , n31292 , n33519 );
and ( n33565 , n31294 , n33521 );
and ( n33566 , n31296 , n33523 );
and ( n33567 , n31298 , n33525 );
and ( n33568 , n31300 , n33527 );
and ( n33569 , n31302 , n33529 );
and ( n33570 , n31304 , n33531 );
or ( n33571 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 );
and ( n33572 , n33554 , n33571 );
xor ( n33573 , n33439 , n33446 );
and ( n33574 , n31240 , n33501 );
and ( n33575 , n31242 , n33503 );
and ( n33576 , n31244 , n33505 );
and ( n33577 , n31246 , n33507 );
and ( n33578 , n31248 , n33509 );
and ( n33579 , n31250 , n33511 );
and ( n33580 , n31252 , n33513 );
and ( n33581 , n31254 , n33515 );
and ( n33582 , n31256 , n33517 );
and ( n33583 , n31258 , n33519 );
and ( n33584 , n31260 , n33521 );
and ( n33585 , n31262 , n33523 );
and ( n33586 , n31264 , n33525 );
and ( n33587 , n31266 , n33527 );
and ( n33588 , n31268 , n33529 );
and ( n33589 , n31270 , n33531 );
or ( n33590 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 );
and ( n33591 , n33573 , n33590 );
xor ( n33592 , n33440 , n33445 );
and ( n33593 , n31206 , n33501 );
and ( n33594 , n31208 , n33503 );
and ( n33595 , n31210 , n33505 );
and ( n33596 , n31212 , n33507 );
and ( n33597 , n31214 , n33509 );
and ( n33598 , n31216 , n33511 );
and ( n33599 , n31218 , n33513 );
and ( n33600 , n31220 , n33515 );
and ( n33601 , n31222 , n33517 );
and ( n33602 , n31224 , n33519 );
and ( n33603 , n31226 , n33521 );
and ( n33604 , n31228 , n33523 );
and ( n33605 , n31230 , n33525 );
and ( n33606 , n31232 , n33527 );
and ( n33607 , n31234 , n33529 );
and ( n33608 , n31236 , n33531 );
or ( n33609 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 );
and ( n33610 , n33592 , n33609 );
xnor ( n33611 , n33441 , n33444 );
and ( n33612 , n31173 , n33501 );
and ( n33613 , n31175 , n33503 );
and ( n33614 , n31177 , n33505 );
and ( n33615 , n31179 , n33507 );
and ( n33616 , n31181 , n33509 );
and ( n33617 , n31183 , n33511 );
and ( n33618 , n31185 , n33513 );
and ( n33619 , n31187 , n33515 );
and ( n33620 , n31189 , n33517 );
and ( n33621 , n31191 , n33519 );
and ( n33622 , n31193 , n33521 );
and ( n33623 , n31195 , n33523 );
and ( n33624 , n31197 , n33525 );
and ( n33625 , n31199 , n33527 );
and ( n33626 , n31201 , n33529 );
and ( n33627 , n31203 , n33531 );
or ( n33628 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 );
and ( n33629 , n33611 , n33628 );
xor ( n33630 , n33442 , n33443 );
and ( n33631 , n31140 , n33501 );
and ( n33632 , n31142 , n33503 );
and ( n33633 , n31144 , n33505 );
and ( n33634 , n31146 , n33507 );
and ( n33635 , n31148 , n33509 );
and ( n33636 , n31150 , n33511 );
and ( n33637 , n31152 , n33513 );
and ( n33638 , n31154 , n33515 );
and ( n33639 , n31156 , n33517 );
and ( n33640 , n31158 , n33519 );
and ( n33641 , n31160 , n33521 );
and ( n33642 , n31162 , n33523 );
and ( n33643 , n31164 , n33525 );
and ( n33644 , n31166 , n33527 );
and ( n33645 , n31168 , n33529 );
and ( n33646 , n31170 , n33531 );
or ( n33647 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 );
and ( n33648 , n33630 , n33647 );
not ( n33649 , n33443 );
and ( n33650 , n31086 , n33501 );
and ( n33651 , n31090 , n33503 );
and ( n33652 , n31094 , n33505 );
and ( n33653 , n31098 , n33507 );
and ( n33654 , n31101 , n33509 );
and ( n33655 , n31105 , n33511 );
and ( n33656 , n31108 , n33513 );
and ( n33657 , n31111 , n33515 );
and ( n33658 , n31114 , n33517 );
and ( n33659 , n31117 , n33519 );
and ( n33660 , n31120 , n33521 );
and ( n33661 , n31123 , n33523 );
and ( n33662 , n31126 , n33525 );
and ( n33663 , n31129 , n33527 );
and ( n33664 , n31132 , n33529 );
and ( n33665 , n31135 , n33531 );
or ( n33666 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 );
and ( n33667 , n33649 , n33666 );
and ( n33668 , n33647 , n33667 );
and ( n33669 , n33630 , n33667 );
or ( n33670 , n33648 , n33668 , n33669 );
and ( n33671 , n33628 , n33670 );
and ( n33672 , n33611 , n33670 );
or ( n33673 , n33629 , n33671 , n33672 );
and ( n33674 , n33609 , n33673 );
and ( n33675 , n33592 , n33673 );
or ( n33676 , n33610 , n33674 , n33675 );
and ( n33677 , n33590 , n33676 );
and ( n33678 , n33573 , n33676 );
or ( n33679 , n33591 , n33677 , n33678 );
and ( n33680 , n33571 , n33679 );
and ( n33681 , n33554 , n33679 );
or ( n33682 , n33572 , n33680 , n33681 );
and ( n33683 , n33552 , n33682 );
and ( n33684 , n33535 , n33682 );
or ( n33685 , n33553 , n33683 , n33684 );
and ( n33686 , n33533 , n33685 );
and ( n33687 , n33478 , n33685 );
or ( n33688 , n33534 , n33686 , n33687 );
and ( n33689 , n33477 , n33688 );
and ( n33690 , n33476 , n33689 );
and ( n33691 , n33475 , n33690 );
and ( n33692 , n33474 , n33691 );
and ( n33693 , n33473 , n33692 );
and ( n33694 , n33472 , n33693 );
and ( n33695 , n33471 , n33694 );
and ( n33696 , n33470 , n33695 );
and ( n33697 , n33469 , n33696 );
and ( n33698 , n33468 , n33697 );
and ( n33699 , n33467 , n33698 );
and ( n33700 , n33466 , n33699 );
and ( n33701 , n33465 , n33700 );
xor ( n33702 , n33464 , n33701 );
and ( n33703 , n33702 , n33419 );
or ( n33704 , n33421 , n33703 );
and ( n33705 , n33704 , n31529 );
not ( n33706 , n31041 );
buf ( n33707 , n31041 );
buf ( n33708 , n31041 );
buf ( n33709 , n31041 );
buf ( n33710 , n31041 );
buf ( n33711 , n31041 );
buf ( n33712 , n31041 );
buf ( n33713 , n31041 );
buf ( n33714 , n31041 );
buf ( n33715 , n31041 );
buf ( n33716 , n31041 );
buf ( n33717 , n31041 );
buf ( n33718 , n31041 );
buf ( n33719 , n31041 );
buf ( n33720 , n31041 );
buf ( n33721 , n31041 );
buf ( n33722 , n31041 );
buf ( n33723 , n31041 );
buf ( n33724 , n31041 );
buf ( n33725 , n31041 );
buf ( n33726 , n31041 );
buf ( n33727 , n31041 );
buf ( n33728 , n31041 );
buf ( n33729 , n31041 );
buf ( n33730 , n31041 );
buf ( n33731 , n31041 );
and ( n33732 , n33415 , n31075 );
or ( n33733 , n31044 , n31046 , n31048 , n31041 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 );
and ( n33734 , n33706 , n33733 );
not ( n33735 , n33734 );
and ( n33736 , n33735 , n31570 );
not ( n33737 , n33533 );
and ( n33738 , n33441 , n33442 );
and ( n33739 , n33440 , n33738 );
and ( n33740 , n33439 , n33739 );
and ( n33741 , n33438 , n33740 );
and ( n33742 , n33437 , n33741 );
and ( n33743 , n33436 , n33742 );
and ( n33744 , n33435 , n33743 );
and ( n33745 , n33434 , n33744 );
and ( n33746 , n33433 , n33745 );
and ( n33747 , n33432 , n33746 );
and ( n33748 , n33431 , n33747 );
and ( n33749 , n33430 , n33748 );
and ( n33750 , n33429 , n33749 );
and ( n33751 , n33428 , n33750 );
and ( n33752 , n33427 , n33751 );
and ( n33753 , n33426 , n33752 );
and ( n33754 , n33425 , n33753 );
and ( n33755 , n33424 , n33754 );
and ( n33756 , n33423 , n33755 );
xor ( n33757 , n33422 , n33756 );
xor ( n33758 , n33423 , n33755 );
xor ( n33759 , n33424 , n33754 );
xor ( n33760 , n33425 , n33753 );
xor ( n33761 , n33426 , n33752 );
xor ( n33762 , n33427 , n33751 );
xor ( n33763 , n33428 , n33750 );
xor ( n33764 , n33429 , n33749 );
xor ( n33765 , n33430 , n33748 );
xor ( n33766 , n33431 , n33747 );
xor ( n33767 , n33432 , n33746 );
xor ( n33768 , n33433 , n33745 );
xor ( n33769 , n33434 , n33744 );
xor ( n33770 , n33435 , n33743 );
xor ( n33771 , n33436 , n33742 );
and ( n33772 , n33771 , n33533 );
xor ( n33773 , n33437 , n33741 );
and ( n33774 , n33773 , n33552 );
xor ( n33775 , n33438 , n33740 );
and ( n33776 , n33775 , n33571 );
xor ( n33777 , n33439 , n33739 );
and ( n33778 , n33777 , n33590 );
xor ( n33779 , n33440 , n33738 );
and ( n33780 , n33779 , n33609 );
xor ( n33781 , n33441 , n33442 );
and ( n33782 , n33781 , n33628 );
not ( n33783 , n33442 );
and ( n33784 , n33783 , n33647 );
and ( n33785 , n33443 , n33666 );
and ( n33786 , n33647 , n33785 );
and ( n33787 , n33783 , n33785 );
or ( n33788 , n33784 , n33786 , n33787 );
and ( n33789 , n33628 , n33788 );
and ( n33790 , n33781 , n33788 );
or ( n33791 , n33782 , n33789 , n33790 );
and ( n33792 , n33609 , n33791 );
and ( n33793 , n33779 , n33791 );
or ( n33794 , n33780 , n33792 , n33793 );
and ( n33795 , n33590 , n33794 );
and ( n33796 , n33777 , n33794 );
or ( n33797 , n33778 , n33795 , n33796 );
and ( n33798 , n33571 , n33797 );
and ( n33799 , n33775 , n33797 );
or ( n33800 , n33776 , n33798 , n33799 );
and ( n33801 , n33552 , n33800 );
and ( n33802 , n33773 , n33800 );
or ( n33803 , n33774 , n33801 , n33802 );
and ( n33804 , n33533 , n33803 );
and ( n33805 , n33771 , n33803 );
or ( n33806 , n33772 , n33804 , n33805 );
and ( n33807 , n33770 , n33806 );
and ( n33808 , n33769 , n33807 );
and ( n33809 , n33768 , n33808 );
and ( n33810 , n33767 , n33809 );
and ( n33811 , n33766 , n33810 );
and ( n33812 , n33765 , n33811 );
and ( n33813 , n33764 , n33812 );
and ( n33814 , n33763 , n33813 );
and ( n33815 , n33762 , n33814 );
and ( n33816 , n33761 , n33815 );
and ( n33817 , n33760 , n33816 );
and ( n33818 , n33759 , n33817 );
and ( n33819 , n33758 , n33818 );
xor ( n33820 , n33757 , n33819 );
and ( n33821 , n33737 , n33820 );
and ( n33822 , n33442 , n33443 );
and ( n33823 , n33441 , n33822 );
and ( n33824 , n33440 , n33823 );
and ( n33825 , n33439 , n33824 );
and ( n33826 , n33438 , n33825 );
and ( n33827 , n33437 , n33826 );
and ( n33828 , n33436 , n33827 );
and ( n33829 , n33435 , n33828 );
and ( n33830 , n33434 , n33829 );
and ( n33831 , n33433 , n33830 );
and ( n33832 , n33432 , n33831 );
and ( n33833 , n33431 , n33832 );
and ( n33834 , n33430 , n33833 );
and ( n33835 , n33429 , n33834 );
and ( n33836 , n33428 , n33835 );
and ( n33837 , n33427 , n33836 );
and ( n33838 , n33426 , n33837 );
and ( n33839 , n33425 , n33838 );
and ( n33840 , n33424 , n33839 );
and ( n33841 , n33423 , n33840 );
xor ( n33842 , n33422 , n33841 );
xor ( n33843 , n33423 , n33840 );
xor ( n33844 , n33424 , n33839 );
xor ( n33845 , n33425 , n33838 );
xor ( n33846 , n33426 , n33837 );
xor ( n33847 , n33427 , n33836 );
xor ( n33848 , n33428 , n33835 );
xor ( n33849 , n33429 , n33834 );
xor ( n33850 , n33430 , n33833 );
xor ( n33851 , n33431 , n33832 );
xor ( n33852 , n33432 , n33831 );
xor ( n33853 , n33433 , n33830 );
xor ( n33854 , n33434 , n33829 );
xor ( n33855 , n33435 , n33828 );
xor ( n33856 , n33436 , n33827 );
not ( n33857 , n33533 );
not ( n33858 , n33857 );
and ( n33859 , n33856 , n33858 );
xor ( n33860 , n33437 , n33826 );
not ( n33861 , n33552 );
not ( n33862 , n33861 );
and ( n33863 , n33860 , n33862 );
xor ( n33864 , n33438 , n33825 );
not ( n33865 , n33571 );
not ( n33866 , n33865 );
and ( n33867 , n33864 , n33866 );
xor ( n33868 , n33439 , n33824 );
not ( n33869 , n33590 );
not ( n33870 , n33869 );
and ( n33871 , n33868 , n33870 );
xor ( n33872 , n33440 , n33823 );
not ( n33873 , n33609 );
not ( n33874 , n33873 );
and ( n33875 , n33872 , n33874 );
xor ( n33876 , n33441 , n33822 );
not ( n33877 , n33628 );
not ( n33878 , n33877 );
and ( n33879 , n33876 , n33878 );
xor ( n33880 , n33442 , n33443 );
not ( n33881 , n33647 );
not ( n33882 , n33881 );
and ( n33883 , n33880 , n33882 );
not ( n33884 , n33443 );
not ( n33885 , n33666 );
not ( n33886 , n33885 );
or ( n33887 , n33884 , n33886 );
and ( n33888 , n33882 , n33887 );
and ( n33889 , n33880 , n33887 );
or ( n33890 , n33883 , n33888 , n33889 );
and ( n33891 , n33878 , n33890 );
and ( n33892 , n33876 , n33890 );
or ( n33893 , n33879 , n33891 , n33892 );
and ( n33894 , n33874 , n33893 );
and ( n33895 , n33872 , n33893 );
or ( n33896 , n33875 , n33894 , n33895 );
and ( n33897 , n33870 , n33896 );
and ( n33898 , n33868 , n33896 );
or ( n33899 , n33871 , n33897 , n33898 );
and ( n33900 , n33866 , n33899 );
and ( n33901 , n33864 , n33899 );
or ( n33902 , n33867 , n33900 , n33901 );
and ( n33903 , n33862 , n33902 );
and ( n33904 , n33860 , n33902 );
or ( n33905 , n33863 , n33903 , n33904 );
and ( n33906 , n33858 , n33905 );
and ( n33907 , n33856 , n33905 );
or ( n33908 , n33859 , n33906 , n33907 );
or ( n33909 , n33855 , n33908 );
or ( n33910 , n33854 , n33909 );
or ( n33911 , n33853 , n33910 );
or ( n33912 , n33852 , n33911 );
or ( n33913 , n33851 , n33912 );
or ( n33914 , n33850 , n33913 );
or ( n33915 , n33849 , n33914 );
or ( n33916 , n33848 , n33915 );
or ( n33917 , n33847 , n33916 );
or ( n33918 , n33846 , n33917 );
or ( n33919 , n33845 , n33918 );
or ( n33920 , n33844 , n33919 );
or ( n33921 , n33843 , n33920 );
xnor ( n33922 , n33842 , n33921 );
and ( n33923 , n33922 , n33533 );
or ( n33924 , n33821 , n33923 );
and ( n33925 , n33924 , n33734 );
or ( n33926 , n33736 , n33925 );
and ( n33927 , n33926 , n31527 );
or ( n33928 , n31525 , n31531 );
or ( n33929 , n33928 , n31534 );
or ( n33930 , n33929 , n31536 );
or ( n33931 , n33930 , n31538 );
or ( n33932 , n33931 , n31521 );
or ( n33933 , n33932 , n31468 );
or ( n33934 , n33933 , n31408 );
or ( n33935 , n33934 , n31373 );
or ( n33936 , n33935 , n31540 );
or ( n33937 , n33936 , n31542 );
or ( n33938 , n33937 , n31544 );
or ( n33939 , n33938 , n31546 );
or ( n33940 , n33939 , n31548 );
or ( n33941 , n33940 , n31550 );
or ( n33942 , n33941 , n31552 );
and ( n33943 , n31570 , n33942 );
or ( n33944 , n33705 , n33927 , n33943 );
and ( n33945 , n33944 , n31557 );
xor ( n33946 , n31570 , n31608 );
and ( n33947 , n33946 , n31643 );
not ( n33948 , n31452 );
and ( n33949 , n33948 , n33946 );
and ( n33950 , n30989 , n31588 );
and ( n33951 , n31587 , n33950 );
and ( n33952 , n31586 , n33951 );
and ( n33953 , n31585 , n33952 );
and ( n33954 , n31584 , n33953 );
and ( n33955 , n31583 , n33954 );
and ( n33956 , n31582 , n33955 );
and ( n33957 , n31581 , n33956 );
and ( n33958 , n31580 , n33957 );
and ( n33959 , n31579 , n33958 );
and ( n33960 , n31578 , n33959 );
and ( n33961 , n31577 , n33960 );
and ( n33962 , n31576 , n33961 );
and ( n33963 , n31575 , n33962 );
and ( n33964 , n31574 , n33963 );
and ( n33965 , n31573 , n33964 );
and ( n33966 , n31572 , n33965 );
and ( n33967 , n31571 , n33966 );
xor ( n33968 , n31570 , n33967 );
and ( n33969 , n33968 , n31452 );
or ( n33970 , n33949 , n33969 );
and ( n33971 , n33970 , n31638 );
buf ( n33972 , RI15b57fc0_867);
nor ( n33973 , n30990 , n30999 , n31002 , n31005 );
and ( n33974 , n33972 , n33973 );
or ( n33975 , n31642 , n31645 );
or ( n33976 , n33975 , n31647 );
or ( n33977 , n33976 , n31649 );
or ( n33978 , n33977 , n31007 );
and ( n33979 , n31570 , n33978 );
or ( n33980 , C0 , n33945 , n33947 , n33971 , n33974 , n33979 );
buf ( n33981 , n33980 );
buf ( n33982 , n33981 );
buf ( n33983 , n30987 );
and ( n33984 , n31574 , n31007 );
not ( n33985 , n31077 );
buf ( n33986 , RI15b57de0_863);
and ( n33987 , n33985 , n33986 );
buf ( n33988 , n33987 );
and ( n33989 , n33988 , n31373 );
not ( n33990 , n31402 );
and ( n33991 , n33990 , n33986 );
buf ( n33992 , n33991 );
and ( n33993 , n33992 , n31408 );
not ( n33994 , n31437 );
and ( n33995 , n33994 , n33986 );
not ( n33996 , n31455 );
buf ( n33997 , RI15b55fe0_799);
and ( n33998 , n33996 , n33997 );
buf ( n33999 , RI15b57d68_862);
buf ( n34000 , RI15b57cf0_861);
buf ( n34001 , RI15b57c78_860);
buf ( n34002 , RI15b57c00_859);
buf ( n34003 , RI15b57b88_858);
buf ( n34004 , RI15b57b10_857);
buf ( n34005 , RI15b57a98_856);
buf ( n34006 , RI15b57a20_855);
buf ( n34007 , RI15b579a8_854);
buf ( n34008 , RI15b57930_853);
buf ( n34009 , RI15b578b8_852);
buf ( n34010 , RI15b57840_851);
buf ( n34011 , RI15b577c8_850);
and ( n34012 , n31079 , n31461 );
and ( n34013 , n34011 , n34012 );
and ( n34014 , n34010 , n34013 );
and ( n34015 , n34009 , n34014 );
and ( n34016 , n34008 , n34015 );
and ( n34017 , n34007 , n34016 );
and ( n34018 , n34006 , n34017 );
and ( n34019 , n34005 , n34018 );
and ( n34020 , n34004 , n34019 );
and ( n34021 , n34003 , n34020 );
and ( n34022 , n34002 , n34021 );
and ( n34023 , n34001 , n34022 );
and ( n34024 , n34000 , n34023 );
and ( n34025 , n33999 , n34024 );
xor ( n34026 , n33986 , n34025 );
and ( n34027 , n34026 , n31455 );
or ( n34028 , n33998 , n34027 );
and ( n34029 , n34028 , n31437 );
or ( n34030 , n33995 , n34029 );
and ( n34031 , n34030 , n31468 );
not ( n34032 , n31497 );
and ( n34033 , n34032 , n33986 );
not ( n34034 , n31454 );
not ( n34035 , n31501 );
and ( n34036 , n34035 , n33997 );
not ( n34037 , n33997 );
buf ( n34038 , RI15b55f68_798);
not ( n34039 , n34038 );
buf ( n34040 , RI15b55ef0_797);
not ( n34041 , n34040 );
buf ( n34042 , RI15b55e78_796);
not ( n34043 , n34042 );
buf ( n34044 , RI15b55e00_795);
not ( n34045 , n34044 );
buf ( n34046 , RI15b55d88_794);
not ( n34047 , n34046 );
buf ( n34048 , RI15b55d10_793);
not ( n34049 , n34048 );
buf ( n34050 , RI15b55c98_792);
not ( n34051 , n34050 );
buf ( n34052 , RI15b55c20_791);
not ( n34053 , n34052 );
buf ( n34054 , RI15b55ba8_790);
not ( n34055 , n34054 );
buf ( n34056 , RI15b55b30_789);
not ( n34057 , n34056 );
buf ( n34058 , RI15b55ab8_788);
not ( n34059 , n34058 );
buf ( n34060 , RI15b55a40_787);
not ( n34061 , n34060 );
buf ( n34062 , RI15b559c8_786);
not ( n34063 , n34062 );
and ( n34064 , n31504 , n31512 );
and ( n34065 , n34063 , n34064 );
and ( n34066 , n34061 , n34065 );
and ( n34067 , n34059 , n34066 );
and ( n34068 , n34057 , n34067 );
and ( n34069 , n34055 , n34068 );
and ( n34070 , n34053 , n34069 );
and ( n34071 , n34051 , n34070 );
and ( n34072 , n34049 , n34071 );
and ( n34073 , n34047 , n34072 );
and ( n34074 , n34045 , n34073 );
and ( n34075 , n34043 , n34074 );
and ( n34076 , n34041 , n34075 );
and ( n34077 , n34039 , n34076 );
xor ( n34078 , n34037 , n34077 );
and ( n34079 , n34078 , n31501 );
or ( n34080 , n34036 , n34079 );
and ( n34081 , n34034 , n34080 );
and ( n34082 , n34026 , n31454 );
or ( n34083 , n34081 , n34082 );
and ( n34084 , n34083 , n31497 );
or ( n34085 , n34033 , n34084 );
and ( n34086 , n34085 , n31521 );
and ( n34087 , n33986 , n31553 );
or ( n34088 , n33989 , n33993 , n34031 , n34086 , n34087 );
and ( n34089 , n34088 , n31557 );
not ( n34090 , n31452 );
not ( n34091 , n31619 );
xor ( n34092 , n31574 , n31604 );
and ( n34093 , n34091 , n34092 );
not ( n34094 , n34092 );
xor ( n34095 , n31575 , n31603 );
not ( n34096 , n34095 );
xor ( n34097 , n31576 , n31602 );
not ( n34098 , n34097 );
xor ( n34099 , n31577 , n31601 );
not ( n34100 , n34099 );
xor ( n34101 , n31578 , n31600 );
not ( n34102 , n34101 );
xor ( n34103 , n31579 , n31599 );
not ( n34104 , n34103 );
xor ( n34105 , n31580 , n31598 );
not ( n34106 , n34105 );
xor ( n34107 , n31581 , n31597 );
not ( n34108 , n34107 );
xor ( n34109 , n31582 , n31596 );
not ( n34110 , n34109 );
xor ( n34111 , n31583 , n31595 );
not ( n34112 , n34111 );
xor ( n34113 , n31584 , n31594 );
not ( n34114 , n34113 );
xor ( n34115 , n31585 , n31593 );
not ( n34116 , n34115 );
xor ( n34117 , n31586 , n31592 );
not ( n34118 , n34117 );
xor ( n34119 , n31587 , n31591 );
not ( n34120 , n34119 );
and ( n34121 , n31623 , n31631 );
and ( n34122 , n34120 , n34121 );
and ( n34123 , n34118 , n34122 );
and ( n34124 , n34116 , n34123 );
and ( n34125 , n34114 , n34124 );
and ( n34126 , n34112 , n34125 );
and ( n34127 , n34110 , n34126 );
and ( n34128 , n34108 , n34127 );
and ( n34129 , n34106 , n34128 );
and ( n34130 , n34104 , n34129 );
and ( n34131 , n34102 , n34130 );
and ( n34132 , n34100 , n34131 );
and ( n34133 , n34098 , n34132 );
and ( n34134 , n34096 , n34133 );
xor ( n34135 , n34094 , n34134 );
and ( n34136 , n34135 , n31619 );
or ( n34137 , n34093 , n34136 );
and ( n34138 , n34090 , n34137 );
and ( n34139 , n33986 , n31452 );
or ( n34140 , n34138 , n34139 );
and ( n34141 , n34140 , n31638 );
buf ( n34142 , n33973 );
and ( n34143 , n33986 , n31650 );
or ( n34144 , C0 , n33984 , n34089 , n34141 , n34142 , n34143 );
buf ( n34145 , n34144 );
buf ( n34146 , n34145 );
buf ( n34147 , n31655 );
buf ( n34148 , n31655 );
buf ( n34149 , n30987 );
not ( n34150 , n32531 );
not ( n34151 , n34150 );
and ( n34152 , n34151 , n32783 );
not ( n34153 , n32542 );
nor ( n34154 , n32546 , n34153 , n32538 , n32534 , n32530 );
not ( n34155 , n34154 );
and ( n34156 , n34155 , n32783 );
and ( n34157 , n32789 , n34154 );
or ( n34158 , n34156 , n34157 );
and ( n34159 , n34158 , n34150 );
or ( n34160 , n34152 , n34159 );
and ( n34161 , n34160 , n33381 );
not ( n34162 , n32546 );
not ( n34163 , n34162 );
buf ( n34164 , n34163 );
not ( n34165 , n34164 );
xor ( n34166 , n32542 , n32546 );
not ( n34167 , n34166 );
buf ( n34168 , n34167 );
buf ( n34169 , n34168 );
not ( n34170 , n34169 );
not ( n34171 , n34170 );
and ( n34172 , n32542 , n32546 );
xor ( n34173 , n32538 , n34172 );
not ( n34174 , n34173 );
buf ( n34175 , n34174 );
buf ( n34176 , n34175 );
not ( n34177 , n34176 );
and ( n34178 , n32538 , n34172 );
xor ( n34179 , n32534 , n34178 );
not ( n34180 , n34179 );
buf ( n34181 , n34180 );
buf ( n34182 , n34181 );
not ( n34183 , n34182 );
nor ( n34184 , n34165 , n34171 , n34177 , n34183 , C0 );
not ( n34185 , n34184 );
not ( n34186 , n34154 );
and ( n34187 , n34186 , n32783 );
buf ( n34188 , RI15b65850_1329);
buf ( n34189 , n34188 );
not ( n34190 , n34189 );
buf ( n34191 , n34190 );
not ( n34192 , n34191 );
buf ( n34193 , RI15b666d8_1360);
not ( n34194 , n34193 );
buf ( n34195 , RI15b658c8_1330);
and ( n34196 , n34194 , n34195 );
not ( n34197 , n34195 );
not ( n34198 , n34188 );
xor ( n34199 , n34197 , n34198 );
and ( n34200 , n34199 , n34193 );
or ( n34201 , n34196 , n34200 );
not ( n34202 , n34201 );
buf ( n34203 , n34202 );
buf ( n34204 , n34203 );
not ( n34205 , n34204 );
or ( n34206 , n34192 , n34205 );
not ( n34207 , n34193 );
buf ( n34208 , RI15b65940_1331);
and ( n34209 , n34207 , n34208 );
not ( n34210 , n34208 );
and ( n34211 , n34197 , n34198 );
xor ( n34212 , n34210 , n34211 );
and ( n34213 , n34212 , n34193 );
or ( n34214 , n34209 , n34213 );
not ( n34215 , n34214 );
buf ( n34216 , n34215 );
buf ( n34217 , n34216 );
not ( n34218 , n34217 );
or ( n34219 , n34206 , n34218 );
not ( n34220 , n34193 );
buf ( n34221 , RI15b659b8_1332);
and ( n34222 , n34220 , n34221 );
not ( n34223 , n34221 );
and ( n34224 , n34210 , n34211 );
xor ( n34225 , n34223 , n34224 );
and ( n34226 , n34225 , n34193 );
or ( n34227 , n34222 , n34226 );
not ( n34228 , n34227 );
buf ( n34229 , n34228 );
buf ( n34230 , n34229 );
not ( n34231 , n34230 );
or ( n34232 , n34219 , n34231 );
not ( n34233 , n34193 );
buf ( n34234 , RI15b65a30_1333);
and ( n34235 , n34233 , n34234 );
not ( n34236 , n34234 );
and ( n34237 , n34223 , n34224 );
xor ( n34238 , n34236 , n34237 );
and ( n34239 , n34238 , n34193 );
or ( n34240 , n34235 , n34239 );
not ( n34241 , n34240 );
buf ( n34242 , n34241 );
buf ( n34243 , n34242 );
not ( n34244 , n34243 );
or ( n34245 , n34232 , n34244 );
not ( n34246 , n34193 );
buf ( n34247 , RI15b65aa8_1334);
and ( n34248 , n34246 , n34247 );
not ( n34249 , n34247 );
and ( n34250 , n34236 , n34237 );
xor ( n34251 , n34249 , n34250 );
and ( n34252 , n34251 , n34193 );
or ( n34253 , n34248 , n34252 );
not ( n34254 , n34253 );
buf ( n34255 , n34254 );
buf ( n34256 , n34255 );
not ( n34257 , n34256 );
or ( n34258 , n34245 , n34257 );
not ( n34259 , n34193 );
buf ( n34260 , RI15b65b20_1335);
and ( n34261 , n34259 , n34260 );
not ( n34262 , n34260 );
and ( n34263 , n34249 , n34250 );
xor ( n34264 , n34262 , n34263 );
and ( n34265 , n34264 , n34193 );
or ( n34266 , n34261 , n34265 );
not ( n34267 , n34266 );
buf ( n34268 , n34267 );
buf ( n34269 , n34268 );
not ( n34270 , n34269 );
or ( n34271 , n34258 , n34270 );
not ( n34272 , n34193 );
buf ( n34273 , RI15b65b98_1336);
and ( n34274 , n34272 , n34273 );
not ( n34275 , n34273 );
and ( n34276 , n34262 , n34263 );
xor ( n34277 , n34275 , n34276 );
and ( n34278 , n34277 , n34193 );
or ( n34279 , n34274 , n34278 );
not ( n34280 , n34279 );
buf ( n34281 , n34280 );
buf ( n34282 , n34281 );
not ( n34283 , n34282 );
or ( n34284 , n34271 , n34283 );
buf ( n34285 , n34284 );
buf ( n34286 , n34285 );
and ( n34287 , n34286 , n34193 );
not ( n34288 , n34287 );
and ( n34289 , n34288 , n34244 );
xor ( n34290 , n34244 , n34193 );
xor ( n34291 , n34231 , n34193 );
xor ( n34292 , n34218 , n34193 );
xor ( n34293 , n34205 , n34193 );
xor ( n34294 , n34192 , n34193 );
and ( n34295 , n34294 , n34193 );
and ( n34296 , n34293 , n34295 );
and ( n34297 , n34292 , n34296 );
and ( n34298 , n34291 , n34297 );
xor ( n34299 , n34290 , n34298 );
and ( n34300 , n34299 , n34287 );
or ( n34301 , n34289 , n34300 );
and ( n34302 , n34301 , n34154 );
or ( n34303 , n34187 , n34302 );
and ( n34304 , n34185 , n34303 );
and ( n34305 , n34301 , n34184 );
or ( n34306 , n34304 , n34305 );
and ( n34307 , n34306 , n33375 );
not ( n34308 , n32968 );
not ( n34309 , n34184 );
not ( n34310 , n34154 );
and ( n34311 , n34310 , n32783 );
and ( n34312 , n34301 , n34154 );
or ( n34313 , n34311 , n34312 );
and ( n34314 , n34309 , n34313 );
and ( n34315 , n34301 , n34184 );
or ( n34316 , n34314 , n34315 );
and ( n34317 , n34308 , n34316 );
not ( n34318 , n34165 );
not ( n34319 , n34318 );
buf ( n34320 , n34319 );
not ( n34321 , n34320 );
not ( n34322 , n34321 );
not ( n34323 , n34322 );
buf ( n34324 , n34323 );
not ( n34325 , n34324 );
xor ( n34326 , n34170 , n34165 );
not ( n34327 , n34326 );
buf ( n34328 , n34327 );
not ( n34329 , n34328 );
xor ( n34330 , n34329 , n34321 );
not ( n34331 , n34330 );
buf ( n34332 , n34331 );
not ( n34333 , n34332 );
not ( n34334 , n34333 );
and ( n34335 , n34170 , n34165 );
xor ( n34336 , n34177 , n34335 );
not ( n34337 , n34336 );
buf ( n34338 , n34337 );
not ( n34339 , n34338 );
and ( n34340 , n34329 , n34321 );
xor ( n34341 , n34339 , n34340 );
not ( n34342 , n34341 );
buf ( n34343 , n34342 );
not ( n34344 , n34343 );
and ( n34345 , n34177 , n34335 );
xor ( n34346 , n34183 , n34345 );
not ( n34347 , n34346 );
buf ( n34348 , n34347 );
not ( n34349 , n34348 );
and ( n34350 , n34339 , n34340 );
xor ( n34351 , n34349 , n34350 );
not ( n34352 , n34351 );
buf ( n34353 , n34352 );
not ( n34354 , n34353 );
nor ( n34355 , n34325 , n34334 , n34344 , n34354 , C0 );
not ( n34356 , n34355 );
not ( n34357 , n34329 );
nor ( n34358 , n34321 , n34357 , n34339 , n34349 , C0 );
not ( n34359 , n34358 );
and ( n34360 , n34359 , n34316 );
not ( n34361 , n34193 );
buf ( n34362 , RI15b65fd0_1345);
and ( n34363 , n34361 , n34362 );
not ( n34364 , n34362 );
buf ( n34365 , RI15b65f58_1344);
not ( n34366 , n34365 );
buf ( n34367 , RI15b65ee0_1343);
not ( n34368 , n34367 );
buf ( n34369 , RI15b65e68_1342);
not ( n34370 , n34369 );
buf ( n34371 , RI15b65df0_1341);
not ( n34372 , n34371 );
buf ( n34373 , RI15b65d78_1340);
not ( n34374 , n34373 );
buf ( n34375 , RI15b65d00_1339);
not ( n34376 , n34375 );
buf ( n34377 , RI15b65c88_1338);
not ( n34378 , n34377 );
buf ( n34379 , RI15b65c10_1337);
not ( n34380 , n34379 );
not ( n34381 , n34273 );
not ( n34382 , n34260 );
not ( n34383 , n34247 );
not ( n34384 , n34234 );
not ( n34385 , n34221 );
not ( n34386 , n34208 );
not ( n34387 , n34195 );
not ( n34388 , n34188 );
and ( n34389 , n34387 , n34388 );
and ( n34390 , n34386 , n34389 );
and ( n34391 , n34385 , n34390 );
and ( n34392 , n34384 , n34391 );
and ( n34393 , n34383 , n34392 );
and ( n34394 , n34382 , n34393 );
and ( n34395 , n34381 , n34394 );
and ( n34396 , n34380 , n34395 );
and ( n34397 , n34378 , n34396 );
and ( n34398 , n34376 , n34397 );
and ( n34399 , n34374 , n34398 );
and ( n34400 , n34372 , n34399 );
and ( n34401 , n34370 , n34400 );
and ( n34402 , n34368 , n34401 );
and ( n34403 , n34366 , n34402 );
xor ( n34404 , n34364 , n34403 );
and ( n34405 , n34404 , n34193 );
or ( n34406 , n34363 , n34405 );
not ( n34407 , n34406 );
buf ( n34408 , n34407 );
buf ( n34409 , n34408 );
not ( n34410 , n34409 );
buf ( n34411 , n34410 );
buf ( n34412 , n34411 );
not ( n34413 , n34412 );
buf ( n34414 , n34413 );
not ( n34415 , n34414 );
not ( n34416 , n34193 );
buf ( n34417 , RI15b66660_1359);
not ( n34418 , n34417 );
buf ( n34419 , RI15b665e8_1358);
not ( n34420 , n34419 );
buf ( n34421 , RI15b66570_1357);
not ( n34422 , n34421 );
buf ( n34423 , RI15b664f8_1356);
not ( n34424 , n34423 );
buf ( n34425 , RI15b66480_1355);
not ( n34426 , n34425 );
buf ( n34427 , RI15b66408_1354);
not ( n34428 , n34427 );
buf ( n34429 , RI15b66390_1353);
not ( n34430 , n34429 );
buf ( n34431 , RI15b66318_1352);
not ( n34432 , n34431 );
buf ( n34433 , RI15b662a0_1351);
not ( n34434 , n34433 );
buf ( n34435 , RI15b66228_1350);
not ( n34436 , n34435 );
buf ( n34437 , RI15b661b0_1349);
not ( n34438 , n34437 );
buf ( n34439 , RI15b66138_1348);
not ( n34440 , n34439 );
buf ( n34441 , RI15b660c0_1347);
not ( n34442 , n34441 );
buf ( n34443 , RI15b66048_1346);
not ( n34444 , n34443 );
and ( n34445 , n34364 , n34403 );
and ( n34446 , n34444 , n34445 );
and ( n34447 , n34442 , n34446 );
and ( n34448 , n34440 , n34447 );
and ( n34449 , n34438 , n34448 );
and ( n34450 , n34436 , n34449 );
and ( n34451 , n34434 , n34450 );
and ( n34452 , n34432 , n34451 );
and ( n34453 , n34430 , n34452 );
and ( n34454 , n34428 , n34453 );
and ( n34455 , n34426 , n34454 );
and ( n34456 , n34424 , n34455 );
and ( n34457 , n34422 , n34456 );
and ( n34458 , n34420 , n34457 );
and ( n34459 , n34418 , n34458 );
xor ( n34460 , n34416 , n34459 );
buf ( n34461 , n34193 );
and ( n34462 , n34460 , n34461 );
buf ( n34463 , n34462 );
not ( n34464 , n34463 );
not ( n34465 , n34464 );
not ( n34466 , n34465 );
not ( n34467 , n34193 );
and ( n34468 , n34467 , n34417 );
xor ( n34469 , n34418 , n34458 );
and ( n34470 , n34469 , n34193 );
or ( n34471 , n34468 , n34470 );
not ( n34472 , n34471 );
buf ( n34473 , n34472 );
buf ( n34474 , n34473 );
not ( n34475 , n34474 );
not ( n34476 , n34475 );
not ( n34477 , n34193 );
and ( n34478 , n34477 , n34419 );
xor ( n34479 , n34420 , n34457 );
and ( n34480 , n34479 , n34193 );
or ( n34481 , n34478 , n34480 );
not ( n34482 , n34481 );
buf ( n34483 , n34482 );
buf ( n34484 , n34483 );
not ( n34485 , n34484 );
not ( n34486 , n34485 );
not ( n34487 , n34193 );
and ( n34488 , n34487 , n34421 );
xor ( n34489 , n34422 , n34456 );
and ( n34490 , n34489 , n34193 );
or ( n34491 , n34488 , n34490 );
not ( n34492 , n34491 );
buf ( n34493 , n34492 );
buf ( n34494 , n34493 );
not ( n34495 , n34494 );
not ( n34496 , n34495 );
not ( n34497 , n34193 );
and ( n34498 , n34497 , n34423 );
xor ( n34499 , n34424 , n34455 );
and ( n34500 , n34499 , n34193 );
or ( n34501 , n34498 , n34500 );
not ( n34502 , n34501 );
buf ( n34503 , n34502 );
buf ( n34504 , n34503 );
not ( n34505 , n34504 );
not ( n34506 , n34505 );
not ( n34507 , n34193 );
and ( n34508 , n34507 , n34425 );
xor ( n34509 , n34426 , n34454 );
and ( n34510 , n34509 , n34193 );
or ( n34511 , n34508 , n34510 );
not ( n34512 , n34511 );
buf ( n34513 , n34512 );
buf ( n34514 , n34513 );
not ( n34515 , n34514 );
not ( n34516 , n34515 );
not ( n34517 , n34193 );
and ( n34518 , n34517 , n34427 );
xor ( n34519 , n34428 , n34453 );
and ( n34520 , n34519 , n34193 );
or ( n34521 , n34518 , n34520 );
not ( n34522 , n34521 );
buf ( n34523 , n34522 );
buf ( n34524 , n34523 );
not ( n34525 , n34524 );
not ( n34526 , n34525 );
not ( n34527 , n34193 );
and ( n34528 , n34527 , n34429 );
xor ( n34529 , n34430 , n34452 );
and ( n34530 , n34529 , n34193 );
or ( n34531 , n34528 , n34530 );
not ( n34532 , n34531 );
buf ( n34533 , n34532 );
buf ( n34534 , n34533 );
not ( n34535 , n34534 );
not ( n34536 , n34535 );
not ( n34537 , n34193 );
and ( n34538 , n34537 , n34431 );
xor ( n34539 , n34432 , n34451 );
and ( n34540 , n34539 , n34193 );
or ( n34541 , n34538 , n34540 );
not ( n34542 , n34541 );
buf ( n34543 , n34542 );
buf ( n34544 , n34543 );
not ( n34545 , n34544 );
not ( n34546 , n34545 );
not ( n34547 , n34193 );
and ( n34548 , n34547 , n34433 );
xor ( n34549 , n34434 , n34450 );
and ( n34550 , n34549 , n34193 );
or ( n34551 , n34548 , n34550 );
not ( n34552 , n34551 );
buf ( n34553 , n34552 );
buf ( n34554 , n34553 );
not ( n34555 , n34554 );
not ( n34556 , n34555 );
not ( n34557 , n34193 );
and ( n34558 , n34557 , n34435 );
xor ( n34559 , n34436 , n34449 );
and ( n34560 , n34559 , n34193 );
or ( n34561 , n34558 , n34560 );
not ( n34562 , n34561 );
buf ( n34563 , n34562 );
buf ( n34564 , n34563 );
not ( n34565 , n34564 );
not ( n34566 , n34565 );
not ( n34567 , n34193 );
and ( n34568 , n34567 , n34437 );
xor ( n34569 , n34438 , n34448 );
and ( n34570 , n34569 , n34193 );
or ( n34571 , n34568 , n34570 );
not ( n34572 , n34571 );
buf ( n34573 , n34572 );
buf ( n34574 , n34573 );
not ( n34575 , n34574 );
not ( n34576 , n34575 );
not ( n34577 , n34193 );
and ( n34578 , n34577 , n34439 );
xor ( n34579 , n34440 , n34447 );
and ( n34580 , n34579 , n34193 );
or ( n34581 , n34578 , n34580 );
not ( n34582 , n34581 );
buf ( n34583 , n34582 );
buf ( n34584 , n34583 );
not ( n34585 , n34584 );
not ( n34586 , n34585 );
not ( n34587 , n34193 );
and ( n34588 , n34587 , n34441 );
xor ( n34589 , n34442 , n34446 );
and ( n34590 , n34589 , n34193 );
or ( n34591 , n34588 , n34590 );
not ( n34592 , n34591 );
buf ( n34593 , n34592 );
buf ( n34594 , n34593 );
not ( n34595 , n34594 );
not ( n34596 , n34595 );
not ( n34597 , n34193 );
and ( n34598 , n34597 , n34443 );
xor ( n34599 , n34444 , n34445 );
and ( n34600 , n34599 , n34193 );
or ( n34601 , n34598 , n34600 );
not ( n34602 , n34601 );
buf ( n34603 , n34602 );
buf ( n34604 , n34603 );
not ( n34605 , n34604 );
not ( n34606 , n34605 );
not ( n34607 , n34410 );
and ( n34608 , n34606 , n34607 );
and ( n34609 , n34596 , n34608 );
and ( n34610 , n34586 , n34609 );
and ( n34611 , n34576 , n34610 );
and ( n34612 , n34566 , n34611 );
and ( n34613 , n34556 , n34612 );
and ( n34614 , n34546 , n34613 );
and ( n34615 , n34536 , n34614 );
and ( n34616 , n34526 , n34615 );
and ( n34617 , n34516 , n34616 );
and ( n34618 , n34506 , n34617 );
and ( n34619 , n34496 , n34618 );
and ( n34620 , n34486 , n34619 );
and ( n34621 , n34476 , n34620 );
and ( n34622 , n34466 , n34621 );
not ( n34623 , n34622 );
and ( n34624 , n34623 , n34193 );
buf ( n34625 , n34624 );
not ( n34626 , n34625 );
not ( n34627 , n34193 );
and ( n34628 , n34627 , n34605 );
xor ( n34629 , n34606 , n34607 );
and ( n34630 , n34629 , n34193 );
or ( n34631 , n34628 , n34630 );
and ( n34632 , n34626 , n34631 );
not ( n34633 , n34631 );
not ( n34634 , n34411 );
xor ( n34635 , n34633 , n34634 );
and ( n34636 , n34635 , n34625 );
or ( n34637 , n34632 , n34636 );
not ( n34638 , n34637 );
buf ( n34639 , n34638 );
buf ( n34640 , n34639 );
not ( n34641 , n34640 );
or ( n34642 , n34415 , n34641 );
not ( n34643 , n34625 );
not ( n34644 , n34193 );
and ( n34645 , n34644 , n34595 );
xor ( n34646 , n34596 , n34608 );
and ( n34647 , n34646 , n34193 );
or ( n34648 , n34645 , n34647 );
and ( n34649 , n34643 , n34648 );
not ( n34650 , n34648 );
and ( n34651 , n34633 , n34634 );
xor ( n34652 , n34650 , n34651 );
and ( n34653 , n34652 , n34625 );
or ( n34654 , n34649 , n34653 );
not ( n34655 , n34654 );
buf ( n34656 , n34655 );
buf ( n34657 , n34656 );
not ( n34658 , n34657 );
or ( n34659 , n34642 , n34658 );
not ( n34660 , n34625 );
not ( n34661 , n34193 );
and ( n34662 , n34661 , n34585 );
xor ( n34663 , n34586 , n34609 );
and ( n34664 , n34663 , n34193 );
or ( n34665 , n34662 , n34664 );
and ( n34666 , n34660 , n34665 );
not ( n34667 , n34665 );
and ( n34668 , n34650 , n34651 );
xor ( n34669 , n34667 , n34668 );
and ( n34670 , n34669 , n34625 );
or ( n34671 , n34666 , n34670 );
not ( n34672 , n34671 );
buf ( n34673 , n34672 );
buf ( n34674 , n34673 );
not ( n34675 , n34674 );
or ( n34676 , n34659 , n34675 );
not ( n34677 , n34625 );
not ( n34678 , n34193 );
and ( n34679 , n34678 , n34575 );
xor ( n34680 , n34576 , n34610 );
and ( n34681 , n34680 , n34193 );
or ( n34682 , n34679 , n34681 );
and ( n34683 , n34677 , n34682 );
not ( n34684 , n34682 );
and ( n34685 , n34667 , n34668 );
xor ( n34686 , n34684 , n34685 );
and ( n34687 , n34686 , n34625 );
or ( n34688 , n34683 , n34687 );
not ( n34689 , n34688 );
buf ( n34690 , n34689 );
buf ( n34691 , n34690 );
not ( n34692 , n34691 );
or ( n34693 , n34676 , n34692 );
not ( n34694 , n34625 );
not ( n34695 , n34193 );
and ( n34696 , n34695 , n34565 );
xor ( n34697 , n34566 , n34611 );
and ( n34698 , n34697 , n34193 );
or ( n34699 , n34696 , n34698 );
and ( n34700 , n34694 , n34699 );
not ( n34701 , n34699 );
and ( n34702 , n34684 , n34685 );
xor ( n34703 , n34701 , n34702 );
and ( n34704 , n34703 , n34625 );
or ( n34705 , n34700 , n34704 );
not ( n34706 , n34705 );
buf ( n34707 , n34706 );
buf ( n34708 , n34707 );
not ( n34709 , n34708 );
or ( n34710 , n34693 , n34709 );
not ( n34711 , n34625 );
not ( n34712 , n34193 );
and ( n34713 , n34712 , n34555 );
xor ( n34714 , n34556 , n34612 );
and ( n34715 , n34714 , n34193 );
or ( n34716 , n34713 , n34715 );
and ( n34717 , n34711 , n34716 );
not ( n34718 , n34716 );
and ( n34719 , n34701 , n34702 );
xor ( n34720 , n34718 , n34719 );
and ( n34721 , n34720 , n34625 );
or ( n34722 , n34717 , n34721 );
not ( n34723 , n34722 );
buf ( n34724 , n34723 );
buf ( n34725 , n34724 );
not ( n34726 , n34725 );
or ( n34727 , n34710 , n34726 );
not ( n34728 , n34625 );
not ( n34729 , n34193 );
and ( n34730 , n34729 , n34545 );
xor ( n34731 , n34546 , n34613 );
and ( n34732 , n34731 , n34193 );
or ( n34733 , n34730 , n34732 );
and ( n34734 , n34728 , n34733 );
not ( n34735 , n34733 );
and ( n34736 , n34718 , n34719 );
xor ( n34737 , n34735 , n34736 );
and ( n34738 , n34737 , n34625 );
or ( n34739 , n34734 , n34738 );
not ( n34740 , n34739 );
buf ( n34741 , n34740 );
buf ( n34742 , n34741 );
not ( n34743 , n34742 );
or ( n34744 , n34727 , n34743 );
buf ( n34745 , n34744 );
buf ( n34746 , n34745 );
and ( n34747 , n34746 , n34625 );
not ( n34748 , n34747 );
and ( n34749 , n34748 , n34692 );
xor ( n34750 , n34692 , n34625 );
xor ( n34751 , n34675 , n34625 );
xor ( n34752 , n34658 , n34625 );
xor ( n34753 , n34641 , n34625 );
xor ( n34754 , n34415 , n34625 );
and ( n34755 , n34754 , n34625 );
and ( n34756 , n34753 , n34755 );
and ( n34757 , n34752 , n34756 );
and ( n34758 , n34751 , n34757 );
xor ( n34759 , n34750 , n34758 );
and ( n34760 , n34759 , n34747 );
or ( n34761 , n34749 , n34760 );
and ( n34762 , n34761 , n34358 );
or ( n34763 , n34360 , n34762 );
and ( n34764 , n34356 , n34763 );
not ( n34765 , n34193 );
and ( n34766 , n34765 , n34429 );
not ( n34767 , n34429 );
not ( n34768 , n34431 );
not ( n34769 , n34433 );
not ( n34770 , n34435 );
not ( n34771 , n34437 );
not ( n34772 , n34439 );
not ( n34773 , n34441 );
not ( n34774 , n34443 );
not ( n34775 , n34362 );
not ( n34776 , n34365 );
not ( n34777 , n34367 );
not ( n34778 , n34369 );
not ( n34779 , n34371 );
not ( n34780 , n34373 );
not ( n34781 , n34375 );
not ( n34782 , n34377 );
not ( n34783 , n34379 );
not ( n34784 , n34273 );
not ( n34785 , n34260 );
not ( n34786 , n34247 );
not ( n34787 , n34234 );
not ( n34788 , n34221 );
not ( n34789 , n34208 );
not ( n34790 , n34195 );
not ( n34791 , n34188 );
and ( n34792 , n34790 , n34791 );
and ( n34793 , n34789 , n34792 );
and ( n34794 , n34788 , n34793 );
and ( n34795 , n34787 , n34794 );
and ( n34796 , n34786 , n34795 );
and ( n34797 , n34785 , n34796 );
and ( n34798 , n34784 , n34797 );
and ( n34799 , n34783 , n34798 );
and ( n34800 , n34782 , n34799 );
and ( n34801 , n34781 , n34800 );
and ( n34802 , n34780 , n34801 );
and ( n34803 , n34779 , n34802 );
and ( n34804 , n34778 , n34803 );
and ( n34805 , n34777 , n34804 );
and ( n34806 , n34776 , n34805 );
and ( n34807 , n34775 , n34806 );
and ( n34808 , n34774 , n34807 );
and ( n34809 , n34773 , n34808 );
and ( n34810 , n34772 , n34809 );
and ( n34811 , n34771 , n34810 );
and ( n34812 , n34770 , n34811 );
and ( n34813 , n34769 , n34812 );
and ( n34814 , n34768 , n34813 );
xor ( n34815 , n34767 , n34814 );
and ( n34816 , n34815 , n34193 );
or ( n34817 , n34766 , n34816 );
not ( n34818 , n34817 );
buf ( n34819 , n34818 );
buf ( n34820 , n34819 );
not ( n34821 , n34820 );
buf ( n34822 , n34821 );
buf ( n34823 , n34822 );
not ( n34824 , n34823 );
buf ( n34825 , n34824 );
not ( n34826 , n34825 );
not ( n34827 , n34193 );
not ( n34828 , n34417 );
not ( n34829 , n34419 );
not ( n34830 , n34421 );
not ( n34831 , n34423 );
not ( n34832 , n34425 );
not ( n34833 , n34427 );
and ( n34834 , n34767 , n34814 );
and ( n34835 , n34833 , n34834 );
and ( n34836 , n34832 , n34835 );
and ( n34837 , n34831 , n34836 );
and ( n34838 , n34830 , n34837 );
and ( n34839 , n34829 , n34838 );
and ( n34840 , n34828 , n34839 );
xor ( n34841 , n34827 , n34840 );
buf ( n34842 , n34193 );
and ( n34843 , n34841 , n34842 );
buf ( n34844 , n34843 );
not ( n34845 , n34844 );
not ( n34846 , n34845 );
not ( n34847 , n34846 );
not ( n34848 , n34193 );
and ( n34849 , n34848 , n34417 );
xor ( n34850 , n34828 , n34839 );
and ( n34851 , n34850 , n34193 );
or ( n34852 , n34849 , n34851 );
not ( n34853 , n34852 );
buf ( n34854 , n34853 );
buf ( n34855 , n34854 );
not ( n34856 , n34855 );
not ( n34857 , n34856 );
not ( n34858 , n34193 );
and ( n34859 , n34858 , n34419 );
xor ( n34860 , n34829 , n34838 );
and ( n34861 , n34860 , n34193 );
or ( n34862 , n34859 , n34861 );
not ( n34863 , n34862 );
buf ( n34864 , n34863 );
buf ( n34865 , n34864 );
not ( n34866 , n34865 );
not ( n34867 , n34866 );
not ( n34868 , n34193 );
and ( n34869 , n34868 , n34421 );
xor ( n34870 , n34830 , n34837 );
and ( n34871 , n34870 , n34193 );
or ( n34872 , n34869 , n34871 );
not ( n34873 , n34872 );
buf ( n34874 , n34873 );
buf ( n34875 , n34874 );
not ( n34876 , n34875 );
not ( n34877 , n34876 );
not ( n34878 , n34193 );
and ( n34879 , n34878 , n34423 );
xor ( n34880 , n34831 , n34836 );
and ( n34881 , n34880 , n34193 );
or ( n34882 , n34879 , n34881 );
not ( n34883 , n34882 );
buf ( n34884 , n34883 );
buf ( n34885 , n34884 );
not ( n34886 , n34885 );
not ( n34887 , n34886 );
not ( n34888 , n34193 );
and ( n34889 , n34888 , n34425 );
xor ( n34890 , n34832 , n34835 );
and ( n34891 , n34890 , n34193 );
or ( n34892 , n34889 , n34891 );
not ( n34893 , n34892 );
buf ( n34894 , n34893 );
buf ( n34895 , n34894 );
not ( n34896 , n34895 );
not ( n34897 , n34896 );
not ( n34898 , n34193 );
and ( n34899 , n34898 , n34427 );
xor ( n34900 , n34833 , n34834 );
and ( n34901 , n34900 , n34193 );
or ( n34902 , n34899 , n34901 );
not ( n34903 , n34902 );
buf ( n34904 , n34903 );
buf ( n34905 , n34904 );
not ( n34906 , n34905 );
not ( n34907 , n34906 );
not ( n34908 , n34821 );
and ( n34909 , n34907 , n34908 );
and ( n34910 , n34897 , n34909 );
and ( n34911 , n34887 , n34910 );
and ( n34912 , n34877 , n34911 );
and ( n34913 , n34867 , n34912 );
and ( n34914 , n34857 , n34913 );
and ( n34915 , n34847 , n34914 );
not ( n34916 , n34915 );
and ( n34917 , n34916 , n34193 );
buf ( n34918 , n34917 );
not ( n34919 , n34918 );
not ( n34920 , n34193 );
and ( n34921 , n34920 , n34906 );
xor ( n34922 , n34907 , n34908 );
and ( n34923 , n34922 , n34193 );
or ( n34924 , n34921 , n34923 );
and ( n34925 , n34919 , n34924 );
not ( n34926 , n34924 );
not ( n34927 , n34822 );
xor ( n34928 , n34926 , n34927 );
and ( n34929 , n34928 , n34918 );
or ( n34930 , n34925 , n34929 );
not ( n34931 , n34930 );
buf ( n34932 , n34931 );
buf ( n34933 , n34932 );
not ( n34934 , n34933 );
or ( n34935 , n34826 , n34934 );
not ( n34936 , n34918 );
not ( n34937 , n34193 );
and ( n34938 , n34937 , n34896 );
xor ( n34939 , n34897 , n34909 );
and ( n34940 , n34939 , n34193 );
or ( n34941 , n34938 , n34940 );
and ( n34942 , n34936 , n34941 );
not ( n34943 , n34941 );
and ( n34944 , n34926 , n34927 );
xor ( n34945 , n34943 , n34944 );
and ( n34946 , n34945 , n34918 );
or ( n34947 , n34942 , n34946 );
not ( n34948 , n34947 );
buf ( n34949 , n34948 );
buf ( n34950 , n34949 );
not ( n34951 , n34950 );
or ( n34952 , n34935 , n34951 );
not ( n34953 , n34918 );
not ( n34954 , n34193 );
and ( n34955 , n34954 , n34886 );
xor ( n34956 , n34887 , n34910 );
and ( n34957 , n34956 , n34193 );
or ( n34958 , n34955 , n34957 );
and ( n34959 , n34953 , n34958 );
not ( n34960 , n34958 );
and ( n34961 , n34943 , n34944 );
xor ( n34962 , n34960 , n34961 );
and ( n34963 , n34962 , n34918 );
or ( n34964 , n34959 , n34963 );
not ( n34965 , n34964 );
buf ( n34966 , n34965 );
buf ( n34967 , n34966 );
not ( n34968 , n34967 );
or ( n34969 , n34952 , n34968 );
not ( n34970 , n34918 );
not ( n34971 , n34193 );
and ( n34972 , n34971 , n34876 );
xor ( n34973 , n34877 , n34911 );
and ( n34974 , n34973 , n34193 );
or ( n34975 , n34972 , n34974 );
and ( n34976 , n34970 , n34975 );
not ( n34977 , n34975 );
and ( n34978 , n34960 , n34961 );
xor ( n34979 , n34977 , n34978 );
and ( n34980 , n34979 , n34918 );
or ( n34981 , n34976 , n34980 );
not ( n34982 , n34981 );
buf ( n34983 , n34982 );
buf ( n34984 , n34983 );
not ( n34985 , n34984 );
or ( n34986 , n34969 , n34985 );
not ( n34987 , n34918 );
not ( n34988 , n34193 );
and ( n34989 , n34988 , n34866 );
xor ( n34990 , n34867 , n34912 );
and ( n34991 , n34990 , n34193 );
or ( n34992 , n34989 , n34991 );
and ( n34993 , n34987 , n34992 );
not ( n34994 , n34992 );
and ( n34995 , n34977 , n34978 );
xor ( n34996 , n34994 , n34995 );
and ( n34997 , n34996 , n34918 );
or ( n34998 , n34993 , n34997 );
not ( n34999 , n34998 );
buf ( n35000 , n34999 );
buf ( n35001 , n35000 );
not ( n35002 , n35001 );
or ( n35003 , n34986 , n35002 );
not ( n35004 , n34918 );
not ( n35005 , n34193 );
and ( n35006 , n35005 , n34856 );
xor ( n35007 , n34857 , n34913 );
and ( n35008 , n35007 , n34193 );
or ( n35009 , n35006 , n35008 );
and ( n35010 , n35004 , n35009 );
not ( n35011 , n35009 );
and ( n35012 , n34994 , n34995 );
xor ( n35013 , n35011 , n35012 );
and ( n35014 , n35013 , n34918 );
or ( n35015 , n35010 , n35014 );
not ( n35016 , n35015 );
buf ( n35017 , n35016 );
buf ( n35018 , n35017 );
not ( n35019 , n35018 );
or ( n35020 , n35003 , n35019 );
xor ( n35021 , n34847 , n34914 );
and ( n35022 , n35021 , n34193 );
buf ( n35023 , n35022 );
not ( n35024 , n35023 );
and ( n35025 , n35011 , n35012 );
xor ( n35026 , n35024 , n35025 );
and ( n35027 , n35026 , n34918 );
buf ( n35028 , n35027 );
not ( n35029 , n35028 );
buf ( n35030 , n35029 );
buf ( n35031 , n35030 );
not ( n35032 , n35031 );
or ( n35033 , n35020 , n35032 );
buf ( n35034 , n35033 );
buf ( n35035 , n35034 );
and ( n35036 , n35035 , n34918 );
not ( n35037 , n35036 );
and ( n35038 , n35037 , n34985 );
xor ( n35039 , n34985 , n34918 );
xor ( n35040 , n34968 , n34918 );
xor ( n35041 , n34951 , n34918 );
xor ( n35042 , n34934 , n34918 );
xor ( n35043 , n34826 , n34918 );
and ( n35044 , n35043 , n34918 );
and ( n35045 , n35042 , n35044 );
and ( n35046 , n35041 , n35045 );
and ( n35047 , n35040 , n35046 );
xor ( n35048 , n35039 , n35047 );
and ( n35049 , n35048 , n35036 );
or ( n35050 , n35038 , n35049 );
and ( n35051 , n35050 , n34355 );
or ( n35052 , n34764 , n35051 );
and ( n35053 , n35052 , n32968 );
or ( n35054 , n34317 , n35053 );
and ( n35055 , n35054 , n33370 );
nor ( n35056 , n32511 , n32520 , n32523 , n32526 );
or ( n35057 , n33372 , n35056 );
or ( n35058 , n35057 , n33373 );
or ( n35059 , n35058 , n33208 );
or ( n35060 , n35059 , n33377 );
or ( n35061 , n35060 , n33379 );
or ( n35062 , n35061 , n32528 );
and ( n35063 , n32783 , n35062 );
or ( n35064 , C0 , n34161 , n34307 , n35055 , n35063 );
buf ( n35065 , n35064 );
buf ( n35066 , n35065 );
not ( n35067 , n34150 );
and ( n35068 , n35067 , n32749 );
not ( n35069 , n34154 );
and ( n35070 , n35069 , n32749 );
and ( n35071 , n32755 , n34154 );
or ( n35072 , n35070 , n35071 );
and ( n35073 , n35072 , n34150 );
or ( n35074 , n35068 , n35073 );
and ( n35075 , n35074 , n33381 );
not ( n35076 , n34184 );
not ( n35077 , n34154 );
and ( n35078 , n35077 , n32749 );
not ( n35079 , n34287 );
and ( n35080 , n35079 , n34231 );
xor ( n35081 , n34291 , n34297 );
and ( n35082 , n35081 , n34287 );
or ( n35083 , n35080 , n35082 );
and ( n35084 , n35083 , n34154 );
or ( n35085 , n35078 , n35084 );
and ( n35086 , n35076 , n35085 );
and ( n35087 , n35083 , n34184 );
or ( n35088 , n35086 , n35087 );
and ( n35089 , n35088 , n33375 );
not ( n35090 , n32968 );
not ( n35091 , n34184 );
not ( n35092 , n34154 );
and ( n35093 , n35092 , n32749 );
and ( n35094 , n35083 , n34154 );
or ( n35095 , n35093 , n35094 );
and ( n35096 , n35091 , n35095 );
and ( n35097 , n35083 , n34184 );
or ( n35098 , n35096 , n35097 );
and ( n35099 , n35090 , n35098 );
not ( n35100 , n34355 );
not ( n35101 , n34358 );
and ( n35102 , n35101 , n35098 );
not ( n35103 , n34747 );
and ( n35104 , n35103 , n34675 );
xor ( n35105 , n34751 , n34757 );
and ( n35106 , n35105 , n34747 );
or ( n35107 , n35104 , n35106 );
and ( n35108 , n35107 , n34358 );
or ( n35109 , n35102 , n35108 );
and ( n35110 , n35100 , n35109 );
not ( n35111 , n35036 );
and ( n35112 , n35111 , n34968 );
xor ( n35113 , n35040 , n35046 );
and ( n35114 , n35113 , n35036 );
or ( n35115 , n35112 , n35114 );
and ( n35116 , n35115 , n34355 );
or ( n35117 , n35110 , n35116 );
and ( n35118 , n35117 , n32968 );
or ( n35119 , n35099 , n35118 );
and ( n35120 , n35119 , n33370 );
and ( n35121 , n32749 , n35062 );
or ( n35122 , C0 , n35075 , n35089 , n35120 , n35121 );
buf ( n35123 , n35122 );
buf ( n35124 , n35123 );
buf ( n35125 , n31655 );
buf ( n35126 , n30987 );
and ( n35127 , n33235 , n32528 );
not ( n35128 , n32598 );
and ( n35129 , n35128 , n32998 );
buf ( n35130 , n35129 );
and ( n35131 , n35130 , n32890 );
not ( n35132 , n32919 );
and ( n35133 , n35132 , n32998 );
buf ( n35134 , n35133 );
and ( n35135 , n35134 , n32924 );
not ( n35136 , n32953 );
and ( n35137 , n35136 , n32998 );
not ( n35138 , n32971 );
and ( n35139 , n35138 , n33121 );
xor ( n35140 , n32998 , n33007 );
and ( n35141 , n35140 , n32971 );
or ( n35142 , n35139 , n35141 );
and ( n35143 , n35142 , n32953 );
or ( n35144 , n35137 , n35143 );
and ( n35145 , n35144 , n33038 );
not ( n35146 , n33067 );
and ( n35147 , n35146 , n32998 );
not ( n35148 , n32970 );
not ( n35149 , n33071 );
and ( n35150 , n35149 , n33121 );
xor ( n35151 , n33122 , n33139 );
and ( n35152 , n35151 , n33071 );
or ( n35153 , n35150 , n35152 );
and ( n35154 , n35148 , n35153 );
and ( n35155 , n35140 , n32970 );
or ( n35156 , n35154 , n35155 );
and ( n35157 , n35156 , n33067 );
or ( n35158 , n35147 , n35157 );
and ( n35159 , n35158 , n33172 );
and ( n35160 , n32998 , n33204 );
or ( n35161 , n35131 , n35135 , n35145 , n35159 , n35160 );
and ( n35162 , n35161 , n33208 );
not ( n35163 , n32968 );
not ( n35164 , n33270 );
and ( n35165 , n35164 , n33321 );
xor ( n35166 , n33322 , n33339 );
and ( n35167 , n35166 , n33270 );
or ( n35168 , n35165 , n35167 );
and ( n35169 , n35163 , n35168 );
and ( n35170 , n32998 , n32968 );
or ( n35171 , n35169 , n35170 );
and ( n35172 , n35171 , n33370 );
buf ( n35173 , n35056 );
and ( n35174 , n32998 , n33382 );
or ( n35175 , C0 , n35127 , n35162 , n35172 , n35173 , n35174 );
buf ( n35176 , n35175 );
buf ( n35177 , n35176 );
buf ( n35178 , n31655 );
buf ( n35179 , n30987 );
buf ( n35180 , n30987 );
buf ( n35181 , n31655 );
buf ( n35182 , RI15b62b50_1233);
and ( n35183 , n35182 , n32500 );
not ( n35184 , n31689 );
buf ( n35185 , n31689 );
buf ( n35186 , n31689 );
buf ( n35187 , n31689 );
buf ( n35188 , n31689 );
buf ( n35189 , n31689 );
buf ( n35190 , n31689 );
buf ( n35191 , n31689 );
buf ( n35192 , n31689 );
buf ( n35193 , n31689 );
buf ( n35194 , n31689 );
buf ( n35195 , n31689 );
buf ( n35196 , n31689 );
buf ( n35197 , n31689 );
buf ( n35198 , n31689 );
buf ( n35199 , n31689 );
buf ( n35200 , n31689 );
buf ( n35201 , n31689 );
buf ( n35202 , n31689 );
buf ( n35203 , n31689 );
buf ( n35204 , n31689 );
buf ( n35205 , n31689 );
buf ( n35206 , n31689 );
buf ( n35207 , n31689 );
buf ( n35208 , n31689 );
buf ( n35209 , n31689 );
or ( n35210 , n31721 , n31692 , n31694 , n31689 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n31723 );
and ( n35211 , n35184 , n35210 );
not ( n35212 , n35211 );
buf ( n35213 , RI15b63a50_1265);
and ( n35214 , n35212 , n35213 );
and ( n35215 , n31751 , n35211 );
or ( n35216 , n35214 , n35215 );
and ( n35217 , n35216 , n32421 );
not ( n35218 , n31689 );
buf ( n35219 , n31689 );
buf ( n35220 , n31689 );
buf ( n35221 , n31689 );
buf ( n35222 , n31689 );
buf ( n35223 , n31689 );
buf ( n35224 , n31689 );
buf ( n35225 , n31689 );
buf ( n35226 , n31689 );
buf ( n35227 , n31689 );
buf ( n35228 , n31689 );
buf ( n35229 , n31689 );
buf ( n35230 , n31689 );
buf ( n35231 , n31689 );
buf ( n35232 , n31689 );
buf ( n35233 , n31689 );
buf ( n35234 , n31689 );
buf ( n35235 , n31689 );
buf ( n35236 , n31689 );
buf ( n35237 , n31689 );
buf ( n35238 , n31689 );
buf ( n35239 , n31689 );
buf ( n35240 , n31689 );
buf ( n35241 , n31689 );
buf ( n35242 , n31689 );
buf ( n35243 , n31689 );
or ( n35244 , n31721 , n31692 , n31694 , n31689 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n31723 );
and ( n35245 , n35218 , n35244 );
not ( n35246 , n35245 );
and ( n35247 , n35246 , n35213 );
and ( n35248 , n31751 , n35245 );
or ( n35249 , n35247 , n35248 );
and ( n35250 , n35249 , n32419 );
not ( n35251 , n31689 );
buf ( n35252 , n31689 );
buf ( n35253 , n31689 );
buf ( n35254 , n31689 );
buf ( n35255 , n31689 );
buf ( n35256 , n31689 );
buf ( n35257 , n31689 );
buf ( n35258 , n31689 );
buf ( n35259 , n31689 );
buf ( n35260 , n31689 );
buf ( n35261 , n31689 );
buf ( n35262 , n31689 );
buf ( n35263 , n31689 );
buf ( n35264 , n31689 );
buf ( n35265 , n31689 );
buf ( n35266 , n31689 );
buf ( n35267 , n31689 );
buf ( n35268 , n31689 );
buf ( n35269 , n31689 );
buf ( n35270 , n31689 );
buf ( n35271 , n31689 );
buf ( n35272 , n31689 );
buf ( n35273 , n31689 );
buf ( n35274 , n31689 );
buf ( n35275 , n31689 );
buf ( n35276 , n31689 );
or ( n35277 , n31721 , n31692 , n31694 , n31689 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n31723 );
and ( n35278 , n35251 , n35277 );
not ( n35279 , n35278 );
and ( n35280 , n35279 , n35213 );
buf ( n35281 , RI15b60be8_1166);
buf ( n35282 , RI15b60c60_1167);
not ( n35283 , n35282 );
buf ( n35284 , RI15b60cd8_1168);
nor ( n35285 , n35281 , n35283 , n35284 );
not ( n35286 , n35281 );
and ( n35287 , n35286 , n35283 , n35284 );
or ( n35288 , n35285 , n35287 );
buf ( n35289 , RI15b66750_1361);
buf ( n35290 , RI15b3fb28_38);
and ( n35291 , n35289 , n35290 );
not ( n35292 , n35291 );
not ( n35293 , n32475 );
and ( n35294 , n35292 , n35293 );
and ( n35295 , n35288 , n35294 );
not ( n35296 , n35295 );
buf ( n35297 , RI15b61c50_1201);
and ( n35298 , n35296 , n35297 );
and ( n35299 , n35213 , n35295 );
or ( n35300 , n35298 , n35299 );
and ( n35301 , n35300 , n35278 );
or ( n35302 , n35280 , n35301 );
and ( n35303 , n35302 , n32417 );
not ( n35304 , n31689 );
buf ( n35305 , n31689 );
buf ( n35306 , n31689 );
buf ( n35307 , n31689 );
buf ( n35308 , n31689 );
buf ( n35309 , n31689 );
buf ( n35310 , n31689 );
buf ( n35311 , n31689 );
buf ( n35312 , n31689 );
buf ( n35313 , n31689 );
buf ( n35314 , n31689 );
buf ( n35315 , n31689 );
buf ( n35316 , n31689 );
buf ( n35317 , n31689 );
buf ( n35318 , n31689 );
buf ( n35319 , n31689 );
buf ( n35320 , n31689 );
buf ( n35321 , n31689 );
buf ( n35322 , n31689 );
buf ( n35323 , n31689 );
buf ( n35324 , n31689 );
buf ( n35325 , n31689 );
buf ( n35326 , n31689 );
buf ( n35327 , n31689 );
buf ( n35328 , n31689 );
buf ( n35329 , n31689 );
or ( n35330 , n31721 , n31692 , n31694 , n31689 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n31723 );
and ( n35331 , n35304 , n35330 );
not ( n35332 , n35331 );
and ( n35333 , n35332 , n35213 );
not ( n35334 , n35294 );
buf ( n35335 , n35297 );
and ( n35336 , n35334 , n35335 );
and ( n35337 , n35213 , n35294 );
or ( n35338 , n35336 , n35337 );
and ( n35339 , n35338 , n35331 );
or ( n35340 , n35333 , n35339 );
and ( n35341 , n35340 , n32415 );
or ( n35342 , n32405 , n32398 );
or ( n35343 , n35342 , n32253 );
or ( n35344 , n35343 , n32406 );
or ( n35345 , n35344 , n32409 );
or ( n35346 , n35345 , n32411 );
or ( n35347 , n35346 , n32413 );
or ( n35348 , n35347 , n32423 );
or ( n35349 , n35348 , n32425 );
or ( n35350 , n35349 , n32427 );
or ( n35351 , n35350 , n32429 );
or ( n35352 , n35351 , n32431 );
or ( n35353 , n35352 , n32433 );
or ( n35354 , n35353 , n32435 );
and ( n35355 , n35213 , n35354 );
or ( n35356 , n35217 , n35250 , n35303 , n35341 , n35355 );
and ( n35357 , n35356 , n32456 );
not ( n35358 , n32475 );
buf ( n35359 , n35182 );
and ( n35360 , n35358 , n35359 );
and ( n35361 , n35213 , n32475 );
or ( n35362 , n35360 , n35361 );
and ( n35363 , n35362 , n32486 );
or ( n35364 , n32493 , n32473 );
or ( n35365 , n35364 , n32494 );
or ( n35366 , n35365 , n32496 );
or ( n35367 , n35366 , n32498 );
and ( n35368 , n35213 , n35367 );
or ( n35369 , C0 , n35183 , n35357 , n35363 , C0 , n35368 );
buf ( n35370 , n35369 );
buf ( n35371 , n35370 );
buf ( n35372 , n30987 );
and ( n35373 , n31560 , n31007 );
not ( n35374 , n31077 );
buf ( n35375 , RI15b58470_877);
and ( n35376 , n35374 , n35375 );
buf ( n35377 , n35376 );
and ( n35378 , n35377 , n31373 );
not ( n35379 , n31402 );
and ( n35380 , n35379 , n35375 );
buf ( n35381 , n35380 );
and ( n35382 , n35381 , n31408 );
not ( n35383 , n31437 );
and ( n35384 , n35383 , n35375 );
not ( n35385 , n31455 );
and ( n35386 , n35385 , n31501 );
buf ( n35387 , RI15b583f8_876);
buf ( n35388 , RI15b58380_875);
buf ( n35389 , RI15b58308_874);
buf ( n35390 , RI15b58290_873);
buf ( n35391 , RI15b58218_872);
buf ( n35392 , RI15b581a0_871);
buf ( n35393 , RI15b58128_870);
buf ( n35394 , RI15b580b0_869);
buf ( n35395 , RI15b58038_868);
buf ( n35396 , RI15b57f48_866);
buf ( n35397 , RI15b57ed0_865);
buf ( n35398 , RI15b57e58_864);
and ( n35399 , n33986 , n34025 );
and ( n35400 , n35398 , n35399 );
and ( n35401 , n35397 , n35400 );
and ( n35402 , n35396 , n35401 );
and ( n35403 , n33972 , n35402 );
and ( n35404 , n35395 , n35403 );
and ( n35405 , n35394 , n35404 );
and ( n35406 , n35393 , n35405 );
and ( n35407 , n35392 , n35406 );
and ( n35408 , n35391 , n35407 );
and ( n35409 , n35390 , n35408 );
and ( n35410 , n35389 , n35409 );
and ( n35411 , n35388 , n35410 );
and ( n35412 , n35387 , n35411 );
xor ( n35413 , n35375 , n35412 );
and ( n35414 , n35413 , n31455 );
or ( n35415 , n35386 , n35414 );
and ( n35416 , n35415 , n31437 );
or ( n35417 , n35384 , n35416 );
and ( n35418 , n35417 , n31468 );
not ( n35419 , n31497 );
and ( n35420 , n35419 , n35375 );
not ( n35421 , n31454 );
not ( n35422 , n31501 );
buf ( n35423 , RI15b565f8_812);
not ( n35424 , n35423 );
buf ( n35425 , RI15b56580_811);
not ( n35426 , n35425 );
buf ( n35427 , RI15b56508_810);
not ( n35428 , n35427 );
buf ( n35429 , RI15b56490_809);
not ( n35430 , n35429 );
buf ( n35431 , RI15b56418_808);
not ( n35432 , n35431 );
buf ( n35433 , RI15b563a0_807);
not ( n35434 , n35433 );
buf ( n35435 , RI15b56328_806);
not ( n35436 , n35435 );
buf ( n35437 , RI15b562b0_805);
not ( n35438 , n35437 );
buf ( n35439 , RI15b56238_804);
not ( n35440 , n35439 );
buf ( n35441 , RI15b561c0_803);
not ( n35442 , n35441 );
buf ( n35443 , RI15b56148_802);
not ( n35444 , n35443 );
buf ( n35445 , RI15b560d0_801);
not ( n35446 , n35445 );
buf ( n35447 , RI15b56058_800);
not ( n35448 , n35447 );
and ( n35449 , n34037 , n34077 );
and ( n35450 , n35448 , n35449 );
and ( n35451 , n35446 , n35450 );
and ( n35452 , n35444 , n35451 );
and ( n35453 , n35442 , n35452 );
and ( n35454 , n35440 , n35453 );
and ( n35455 , n35438 , n35454 );
and ( n35456 , n35436 , n35455 );
and ( n35457 , n35434 , n35456 );
and ( n35458 , n35432 , n35457 );
and ( n35459 , n35430 , n35458 );
and ( n35460 , n35428 , n35459 );
and ( n35461 , n35426 , n35460 );
and ( n35462 , n35424 , n35461 );
xor ( n35463 , n35422 , n35462 );
buf ( n35464 , n31501 );
and ( n35465 , n35463 , n35464 );
buf ( n35466 , n35465 );
and ( n35467 , n35421 , n35466 );
and ( n35468 , n35413 , n31454 );
or ( n35469 , n35467 , n35468 );
and ( n35470 , n35469 , n31497 );
or ( n35471 , n35420 , n35470 );
and ( n35472 , n35471 , n31521 );
and ( n35473 , n35375 , n31553 );
or ( n35474 , n35378 , n35382 , n35418 , n35472 , n35473 );
and ( n35475 , n35474 , n31557 );
not ( n35476 , n31452 );
not ( n35477 , n31619 );
xor ( n35478 , n31561 , n31617 );
not ( n35479 , n35478 );
xor ( n35480 , n31562 , n31616 );
not ( n35481 , n35480 );
xor ( n35482 , n31563 , n31615 );
not ( n35483 , n35482 );
xor ( n35484 , n31564 , n31614 );
not ( n35485 , n35484 );
xor ( n35486 , n31565 , n31613 );
not ( n35487 , n35486 );
xor ( n35488 , n31566 , n31612 );
not ( n35489 , n35488 );
xor ( n35490 , n31567 , n31611 );
not ( n35491 , n35490 );
xor ( n35492 , n31568 , n31610 );
not ( n35493 , n35492 );
xor ( n35494 , n31569 , n31609 );
not ( n35495 , n35494 );
not ( n35496 , n33946 );
xor ( n35497 , n31571 , n31607 );
not ( n35498 , n35497 );
xor ( n35499 , n31572 , n31606 );
not ( n35500 , n35499 );
xor ( n35501 , n31573 , n31605 );
not ( n35502 , n35501 );
and ( n35503 , n34094 , n34134 );
and ( n35504 , n35502 , n35503 );
and ( n35505 , n35500 , n35504 );
and ( n35506 , n35498 , n35505 );
and ( n35507 , n35496 , n35506 );
and ( n35508 , n35495 , n35507 );
and ( n35509 , n35493 , n35508 );
and ( n35510 , n35491 , n35509 );
and ( n35511 , n35489 , n35510 );
and ( n35512 , n35487 , n35511 );
and ( n35513 , n35485 , n35512 );
and ( n35514 , n35483 , n35513 );
and ( n35515 , n35481 , n35514 );
and ( n35516 , n35479 , n35515 );
xor ( n35517 , n35477 , n35516 );
buf ( n35518 , n31619 );
and ( n35519 , n35517 , n35518 );
buf ( n35520 , n35519 );
and ( n35521 , n35476 , n35520 );
and ( n35522 , n35375 , n31452 );
or ( n35523 , n35521 , n35522 );
and ( n35524 , n35523 , n31638 );
and ( n35525 , n35375 , n31650 );
or ( n35526 , C0 , n35373 , n35475 , n35524 , C0 , n35525 );
buf ( n35527 , n35526 );
buf ( n35528 , n35527 );
buf ( n35529 , RI15b605d0_1153);
buf ( n35530 , RI15b60648_1154);
not ( n35531 , n35530 );
nand ( n35532 , n35529 , n35531 );
buf ( n35533 , RI15b54168_734);
buf ( n35534 , RI15b541e0_735);
not ( n35535 , n35534 );
nand ( n35536 , n35533 , n35535 );
and ( n35537 , n35532 , n35536 );
buf ( n35538 , RI15b47d00_315);
buf ( n35539 , RI15b47d78_316);
not ( n35540 , n35539 );
nand ( n35541 , n35538 , n35540 );
and ( n35542 , n35537 , n35541 );
not ( n35543 , n35542 );
buf ( n35544 , RI15b51558_640);
and ( n35545 , n35543 , n35544 );
buf ( n35546 , RI15b450f0_221);
and ( n35547 , n35546 , n35542 );
or ( n35548 , n35545 , n35547 );
buf ( n35549 , n35548 );
buf ( n35550 , n35549 );
buf ( n35551 , n31655 );
buf ( n35552 , n30987 );
not ( n35553 , n33419 );
and ( n35554 , n35553 , n31584 );
xor ( n35555 , n33478 , n33533 );
xor ( n35556 , n35555 , n33685 );
and ( n35557 , n35556 , n33419 );
or ( n35558 , n35554 , n35557 );
and ( n35559 , n35558 , n31529 );
not ( n35560 , n33734 );
and ( n35561 , n35560 , n31584 );
not ( n35562 , n33533 );
xor ( n35563 , n33771 , n33533 );
xor ( n35564 , n35563 , n33803 );
and ( n35565 , n35562 , n35564 );
xor ( n35566 , n33856 , n33858 );
xor ( n35567 , n35566 , n33905 );
and ( n35568 , n35567 , n33533 );
or ( n35569 , n35565 , n35568 );
and ( n35570 , n35569 , n33734 );
or ( n35571 , n35561 , n35570 );
and ( n35572 , n35571 , n31527 );
and ( n35573 , n31584 , n33942 );
or ( n35574 , n35559 , n35572 , n35573 );
and ( n35575 , n35574 , n31557 );
and ( n35576 , n34113 , n31643 );
not ( n35577 , n31452 );
and ( n35578 , n35577 , n34113 );
xor ( n35579 , n31584 , n33953 );
and ( n35580 , n35579 , n31452 );
or ( n35581 , n35578 , n35580 );
and ( n35582 , n35581 , n31638 );
and ( n35583 , n34008 , n33973 );
and ( n35584 , n31584 , n33978 );
or ( n35585 , C0 , n35575 , n35576 , n35582 , n35583 , n35584 );
buf ( n35586 , n35585 );
buf ( n35587 , n35586 );
buf ( n35588 , n31655 );
buf ( n35589 , n30987 );
and ( n35590 , n33211 , n32528 );
not ( n35591 , n32598 );
buf ( n35592 , RI15b4c008_458);
and ( n35593 , n35591 , n35592 );
buf ( n35594 , n35593 );
and ( n35595 , n35594 , n32890 );
not ( n35596 , n32919 );
and ( n35597 , n35596 , n35592 );
buf ( n35598 , n35597 );
and ( n35599 , n35598 , n32924 );
not ( n35600 , n32953 );
and ( n35601 , n35600 , n35592 );
not ( n35602 , n32971 );
and ( n35603 , n35602 , n33071 );
and ( n35604 , n32600 , n33031 );
xor ( n35605 , n35592 , n35604 );
and ( n35606 , n35605 , n32971 );
or ( n35607 , n35603 , n35606 );
and ( n35608 , n35607 , n32953 );
or ( n35609 , n35601 , n35608 );
and ( n35610 , n35609 , n33038 );
not ( n35611 , n33067 );
and ( n35612 , n35611 , n35592 );
not ( n35613 , n32970 );
not ( n35614 , n33071 );
and ( n35615 , n33074 , n33163 );
xor ( n35616 , n35614 , n35615 );
buf ( n35617 , n33071 );
and ( n35618 , n35616 , n35617 );
buf ( n35619 , n35618 );
and ( n35620 , n35613 , n35619 );
and ( n35621 , n35605 , n32970 );
or ( n35622 , n35620 , n35621 );
and ( n35623 , n35622 , n33067 );
or ( n35624 , n35612 , n35623 );
and ( n35625 , n35624 , n33172 );
and ( n35626 , n35592 , n33204 );
or ( n35627 , n35595 , n35599 , n35610 , n35625 , n35626 );
and ( n35628 , n35627 , n33208 );
not ( n35629 , n32968 );
not ( n35630 , n33270 );
and ( n35631 , n33274 , n33363 );
xor ( n35632 , n35630 , n35631 );
buf ( n35633 , n33270 );
and ( n35634 , n35632 , n35633 );
buf ( n35635 , n35634 );
and ( n35636 , n35629 , n35635 );
and ( n35637 , n35592 , n32968 );
or ( n35638 , n35636 , n35637 );
and ( n35639 , n35638 , n33370 );
and ( n35640 , n35592 , n33382 );
or ( n35641 , C0 , n35590 , n35628 , n35639 , C0 , n35640 );
buf ( n35642 , n35641 );
buf ( n35643 , n35642 );
buf ( n35644 , n30987 );
buf ( n35645 , n31655 );
not ( n35646 , n31728 );
and ( n35647 , n35646 , n32458 );
xor ( n35648 , n31749 , n31823 );
xor ( n35649 , n35648 , n32087 );
and ( n35650 , n35649 , n31728 );
or ( n35651 , n35647 , n35650 );
and ( n35652 , n35651 , n32253 );
not ( n35653 , n32283 );
and ( n35654 , n35653 , n32458 );
not ( n35655 , n31823 );
xor ( n35656 , n32294 , n31823 );
xor ( n35657 , n35656 , n32326 );
and ( n35658 , n35655 , n35657 );
xor ( n35659 , n32340 , n32342 );
xor ( n35660 , n35659 , n32389 );
and ( n35661 , n35660 , n31823 );
or ( n35662 , n35658 , n35661 );
and ( n35663 , n35662 , n32283 );
or ( n35664 , n35654 , n35663 );
and ( n35665 , n35664 , n32398 );
and ( n35666 , n32458 , n32436 );
or ( n35667 , n35652 , n35665 , n35666 );
and ( n35668 , n35667 , n32456 );
xor ( n35669 , n32458 , n32469 );
and ( n35670 , n35669 , n32473 );
not ( n35671 , n32475 );
and ( n35672 , n35671 , n35669 );
xor ( n35673 , n32458 , n32481 );
and ( n35674 , n35673 , n32475 );
or ( n35675 , n35672 , n35674 );
and ( n35676 , n35675 , n32486 );
buf ( n35677 , RI15b63d98_1272);
and ( n35678 , n35677 , n32489 );
and ( n35679 , n32458 , n32501 );
or ( n35680 , C0 , n35668 , n35670 , n35676 , n35678 , n35679 );
buf ( n35681 , n35680 );
buf ( n35682 , n35681 );
buf ( n35683 , n31655 );
not ( n35684 , n35375 );
and ( n35685 , n35684 , n31460 );
not ( n35686 , n31460 );
buf ( n35687 , RI15b575e8_846);
not ( n35688 , n35687 );
xor ( n35689 , n35686 , n35688 );
and ( n35690 , n35689 , n35375 );
or ( n35691 , n35685 , n35690 );
not ( n35692 , n35691 );
buf ( n35693 , n35692 );
buf ( n35694 , n35693 );
not ( n35695 , n35694 );
buf ( n35696 , n35695 );
buf ( n35697 , n35696 );
not ( n35698 , n35697 );
buf ( n35699 , n35698 );
not ( n35700 , n35699 );
not ( n35701 , n35375 );
not ( n35702 , n35387 );
not ( n35703 , n35388 );
not ( n35704 , n35389 );
not ( n35705 , n35390 );
not ( n35706 , n35391 );
not ( n35707 , n35392 );
not ( n35708 , n35393 );
not ( n35709 , n35394 );
not ( n35710 , n35395 );
not ( n35711 , n33972 );
not ( n35712 , n35396 );
not ( n35713 , n35397 );
not ( n35714 , n35398 );
not ( n35715 , n33986 );
not ( n35716 , n33999 );
not ( n35717 , n34000 );
not ( n35718 , n34001 );
not ( n35719 , n34002 );
not ( n35720 , n34003 );
not ( n35721 , n34004 );
not ( n35722 , n34005 );
not ( n35723 , n34006 );
not ( n35724 , n34007 );
not ( n35725 , n34008 );
not ( n35726 , n34009 );
not ( n35727 , n34010 );
not ( n35728 , n34011 );
not ( n35729 , n31079 );
not ( n35730 , n31459 );
and ( n35731 , n35686 , n35688 );
and ( n35732 , n35730 , n35731 );
and ( n35733 , n35729 , n35732 );
and ( n35734 , n35728 , n35733 );
and ( n35735 , n35727 , n35734 );
and ( n35736 , n35726 , n35735 );
and ( n35737 , n35725 , n35736 );
and ( n35738 , n35724 , n35737 );
and ( n35739 , n35723 , n35738 );
and ( n35740 , n35722 , n35739 );
and ( n35741 , n35721 , n35740 );
and ( n35742 , n35720 , n35741 );
and ( n35743 , n35719 , n35742 );
and ( n35744 , n35718 , n35743 );
and ( n35745 , n35717 , n35744 );
and ( n35746 , n35716 , n35745 );
and ( n35747 , n35715 , n35746 );
and ( n35748 , n35714 , n35747 );
and ( n35749 , n35713 , n35748 );
and ( n35750 , n35712 , n35749 );
and ( n35751 , n35711 , n35750 );
and ( n35752 , n35710 , n35751 );
and ( n35753 , n35709 , n35752 );
and ( n35754 , n35708 , n35753 );
and ( n35755 , n35707 , n35754 );
and ( n35756 , n35706 , n35755 );
and ( n35757 , n35705 , n35756 );
and ( n35758 , n35704 , n35757 );
and ( n35759 , n35703 , n35758 );
and ( n35760 , n35702 , n35759 );
xor ( n35761 , n35701 , n35760 );
buf ( n35762 , n35375 );
and ( n35763 , n35761 , n35762 );
buf ( n35764 , n35763 );
not ( n35765 , n35764 );
not ( n35766 , n35765 );
not ( n35767 , n35766 );
not ( n35768 , n35375 );
and ( n35769 , n35768 , n35387 );
xor ( n35770 , n35702 , n35759 );
and ( n35771 , n35770 , n35375 );
or ( n35772 , n35769 , n35771 );
not ( n35773 , n35772 );
buf ( n35774 , n35773 );
buf ( n35775 , n35774 );
not ( n35776 , n35775 );
not ( n35777 , n35776 );
not ( n35778 , n35375 );
and ( n35779 , n35778 , n35388 );
xor ( n35780 , n35703 , n35758 );
and ( n35781 , n35780 , n35375 );
or ( n35782 , n35779 , n35781 );
not ( n35783 , n35782 );
buf ( n35784 , n35783 );
buf ( n35785 , n35784 );
not ( n35786 , n35785 );
not ( n35787 , n35786 );
not ( n35788 , n35375 );
and ( n35789 , n35788 , n35389 );
xor ( n35790 , n35704 , n35757 );
and ( n35791 , n35790 , n35375 );
or ( n35792 , n35789 , n35791 );
not ( n35793 , n35792 );
buf ( n35794 , n35793 );
buf ( n35795 , n35794 );
not ( n35796 , n35795 );
not ( n35797 , n35796 );
not ( n35798 , n35375 );
and ( n35799 , n35798 , n35390 );
xor ( n35800 , n35705 , n35756 );
and ( n35801 , n35800 , n35375 );
or ( n35802 , n35799 , n35801 );
not ( n35803 , n35802 );
buf ( n35804 , n35803 );
buf ( n35805 , n35804 );
not ( n35806 , n35805 );
not ( n35807 , n35806 );
not ( n35808 , n35375 );
and ( n35809 , n35808 , n35391 );
xor ( n35810 , n35706 , n35755 );
and ( n35811 , n35810 , n35375 );
or ( n35812 , n35809 , n35811 );
not ( n35813 , n35812 );
buf ( n35814 , n35813 );
buf ( n35815 , n35814 );
not ( n35816 , n35815 );
not ( n35817 , n35816 );
not ( n35818 , n35375 );
and ( n35819 , n35818 , n35392 );
xor ( n35820 , n35707 , n35754 );
and ( n35821 , n35820 , n35375 );
or ( n35822 , n35819 , n35821 );
not ( n35823 , n35822 );
buf ( n35824 , n35823 );
buf ( n35825 , n35824 );
not ( n35826 , n35825 );
not ( n35827 , n35826 );
not ( n35828 , n35375 );
and ( n35829 , n35828 , n35393 );
xor ( n35830 , n35708 , n35753 );
and ( n35831 , n35830 , n35375 );
or ( n35832 , n35829 , n35831 );
not ( n35833 , n35832 );
buf ( n35834 , n35833 );
buf ( n35835 , n35834 );
not ( n35836 , n35835 );
not ( n35837 , n35836 );
not ( n35838 , n35375 );
and ( n35839 , n35838 , n35394 );
xor ( n35840 , n35709 , n35752 );
and ( n35841 , n35840 , n35375 );
or ( n35842 , n35839 , n35841 );
not ( n35843 , n35842 );
buf ( n35844 , n35843 );
buf ( n35845 , n35844 );
not ( n35846 , n35845 );
not ( n35847 , n35846 );
not ( n35848 , n35375 );
and ( n35849 , n35848 , n35395 );
xor ( n35850 , n35710 , n35751 );
and ( n35851 , n35850 , n35375 );
or ( n35852 , n35849 , n35851 );
not ( n35853 , n35852 );
buf ( n35854 , n35853 );
buf ( n35855 , n35854 );
not ( n35856 , n35855 );
not ( n35857 , n35856 );
not ( n35858 , n35375 );
and ( n35859 , n35858 , n33972 );
xor ( n35860 , n35711 , n35750 );
and ( n35861 , n35860 , n35375 );
or ( n35862 , n35859 , n35861 );
not ( n35863 , n35862 );
buf ( n35864 , n35863 );
buf ( n35865 , n35864 );
not ( n35866 , n35865 );
not ( n35867 , n35866 );
not ( n35868 , n35375 );
and ( n35869 , n35868 , n35396 );
xor ( n35870 , n35712 , n35749 );
and ( n35871 , n35870 , n35375 );
or ( n35872 , n35869 , n35871 );
not ( n35873 , n35872 );
buf ( n35874 , n35873 );
buf ( n35875 , n35874 );
not ( n35876 , n35875 );
not ( n35877 , n35876 );
not ( n35878 , n35375 );
and ( n35879 , n35878 , n35397 );
xor ( n35880 , n35713 , n35748 );
and ( n35881 , n35880 , n35375 );
or ( n35882 , n35879 , n35881 );
not ( n35883 , n35882 );
buf ( n35884 , n35883 );
buf ( n35885 , n35884 );
not ( n35886 , n35885 );
not ( n35887 , n35886 );
not ( n35888 , n35375 );
and ( n35889 , n35888 , n35398 );
xor ( n35890 , n35714 , n35747 );
and ( n35891 , n35890 , n35375 );
or ( n35892 , n35889 , n35891 );
not ( n35893 , n35892 );
buf ( n35894 , n35893 );
buf ( n35895 , n35894 );
not ( n35896 , n35895 );
not ( n35897 , n35896 );
not ( n35898 , n35375 );
and ( n35899 , n35898 , n33986 );
xor ( n35900 , n35715 , n35746 );
and ( n35901 , n35900 , n35375 );
or ( n35902 , n35899 , n35901 );
not ( n35903 , n35902 );
buf ( n35904 , n35903 );
buf ( n35905 , n35904 );
not ( n35906 , n35905 );
not ( n35907 , n35906 );
not ( n35908 , n35375 );
and ( n35909 , n35908 , n33999 );
xor ( n35910 , n35716 , n35745 );
and ( n35911 , n35910 , n35375 );
or ( n35912 , n35909 , n35911 );
not ( n35913 , n35912 );
buf ( n35914 , n35913 );
buf ( n35915 , n35914 );
not ( n35916 , n35915 );
not ( n35917 , n35916 );
not ( n35918 , n35375 );
and ( n35919 , n35918 , n34000 );
xor ( n35920 , n35717 , n35744 );
and ( n35921 , n35920 , n35375 );
or ( n35922 , n35919 , n35921 );
not ( n35923 , n35922 );
buf ( n35924 , n35923 );
buf ( n35925 , n35924 );
not ( n35926 , n35925 );
not ( n35927 , n35926 );
not ( n35928 , n35375 );
and ( n35929 , n35928 , n34001 );
xor ( n35930 , n35718 , n35743 );
and ( n35931 , n35930 , n35375 );
or ( n35932 , n35929 , n35931 );
not ( n35933 , n35932 );
buf ( n35934 , n35933 );
buf ( n35935 , n35934 );
not ( n35936 , n35935 );
not ( n35937 , n35936 );
not ( n35938 , n35375 );
and ( n35939 , n35938 , n34002 );
xor ( n35940 , n35719 , n35742 );
and ( n35941 , n35940 , n35375 );
or ( n35942 , n35939 , n35941 );
not ( n35943 , n35942 );
buf ( n35944 , n35943 );
buf ( n35945 , n35944 );
not ( n35946 , n35945 );
not ( n35947 , n35946 );
not ( n35948 , n35375 );
and ( n35949 , n35948 , n34003 );
xor ( n35950 , n35720 , n35741 );
and ( n35951 , n35950 , n35375 );
or ( n35952 , n35949 , n35951 );
not ( n35953 , n35952 );
buf ( n35954 , n35953 );
buf ( n35955 , n35954 );
not ( n35956 , n35955 );
not ( n35957 , n35956 );
not ( n35958 , n35375 );
and ( n35959 , n35958 , n34004 );
xor ( n35960 , n35721 , n35740 );
and ( n35961 , n35960 , n35375 );
or ( n35962 , n35959 , n35961 );
not ( n35963 , n35962 );
buf ( n35964 , n35963 );
buf ( n35965 , n35964 );
not ( n35966 , n35965 );
not ( n35967 , n35966 );
not ( n35968 , n35375 );
and ( n35969 , n35968 , n34005 );
xor ( n35970 , n35722 , n35739 );
and ( n35971 , n35970 , n35375 );
or ( n35972 , n35969 , n35971 );
not ( n35973 , n35972 );
buf ( n35974 , n35973 );
buf ( n35975 , n35974 );
not ( n35976 , n35975 );
not ( n35977 , n35976 );
not ( n35978 , n35375 );
and ( n35979 , n35978 , n34006 );
xor ( n35980 , n35723 , n35738 );
and ( n35981 , n35980 , n35375 );
or ( n35982 , n35979 , n35981 );
not ( n35983 , n35982 );
buf ( n35984 , n35983 );
buf ( n35985 , n35984 );
not ( n35986 , n35985 );
not ( n35987 , n35986 );
not ( n35988 , n35375 );
and ( n35989 , n35988 , n34007 );
xor ( n35990 , n35724 , n35737 );
and ( n35991 , n35990 , n35375 );
or ( n35992 , n35989 , n35991 );
not ( n35993 , n35992 );
buf ( n35994 , n35993 );
buf ( n35995 , n35994 );
not ( n35996 , n35995 );
not ( n35997 , n35996 );
not ( n35998 , n35375 );
and ( n35999 , n35998 , n34008 );
xor ( n36000 , n35725 , n35736 );
and ( n36001 , n36000 , n35375 );
or ( n36002 , n35999 , n36001 );
not ( n36003 , n36002 );
buf ( n36004 , n36003 );
buf ( n36005 , n36004 );
not ( n36006 , n36005 );
not ( n36007 , n36006 );
not ( n36008 , n35375 );
and ( n36009 , n36008 , n34009 );
xor ( n36010 , n35726 , n35735 );
and ( n36011 , n36010 , n35375 );
or ( n36012 , n36009 , n36011 );
not ( n36013 , n36012 );
buf ( n36014 , n36013 );
buf ( n36015 , n36014 );
not ( n36016 , n36015 );
not ( n36017 , n36016 );
not ( n36018 , n35375 );
and ( n36019 , n36018 , n34010 );
xor ( n36020 , n35727 , n35734 );
and ( n36021 , n36020 , n35375 );
or ( n36022 , n36019 , n36021 );
not ( n36023 , n36022 );
buf ( n36024 , n36023 );
buf ( n36025 , n36024 );
not ( n36026 , n36025 );
not ( n36027 , n36026 );
not ( n36028 , n35375 );
and ( n36029 , n36028 , n34011 );
xor ( n36030 , n35728 , n35733 );
and ( n36031 , n36030 , n35375 );
or ( n36032 , n36029 , n36031 );
not ( n36033 , n36032 );
buf ( n36034 , n36033 );
buf ( n36035 , n36034 );
not ( n36036 , n36035 );
not ( n36037 , n36036 );
not ( n36038 , n35375 );
and ( n36039 , n36038 , n31079 );
xor ( n36040 , n35729 , n35732 );
and ( n36041 , n36040 , n35375 );
or ( n36042 , n36039 , n36041 );
not ( n36043 , n36042 );
buf ( n36044 , n36043 );
buf ( n36045 , n36044 );
not ( n36046 , n36045 );
not ( n36047 , n36046 );
not ( n36048 , n35375 );
and ( n36049 , n36048 , n31459 );
xor ( n36050 , n35730 , n35731 );
and ( n36051 , n36050 , n35375 );
or ( n36052 , n36049 , n36051 );
not ( n36053 , n36052 );
buf ( n36054 , n36053 );
buf ( n36055 , n36054 );
not ( n36056 , n36055 );
not ( n36057 , n36056 );
not ( n36058 , n35695 );
and ( n36059 , n36057 , n36058 );
and ( n36060 , n36047 , n36059 );
and ( n36061 , n36037 , n36060 );
and ( n36062 , n36027 , n36061 );
and ( n36063 , n36017 , n36062 );
and ( n36064 , n36007 , n36063 );
and ( n36065 , n35997 , n36064 );
and ( n36066 , n35987 , n36065 );
and ( n36067 , n35977 , n36066 );
and ( n36068 , n35967 , n36067 );
and ( n36069 , n35957 , n36068 );
and ( n36070 , n35947 , n36069 );
and ( n36071 , n35937 , n36070 );
and ( n36072 , n35927 , n36071 );
and ( n36073 , n35917 , n36072 );
and ( n36074 , n35907 , n36073 );
and ( n36075 , n35897 , n36074 );
and ( n36076 , n35887 , n36075 );
and ( n36077 , n35877 , n36076 );
and ( n36078 , n35867 , n36077 );
and ( n36079 , n35857 , n36078 );
and ( n36080 , n35847 , n36079 );
and ( n36081 , n35837 , n36080 );
and ( n36082 , n35827 , n36081 );
and ( n36083 , n35817 , n36082 );
and ( n36084 , n35807 , n36083 );
and ( n36085 , n35797 , n36084 );
and ( n36086 , n35787 , n36085 );
and ( n36087 , n35777 , n36086 );
and ( n36088 , n35767 , n36087 );
not ( n36089 , n36088 );
and ( n36090 , n36089 , n35375 );
buf ( n36091 , n36090 );
not ( n36092 , n36091 );
not ( n36093 , n35375 );
and ( n36094 , n36093 , n36056 );
xor ( n36095 , n36057 , n36058 );
and ( n36096 , n36095 , n35375 );
or ( n36097 , n36094 , n36096 );
and ( n36098 , n36092 , n36097 );
not ( n36099 , n36097 );
not ( n36100 , n35696 );
xor ( n36101 , n36099 , n36100 );
and ( n36102 , n36101 , n36091 );
or ( n36103 , n36098 , n36102 );
not ( n36104 , n36103 );
buf ( n36105 , n36104 );
buf ( n36106 , n36105 );
not ( n36107 , n36106 );
or ( n36108 , n35700 , n36107 );
not ( n36109 , n36091 );
not ( n36110 , n35375 );
and ( n36111 , n36110 , n36046 );
xor ( n36112 , n36047 , n36059 );
and ( n36113 , n36112 , n35375 );
or ( n36114 , n36111 , n36113 );
and ( n36115 , n36109 , n36114 );
not ( n36116 , n36114 );
and ( n36117 , n36099 , n36100 );
xor ( n36118 , n36116 , n36117 );
and ( n36119 , n36118 , n36091 );
or ( n36120 , n36115 , n36119 );
not ( n36121 , n36120 );
buf ( n36122 , n36121 );
buf ( n36123 , n36122 );
not ( n36124 , n36123 );
or ( n36125 , n36108 , n36124 );
not ( n36126 , n36091 );
not ( n36127 , n35375 );
and ( n36128 , n36127 , n36036 );
xor ( n36129 , n36037 , n36060 );
and ( n36130 , n36129 , n35375 );
or ( n36131 , n36128 , n36130 );
and ( n36132 , n36126 , n36131 );
not ( n36133 , n36131 );
and ( n36134 , n36116 , n36117 );
xor ( n36135 , n36133 , n36134 );
and ( n36136 , n36135 , n36091 );
or ( n36137 , n36132 , n36136 );
not ( n36138 , n36137 );
buf ( n36139 , n36138 );
buf ( n36140 , n36139 );
not ( n36141 , n36140 );
or ( n36142 , n36125 , n36141 );
not ( n36143 , n36091 );
not ( n36144 , n35375 );
and ( n36145 , n36144 , n36026 );
xor ( n36146 , n36027 , n36061 );
and ( n36147 , n36146 , n35375 );
or ( n36148 , n36145 , n36147 );
and ( n36149 , n36143 , n36148 );
not ( n36150 , n36148 );
and ( n36151 , n36133 , n36134 );
xor ( n36152 , n36150 , n36151 );
and ( n36153 , n36152 , n36091 );
or ( n36154 , n36149 , n36153 );
not ( n36155 , n36154 );
buf ( n36156 , n36155 );
buf ( n36157 , n36156 );
not ( n36158 , n36157 );
or ( n36159 , n36142 , n36158 );
not ( n36160 , n36091 );
not ( n36161 , n35375 );
and ( n36162 , n36161 , n36016 );
xor ( n36163 , n36017 , n36062 );
and ( n36164 , n36163 , n35375 );
or ( n36165 , n36162 , n36164 );
and ( n36166 , n36160 , n36165 );
not ( n36167 , n36165 );
and ( n36168 , n36150 , n36151 );
xor ( n36169 , n36167 , n36168 );
and ( n36170 , n36169 , n36091 );
or ( n36171 , n36166 , n36170 );
not ( n36172 , n36171 );
buf ( n36173 , n36172 );
buf ( n36174 , n36173 );
not ( n36175 , n36174 );
or ( n36176 , n36159 , n36175 );
not ( n36177 , n36091 );
not ( n36178 , n35375 );
and ( n36179 , n36178 , n36006 );
xor ( n36180 , n36007 , n36063 );
and ( n36181 , n36180 , n35375 );
or ( n36182 , n36179 , n36181 );
and ( n36183 , n36177 , n36182 );
not ( n36184 , n36182 );
and ( n36185 , n36167 , n36168 );
xor ( n36186 , n36184 , n36185 );
and ( n36187 , n36186 , n36091 );
or ( n36188 , n36183 , n36187 );
not ( n36189 , n36188 );
buf ( n36190 , n36189 );
buf ( n36191 , n36190 );
not ( n36192 , n36191 );
or ( n36193 , n36176 , n36192 );
not ( n36194 , n36091 );
not ( n36195 , n35375 );
and ( n36196 , n36195 , n35996 );
xor ( n36197 , n35997 , n36064 );
and ( n36198 , n36197 , n35375 );
or ( n36199 , n36196 , n36198 );
and ( n36200 , n36194 , n36199 );
not ( n36201 , n36199 );
and ( n36202 , n36184 , n36185 );
xor ( n36203 , n36201 , n36202 );
and ( n36204 , n36203 , n36091 );
or ( n36205 , n36200 , n36204 );
not ( n36206 , n36205 );
buf ( n36207 , n36206 );
buf ( n36208 , n36207 );
not ( n36209 , n36208 );
or ( n36210 , n36193 , n36209 );
not ( n36211 , n36091 );
not ( n36212 , n35375 );
and ( n36213 , n36212 , n35986 );
xor ( n36214 , n35987 , n36065 );
and ( n36215 , n36214 , n35375 );
or ( n36216 , n36213 , n36215 );
and ( n36217 , n36211 , n36216 );
not ( n36218 , n36216 );
and ( n36219 , n36201 , n36202 );
xor ( n36220 , n36218 , n36219 );
and ( n36221 , n36220 , n36091 );
or ( n36222 , n36217 , n36221 );
not ( n36223 , n36222 );
buf ( n36224 , n36223 );
buf ( n36225 , n36224 );
not ( n36226 , n36225 );
or ( n36227 , n36210 , n36226 );
not ( n36228 , n36091 );
not ( n36229 , n35375 );
and ( n36230 , n36229 , n35976 );
xor ( n36231 , n35977 , n36066 );
and ( n36232 , n36231 , n35375 );
or ( n36233 , n36230 , n36232 );
and ( n36234 , n36228 , n36233 );
not ( n36235 , n36233 );
and ( n36236 , n36218 , n36219 );
xor ( n36237 , n36235 , n36236 );
and ( n36238 , n36237 , n36091 );
or ( n36239 , n36234 , n36238 );
not ( n36240 , n36239 );
buf ( n36241 , n36240 );
buf ( n36242 , n36241 );
not ( n36243 , n36242 );
or ( n36244 , n36227 , n36243 );
not ( n36245 , n36091 );
not ( n36246 , n35375 );
and ( n36247 , n36246 , n35966 );
xor ( n36248 , n35967 , n36067 );
and ( n36249 , n36248 , n35375 );
or ( n36250 , n36247 , n36249 );
and ( n36251 , n36245 , n36250 );
not ( n36252 , n36250 );
and ( n36253 , n36235 , n36236 );
xor ( n36254 , n36252 , n36253 );
and ( n36255 , n36254 , n36091 );
or ( n36256 , n36251 , n36255 );
not ( n36257 , n36256 );
buf ( n36258 , n36257 );
buf ( n36259 , n36258 );
not ( n36260 , n36259 );
or ( n36261 , n36244 , n36260 );
not ( n36262 , n36091 );
not ( n36263 , n35375 );
and ( n36264 , n36263 , n35956 );
xor ( n36265 , n35957 , n36068 );
and ( n36266 , n36265 , n35375 );
or ( n36267 , n36264 , n36266 );
and ( n36268 , n36262 , n36267 );
not ( n36269 , n36267 );
and ( n36270 , n36252 , n36253 );
xor ( n36271 , n36269 , n36270 );
and ( n36272 , n36271 , n36091 );
or ( n36273 , n36268 , n36272 );
not ( n36274 , n36273 );
buf ( n36275 , n36274 );
buf ( n36276 , n36275 );
not ( n36277 , n36276 );
or ( n36278 , n36261 , n36277 );
not ( n36279 , n36091 );
not ( n36280 , n35375 );
and ( n36281 , n36280 , n35946 );
xor ( n36282 , n35947 , n36069 );
and ( n36283 , n36282 , n35375 );
or ( n36284 , n36281 , n36283 );
and ( n36285 , n36279 , n36284 );
not ( n36286 , n36284 );
and ( n36287 , n36269 , n36270 );
xor ( n36288 , n36286 , n36287 );
and ( n36289 , n36288 , n36091 );
or ( n36290 , n36285 , n36289 );
not ( n36291 , n36290 );
buf ( n36292 , n36291 );
buf ( n36293 , n36292 );
not ( n36294 , n36293 );
or ( n36295 , n36278 , n36294 );
not ( n36296 , n36091 );
not ( n36297 , n35375 );
and ( n36298 , n36297 , n35936 );
xor ( n36299 , n35937 , n36070 );
and ( n36300 , n36299 , n35375 );
or ( n36301 , n36298 , n36300 );
and ( n36302 , n36296 , n36301 );
not ( n36303 , n36301 );
and ( n36304 , n36286 , n36287 );
xor ( n36305 , n36303 , n36304 );
and ( n36306 , n36305 , n36091 );
or ( n36307 , n36302 , n36306 );
not ( n36308 , n36307 );
buf ( n36309 , n36308 );
buf ( n36310 , n36309 );
not ( n36311 , n36310 );
or ( n36312 , n36295 , n36311 );
not ( n36313 , n36091 );
not ( n36314 , n35375 );
and ( n36315 , n36314 , n35926 );
xor ( n36316 , n35927 , n36071 );
and ( n36317 , n36316 , n35375 );
or ( n36318 , n36315 , n36317 );
and ( n36319 , n36313 , n36318 );
not ( n36320 , n36318 );
and ( n36321 , n36303 , n36304 );
xor ( n36322 , n36320 , n36321 );
and ( n36323 , n36322 , n36091 );
or ( n36324 , n36319 , n36323 );
not ( n36325 , n36324 );
buf ( n36326 , n36325 );
buf ( n36327 , n36326 );
not ( n36328 , n36327 );
or ( n36329 , n36312 , n36328 );
not ( n36330 , n36091 );
not ( n36331 , n35375 );
and ( n36332 , n36331 , n35916 );
xor ( n36333 , n35917 , n36072 );
and ( n36334 , n36333 , n35375 );
or ( n36335 , n36332 , n36334 );
and ( n36336 , n36330 , n36335 );
not ( n36337 , n36335 );
and ( n36338 , n36320 , n36321 );
xor ( n36339 , n36337 , n36338 );
and ( n36340 , n36339 , n36091 );
or ( n36341 , n36336 , n36340 );
not ( n36342 , n36341 );
buf ( n36343 , n36342 );
buf ( n36344 , n36343 );
not ( n36345 , n36344 );
or ( n36346 , n36329 , n36345 );
not ( n36347 , n36091 );
not ( n36348 , n35375 );
and ( n36349 , n36348 , n35906 );
xor ( n36350 , n35907 , n36073 );
and ( n36351 , n36350 , n35375 );
or ( n36352 , n36349 , n36351 );
and ( n36353 , n36347 , n36352 );
not ( n36354 , n36352 );
and ( n36355 , n36337 , n36338 );
xor ( n36356 , n36354 , n36355 );
and ( n36357 , n36356 , n36091 );
or ( n36358 , n36353 , n36357 );
not ( n36359 , n36358 );
buf ( n36360 , n36359 );
buf ( n36361 , n36360 );
not ( n36362 , n36361 );
or ( n36363 , n36346 , n36362 );
not ( n36364 , n36091 );
not ( n36365 , n35375 );
and ( n36366 , n36365 , n35896 );
xor ( n36367 , n35897 , n36074 );
and ( n36368 , n36367 , n35375 );
or ( n36369 , n36366 , n36368 );
and ( n36370 , n36364 , n36369 );
not ( n36371 , n36369 );
and ( n36372 , n36354 , n36355 );
xor ( n36373 , n36371 , n36372 );
and ( n36374 , n36373 , n36091 );
or ( n36375 , n36370 , n36374 );
not ( n36376 , n36375 );
buf ( n36377 , n36376 );
buf ( n36378 , n36377 );
not ( n36379 , n36378 );
or ( n36380 , n36363 , n36379 );
not ( n36381 , n36091 );
not ( n36382 , n35375 );
and ( n36383 , n36382 , n35886 );
xor ( n36384 , n35887 , n36075 );
and ( n36385 , n36384 , n35375 );
or ( n36386 , n36383 , n36385 );
and ( n36387 , n36381 , n36386 );
not ( n36388 , n36386 );
and ( n36389 , n36371 , n36372 );
xor ( n36390 , n36388 , n36389 );
and ( n36391 , n36390 , n36091 );
or ( n36392 , n36387 , n36391 );
not ( n36393 , n36392 );
buf ( n36394 , n36393 );
buf ( n36395 , n36394 );
not ( n36396 , n36395 );
or ( n36397 , n36380 , n36396 );
not ( n36398 , n36091 );
not ( n36399 , n35375 );
and ( n36400 , n36399 , n35876 );
xor ( n36401 , n35877 , n36076 );
and ( n36402 , n36401 , n35375 );
or ( n36403 , n36400 , n36402 );
and ( n36404 , n36398 , n36403 );
not ( n36405 , n36403 );
and ( n36406 , n36388 , n36389 );
xor ( n36407 , n36405 , n36406 );
and ( n36408 , n36407 , n36091 );
or ( n36409 , n36404 , n36408 );
not ( n36410 , n36409 );
buf ( n36411 , n36410 );
buf ( n36412 , n36411 );
not ( n36413 , n36412 );
or ( n36414 , n36397 , n36413 );
not ( n36415 , n36091 );
not ( n36416 , n35375 );
and ( n36417 , n36416 , n35866 );
xor ( n36418 , n35867 , n36077 );
and ( n36419 , n36418 , n35375 );
or ( n36420 , n36417 , n36419 );
and ( n36421 , n36415 , n36420 );
not ( n36422 , n36420 );
and ( n36423 , n36405 , n36406 );
xor ( n36424 , n36422 , n36423 );
and ( n36425 , n36424 , n36091 );
or ( n36426 , n36421 , n36425 );
not ( n36427 , n36426 );
buf ( n36428 , n36427 );
buf ( n36429 , n36428 );
not ( n36430 , n36429 );
or ( n36431 , n36414 , n36430 );
not ( n36432 , n36091 );
not ( n36433 , n35375 );
and ( n36434 , n36433 , n35856 );
xor ( n36435 , n35857 , n36078 );
and ( n36436 , n36435 , n35375 );
or ( n36437 , n36434 , n36436 );
and ( n36438 , n36432 , n36437 );
not ( n36439 , n36437 );
and ( n36440 , n36422 , n36423 );
xor ( n36441 , n36439 , n36440 );
and ( n36442 , n36441 , n36091 );
or ( n36443 , n36438 , n36442 );
not ( n36444 , n36443 );
buf ( n36445 , n36444 );
buf ( n36446 , n36445 );
not ( n36447 , n36446 );
or ( n36448 , n36431 , n36447 );
not ( n36449 , n36091 );
not ( n36450 , n35375 );
and ( n36451 , n36450 , n35846 );
xor ( n36452 , n35847 , n36079 );
and ( n36453 , n36452 , n35375 );
or ( n36454 , n36451 , n36453 );
and ( n36455 , n36449 , n36454 );
not ( n36456 , n36454 );
and ( n36457 , n36439 , n36440 );
xor ( n36458 , n36456 , n36457 );
and ( n36459 , n36458 , n36091 );
or ( n36460 , n36455 , n36459 );
not ( n36461 , n36460 );
buf ( n36462 , n36461 );
buf ( n36463 , n36462 );
not ( n36464 , n36463 );
or ( n36465 , n36448 , n36464 );
not ( n36466 , n36091 );
not ( n36467 , n35375 );
and ( n36468 , n36467 , n35836 );
xor ( n36469 , n35837 , n36080 );
and ( n36470 , n36469 , n35375 );
or ( n36471 , n36468 , n36470 );
and ( n36472 , n36466 , n36471 );
not ( n36473 , n36471 );
and ( n36474 , n36456 , n36457 );
xor ( n36475 , n36473 , n36474 );
and ( n36476 , n36475 , n36091 );
or ( n36477 , n36472 , n36476 );
not ( n36478 , n36477 );
buf ( n36479 , n36478 );
buf ( n36480 , n36479 );
not ( n36481 , n36480 );
or ( n36482 , n36465 , n36481 );
not ( n36483 , n36091 );
not ( n36484 , n35375 );
and ( n36485 , n36484 , n35826 );
xor ( n36486 , n35827 , n36081 );
and ( n36487 , n36486 , n35375 );
or ( n36488 , n36485 , n36487 );
and ( n36489 , n36483 , n36488 );
not ( n36490 , n36488 );
and ( n36491 , n36473 , n36474 );
xor ( n36492 , n36490 , n36491 );
and ( n36493 , n36492 , n36091 );
or ( n36494 , n36489 , n36493 );
not ( n36495 , n36494 );
buf ( n36496 , n36495 );
buf ( n36497 , n36496 );
not ( n36498 , n36497 );
or ( n36499 , n36482 , n36498 );
not ( n36500 , n36091 );
not ( n36501 , n35375 );
and ( n36502 , n36501 , n35816 );
xor ( n36503 , n35817 , n36082 );
and ( n36504 , n36503 , n35375 );
or ( n36505 , n36502 , n36504 );
and ( n36506 , n36500 , n36505 );
not ( n36507 , n36505 );
and ( n36508 , n36490 , n36491 );
xor ( n36509 , n36507 , n36508 );
and ( n36510 , n36509 , n36091 );
or ( n36511 , n36506 , n36510 );
not ( n36512 , n36511 );
buf ( n36513 , n36512 );
buf ( n36514 , n36513 );
not ( n36515 , n36514 );
or ( n36516 , n36499 , n36515 );
not ( n36517 , n36091 );
not ( n36518 , n35375 );
and ( n36519 , n36518 , n35806 );
xor ( n36520 , n35807 , n36083 );
and ( n36521 , n36520 , n35375 );
or ( n36522 , n36519 , n36521 );
and ( n36523 , n36517 , n36522 );
not ( n36524 , n36522 );
and ( n36525 , n36507 , n36508 );
xor ( n36526 , n36524 , n36525 );
and ( n36527 , n36526 , n36091 );
or ( n36528 , n36523 , n36527 );
not ( n36529 , n36528 );
buf ( n36530 , n36529 );
buf ( n36531 , n36530 );
not ( n36532 , n36531 );
or ( n36533 , n36516 , n36532 );
not ( n36534 , n36091 );
not ( n36535 , n35375 );
and ( n36536 , n36535 , n35796 );
xor ( n36537 , n35797 , n36084 );
and ( n36538 , n36537 , n35375 );
or ( n36539 , n36536 , n36538 );
and ( n36540 , n36534 , n36539 );
not ( n36541 , n36539 );
and ( n36542 , n36524 , n36525 );
xor ( n36543 , n36541 , n36542 );
and ( n36544 , n36543 , n36091 );
or ( n36545 , n36540 , n36544 );
not ( n36546 , n36545 );
buf ( n36547 , n36546 );
buf ( n36548 , n36547 );
not ( n36549 , n36548 );
or ( n36550 , n36533 , n36549 );
not ( n36551 , n36091 );
not ( n36552 , n35375 );
and ( n36553 , n36552 , n35786 );
xor ( n36554 , n35787 , n36085 );
and ( n36555 , n36554 , n35375 );
or ( n36556 , n36553 , n36555 );
and ( n36557 , n36551 , n36556 );
not ( n36558 , n36556 );
and ( n36559 , n36541 , n36542 );
xor ( n36560 , n36558 , n36559 );
and ( n36561 , n36560 , n36091 );
or ( n36562 , n36557 , n36561 );
not ( n36563 , n36562 );
buf ( n36564 , n36563 );
buf ( n36565 , n36564 );
not ( n36566 , n36565 );
or ( n36567 , n36550 , n36566 );
not ( n36568 , n36091 );
not ( n36569 , n35375 );
and ( n36570 , n36569 , n35776 );
xor ( n36571 , n35777 , n36086 );
and ( n36572 , n36571 , n35375 );
or ( n36573 , n36570 , n36572 );
and ( n36574 , n36568 , n36573 );
not ( n36575 , n36573 );
and ( n36576 , n36558 , n36559 );
xor ( n36577 , n36575 , n36576 );
and ( n36578 , n36577 , n36091 );
or ( n36579 , n36574 , n36578 );
not ( n36580 , n36579 );
buf ( n36581 , n36580 );
buf ( n36582 , n36581 );
not ( n36583 , n36582 );
or ( n36584 , n36567 , n36583 );
buf ( n36585 , n36584 );
buf ( n36586 , n36585 );
and ( n36587 , n36586 , n36091 );
not ( n36588 , n36587 );
and ( n36589 , n36588 , n36107 );
xor ( n36590 , n36107 , n36091 );
xor ( n36591 , n35700 , n36091 );
and ( n36592 , n36591 , n36091 );
xor ( n36593 , n36590 , n36592 );
and ( n36594 , n36593 , n36587 );
or ( n36595 , n36589 , n36594 );
and ( n36596 , n31445 , n31441 , n31443 );
and ( n36597 , n36595 , n36596 );
not ( n36598 , n35375 );
and ( n36599 , n36598 , n31459 );
not ( n36600 , n31459 );
not ( n36601 , n31460 );
not ( n36602 , n35687 );
and ( n36603 , n36601 , n36602 );
xor ( n36604 , n36600 , n36603 );
and ( n36605 , n36604 , n35375 );
or ( n36606 , n36599 , n36605 );
not ( n36607 , n36606 );
buf ( n36608 , n36607 );
buf ( n36609 , n36608 );
not ( n36610 , n36609 );
buf ( n36611 , n36610 );
buf ( n36612 , n36611 );
not ( n36613 , n36612 );
buf ( n36614 , n36613 );
not ( n36615 , n36614 );
not ( n36616 , n35375 );
not ( n36617 , n35387 );
not ( n36618 , n35388 );
not ( n36619 , n35389 );
not ( n36620 , n35390 );
not ( n36621 , n35391 );
not ( n36622 , n35392 );
not ( n36623 , n35393 );
not ( n36624 , n35394 );
not ( n36625 , n35395 );
not ( n36626 , n33972 );
not ( n36627 , n35396 );
not ( n36628 , n35397 );
not ( n36629 , n35398 );
not ( n36630 , n33986 );
not ( n36631 , n33999 );
not ( n36632 , n34000 );
not ( n36633 , n34001 );
not ( n36634 , n34002 );
not ( n36635 , n34003 );
not ( n36636 , n34004 );
not ( n36637 , n34005 );
not ( n36638 , n34006 );
not ( n36639 , n34007 );
not ( n36640 , n34008 );
not ( n36641 , n34009 );
not ( n36642 , n34010 );
not ( n36643 , n34011 );
not ( n36644 , n31079 );
and ( n36645 , n36600 , n36603 );
and ( n36646 , n36644 , n36645 );
and ( n36647 , n36643 , n36646 );
and ( n36648 , n36642 , n36647 );
and ( n36649 , n36641 , n36648 );
and ( n36650 , n36640 , n36649 );
and ( n36651 , n36639 , n36650 );
and ( n36652 , n36638 , n36651 );
and ( n36653 , n36637 , n36652 );
and ( n36654 , n36636 , n36653 );
and ( n36655 , n36635 , n36654 );
and ( n36656 , n36634 , n36655 );
and ( n36657 , n36633 , n36656 );
and ( n36658 , n36632 , n36657 );
and ( n36659 , n36631 , n36658 );
and ( n36660 , n36630 , n36659 );
and ( n36661 , n36629 , n36660 );
and ( n36662 , n36628 , n36661 );
and ( n36663 , n36627 , n36662 );
and ( n36664 , n36626 , n36663 );
and ( n36665 , n36625 , n36664 );
and ( n36666 , n36624 , n36665 );
and ( n36667 , n36623 , n36666 );
and ( n36668 , n36622 , n36667 );
and ( n36669 , n36621 , n36668 );
and ( n36670 , n36620 , n36669 );
and ( n36671 , n36619 , n36670 );
and ( n36672 , n36618 , n36671 );
and ( n36673 , n36617 , n36672 );
xor ( n36674 , n36616 , n36673 );
buf ( n36675 , n35375 );
and ( n36676 , n36674 , n36675 );
buf ( n36677 , n36676 );
not ( n36678 , n36677 );
not ( n36679 , n36678 );
not ( n36680 , n36679 );
not ( n36681 , n35375 );
and ( n36682 , n36681 , n35387 );
xor ( n36683 , n36617 , n36672 );
and ( n36684 , n36683 , n35375 );
or ( n36685 , n36682 , n36684 );
not ( n36686 , n36685 );
buf ( n36687 , n36686 );
buf ( n36688 , n36687 );
not ( n36689 , n36688 );
not ( n36690 , n36689 );
not ( n36691 , n35375 );
and ( n36692 , n36691 , n35388 );
xor ( n36693 , n36618 , n36671 );
and ( n36694 , n36693 , n35375 );
or ( n36695 , n36692 , n36694 );
not ( n36696 , n36695 );
buf ( n36697 , n36696 );
buf ( n36698 , n36697 );
not ( n36699 , n36698 );
not ( n36700 , n36699 );
not ( n36701 , n35375 );
and ( n36702 , n36701 , n35389 );
xor ( n36703 , n36619 , n36670 );
and ( n36704 , n36703 , n35375 );
or ( n36705 , n36702 , n36704 );
not ( n36706 , n36705 );
buf ( n36707 , n36706 );
buf ( n36708 , n36707 );
not ( n36709 , n36708 );
not ( n36710 , n36709 );
not ( n36711 , n35375 );
and ( n36712 , n36711 , n35390 );
xor ( n36713 , n36620 , n36669 );
and ( n36714 , n36713 , n35375 );
or ( n36715 , n36712 , n36714 );
not ( n36716 , n36715 );
buf ( n36717 , n36716 );
buf ( n36718 , n36717 );
not ( n36719 , n36718 );
not ( n36720 , n36719 );
not ( n36721 , n35375 );
and ( n36722 , n36721 , n35391 );
xor ( n36723 , n36621 , n36668 );
and ( n36724 , n36723 , n35375 );
or ( n36725 , n36722 , n36724 );
not ( n36726 , n36725 );
buf ( n36727 , n36726 );
buf ( n36728 , n36727 );
not ( n36729 , n36728 );
not ( n36730 , n36729 );
not ( n36731 , n35375 );
and ( n36732 , n36731 , n35392 );
xor ( n36733 , n36622 , n36667 );
and ( n36734 , n36733 , n35375 );
or ( n36735 , n36732 , n36734 );
not ( n36736 , n36735 );
buf ( n36737 , n36736 );
buf ( n36738 , n36737 );
not ( n36739 , n36738 );
not ( n36740 , n36739 );
not ( n36741 , n35375 );
and ( n36742 , n36741 , n35393 );
xor ( n36743 , n36623 , n36666 );
and ( n36744 , n36743 , n35375 );
or ( n36745 , n36742 , n36744 );
not ( n36746 , n36745 );
buf ( n36747 , n36746 );
buf ( n36748 , n36747 );
not ( n36749 , n36748 );
not ( n36750 , n36749 );
not ( n36751 , n35375 );
and ( n36752 , n36751 , n35394 );
xor ( n36753 , n36624 , n36665 );
and ( n36754 , n36753 , n35375 );
or ( n36755 , n36752 , n36754 );
not ( n36756 , n36755 );
buf ( n36757 , n36756 );
buf ( n36758 , n36757 );
not ( n36759 , n36758 );
not ( n36760 , n36759 );
not ( n36761 , n35375 );
and ( n36762 , n36761 , n35395 );
xor ( n36763 , n36625 , n36664 );
and ( n36764 , n36763 , n35375 );
or ( n36765 , n36762 , n36764 );
not ( n36766 , n36765 );
buf ( n36767 , n36766 );
buf ( n36768 , n36767 );
not ( n36769 , n36768 );
not ( n36770 , n36769 );
not ( n36771 , n35375 );
and ( n36772 , n36771 , n33972 );
xor ( n36773 , n36626 , n36663 );
and ( n36774 , n36773 , n35375 );
or ( n36775 , n36772 , n36774 );
not ( n36776 , n36775 );
buf ( n36777 , n36776 );
buf ( n36778 , n36777 );
not ( n36779 , n36778 );
not ( n36780 , n36779 );
not ( n36781 , n35375 );
and ( n36782 , n36781 , n35396 );
xor ( n36783 , n36627 , n36662 );
and ( n36784 , n36783 , n35375 );
or ( n36785 , n36782 , n36784 );
not ( n36786 , n36785 );
buf ( n36787 , n36786 );
buf ( n36788 , n36787 );
not ( n36789 , n36788 );
not ( n36790 , n36789 );
not ( n36791 , n35375 );
and ( n36792 , n36791 , n35397 );
xor ( n36793 , n36628 , n36661 );
and ( n36794 , n36793 , n35375 );
or ( n36795 , n36792 , n36794 );
not ( n36796 , n36795 );
buf ( n36797 , n36796 );
buf ( n36798 , n36797 );
not ( n36799 , n36798 );
not ( n36800 , n36799 );
not ( n36801 , n35375 );
and ( n36802 , n36801 , n35398 );
xor ( n36803 , n36629 , n36660 );
and ( n36804 , n36803 , n35375 );
or ( n36805 , n36802 , n36804 );
not ( n36806 , n36805 );
buf ( n36807 , n36806 );
buf ( n36808 , n36807 );
not ( n36809 , n36808 );
not ( n36810 , n36809 );
not ( n36811 , n35375 );
and ( n36812 , n36811 , n33986 );
xor ( n36813 , n36630 , n36659 );
and ( n36814 , n36813 , n35375 );
or ( n36815 , n36812 , n36814 );
not ( n36816 , n36815 );
buf ( n36817 , n36816 );
buf ( n36818 , n36817 );
not ( n36819 , n36818 );
not ( n36820 , n36819 );
not ( n36821 , n35375 );
and ( n36822 , n36821 , n33999 );
xor ( n36823 , n36631 , n36658 );
and ( n36824 , n36823 , n35375 );
or ( n36825 , n36822 , n36824 );
not ( n36826 , n36825 );
buf ( n36827 , n36826 );
buf ( n36828 , n36827 );
not ( n36829 , n36828 );
not ( n36830 , n36829 );
not ( n36831 , n35375 );
and ( n36832 , n36831 , n34000 );
xor ( n36833 , n36632 , n36657 );
and ( n36834 , n36833 , n35375 );
or ( n36835 , n36832 , n36834 );
not ( n36836 , n36835 );
buf ( n36837 , n36836 );
buf ( n36838 , n36837 );
not ( n36839 , n36838 );
not ( n36840 , n36839 );
not ( n36841 , n35375 );
and ( n36842 , n36841 , n34001 );
xor ( n36843 , n36633 , n36656 );
and ( n36844 , n36843 , n35375 );
or ( n36845 , n36842 , n36844 );
not ( n36846 , n36845 );
buf ( n36847 , n36846 );
buf ( n36848 , n36847 );
not ( n36849 , n36848 );
not ( n36850 , n36849 );
not ( n36851 , n35375 );
and ( n36852 , n36851 , n34002 );
xor ( n36853 , n36634 , n36655 );
and ( n36854 , n36853 , n35375 );
or ( n36855 , n36852 , n36854 );
not ( n36856 , n36855 );
buf ( n36857 , n36856 );
buf ( n36858 , n36857 );
not ( n36859 , n36858 );
not ( n36860 , n36859 );
not ( n36861 , n35375 );
and ( n36862 , n36861 , n34003 );
xor ( n36863 , n36635 , n36654 );
and ( n36864 , n36863 , n35375 );
or ( n36865 , n36862 , n36864 );
not ( n36866 , n36865 );
buf ( n36867 , n36866 );
buf ( n36868 , n36867 );
not ( n36869 , n36868 );
not ( n36870 , n36869 );
not ( n36871 , n35375 );
and ( n36872 , n36871 , n34004 );
xor ( n36873 , n36636 , n36653 );
and ( n36874 , n36873 , n35375 );
or ( n36875 , n36872 , n36874 );
not ( n36876 , n36875 );
buf ( n36877 , n36876 );
buf ( n36878 , n36877 );
not ( n36879 , n36878 );
not ( n36880 , n36879 );
not ( n36881 , n35375 );
and ( n36882 , n36881 , n34005 );
xor ( n36883 , n36637 , n36652 );
and ( n36884 , n36883 , n35375 );
or ( n36885 , n36882 , n36884 );
not ( n36886 , n36885 );
buf ( n36887 , n36886 );
buf ( n36888 , n36887 );
not ( n36889 , n36888 );
not ( n36890 , n36889 );
not ( n36891 , n35375 );
and ( n36892 , n36891 , n34006 );
xor ( n36893 , n36638 , n36651 );
and ( n36894 , n36893 , n35375 );
or ( n36895 , n36892 , n36894 );
not ( n36896 , n36895 );
buf ( n36897 , n36896 );
buf ( n36898 , n36897 );
not ( n36899 , n36898 );
not ( n36900 , n36899 );
not ( n36901 , n35375 );
and ( n36902 , n36901 , n34007 );
xor ( n36903 , n36639 , n36650 );
and ( n36904 , n36903 , n35375 );
or ( n36905 , n36902 , n36904 );
not ( n36906 , n36905 );
buf ( n36907 , n36906 );
buf ( n36908 , n36907 );
not ( n36909 , n36908 );
not ( n36910 , n36909 );
not ( n36911 , n35375 );
and ( n36912 , n36911 , n34008 );
xor ( n36913 , n36640 , n36649 );
and ( n36914 , n36913 , n35375 );
or ( n36915 , n36912 , n36914 );
not ( n36916 , n36915 );
buf ( n36917 , n36916 );
buf ( n36918 , n36917 );
not ( n36919 , n36918 );
not ( n36920 , n36919 );
not ( n36921 , n35375 );
and ( n36922 , n36921 , n34009 );
xor ( n36923 , n36641 , n36648 );
and ( n36924 , n36923 , n35375 );
or ( n36925 , n36922 , n36924 );
not ( n36926 , n36925 );
buf ( n36927 , n36926 );
buf ( n36928 , n36927 );
not ( n36929 , n36928 );
not ( n36930 , n36929 );
not ( n36931 , n35375 );
and ( n36932 , n36931 , n34010 );
xor ( n36933 , n36642 , n36647 );
and ( n36934 , n36933 , n35375 );
or ( n36935 , n36932 , n36934 );
not ( n36936 , n36935 );
buf ( n36937 , n36936 );
buf ( n36938 , n36937 );
not ( n36939 , n36938 );
not ( n36940 , n36939 );
not ( n36941 , n35375 );
and ( n36942 , n36941 , n34011 );
xor ( n36943 , n36643 , n36646 );
and ( n36944 , n36943 , n35375 );
or ( n36945 , n36942 , n36944 );
not ( n36946 , n36945 );
buf ( n36947 , n36946 );
buf ( n36948 , n36947 );
not ( n36949 , n36948 );
not ( n36950 , n36949 );
not ( n36951 , n35375 );
and ( n36952 , n36951 , n31079 );
xor ( n36953 , n36644 , n36645 );
and ( n36954 , n36953 , n35375 );
or ( n36955 , n36952 , n36954 );
not ( n36956 , n36955 );
buf ( n36957 , n36956 );
buf ( n36958 , n36957 );
not ( n36959 , n36958 );
not ( n36960 , n36959 );
not ( n36961 , n36610 );
and ( n36962 , n36960 , n36961 );
and ( n36963 , n36950 , n36962 );
and ( n36964 , n36940 , n36963 );
and ( n36965 , n36930 , n36964 );
and ( n36966 , n36920 , n36965 );
and ( n36967 , n36910 , n36966 );
and ( n36968 , n36900 , n36967 );
and ( n36969 , n36890 , n36968 );
and ( n36970 , n36880 , n36969 );
and ( n36971 , n36870 , n36970 );
and ( n36972 , n36860 , n36971 );
and ( n36973 , n36850 , n36972 );
and ( n36974 , n36840 , n36973 );
and ( n36975 , n36830 , n36974 );
and ( n36976 , n36820 , n36975 );
and ( n36977 , n36810 , n36976 );
and ( n36978 , n36800 , n36977 );
and ( n36979 , n36790 , n36978 );
and ( n36980 , n36780 , n36979 );
and ( n36981 , n36770 , n36980 );
and ( n36982 , n36760 , n36981 );
and ( n36983 , n36750 , n36982 );
and ( n36984 , n36740 , n36983 );
and ( n36985 , n36730 , n36984 );
and ( n36986 , n36720 , n36985 );
and ( n36987 , n36710 , n36986 );
and ( n36988 , n36700 , n36987 );
and ( n36989 , n36690 , n36988 );
and ( n36990 , n36680 , n36989 );
not ( n36991 , n36990 );
and ( n36992 , n36991 , n35375 );
buf ( n36993 , n36992 );
not ( n36994 , n36993 );
not ( n36995 , n35375 );
and ( n36996 , n36995 , n36959 );
xor ( n36997 , n36960 , n36961 );
and ( n36998 , n36997 , n35375 );
or ( n36999 , n36996 , n36998 );
and ( n37000 , n36994 , n36999 );
not ( n37001 , n36999 );
not ( n37002 , n36611 );
xor ( n37003 , n37001 , n37002 );
and ( n37004 , n37003 , n36993 );
or ( n37005 , n37000 , n37004 );
not ( n37006 , n37005 );
buf ( n37007 , n37006 );
buf ( n37008 , n37007 );
not ( n37009 , n37008 );
or ( n37010 , n36615 , n37009 );
not ( n37011 , n36993 );
not ( n37012 , n35375 );
and ( n37013 , n37012 , n36949 );
xor ( n37014 , n36950 , n36962 );
and ( n37015 , n37014 , n35375 );
or ( n37016 , n37013 , n37015 );
and ( n37017 , n37011 , n37016 );
not ( n37018 , n37016 );
and ( n37019 , n37001 , n37002 );
xor ( n37020 , n37018 , n37019 );
and ( n37021 , n37020 , n36993 );
or ( n37022 , n37017 , n37021 );
not ( n37023 , n37022 );
buf ( n37024 , n37023 );
buf ( n37025 , n37024 );
not ( n37026 , n37025 );
or ( n37027 , n37010 , n37026 );
not ( n37028 , n36993 );
not ( n37029 , n35375 );
and ( n37030 , n37029 , n36939 );
xor ( n37031 , n36940 , n36963 );
and ( n37032 , n37031 , n35375 );
or ( n37033 , n37030 , n37032 );
and ( n37034 , n37028 , n37033 );
not ( n37035 , n37033 );
and ( n37036 , n37018 , n37019 );
xor ( n37037 , n37035 , n37036 );
and ( n37038 , n37037 , n36993 );
or ( n37039 , n37034 , n37038 );
not ( n37040 , n37039 );
buf ( n37041 , n37040 );
buf ( n37042 , n37041 );
not ( n37043 , n37042 );
or ( n37044 , n37027 , n37043 );
not ( n37045 , n36993 );
not ( n37046 , n35375 );
and ( n37047 , n37046 , n36929 );
xor ( n37048 , n36930 , n36964 );
and ( n37049 , n37048 , n35375 );
or ( n37050 , n37047 , n37049 );
and ( n37051 , n37045 , n37050 );
not ( n37052 , n37050 );
and ( n37053 , n37035 , n37036 );
xor ( n37054 , n37052 , n37053 );
and ( n37055 , n37054 , n36993 );
or ( n37056 , n37051 , n37055 );
not ( n37057 , n37056 );
buf ( n37058 , n37057 );
buf ( n37059 , n37058 );
not ( n37060 , n37059 );
or ( n37061 , n37044 , n37060 );
not ( n37062 , n36993 );
not ( n37063 , n35375 );
and ( n37064 , n37063 , n36919 );
xor ( n37065 , n36920 , n36965 );
and ( n37066 , n37065 , n35375 );
or ( n37067 , n37064 , n37066 );
and ( n37068 , n37062 , n37067 );
not ( n37069 , n37067 );
and ( n37070 , n37052 , n37053 );
xor ( n37071 , n37069 , n37070 );
and ( n37072 , n37071 , n36993 );
or ( n37073 , n37068 , n37072 );
not ( n37074 , n37073 );
buf ( n37075 , n37074 );
buf ( n37076 , n37075 );
not ( n37077 , n37076 );
or ( n37078 , n37061 , n37077 );
not ( n37079 , n36993 );
not ( n37080 , n35375 );
and ( n37081 , n37080 , n36909 );
xor ( n37082 , n36910 , n36966 );
and ( n37083 , n37082 , n35375 );
or ( n37084 , n37081 , n37083 );
and ( n37085 , n37079 , n37084 );
not ( n37086 , n37084 );
and ( n37087 , n37069 , n37070 );
xor ( n37088 , n37086 , n37087 );
and ( n37089 , n37088 , n36993 );
or ( n37090 , n37085 , n37089 );
not ( n37091 , n37090 );
buf ( n37092 , n37091 );
buf ( n37093 , n37092 );
not ( n37094 , n37093 );
or ( n37095 , n37078 , n37094 );
not ( n37096 , n36993 );
not ( n37097 , n35375 );
and ( n37098 , n37097 , n36899 );
xor ( n37099 , n36900 , n36967 );
and ( n37100 , n37099 , n35375 );
or ( n37101 , n37098 , n37100 );
and ( n37102 , n37096 , n37101 );
not ( n37103 , n37101 );
and ( n37104 , n37086 , n37087 );
xor ( n37105 , n37103 , n37104 );
and ( n37106 , n37105 , n36993 );
or ( n37107 , n37102 , n37106 );
not ( n37108 , n37107 );
buf ( n37109 , n37108 );
buf ( n37110 , n37109 );
not ( n37111 , n37110 );
or ( n37112 , n37095 , n37111 );
not ( n37113 , n36993 );
not ( n37114 , n35375 );
and ( n37115 , n37114 , n36889 );
xor ( n37116 , n36890 , n36968 );
and ( n37117 , n37116 , n35375 );
or ( n37118 , n37115 , n37117 );
and ( n37119 , n37113 , n37118 );
not ( n37120 , n37118 );
and ( n37121 , n37103 , n37104 );
xor ( n37122 , n37120 , n37121 );
and ( n37123 , n37122 , n36993 );
or ( n37124 , n37119 , n37123 );
not ( n37125 , n37124 );
buf ( n37126 , n37125 );
buf ( n37127 , n37126 );
not ( n37128 , n37127 );
or ( n37129 , n37112 , n37128 );
not ( n37130 , n36993 );
not ( n37131 , n35375 );
and ( n37132 , n37131 , n36879 );
xor ( n37133 , n36880 , n36969 );
and ( n37134 , n37133 , n35375 );
or ( n37135 , n37132 , n37134 );
and ( n37136 , n37130 , n37135 );
not ( n37137 , n37135 );
and ( n37138 , n37120 , n37121 );
xor ( n37139 , n37137 , n37138 );
and ( n37140 , n37139 , n36993 );
or ( n37141 , n37136 , n37140 );
not ( n37142 , n37141 );
buf ( n37143 , n37142 );
buf ( n37144 , n37143 );
not ( n37145 , n37144 );
or ( n37146 , n37129 , n37145 );
not ( n37147 , n36993 );
not ( n37148 , n35375 );
and ( n37149 , n37148 , n36869 );
xor ( n37150 , n36870 , n36970 );
and ( n37151 , n37150 , n35375 );
or ( n37152 , n37149 , n37151 );
and ( n37153 , n37147 , n37152 );
not ( n37154 , n37152 );
and ( n37155 , n37137 , n37138 );
xor ( n37156 , n37154 , n37155 );
and ( n37157 , n37156 , n36993 );
or ( n37158 , n37153 , n37157 );
not ( n37159 , n37158 );
buf ( n37160 , n37159 );
buf ( n37161 , n37160 );
not ( n37162 , n37161 );
or ( n37163 , n37146 , n37162 );
not ( n37164 , n36993 );
not ( n37165 , n35375 );
and ( n37166 , n37165 , n36859 );
xor ( n37167 , n36860 , n36971 );
and ( n37168 , n37167 , n35375 );
or ( n37169 , n37166 , n37168 );
and ( n37170 , n37164 , n37169 );
not ( n37171 , n37169 );
and ( n37172 , n37154 , n37155 );
xor ( n37173 , n37171 , n37172 );
and ( n37174 , n37173 , n36993 );
or ( n37175 , n37170 , n37174 );
not ( n37176 , n37175 );
buf ( n37177 , n37176 );
buf ( n37178 , n37177 );
not ( n37179 , n37178 );
or ( n37180 , n37163 , n37179 );
not ( n37181 , n36993 );
not ( n37182 , n35375 );
and ( n37183 , n37182 , n36849 );
xor ( n37184 , n36850 , n36972 );
and ( n37185 , n37184 , n35375 );
or ( n37186 , n37183 , n37185 );
and ( n37187 , n37181 , n37186 );
not ( n37188 , n37186 );
and ( n37189 , n37171 , n37172 );
xor ( n37190 , n37188 , n37189 );
and ( n37191 , n37190 , n36993 );
or ( n37192 , n37187 , n37191 );
not ( n37193 , n37192 );
buf ( n37194 , n37193 );
buf ( n37195 , n37194 );
not ( n37196 , n37195 );
or ( n37197 , n37180 , n37196 );
not ( n37198 , n36993 );
not ( n37199 , n35375 );
and ( n37200 , n37199 , n36839 );
xor ( n37201 , n36840 , n36973 );
and ( n37202 , n37201 , n35375 );
or ( n37203 , n37200 , n37202 );
and ( n37204 , n37198 , n37203 );
not ( n37205 , n37203 );
and ( n37206 , n37188 , n37189 );
xor ( n37207 , n37205 , n37206 );
and ( n37208 , n37207 , n36993 );
or ( n37209 , n37204 , n37208 );
not ( n37210 , n37209 );
buf ( n37211 , n37210 );
buf ( n37212 , n37211 );
not ( n37213 , n37212 );
or ( n37214 , n37197 , n37213 );
not ( n37215 , n36993 );
not ( n37216 , n35375 );
and ( n37217 , n37216 , n36829 );
xor ( n37218 , n36830 , n36974 );
and ( n37219 , n37218 , n35375 );
or ( n37220 , n37217 , n37219 );
and ( n37221 , n37215 , n37220 );
not ( n37222 , n37220 );
and ( n37223 , n37205 , n37206 );
xor ( n37224 , n37222 , n37223 );
and ( n37225 , n37224 , n36993 );
or ( n37226 , n37221 , n37225 );
not ( n37227 , n37226 );
buf ( n37228 , n37227 );
buf ( n37229 , n37228 );
not ( n37230 , n37229 );
or ( n37231 , n37214 , n37230 );
not ( n37232 , n36993 );
not ( n37233 , n35375 );
and ( n37234 , n37233 , n36819 );
xor ( n37235 , n36820 , n36975 );
and ( n37236 , n37235 , n35375 );
or ( n37237 , n37234 , n37236 );
and ( n37238 , n37232 , n37237 );
not ( n37239 , n37237 );
and ( n37240 , n37222 , n37223 );
xor ( n37241 , n37239 , n37240 );
and ( n37242 , n37241 , n36993 );
or ( n37243 , n37238 , n37242 );
not ( n37244 , n37243 );
buf ( n37245 , n37244 );
buf ( n37246 , n37245 );
not ( n37247 , n37246 );
or ( n37248 , n37231 , n37247 );
not ( n37249 , n36993 );
not ( n37250 , n35375 );
and ( n37251 , n37250 , n36809 );
xor ( n37252 , n36810 , n36976 );
and ( n37253 , n37252 , n35375 );
or ( n37254 , n37251 , n37253 );
and ( n37255 , n37249 , n37254 );
not ( n37256 , n37254 );
and ( n37257 , n37239 , n37240 );
xor ( n37258 , n37256 , n37257 );
and ( n37259 , n37258 , n36993 );
or ( n37260 , n37255 , n37259 );
not ( n37261 , n37260 );
buf ( n37262 , n37261 );
buf ( n37263 , n37262 );
not ( n37264 , n37263 );
or ( n37265 , n37248 , n37264 );
not ( n37266 , n36993 );
not ( n37267 , n35375 );
and ( n37268 , n37267 , n36799 );
xor ( n37269 , n36800 , n36977 );
and ( n37270 , n37269 , n35375 );
or ( n37271 , n37268 , n37270 );
and ( n37272 , n37266 , n37271 );
not ( n37273 , n37271 );
and ( n37274 , n37256 , n37257 );
xor ( n37275 , n37273 , n37274 );
and ( n37276 , n37275 , n36993 );
or ( n37277 , n37272 , n37276 );
not ( n37278 , n37277 );
buf ( n37279 , n37278 );
buf ( n37280 , n37279 );
not ( n37281 , n37280 );
or ( n37282 , n37265 , n37281 );
not ( n37283 , n36993 );
not ( n37284 , n35375 );
and ( n37285 , n37284 , n36789 );
xor ( n37286 , n36790 , n36978 );
and ( n37287 , n37286 , n35375 );
or ( n37288 , n37285 , n37287 );
and ( n37289 , n37283 , n37288 );
not ( n37290 , n37288 );
and ( n37291 , n37273 , n37274 );
xor ( n37292 , n37290 , n37291 );
and ( n37293 , n37292 , n36993 );
or ( n37294 , n37289 , n37293 );
not ( n37295 , n37294 );
buf ( n37296 , n37295 );
buf ( n37297 , n37296 );
not ( n37298 , n37297 );
or ( n37299 , n37282 , n37298 );
not ( n37300 , n36993 );
not ( n37301 , n35375 );
and ( n37302 , n37301 , n36779 );
xor ( n37303 , n36780 , n36979 );
and ( n37304 , n37303 , n35375 );
or ( n37305 , n37302 , n37304 );
and ( n37306 , n37300 , n37305 );
not ( n37307 , n37305 );
and ( n37308 , n37290 , n37291 );
xor ( n37309 , n37307 , n37308 );
and ( n37310 , n37309 , n36993 );
or ( n37311 , n37306 , n37310 );
not ( n37312 , n37311 );
buf ( n37313 , n37312 );
buf ( n37314 , n37313 );
not ( n37315 , n37314 );
or ( n37316 , n37299 , n37315 );
not ( n37317 , n36993 );
not ( n37318 , n35375 );
and ( n37319 , n37318 , n36769 );
xor ( n37320 , n36770 , n36980 );
and ( n37321 , n37320 , n35375 );
or ( n37322 , n37319 , n37321 );
and ( n37323 , n37317 , n37322 );
not ( n37324 , n37322 );
and ( n37325 , n37307 , n37308 );
xor ( n37326 , n37324 , n37325 );
and ( n37327 , n37326 , n36993 );
or ( n37328 , n37323 , n37327 );
not ( n37329 , n37328 );
buf ( n37330 , n37329 );
buf ( n37331 , n37330 );
not ( n37332 , n37331 );
or ( n37333 , n37316 , n37332 );
not ( n37334 , n36993 );
not ( n37335 , n35375 );
and ( n37336 , n37335 , n36759 );
xor ( n37337 , n36760 , n36981 );
and ( n37338 , n37337 , n35375 );
or ( n37339 , n37336 , n37338 );
and ( n37340 , n37334 , n37339 );
not ( n37341 , n37339 );
and ( n37342 , n37324 , n37325 );
xor ( n37343 , n37341 , n37342 );
and ( n37344 , n37343 , n36993 );
or ( n37345 , n37340 , n37344 );
not ( n37346 , n37345 );
buf ( n37347 , n37346 );
buf ( n37348 , n37347 );
not ( n37349 , n37348 );
or ( n37350 , n37333 , n37349 );
not ( n37351 , n36993 );
not ( n37352 , n35375 );
and ( n37353 , n37352 , n36749 );
xor ( n37354 , n36750 , n36982 );
and ( n37355 , n37354 , n35375 );
or ( n37356 , n37353 , n37355 );
and ( n37357 , n37351 , n37356 );
not ( n37358 , n37356 );
and ( n37359 , n37341 , n37342 );
xor ( n37360 , n37358 , n37359 );
and ( n37361 , n37360 , n36993 );
or ( n37362 , n37357 , n37361 );
not ( n37363 , n37362 );
buf ( n37364 , n37363 );
buf ( n37365 , n37364 );
not ( n37366 , n37365 );
or ( n37367 , n37350 , n37366 );
not ( n37368 , n36993 );
not ( n37369 , n35375 );
and ( n37370 , n37369 , n36739 );
xor ( n37371 , n36740 , n36983 );
and ( n37372 , n37371 , n35375 );
or ( n37373 , n37370 , n37372 );
and ( n37374 , n37368 , n37373 );
not ( n37375 , n37373 );
and ( n37376 , n37358 , n37359 );
xor ( n37377 , n37375 , n37376 );
and ( n37378 , n37377 , n36993 );
or ( n37379 , n37374 , n37378 );
not ( n37380 , n37379 );
buf ( n37381 , n37380 );
buf ( n37382 , n37381 );
not ( n37383 , n37382 );
or ( n37384 , n37367 , n37383 );
not ( n37385 , n36993 );
not ( n37386 , n35375 );
and ( n37387 , n37386 , n36729 );
xor ( n37388 , n36730 , n36984 );
and ( n37389 , n37388 , n35375 );
or ( n37390 , n37387 , n37389 );
and ( n37391 , n37385 , n37390 );
not ( n37392 , n37390 );
and ( n37393 , n37375 , n37376 );
xor ( n37394 , n37392 , n37393 );
and ( n37395 , n37394 , n36993 );
or ( n37396 , n37391 , n37395 );
not ( n37397 , n37396 );
buf ( n37398 , n37397 );
buf ( n37399 , n37398 );
not ( n37400 , n37399 );
or ( n37401 , n37384 , n37400 );
not ( n37402 , n36993 );
not ( n37403 , n35375 );
and ( n37404 , n37403 , n36719 );
xor ( n37405 , n36720 , n36985 );
and ( n37406 , n37405 , n35375 );
or ( n37407 , n37404 , n37406 );
and ( n37408 , n37402 , n37407 );
not ( n37409 , n37407 );
and ( n37410 , n37392 , n37393 );
xor ( n37411 , n37409 , n37410 );
and ( n37412 , n37411 , n36993 );
or ( n37413 , n37408 , n37412 );
not ( n37414 , n37413 );
buf ( n37415 , n37414 );
buf ( n37416 , n37415 );
not ( n37417 , n37416 );
or ( n37418 , n37401 , n37417 );
not ( n37419 , n36993 );
not ( n37420 , n35375 );
and ( n37421 , n37420 , n36709 );
xor ( n37422 , n36710 , n36986 );
and ( n37423 , n37422 , n35375 );
or ( n37424 , n37421 , n37423 );
and ( n37425 , n37419 , n37424 );
not ( n37426 , n37424 );
and ( n37427 , n37409 , n37410 );
xor ( n37428 , n37426 , n37427 );
and ( n37429 , n37428 , n36993 );
or ( n37430 , n37425 , n37429 );
not ( n37431 , n37430 );
buf ( n37432 , n37431 );
buf ( n37433 , n37432 );
not ( n37434 , n37433 );
or ( n37435 , n37418 , n37434 );
not ( n37436 , n36993 );
not ( n37437 , n35375 );
and ( n37438 , n37437 , n36699 );
xor ( n37439 , n36700 , n36987 );
and ( n37440 , n37439 , n35375 );
or ( n37441 , n37438 , n37440 );
and ( n37442 , n37436 , n37441 );
not ( n37443 , n37441 );
and ( n37444 , n37426 , n37427 );
xor ( n37445 , n37443 , n37444 );
and ( n37446 , n37445 , n36993 );
or ( n37447 , n37442 , n37446 );
not ( n37448 , n37447 );
buf ( n37449 , n37448 );
buf ( n37450 , n37449 );
not ( n37451 , n37450 );
or ( n37452 , n37435 , n37451 );
not ( n37453 , n36993 );
not ( n37454 , n35375 );
and ( n37455 , n37454 , n36689 );
xor ( n37456 , n36690 , n36988 );
and ( n37457 , n37456 , n35375 );
or ( n37458 , n37455 , n37457 );
and ( n37459 , n37453 , n37458 );
not ( n37460 , n37458 );
and ( n37461 , n37443 , n37444 );
xor ( n37462 , n37460 , n37461 );
and ( n37463 , n37462 , n36993 );
or ( n37464 , n37459 , n37463 );
not ( n37465 , n37464 );
buf ( n37466 , n37465 );
buf ( n37467 , n37466 );
not ( n37468 , n37467 );
or ( n37469 , n37452 , n37468 );
xor ( n37470 , n36680 , n36989 );
and ( n37471 , n37470 , n35375 );
buf ( n37472 , n37471 );
not ( n37473 , n37472 );
and ( n37474 , n37460 , n37461 );
xor ( n37475 , n37473 , n37474 );
and ( n37476 , n37475 , n36993 );
buf ( n37477 , n37476 );
not ( n37478 , n37477 );
buf ( n37479 , n37478 );
buf ( n37480 , n37479 );
not ( n37481 , n37480 );
or ( n37482 , n37469 , n37481 );
buf ( n37483 , n37482 );
buf ( n37484 , n37483 );
and ( n37485 , n37484 , n36993 );
not ( n37486 , n37485 );
and ( n37487 , n37486 , n37009 );
xor ( n37488 , n37009 , n36993 );
xor ( n37489 , n36615 , n36993 );
and ( n37490 , n37489 , n36993 );
xor ( n37491 , n37488 , n37490 );
and ( n37492 , n37491 , n37485 );
or ( n37493 , n37487 , n37492 );
nor ( n37494 , n31440 , n31442 , n31443 );
and ( n37495 , n37493 , n37494 );
nor ( n37496 , n31445 , n31441 , n31443 );
nor ( n37497 , n31440 , n31441 , n31443 );
or ( n37498 , n37496 , n37497 );
nor ( n37499 , n31445 , n31442 , n31443 );
or ( n37500 , n37498 , n37499 );
and ( n37501 , n31445 , n31442 , n31443 );
or ( n37502 , n37500 , n37501 );
and ( n37503 , n31440 , n31442 , n31443 );
or ( n37504 , n37502 , n37503 );
and ( n37505 , n31440 , n31441 , n31443 );
or ( n37506 , n37504 , n37505 );
and ( n37507 , n35544 , n37506 );
or ( n37508 , n36597 , n37495 , n37507 );
buf ( n37509 , n37508 );
buf ( n37510 , n37509 );
buf ( n37511 , n30987 );
buf ( n37512 , RI15b648d8_1296);
not ( n37513 , n37512 );
buf ( n37514 , RI15b63ac8_1266);
and ( n37515 , n37513 , n37514 );
not ( n37516 , n37514 );
not ( n37517 , n35213 );
xor ( n37518 , n37516 , n37517 );
and ( n37519 , n37518 , n37512 );
or ( n37520 , n37515 , n37519 );
not ( n37521 , n37520 );
buf ( n37522 , n37521 );
buf ( n37523 , n37522 );
not ( n37524 , n37523 );
buf ( n37525 , n37524 );
buf ( n37526 , n37525 );
not ( n37527 , n37526 );
buf ( n37528 , n37527 );
not ( n37529 , n37528 );
not ( n37530 , n37512 );
buf ( n37531 , RI15b64860_1295);
not ( n37532 , n37531 );
buf ( n37533 , RI15b647e8_1294);
not ( n37534 , n37533 );
buf ( n37535 , RI15b64770_1293);
not ( n37536 , n37535 );
buf ( n37537 , RI15b646f8_1292);
not ( n37538 , n37537 );
buf ( n37539 , RI15b64680_1291);
not ( n37540 , n37539 );
buf ( n37541 , RI15b64608_1290);
not ( n37542 , n37541 );
buf ( n37543 , RI15b64590_1289);
not ( n37544 , n37543 );
buf ( n37545 , RI15b64518_1288);
not ( n37546 , n37545 );
buf ( n37547 , RI15b644a0_1287);
not ( n37548 , n37547 );
buf ( n37549 , RI15b64428_1286);
not ( n37550 , n37549 );
buf ( n37551 , RI15b643b0_1285);
not ( n37552 , n37551 );
buf ( n37553 , RI15b64338_1284);
not ( n37554 , n37553 );
buf ( n37555 , RI15b642c0_1283);
not ( n37556 , n37555 );
buf ( n37557 , RI15b64248_1282);
not ( n37558 , n37557 );
buf ( n37559 , RI15b641d0_1281);
not ( n37560 , n37559 );
buf ( n37561 , RI15b64158_1280);
not ( n37562 , n37561 );
buf ( n37563 , RI15b640e0_1279);
not ( n37564 , n37563 );
buf ( n37565 , RI15b64068_1278);
not ( n37566 , n37565 );
buf ( n37567 , RI15b63ff0_1277);
not ( n37568 , n37567 );
buf ( n37569 , RI15b63f78_1276);
not ( n37570 , n37569 );
buf ( n37571 , RI15b63f00_1275);
not ( n37572 , n37571 );
buf ( n37573 , RI15b63e88_1274);
not ( n37574 , n37573 );
not ( n37575 , n32488 );
not ( n37576 , n35677 );
buf ( n37577 , RI15b63d20_1271);
not ( n37578 , n37577 );
buf ( n37579 , RI15b63ca8_1270);
not ( n37580 , n37579 );
buf ( n37581 , RI15b63c30_1269);
not ( n37582 , n37581 );
buf ( n37583 , RI15b63bb8_1268);
not ( n37584 , n37583 );
buf ( n37585 , RI15b63b40_1267);
not ( n37586 , n37585 );
and ( n37587 , n37516 , n37517 );
and ( n37588 , n37586 , n37587 );
and ( n37589 , n37584 , n37588 );
and ( n37590 , n37582 , n37589 );
and ( n37591 , n37580 , n37590 );
and ( n37592 , n37578 , n37591 );
and ( n37593 , n37576 , n37592 );
and ( n37594 , n37575 , n37593 );
and ( n37595 , n37574 , n37594 );
and ( n37596 , n37572 , n37595 );
and ( n37597 , n37570 , n37596 );
and ( n37598 , n37568 , n37597 );
and ( n37599 , n37566 , n37598 );
and ( n37600 , n37564 , n37599 );
and ( n37601 , n37562 , n37600 );
and ( n37602 , n37560 , n37601 );
and ( n37603 , n37558 , n37602 );
and ( n37604 , n37556 , n37603 );
and ( n37605 , n37554 , n37604 );
and ( n37606 , n37552 , n37605 );
and ( n37607 , n37550 , n37606 );
and ( n37608 , n37548 , n37607 );
and ( n37609 , n37546 , n37608 );
and ( n37610 , n37544 , n37609 );
and ( n37611 , n37542 , n37610 );
and ( n37612 , n37540 , n37611 );
and ( n37613 , n37538 , n37612 );
and ( n37614 , n37536 , n37613 );
and ( n37615 , n37534 , n37614 );
and ( n37616 , n37532 , n37615 );
xor ( n37617 , n37530 , n37616 );
buf ( n37618 , n37512 );
and ( n37619 , n37617 , n37618 );
buf ( n37620 , n37619 );
not ( n37621 , n37620 );
not ( n37622 , n37621 );
not ( n37623 , n37622 );
not ( n37624 , n37512 );
and ( n37625 , n37624 , n37531 );
xor ( n37626 , n37532 , n37615 );
and ( n37627 , n37626 , n37512 );
or ( n37628 , n37625 , n37627 );
not ( n37629 , n37628 );
buf ( n37630 , n37629 );
buf ( n37631 , n37630 );
not ( n37632 , n37631 );
not ( n37633 , n37632 );
not ( n37634 , n37512 );
and ( n37635 , n37634 , n37533 );
xor ( n37636 , n37534 , n37614 );
and ( n37637 , n37636 , n37512 );
or ( n37638 , n37635 , n37637 );
not ( n37639 , n37638 );
buf ( n37640 , n37639 );
buf ( n37641 , n37640 );
not ( n37642 , n37641 );
not ( n37643 , n37642 );
not ( n37644 , n37512 );
and ( n37645 , n37644 , n37535 );
xor ( n37646 , n37536 , n37613 );
and ( n37647 , n37646 , n37512 );
or ( n37648 , n37645 , n37647 );
not ( n37649 , n37648 );
buf ( n37650 , n37649 );
buf ( n37651 , n37650 );
not ( n37652 , n37651 );
not ( n37653 , n37652 );
not ( n37654 , n37512 );
and ( n37655 , n37654 , n37537 );
xor ( n37656 , n37538 , n37612 );
and ( n37657 , n37656 , n37512 );
or ( n37658 , n37655 , n37657 );
not ( n37659 , n37658 );
buf ( n37660 , n37659 );
buf ( n37661 , n37660 );
not ( n37662 , n37661 );
not ( n37663 , n37662 );
not ( n37664 , n37512 );
and ( n37665 , n37664 , n37539 );
xor ( n37666 , n37540 , n37611 );
and ( n37667 , n37666 , n37512 );
or ( n37668 , n37665 , n37667 );
not ( n37669 , n37668 );
buf ( n37670 , n37669 );
buf ( n37671 , n37670 );
not ( n37672 , n37671 );
not ( n37673 , n37672 );
not ( n37674 , n37512 );
and ( n37675 , n37674 , n37541 );
xor ( n37676 , n37542 , n37610 );
and ( n37677 , n37676 , n37512 );
or ( n37678 , n37675 , n37677 );
not ( n37679 , n37678 );
buf ( n37680 , n37679 );
buf ( n37681 , n37680 );
not ( n37682 , n37681 );
not ( n37683 , n37682 );
not ( n37684 , n37512 );
and ( n37685 , n37684 , n37543 );
xor ( n37686 , n37544 , n37609 );
and ( n37687 , n37686 , n37512 );
or ( n37688 , n37685 , n37687 );
not ( n37689 , n37688 );
buf ( n37690 , n37689 );
buf ( n37691 , n37690 );
not ( n37692 , n37691 );
not ( n37693 , n37692 );
not ( n37694 , n37512 );
and ( n37695 , n37694 , n37545 );
xor ( n37696 , n37546 , n37608 );
and ( n37697 , n37696 , n37512 );
or ( n37698 , n37695 , n37697 );
not ( n37699 , n37698 );
buf ( n37700 , n37699 );
buf ( n37701 , n37700 );
not ( n37702 , n37701 );
not ( n37703 , n37702 );
not ( n37704 , n37512 );
and ( n37705 , n37704 , n37547 );
xor ( n37706 , n37548 , n37607 );
and ( n37707 , n37706 , n37512 );
or ( n37708 , n37705 , n37707 );
not ( n37709 , n37708 );
buf ( n37710 , n37709 );
buf ( n37711 , n37710 );
not ( n37712 , n37711 );
not ( n37713 , n37712 );
not ( n37714 , n37512 );
and ( n37715 , n37714 , n37549 );
xor ( n37716 , n37550 , n37606 );
and ( n37717 , n37716 , n37512 );
or ( n37718 , n37715 , n37717 );
not ( n37719 , n37718 );
buf ( n37720 , n37719 );
buf ( n37721 , n37720 );
not ( n37722 , n37721 );
not ( n37723 , n37722 );
not ( n37724 , n37512 );
and ( n37725 , n37724 , n37551 );
xor ( n37726 , n37552 , n37605 );
and ( n37727 , n37726 , n37512 );
or ( n37728 , n37725 , n37727 );
not ( n37729 , n37728 );
buf ( n37730 , n37729 );
buf ( n37731 , n37730 );
not ( n37732 , n37731 );
not ( n37733 , n37732 );
not ( n37734 , n37512 );
and ( n37735 , n37734 , n37553 );
xor ( n37736 , n37554 , n37604 );
and ( n37737 , n37736 , n37512 );
or ( n37738 , n37735 , n37737 );
not ( n37739 , n37738 );
buf ( n37740 , n37739 );
buf ( n37741 , n37740 );
not ( n37742 , n37741 );
not ( n37743 , n37742 );
not ( n37744 , n37512 );
and ( n37745 , n37744 , n37555 );
xor ( n37746 , n37556 , n37603 );
and ( n37747 , n37746 , n37512 );
or ( n37748 , n37745 , n37747 );
not ( n37749 , n37748 );
buf ( n37750 , n37749 );
buf ( n37751 , n37750 );
not ( n37752 , n37751 );
not ( n37753 , n37752 );
not ( n37754 , n37512 );
and ( n37755 , n37754 , n37557 );
xor ( n37756 , n37558 , n37602 );
and ( n37757 , n37756 , n37512 );
or ( n37758 , n37755 , n37757 );
not ( n37759 , n37758 );
buf ( n37760 , n37759 );
buf ( n37761 , n37760 );
not ( n37762 , n37761 );
not ( n37763 , n37762 );
not ( n37764 , n37512 );
and ( n37765 , n37764 , n37559 );
xor ( n37766 , n37560 , n37601 );
and ( n37767 , n37766 , n37512 );
or ( n37768 , n37765 , n37767 );
not ( n37769 , n37768 );
buf ( n37770 , n37769 );
buf ( n37771 , n37770 );
not ( n37772 , n37771 );
not ( n37773 , n37772 );
not ( n37774 , n37512 );
and ( n37775 , n37774 , n37561 );
xor ( n37776 , n37562 , n37600 );
and ( n37777 , n37776 , n37512 );
or ( n37778 , n37775 , n37777 );
not ( n37779 , n37778 );
buf ( n37780 , n37779 );
buf ( n37781 , n37780 );
not ( n37782 , n37781 );
not ( n37783 , n37782 );
not ( n37784 , n37512 );
and ( n37785 , n37784 , n37563 );
xor ( n37786 , n37564 , n37599 );
and ( n37787 , n37786 , n37512 );
or ( n37788 , n37785 , n37787 );
not ( n37789 , n37788 );
buf ( n37790 , n37789 );
buf ( n37791 , n37790 );
not ( n37792 , n37791 );
not ( n37793 , n37792 );
not ( n37794 , n37512 );
and ( n37795 , n37794 , n37565 );
xor ( n37796 , n37566 , n37598 );
and ( n37797 , n37796 , n37512 );
or ( n37798 , n37795 , n37797 );
not ( n37799 , n37798 );
buf ( n37800 , n37799 );
buf ( n37801 , n37800 );
not ( n37802 , n37801 );
not ( n37803 , n37802 );
not ( n37804 , n37512 );
and ( n37805 , n37804 , n37567 );
xor ( n37806 , n37568 , n37597 );
and ( n37807 , n37806 , n37512 );
or ( n37808 , n37805 , n37807 );
not ( n37809 , n37808 );
buf ( n37810 , n37809 );
buf ( n37811 , n37810 );
not ( n37812 , n37811 );
not ( n37813 , n37812 );
not ( n37814 , n37512 );
and ( n37815 , n37814 , n37569 );
xor ( n37816 , n37570 , n37596 );
and ( n37817 , n37816 , n37512 );
or ( n37818 , n37815 , n37817 );
not ( n37819 , n37818 );
buf ( n37820 , n37819 );
buf ( n37821 , n37820 );
not ( n37822 , n37821 );
not ( n37823 , n37822 );
not ( n37824 , n37512 );
and ( n37825 , n37824 , n37571 );
xor ( n37826 , n37572 , n37595 );
and ( n37827 , n37826 , n37512 );
or ( n37828 , n37825 , n37827 );
not ( n37829 , n37828 );
buf ( n37830 , n37829 );
buf ( n37831 , n37830 );
not ( n37832 , n37831 );
not ( n37833 , n37832 );
not ( n37834 , n37512 );
and ( n37835 , n37834 , n37573 );
xor ( n37836 , n37574 , n37594 );
and ( n37837 , n37836 , n37512 );
or ( n37838 , n37835 , n37837 );
not ( n37839 , n37838 );
buf ( n37840 , n37839 );
buf ( n37841 , n37840 );
not ( n37842 , n37841 );
not ( n37843 , n37842 );
not ( n37844 , n37512 );
and ( n37845 , n37844 , n32488 );
xor ( n37846 , n37575 , n37593 );
and ( n37847 , n37846 , n37512 );
or ( n37848 , n37845 , n37847 );
not ( n37849 , n37848 );
buf ( n37850 , n37849 );
buf ( n37851 , n37850 );
not ( n37852 , n37851 );
not ( n37853 , n37852 );
not ( n37854 , n37512 );
and ( n37855 , n37854 , n35677 );
xor ( n37856 , n37576 , n37592 );
and ( n37857 , n37856 , n37512 );
or ( n37858 , n37855 , n37857 );
not ( n37859 , n37858 );
buf ( n37860 , n37859 );
buf ( n37861 , n37860 );
not ( n37862 , n37861 );
not ( n37863 , n37862 );
not ( n37864 , n37512 );
and ( n37865 , n37864 , n37577 );
xor ( n37866 , n37578 , n37591 );
and ( n37867 , n37866 , n37512 );
or ( n37868 , n37865 , n37867 );
not ( n37869 , n37868 );
buf ( n37870 , n37869 );
buf ( n37871 , n37870 );
not ( n37872 , n37871 );
not ( n37873 , n37872 );
not ( n37874 , n37512 );
and ( n37875 , n37874 , n37579 );
xor ( n37876 , n37580 , n37590 );
and ( n37877 , n37876 , n37512 );
or ( n37878 , n37875 , n37877 );
not ( n37879 , n37878 );
buf ( n37880 , n37879 );
buf ( n37881 , n37880 );
not ( n37882 , n37881 );
not ( n37883 , n37882 );
not ( n37884 , n37512 );
and ( n37885 , n37884 , n37581 );
xor ( n37886 , n37582 , n37589 );
and ( n37887 , n37886 , n37512 );
or ( n37888 , n37885 , n37887 );
not ( n37889 , n37888 );
buf ( n37890 , n37889 );
buf ( n37891 , n37890 );
not ( n37892 , n37891 );
not ( n37893 , n37892 );
not ( n37894 , n37512 );
and ( n37895 , n37894 , n37583 );
xor ( n37896 , n37584 , n37588 );
and ( n37897 , n37896 , n37512 );
or ( n37898 , n37895 , n37897 );
not ( n37899 , n37898 );
buf ( n37900 , n37899 );
buf ( n37901 , n37900 );
not ( n37902 , n37901 );
not ( n37903 , n37902 );
not ( n37904 , n37512 );
and ( n37905 , n37904 , n37585 );
xor ( n37906 , n37586 , n37587 );
and ( n37907 , n37906 , n37512 );
or ( n37908 , n37905 , n37907 );
not ( n37909 , n37908 );
buf ( n37910 , n37909 );
buf ( n37911 , n37910 );
not ( n37912 , n37911 );
not ( n37913 , n37912 );
not ( n37914 , n37524 );
and ( n37915 , n37913 , n37914 );
and ( n37916 , n37903 , n37915 );
and ( n37917 , n37893 , n37916 );
and ( n37918 , n37883 , n37917 );
and ( n37919 , n37873 , n37918 );
and ( n37920 , n37863 , n37919 );
and ( n37921 , n37853 , n37920 );
and ( n37922 , n37843 , n37921 );
and ( n37923 , n37833 , n37922 );
and ( n37924 , n37823 , n37923 );
and ( n37925 , n37813 , n37924 );
and ( n37926 , n37803 , n37925 );
and ( n37927 , n37793 , n37926 );
and ( n37928 , n37783 , n37927 );
and ( n37929 , n37773 , n37928 );
and ( n37930 , n37763 , n37929 );
and ( n37931 , n37753 , n37930 );
and ( n37932 , n37743 , n37931 );
and ( n37933 , n37733 , n37932 );
and ( n37934 , n37723 , n37933 );
and ( n37935 , n37713 , n37934 );
and ( n37936 , n37703 , n37935 );
and ( n37937 , n37693 , n37936 );
and ( n37938 , n37683 , n37937 );
and ( n37939 , n37673 , n37938 );
and ( n37940 , n37663 , n37939 );
and ( n37941 , n37653 , n37940 );
and ( n37942 , n37643 , n37941 );
and ( n37943 , n37633 , n37942 );
and ( n37944 , n37623 , n37943 );
not ( n37945 , n37944 );
and ( n37946 , n37945 , n37512 );
buf ( n37947 , n37946 );
not ( n37948 , n37947 );
not ( n37949 , n37512 );
and ( n37950 , n37949 , n37912 );
xor ( n37951 , n37913 , n37914 );
and ( n37952 , n37951 , n37512 );
or ( n37953 , n37950 , n37952 );
and ( n37954 , n37948 , n37953 );
not ( n37955 , n37953 );
not ( n37956 , n37525 );
xor ( n37957 , n37955 , n37956 );
and ( n37958 , n37957 , n37947 );
or ( n37959 , n37954 , n37958 );
not ( n37960 , n37959 );
buf ( n37961 , n37960 );
buf ( n37962 , n37961 );
not ( n37963 , n37962 );
or ( n37964 , n37529 , n37963 );
not ( n37965 , n37947 );
not ( n37966 , n37512 );
and ( n37967 , n37966 , n37902 );
xor ( n37968 , n37903 , n37915 );
and ( n37969 , n37968 , n37512 );
or ( n37970 , n37967 , n37969 );
and ( n37971 , n37965 , n37970 );
not ( n37972 , n37970 );
and ( n37973 , n37955 , n37956 );
xor ( n37974 , n37972 , n37973 );
and ( n37975 , n37974 , n37947 );
or ( n37976 , n37971 , n37975 );
not ( n37977 , n37976 );
buf ( n37978 , n37977 );
buf ( n37979 , n37978 );
not ( n37980 , n37979 );
or ( n37981 , n37964 , n37980 );
not ( n37982 , n37947 );
not ( n37983 , n37512 );
and ( n37984 , n37983 , n37892 );
xor ( n37985 , n37893 , n37916 );
and ( n37986 , n37985 , n37512 );
or ( n37987 , n37984 , n37986 );
and ( n37988 , n37982 , n37987 );
not ( n37989 , n37987 );
and ( n37990 , n37972 , n37973 );
xor ( n37991 , n37989 , n37990 );
and ( n37992 , n37991 , n37947 );
or ( n37993 , n37988 , n37992 );
not ( n37994 , n37993 );
buf ( n37995 , n37994 );
buf ( n37996 , n37995 );
not ( n37997 , n37996 );
or ( n37998 , n37981 , n37997 );
not ( n37999 , n37947 );
not ( n38000 , n37512 );
and ( n38001 , n38000 , n37882 );
xor ( n38002 , n37883 , n37917 );
and ( n38003 , n38002 , n37512 );
or ( n38004 , n38001 , n38003 );
and ( n38005 , n37999 , n38004 );
not ( n38006 , n38004 );
and ( n38007 , n37989 , n37990 );
xor ( n38008 , n38006 , n38007 );
and ( n38009 , n38008 , n37947 );
or ( n38010 , n38005 , n38009 );
not ( n38011 , n38010 );
buf ( n38012 , n38011 );
buf ( n38013 , n38012 );
not ( n38014 , n38013 );
or ( n38015 , n37998 , n38014 );
not ( n38016 , n37947 );
not ( n38017 , n37512 );
and ( n38018 , n38017 , n37872 );
xor ( n38019 , n37873 , n37918 );
and ( n38020 , n38019 , n37512 );
or ( n38021 , n38018 , n38020 );
and ( n38022 , n38016 , n38021 );
not ( n38023 , n38021 );
and ( n38024 , n38006 , n38007 );
xor ( n38025 , n38023 , n38024 );
and ( n38026 , n38025 , n37947 );
or ( n38027 , n38022 , n38026 );
not ( n38028 , n38027 );
buf ( n38029 , n38028 );
buf ( n38030 , n38029 );
not ( n38031 , n38030 );
or ( n38032 , n38015 , n38031 );
not ( n38033 , n37947 );
not ( n38034 , n37512 );
and ( n38035 , n38034 , n37862 );
xor ( n38036 , n37863 , n37919 );
and ( n38037 , n38036 , n37512 );
or ( n38038 , n38035 , n38037 );
and ( n38039 , n38033 , n38038 );
not ( n38040 , n38038 );
and ( n38041 , n38023 , n38024 );
xor ( n38042 , n38040 , n38041 );
and ( n38043 , n38042 , n37947 );
or ( n38044 , n38039 , n38043 );
not ( n38045 , n38044 );
buf ( n38046 , n38045 );
buf ( n38047 , n38046 );
not ( n38048 , n38047 );
or ( n38049 , n38032 , n38048 );
not ( n38050 , n37947 );
not ( n38051 , n37512 );
and ( n38052 , n38051 , n37852 );
xor ( n38053 , n37853 , n37920 );
and ( n38054 , n38053 , n37512 );
or ( n38055 , n38052 , n38054 );
and ( n38056 , n38050 , n38055 );
not ( n38057 , n38055 );
and ( n38058 , n38040 , n38041 );
xor ( n38059 , n38057 , n38058 );
and ( n38060 , n38059 , n37947 );
or ( n38061 , n38056 , n38060 );
not ( n38062 , n38061 );
buf ( n38063 , n38062 );
buf ( n38064 , n38063 );
not ( n38065 , n38064 );
or ( n38066 , n38049 , n38065 );
not ( n38067 , n37947 );
not ( n38068 , n37512 );
and ( n38069 , n38068 , n37842 );
xor ( n38070 , n37843 , n37921 );
and ( n38071 , n38070 , n37512 );
or ( n38072 , n38069 , n38071 );
and ( n38073 , n38067 , n38072 );
not ( n38074 , n38072 );
and ( n38075 , n38057 , n38058 );
xor ( n38076 , n38074 , n38075 );
and ( n38077 , n38076 , n37947 );
or ( n38078 , n38073 , n38077 );
not ( n38079 , n38078 );
buf ( n38080 , n38079 );
buf ( n38081 , n38080 );
not ( n38082 , n38081 );
or ( n38083 , n38066 , n38082 );
not ( n38084 , n37947 );
not ( n38085 , n37512 );
and ( n38086 , n38085 , n37832 );
xor ( n38087 , n37833 , n37922 );
and ( n38088 , n38087 , n37512 );
or ( n38089 , n38086 , n38088 );
and ( n38090 , n38084 , n38089 );
not ( n38091 , n38089 );
and ( n38092 , n38074 , n38075 );
xor ( n38093 , n38091 , n38092 );
and ( n38094 , n38093 , n37947 );
or ( n38095 , n38090 , n38094 );
not ( n38096 , n38095 );
buf ( n38097 , n38096 );
buf ( n38098 , n38097 );
not ( n38099 , n38098 );
or ( n38100 , n38083 , n38099 );
not ( n38101 , n37947 );
not ( n38102 , n37512 );
and ( n38103 , n38102 , n37822 );
xor ( n38104 , n37823 , n37923 );
and ( n38105 , n38104 , n37512 );
or ( n38106 , n38103 , n38105 );
and ( n38107 , n38101 , n38106 );
not ( n38108 , n38106 );
and ( n38109 , n38091 , n38092 );
xor ( n38110 , n38108 , n38109 );
and ( n38111 , n38110 , n37947 );
or ( n38112 , n38107 , n38111 );
not ( n38113 , n38112 );
buf ( n38114 , n38113 );
buf ( n38115 , n38114 );
not ( n38116 , n38115 );
or ( n38117 , n38100 , n38116 );
not ( n38118 , n37947 );
not ( n38119 , n37512 );
and ( n38120 , n38119 , n37812 );
xor ( n38121 , n37813 , n37924 );
and ( n38122 , n38121 , n37512 );
or ( n38123 , n38120 , n38122 );
and ( n38124 , n38118 , n38123 );
not ( n38125 , n38123 );
and ( n38126 , n38108 , n38109 );
xor ( n38127 , n38125 , n38126 );
and ( n38128 , n38127 , n37947 );
or ( n38129 , n38124 , n38128 );
not ( n38130 , n38129 );
buf ( n38131 , n38130 );
buf ( n38132 , n38131 );
not ( n38133 , n38132 );
or ( n38134 , n38117 , n38133 );
not ( n38135 , n37947 );
not ( n38136 , n37512 );
and ( n38137 , n38136 , n37802 );
xor ( n38138 , n37803 , n37925 );
and ( n38139 , n38138 , n37512 );
or ( n38140 , n38137 , n38139 );
and ( n38141 , n38135 , n38140 );
not ( n38142 , n38140 );
and ( n38143 , n38125 , n38126 );
xor ( n38144 , n38142 , n38143 );
and ( n38145 , n38144 , n37947 );
or ( n38146 , n38141 , n38145 );
not ( n38147 , n38146 );
buf ( n38148 , n38147 );
buf ( n38149 , n38148 );
not ( n38150 , n38149 );
or ( n38151 , n38134 , n38150 );
not ( n38152 , n37947 );
not ( n38153 , n37512 );
and ( n38154 , n38153 , n37792 );
xor ( n38155 , n37793 , n37926 );
and ( n38156 , n38155 , n37512 );
or ( n38157 , n38154 , n38156 );
and ( n38158 , n38152 , n38157 );
not ( n38159 , n38157 );
and ( n38160 , n38142 , n38143 );
xor ( n38161 , n38159 , n38160 );
and ( n38162 , n38161 , n37947 );
or ( n38163 , n38158 , n38162 );
not ( n38164 , n38163 );
buf ( n38165 , n38164 );
buf ( n38166 , n38165 );
not ( n38167 , n38166 );
or ( n38168 , n38151 , n38167 );
not ( n38169 , n37947 );
not ( n38170 , n37512 );
and ( n38171 , n38170 , n37782 );
xor ( n38172 , n37783 , n37927 );
and ( n38173 , n38172 , n37512 );
or ( n38174 , n38171 , n38173 );
and ( n38175 , n38169 , n38174 );
not ( n38176 , n38174 );
and ( n38177 , n38159 , n38160 );
xor ( n38178 , n38176 , n38177 );
and ( n38179 , n38178 , n37947 );
or ( n38180 , n38175 , n38179 );
not ( n38181 , n38180 );
buf ( n38182 , n38181 );
buf ( n38183 , n38182 );
not ( n38184 , n38183 );
or ( n38185 , n38168 , n38184 );
not ( n38186 , n37947 );
not ( n38187 , n37512 );
and ( n38188 , n38187 , n37772 );
xor ( n38189 , n37773 , n37928 );
and ( n38190 , n38189 , n37512 );
or ( n38191 , n38188 , n38190 );
and ( n38192 , n38186 , n38191 );
not ( n38193 , n38191 );
and ( n38194 , n38176 , n38177 );
xor ( n38195 , n38193 , n38194 );
and ( n38196 , n38195 , n37947 );
or ( n38197 , n38192 , n38196 );
not ( n38198 , n38197 );
buf ( n38199 , n38198 );
buf ( n38200 , n38199 );
not ( n38201 , n38200 );
or ( n38202 , n38185 , n38201 );
not ( n38203 , n37947 );
not ( n38204 , n37512 );
and ( n38205 , n38204 , n37762 );
xor ( n38206 , n37763 , n37929 );
and ( n38207 , n38206 , n37512 );
or ( n38208 , n38205 , n38207 );
and ( n38209 , n38203 , n38208 );
not ( n38210 , n38208 );
and ( n38211 , n38193 , n38194 );
xor ( n38212 , n38210 , n38211 );
and ( n38213 , n38212 , n37947 );
or ( n38214 , n38209 , n38213 );
not ( n38215 , n38214 );
buf ( n38216 , n38215 );
buf ( n38217 , n38216 );
not ( n38218 , n38217 );
or ( n38219 , n38202 , n38218 );
not ( n38220 , n37947 );
not ( n38221 , n37512 );
and ( n38222 , n38221 , n37752 );
xor ( n38223 , n37753 , n37930 );
and ( n38224 , n38223 , n37512 );
or ( n38225 , n38222 , n38224 );
and ( n38226 , n38220 , n38225 );
not ( n38227 , n38225 );
and ( n38228 , n38210 , n38211 );
xor ( n38229 , n38227 , n38228 );
and ( n38230 , n38229 , n37947 );
or ( n38231 , n38226 , n38230 );
not ( n38232 , n38231 );
buf ( n38233 , n38232 );
buf ( n38234 , n38233 );
not ( n38235 , n38234 );
or ( n38236 , n38219 , n38235 );
not ( n38237 , n37947 );
not ( n38238 , n37512 );
and ( n38239 , n38238 , n37742 );
xor ( n38240 , n37743 , n37931 );
and ( n38241 , n38240 , n37512 );
or ( n38242 , n38239 , n38241 );
and ( n38243 , n38237 , n38242 );
not ( n38244 , n38242 );
and ( n38245 , n38227 , n38228 );
xor ( n38246 , n38244 , n38245 );
and ( n38247 , n38246 , n37947 );
or ( n38248 , n38243 , n38247 );
not ( n38249 , n38248 );
buf ( n38250 , n38249 );
buf ( n38251 , n38250 );
not ( n38252 , n38251 );
or ( n38253 , n38236 , n38252 );
not ( n38254 , n37947 );
not ( n38255 , n37512 );
and ( n38256 , n38255 , n37732 );
xor ( n38257 , n37733 , n37932 );
and ( n38258 , n38257 , n37512 );
or ( n38259 , n38256 , n38258 );
and ( n38260 , n38254 , n38259 );
not ( n38261 , n38259 );
and ( n38262 , n38244 , n38245 );
xor ( n38263 , n38261 , n38262 );
and ( n38264 , n38263 , n37947 );
or ( n38265 , n38260 , n38264 );
not ( n38266 , n38265 );
buf ( n38267 , n38266 );
buf ( n38268 , n38267 );
not ( n38269 , n38268 );
or ( n38270 , n38253 , n38269 );
not ( n38271 , n37947 );
not ( n38272 , n37512 );
and ( n38273 , n38272 , n37722 );
xor ( n38274 , n37723 , n37933 );
and ( n38275 , n38274 , n37512 );
or ( n38276 , n38273 , n38275 );
and ( n38277 , n38271 , n38276 );
not ( n38278 , n38276 );
and ( n38279 , n38261 , n38262 );
xor ( n38280 , n38278 , n38279 );
and ( n38281 , n38280 , n37947 );
or ( n38282 , n38277 , n38281 );
not ( n38283 , n38282 );
buf ( n38284 , n38283 );
buf ( n38285 , n38284 );
not ( n38286 , n38285 );
or ( n38287 , n38270 , n38286 );
not ( n38288 , n37947 );
not ( n38289 , n37512 );
and ( n38290 , n38289 , n37712 );
xor ( n38291 , n37713 , n37934 );
and ( n38292 , n38291 , n37512 );
or ( n38293 , n38290 , n38292 );
and ( n38294 , n38288 , n38293 );
not ( n38295 , n38293 );
and ( n38296 , n38278 , n38279 );
xor ( n38297 , n38295 , n38296 );
and ( n38298 , n38297 , n37947 );
or ( n38299 , n38294 , n38298 );
not ( n38300 , n38299 );
buf ( n38301 , n38300 );
buf ( n38302 , n38301 );
not ( n38303 , n38302 );
or ( n38304 , n38287 , n38303 );
not ( n38305 , n37947 );
not ( n38306 , n37512 );
and ( n38307 , n38306 , n37702 );
xor ( n38308 , n37703 , n37935 );
and ( n38309 , n38308 , n37512 );
or ( n38310 , n38307 , n38309 );
and ( n38311 , n38305 , n38310 );
not ( n38312 , n38310 );
and ( n38313 , n38295 , n38296 );
xor ( n38314 , n38312 , n38313 );
and ( n38315 , n38314 , n37947 );
or ( n38316 , n38311 , n38315 );
not ( n38317 , n38316 );
buf ( n38318 , n38317 );
buf ( n38319 , n38318 );
not ( n38320 , n38319 );
or ( n38321 , n38304 , n38320 );
not ( n38322 , n37947 );
not ( n38323 , n37512 );
and ( n38324 , n38323 , n37692 );
xor ( n38325 , n37693 , n37936 );
and ( n38326 , n38325 , n37512 );
or ( n38327 , n38324 , n38326 );
and ( n38328 , n38322 , n38327 );
not ( n38329 , n38327 );
and ( n38330 , n38312 , n38313 );
xor ( n38331 , n38329 , n38330 );
and ( n38332 , n38331 , n37947 );
or ( n38333 , n38328 , n38332 );
not ( n38334 , n38333 );
buf ( n38335 , n38334 );
buf ( n38336 , n38335 );
not ( n38337 , n38336 );
or ( n38338 , n38321 , n38337 );
not ( n38339 , n37947 );
not ( n38340 , n37512 );
and ( n38341 , n38340 , n37682 );
xor ( n38342 , n37683 , n37937 );
and ( n38343 , n38342 , n37512 );
or ( n38344 , n38341 , n38343 );
and ( n38345 , n38339 , n38344 );
not ( n38346 , n38344 );
and ( n38347 , n38329 , n38330 );
xor ( n38348 , n38346 , n38347 );
and ( n38349 , n38348 , n37947 );
or ( n38350 , n38345 , n38349 );
not ( n38351 , n38350 );
buf ( n38352 , n38351 );
buf ( n38353 , n38352 );
not ( n38354 , n38353 );
or ( n38355 , n38338 , n38354 );
not ( n38356 , n37947 );
not ( n38357 , n37512 );
and ( n38358 , n38357 , n37672 );
xor ( n38359 , n37673 , n37938 );
and ( n38360 , n38359 , n37512 );
or ( n38361 , n38358 , n38360 );
and ( n38362 , n38356 , n38361 );
not ( n38363 , n38361 );
and ( n38364 , n38346 , n38347 );
xor ( n38365 , n38363 , n38364 );
and ( n38366 , n38365 , n37947 );
or ( n38367 , n38362 , n38366 );
not ( n38368 , n38367 );
buf ( n38369 , n38368 );
buf ( n38370 , n38369 );
not ( n38371 , n38370 );
or ( n38372 , n38355 , n38371 );
not ( n38373 , n37947 );
not ( n38374 , n37512 );
and ( n38375 , n38374 , n37662 );
xor ( n38376 , n37663 , n37939 );
and ( n38377 , n38376 , n37512 );
or ( n38378 , n38375 , n38377 );
and ( n38379 , n38373 , n38378 );
not ( n38380 , n38378 );
and ( n38381 , n38363 , n38364 );
xor ( n38382 , n38380 , n38381 );
and ( n38383 , n38382 , n37947 );
or ( n38384 , n38379 , n38383 );
not ( n38385 , n38384 );
buf ( n38386 , n38385 );
buf ( n38387 , n38386 );
not ( n38388 , n38387 );
or ( n38389 , n38372 , n38388 );
not ( n38390 , n37947 );
not ( n38391 , n37512 );
and ( n38392 , n38391 , n37652 );
xor ( n38393 , n37653 , n37940 );
and ( n38394 , n38393 , n37512 );
or ( n38395 , n38392 , n38394 );
and ( n38396 , n38390 , n38395 );
not ( n38397 , n38395 );
and ( n38398 , n38380 , n38381 );
xor ( n38399 , n38397 , n38398 );
and ( n38400 , n38399 , n37947 );
or ( n38401 , n38396 , n38400 );
not ( n38402 , n38401 );
buf ( n38403 , n38402 );
buf ( n38404 , n38403 );
not ( n38405 , n38404 );
or ( n38406 , n38389 , n38405 );
not ( n38407 , n37947 );
not ( n38408 , n37512 );
and ( n38409 , n38408 , n37642 );
xor ( n38410 , n37643 , n37941 );
and ( n38411 , n38410 , n37512 );
or ( n38412 , n38409 , n38411 );
and ( n38413 , n38407 , n38412 );
not ( n38414 , n38412 );
and ( n38415 , n38397 , n38398 );
xor ( n38416 , n38414 , n38415 );
and ( n38417 , n38416 , n37947 );
or ( n38418 , n38413 , n38417 );
not ( n38419 , n38418 );
buf ( n38420 , n38419 );
buf ( n38421 , n38420 );
not ( n38422 , n38421 );
or ( n38423 , n38406 , n38422 );
not ( n38424 , n37947 );
not ( n38425 , n37512 );
and ( n38426 , n38425 , n37632 );
xor ( n38427 , n37633 , n37942 );
and ( n38428 , n38427 , n37512 );
or ( n38429 , n38426 , n38428 );
and ( n38430 , n38424 , n38429 );
not ( n38431 , n38429 );
and ( n38432 , n38414 , n38415 );
xor ( n38433 , n38431 , n38432 );
and ( n38434 , n38433 , n37947 );
or ( n38435 , n38430 , n38434 );
not ( n38436 , n38435 );
buf ( n38437 , n38436 );
buf ( n38438 , n38437 );
not ( n38439 , n38438 );
or ( n38440 , n38423 , n38439 );
buf ( n38441 , n38440 );
buf ( n38442 , n38441 );
and ( n38443 , n38442 , n37947 );
not ( n38444 , n38443 );
and ( n38445 , n38444 , n37529 );
xor ( n38446 , n37529 , n37947 );
xor ( n38447 , n38446 , n37947 );
and ( n38448 , n38447 , n38443 );
or ( n38449 , n38445 , n38448 );
and ( n38450 , n35286 , n35282 , n35284 );
and ( n38451 , n38449 , n38450 );
not ( n38452 , n37512 );
and ( n38453 , n38452 , n37585 );
not ( n38454 , n37585 );
not ( n38455 , n37514 );
not ( n38456 , n35213 );
and ( n38457 , n38455 , n38456 );
xor ( n38458 , n38454 , n38457 );
and ( n38459 , n38458 , n37512 );
or ( n38460 , n38453 , n38459 );
not ( n38461 , n38460 );
buf ( n38462 , n38461 );
buf ( n38463 , n38462 );
not ( n38464 , n38463 );
buf ( n38465 , n38464 );
buf ( n38466 , n38465 );
not ( n38467 , n38466 );
buf ( n38468 , n38467 );
not ( n38469 , n38468 );
not ( n38470 , n37512 );
not ( n38471 , n37531 );
not ( n38472 , n37533 );
not ( n38473 , n37535 );
not ( n38474 , n37537 );
not ( n38475 , n37539 );
not ( n38476 , n37541 );
not ( n38477 , n37543 );
not ( n38478 , n37545 );
not ( n38479 , n37547 );
not ( n38480 , n37549 );
not ( n38481 , n37551 );
not ( n38482 , n37553 );
not ( n38483 , n37555 );
not ( n38484 , n37557 );
not ( n38485 , n37559 );
not ( n38486 , n37561 );
not ( n38487 , n37563 );
not ( n38488 , n37565 );
not ( n38489 , n37567 );
not ( n38490 , n37569 );
not ( n38491 , n37571 );
not ( n38492 , n37573 );
not ( n38493 , n32488 );
not ( n38494 , n35677 );
not ( n38495 , n37577 );
not ( n38496 , n37579 );
not ( n38497 , n37581 );
not ( n38498 , n37583 );
and ( n38499 , n38454 , n38457 );
and ( n38500 , n38498 , n38499 );
and ( n38501 , n38497 , n38500 );
and ( n38502 , n38496 , n38501 );
and ( n38503 , n38495 , n38502 );
and ( n38504 , n38494 , n38503 );
and ( n38505 , n38493 , n38504 );
and ( n38506 , n38492 , n38505 );
and ( n38507 , n38491 , n38506 );
and ( n38508 , n38490 , n38507 );
and ( n38509 , n38489 , n38508 );
and ( n38510 , n38488 , n38509 );
and ( n38511 , n38487 , n38510 );
and ( n38512 , n38486 , n38511 );
and ( n38513 , n38485 , n38512 );
and ( n38514 , n38484 , n38513 );
and ( n38515 , n38483 , n38514 );
and ( n38516 , n38482 , n38515 );
and ( n38517 , n38481 , n38516 );
and ( n38518 , n38480 , n38517 );
and ( n38519 , n38479 , n38518 );
and ( n38520 , n38478 , n38519 );
and ( n38521 , n38477 , n38520 );
and ( n38522 , n38476 , n38521 );
and ( n38523 , n38475 , n38522 );
and ( n38524 , n38474 , n38523 );
and ( n38525 , n38473 , n38524 );
and ( n38526 , n38472 , n38525 );
and ( n38527 , n38471 , n38526 );
xor ( n38528 , n38470 , n38527 );
buf ( n38529 , n37512 );
and ( n38530 , n38528 , n38529 );
buf ( n38531 , n38530 );
not ( n38532 , n38531 );
not ( n38533 , n38532 );
not ( n38534 , n38533 );
not ( n38535 , n37512 );
and ( n38536 , n38535 , n37531 );
xor ( n38537 , n38471 , n38526 );
and ( n38538 , n38537 , n37512 );
or ( n38539 , n38536 , n38538 );
not ( n38540 , n38539 );
buf ( n38541 , n38540 );
buf ( n38542 , n38541 );
not ( n38543 , n38542 );
not ( n38544 , n38543 );
not ( n38545 , n37512 );
and ( n38546 , n38545 , n37533 );
xor ( n38547 , n38472 , n38525 );
and ( n38548 , n38547 , n37512 );
or ( n38549 , n38546 , n38548 );
not ( n38550 , n38549 );
buf ( n38551 , n38550 );
buf ( n38552 , n38551 );
not ( n38553 , n38552 );
not ( n38554 , n38553 );
not ( n38555 , n37512 );
and ( n38556 , n38555 , n37535 );
xor ( n38557 , n38473 , n38524 );
and ( n38558 , n38557 , n37512 );
or ( n38559 , n38556 , n38558 );
not ( n38560 , n38559 );
buf ( n38561 , n38560 );
buf ( n38562 , n38561 );
not ( n38563 , n38562 );
not ( n38564 , n38563 );
not ( n38565 , n37512 );
and ( n38566 , n38565 , n37537 );
xor ( n38567 , n38474 , n38523 );
and ( n38568 , n38567 , n37512 );
or ( n38569 , n38566 , n38568 );
not ( n38570 , n38569 );
buf ( n38571 , n38570 );
buf ( n38572 , n38571 );
not ( n38573 , n38572 );
not ( n38574 , n38573 );
not ( n38575 , n37512 );
and ( n38576 , n38575 , n37539 );
xor ( n38577 , n38475 , n38522 );
and ( n38578 , n38577 , n37512 );
or ( n38579 , n38576 , n38578 );
not ( n38580 , n38579 );
buf ( n38581 , n38580 );
buf ( n38582 , n38581 );
not ( n38583 , n38582 );
not ( n38584 , n38583 );
not ( n38585 , n37512 );
and ( n38586 , n38585 , n37541 );
xor ( n38587 , n38476 , n38521 );
and ( n38588 , n38587 , n37512 );
or ( n38589 , n38586 , n38588 );
not ( n38590 , n38589 );
buf ( n38591 , n38590 );
buf ( n38592 , n38591 );
not ( n38593 , n38592 );
not ( n38594 , n38593 );
not ( n38595 , n37512 );
and ( n38596 , n38595 , n37543 );
xor ( n38597 , n38477 , n38520 );
and ( n38598 , n38597 , n37512 );
or ( n38599 , n38596 , n38598 );
not ( n38600 , n38599 );
buf ( n38601 , n38600 );
buf ( n38602 , n38601 );
not ( n38603 , n38602 );
not ( n38604 , n38603 );
not ( n38605 , n37512 );
and ( n38606 , n38605 , n37545 );
xor ( n38607 , n38478 , n38519 );
and ( n38608 , n38607 , n37512 );
or ( n38609 , n38606 , n38608 );
not ( n38610 , n38609 );
buf ( n38611 , n38610 );
buf ( n38612 , n38611 );
not ( n38613 , n38612 );
not ( n38614 , n38613 );
not ( n38615 , n37512 );
and ( n38616 , n38615 , n37547 );
xor ( n38617 , n38479 , n38518 );
and ( n38618 , n38617 , n37512 );
or ( n38619 , n38616 , n38618 );
not ( n38620 , n38619 );
buf ( n38621 , n38620 );
buf ( n38622 , n38621 );
not ( n38623 , n38622 );
not ( n38624 , n38623 );
not ( n38625 , n37512 );
and ( n38626 , n38625 , n37549 );
xor ( n38627 , n38480 , n38517 );
and ( n38628 , n38627 , n37512 );
or ( n38629 , n38626 , n38628 );
not ( n38630 , n38629 );
buf ( n38631 , n38630 );
buf ( n38632 , n38631 );
not ( n38633 , n38632 );
not ( n38634 , n38633 );
not ( n38635 , n37512 );
and ( n38636 , n38635 , n37551 );
xor ( n38637 , n38481 , n38516 );
and ( n38638 , n38637 , n37512 );
or ( n38639 , n38636 , n38638 );
not ( n38640 , n38639 );
buf ( n38641 , n38640 );
buf ( n38642 , n38641 );
not ( n38643 , n38642 );
not ( n38644 , n38643 );
not ( n38645 , n37512 );
and ( n38646 , n38645 , n37553 );
xor ( n38647 , n38482 , n38515 );
and ( n38648 , n38647 , n37512 );
or ( n38649 , n38646 , n38648 );
not ( n38650 , n38649 );
buf ( n38651 , n38650 );
buf ( n38652 , n38651 );
not ( n38653 , n38652 );
not ( n38654 , n38653 );
not ( n38655 , n37512 );
and ( n38656 , n38655 , n37555 );
xor ( n38657 , n38483 , n38514 );
and ( n38658 , n38657 , n37512 );
or ( n38659 , n38656 , n38658 );
not ( n38660 , n38659 );
buf ( n38661 , n38660 );
buf ( n38662 , n38661 );
not ( n38663 , n38662 );
not ( n38664 , n38663 );
not ( n38665 , n37512 );
and ( n38666 , n38665 , n37557 );
xor ( n38667 , n38484 , n38513 );
and ( n38668 , n38667 , n37512 );
or ( n38669 , n38666 , n38668 );
not ( n38670 , n38669 );
buf ( n38671 , n38670 );
buf ( n38672 , n38671 );
not ( n38673 , n38672 );
not ( n38674 , n38673 );
not ( n38675 , n37512 );
and ( n38676 , n38675 , n37559 );
xor ( n38677 , n38485 , n38512 );
and ( n38678 , n38677 , n37512 );
or ( n38679 , n38676 , n38678 );
not ( n38680 , n38679 );
buf ( n38681 , n38680 );
buf ( n38682 , n38681 );
not ( n38683 , n38682 );
not ( n38684 , n38683 );
not ( n38685 , n37512 );
and ( n38686 , n38685 , n37561 );
xor ( n38687 , n38486 , n38511 );
and ( n38688 , n38687 , n37512 );
or ( n38689 , n38686 , n38688 );
not ( n38690 , n38689 );
buf ( n38691 , n38690 );
buf ( n38692 , n38691 );
not ( n38693 , n38692 );
not ( n38694 , n38693 );
not ( n38695 , n37512 );
and ( n38696 , n38695 , n37563 );
xor ( n38697 , n38487 , n38510 );
and ( n38698 , n38697 , n37512 );
or ( n38699 , n38696 , n38698 );
not ( n38700 , n38699 );
buf ( n38701 , n38700 );
buf ( n38702 , n38701 );
not ( n38703 , n38702 );
not ( n38704 , n38703 );
not ( n38705 , n37512 );
and ( n38706 , n38705 , n37565 );
xor ( n38707 , n38488 , n38509 );
and ( n38708 , n38707 , n37512 );
or ( n38709 , n38706 , n38708 );
not ( n38710 , n38709 );
buf ( n38711 , n38710 );
buf ( n38712 , n38711 );
not ( n38713 , n38712 );
not ( n38714 , n38713 );
not ( n38715 , n37512 );
and ( n38716 , n38715 , n37567 );
xor ( n38717 , n38489 , n38508 );
and ( n38718 , n38717 , n37512 );
or ( n38719 , n38716 , n38718 );
not ( n38720 , n38719 );
buf ( n38721 , n38720 );
buf ( n38722 , n38721 );
not ( n38723 , n38722 );
not ( n38724 , n38723 );
not ( n38725 , n37512 );
and ( n38726 , n38725 , n37569 );
xor ( n38727 , n38490 , n38507 );
and ( n38728 , n38727 , n37512 );
or ( n38729 , n38726 , n38728 );
not ( n38730 , n38729 );
buf ( n38731 , n38730 );
buf ( n38732 , n38731 );
not ( n38733 , n38732 );
not ( n38734 , n38733 );
not ( n38735 , n37512 );
and ( n38736 , n38735 , n37571 );
xor ( n38737 , n38491 , n38506 );
and ( n38738 , n38737 , n37512 );
or ( n38739 , n38736 , n38738 );
not ( n38740 , n38739 );
buf ( n38741 , n38740 );
buf ( n38742 , n38741 );
not ( n38743 , n38742 );
not ( n38744 , n38743 );
not ( n38745 , n37512 );
and ( n38746 , n38745 , n37573 );
xor ( n38747 , n38492 , n38505 );
and ( n38748 , n38747 , n37512 );
or ( n38749 , n38746 , n38748 );
not ( n38750 , n38749 );
buf ( n38751 , n38750 );
buf ( n38752 , n38751 );
not ( n38753 , n38752 );
not ( n38754 , n38753 );
not ( n38755 , n37512 );
and ( n38756 , n38755 , n32488 );
xor ( n38757 , n38493 , n38504 );
and ( n38758 , n38757 , n37512 );
or ( n38759 , n38756 , n38758 );
not ( n38760 , n38759 );
buf ( n38761 , n38760 );
buf ( n38762 , n38761 );
not ( n38763 , n38762 );
not ( n38764 , n38763 );
not ( n38765 , n37512 );
and ( n38766 , n38765 , n35677 );
xor ( n38767 , n38494 , n38503 );
and ( n38768 , n38767 , n37512 );
or ( n38769 , n38766 , n38768 );
not ( n38770 , n38769 );
buf ( n38771 , n38770 );
buf ( n38772 , n38771 );
not ( n38773 , n38772 );
not ( n38774 , n38773 );
not ( n38775 , n37512 );
and ( n38776 , n38775 , n37577 );
xor ( n38777 , n38495 , n38502 );
and ( n38778 , n38777 , n37512 );
or ( n38779 , n38776 , n38778 );
not ( n38780 , n38779 );
buf ( n38781 , n38780 );
buf ( n38782 , n38781 );
not ( n38783 , n38782 );
not ( n38784 , n38783 );
not ( n38785 , n37512 );
and ( n38786 , n38785 , n37579 );
xor ( n38787 , n38496 , n38501 );
and ( n38788 , n38787 , n37512 );
or ( n38789 , n38786 , n38788 );
not ( n38790 , n38789 );
buf ( n38791 , n38790 );
buf ( n38792 , n38791 );
not ( n38793 , n38792 );
not ( n38794 , n38793 );
not ( n38795 , n37512 );
and ( n38796 , n38795 , n37581 );
xor ( n38797 , n38497 , n38500 );
and ( n38798 , n38797 , n37512 );
or ( n38799 , n38796 , n38798 );
not ( n38800 , n38799 );
buf ( n38801 , n38800 );
buf ( n38802 , n38801 );
not ( n38803 , n38802 );
not ( n38804 , n38803 );
not ( n38805 , n37512 );
and ( n38806 , n38805 , n37583 );
xor ( n38807 , n38498 , n38499 );
and ( n38808 , n38807 , n37512 );
or ( n38809 , n38806 , n38808 );
not ( n38810 , n38809 );
buf ( n38811 , n38810 );
buf ( n38812 , n38811 );
not ( n38813 , n38812 );
not ( n38814 , n38813 );
not ( n38815 , n38464 );
and ( n38816 , n38814 , n38815 );
and ( n38817 , n38804 , n38816 );
and ( n38818 , n38794 , n38817 );
and ( n38819 , n38784 , n38818 );
and ( n38820 , n38774 , n38819 );
and ( n38821 , n38764 , n38820 );
and ( n38822 , n38754 , n38821 );
and ( n38823 , n38744 , n38822 );
and ( n38824 , n38734 , n38823 );
and ( n38825 , n38724 , n38824 );
and ( n38826 , n38714 , n38825 );
and ( n38827 , n38704 , n38826 );
and ( n38828 , n38694 , n38827 );
and ( n38829 , n38684 , n38828 );
and ( n38830 , n38674 , n38829 );
and ( n38831 , n38664 , n38830 );
and ( n38832 , n38654 , n38831 );
and ( n38833 , n38644 , n38832 );
and ( n38834 , n38634 , n38833 );
and ( n38835 , n38624 , n38834 );
and ( n38836 , n38614 , n38835 );
and ( n38837 , n38604 , n38836 );
and ( n38838 , n38594 , n38837 );
and ( n38839 , n38584 , n38838 );
and ( n38840 , n38574 , n38839 );
and ( n38841 , n38564 , n38840 );
and ( n38842 , n38554 , n38841 );
and ( n38843 , n38544 , n38842 );
and ( n38844 , n38534 , n38843 );
not ( n38845 , n38844 );
and ( n38846 , n38845 , n37512 );
buf ( n38847 , n38846 );
not ( n38848 , n38847 );
not ( n38849 , n37512 );
and ( n38850 , n38849 , n38813 );
xor ( n38851 , n38814 , n38815 );
and ( n38852 , n38851 , n37512 );
or ( n38853 , n38850 , n38852 );
and ( n38854 , n38848 , n38853 );
not ( n38855 , n38853 );
not ( n38856 , n38465 );
xor ( n38857 , n38855 , n38856 );
and ( n38858 , n38857 , n38847 );
or ( n38859 , n38854 , n38858 );
not ( n38860 , n38859 );
buf ( n38861 , n38860 );
buf ( n38862 , n38861 );
not ( n38863 , n38862 );
or ( n38864 , n38469 , n38863 );
not ( n38865 , n38847 );
not ( n38866 , n37512 );
and ( n38867 , n38866 , n38803 );
xor ( n38868 , n38804 , n38816 );
and ( n38869 , n38868 , n37512 );
or ( n38870 , n38867 , n38869 );
and ( n38871 , n38865 , n38870 );
not ( n38872 , n38870 );
and ( n38873 , n38855 , n38856 );
xor ( n38874 , n38872 , n38873 );
and ( n38875 , n38874 , n38847 );
or ( n38876 , n38871 , n38875 );
not ( n38877 , n38876 );
buf ( n38878 , n38877 );
buf ( n38879 , n38878 );
not ( n38880 , n38879 );
or ( n38881 , n38864 , n38880 );
not ( n38882 , n38847 );
not ( n38883 , n37512 );
and ( n38884 , n38883 , n38793 );
xor ( n38885 , n38794 , n38817 );
and ( n38886 , n38885 , n37512 );
or ( n38887 , n38884 , n38886 );
and ( n38888 , n38882 , n38887 );
not ( n38889 , n38887 );
and ( n38890 , n38872 , n38873 );
xor ( n38891 , n38889 , n38890 );
and ( n38892 , n38891 , n38847 );
or ( n38893 , n38888 , n38892 );
not ( n38894 , n38893 );
buf ( n38895 , n38894 );
buf ( n38896 , n38895 );
not ( n38897 , n38896 );
or ( n38898 , n38881 , n38897 );
not ( n38899 , n38847 );
not ( n38900 , n37512 );
and ( n38901 , n38900 , n38783 );
xor ( n38902 , n38784 , n38818 );
and ( n38903 , n38902 , n37512 );
or ( n38904 , n38901 , n38903 );
and ( n38905 , n38899 , n38904 );
not ( n38906 , n38904 );
and ( n38907 , n38889 , n38890 );
xor ( n38908 , n38906 , n38907 );
and ( n38909 , n38908 , n38847 );
or ( n38910 , n38905 , n38909 );
not ( n38911 , n38910 );
buf ( n38912 , n38911 );
buf ( n38913 , n38912 );
not ( n38914 , n38913 );
or ( n38915 , n38898 , n38914 );
not ( n38916 , n38847 );
not ( n38917 , n37512 );
and ( n38918 , n38917 , n38773 );
xor ( n38919 , n38774 , n38819 );
and ( n38920 , n38919 , n37512 );
or ( n38921 , n38918 , n38920 );
and ( n38922 , n38916 , n38921 );
not ( n38923 , n38921 );
and ( n38924 , n38906 , n38907 );
xor ( n38925 , n38923 , n38924 );
and ( n38926 , n38925 , n38847 );
or ( n38927 , n38922 , n38926 );
not ( n38928 , n38927 );
buf ( n38929 , n38928 );
buf ( n38930 , n38929 );
not ( n38931 , n38930 );
or ( n38932 , n38915 , n38931 );
not ( n38933 , n38847 );
not ( n38934 , n37512 );
and ( n38935 , n38934 , n38763 );
xor ( n38936 , n38764 , n38820 );
and ( n38937 , n38936 , n37512 );
or ( n38938 , n38935 , n38937 );
and ( n38939 , n38933 , n38938 );
not ( n38940 , n38938 );
and ( n38941 , n38923 , n38924 );
xor ( n38942 , n38940 , n38941 );
and ( n38943 , n38942 , n38847 );
or ( n38944 , n38939 , n38943 );
not ( n38945 , n38944 );
buf ( n38946 , n38945 );
buf ( n38947 , n38946 );
not ( n38948 , n38947 );
or ( n38949 , n38932 , n38948 );
not ( n38950 , n38847 );
not ( n38951 , n37512 );
and ( n38952 , n38951 , n38753 );
xor ( n38953 , n38754 , n38821 );
and ( n38954 , n38953 , n37512 );
or ( n38955 , n38952 , n38954 );
and ( n38956 , n38950 , n38955 );
not ( n38957 , n38955 );
and ( n38958 , n38940 , n38941 );
xor ( n38959 , n38957 , n38958 );
and ( n38960 , n38959 , n38847 );
or ( n38961 , n38956 , n38960 );
not ( n38962 , n38961 );
buf ( n38963 , n38962 );
buf ( n38964 , n38963 );
not ( n38965 , n38964 );
or ( n38966 , n38949 , n38965 );
not ( n38967 , n38847 );
not ( n38968 , n37512 );
and ( n38969 , n38968 , n38743 );
xor ( n38970 , n38744 , n38822 );
and ( n38971 , n38970 , n37512 );
or ( n38972 , n38969 , n38971 );
and ( n38973 , n38967 , n38972 );
not ( n38974 , n38972 );
and ( n38975 , n38957 , n38958 );
xor ( n38976 , n38974 , n38975 );
and ( n38977 , n38976 , n38847 );
or ( n38978 , n38973 , n38977 );
not ( n38979 , n38978 );
buf ( n38980 , n38979 );
buf ( n38981 , n38980 );
not ( n38982 , n38981 );
or ( n38983 , n38966 , n38982 );
not ( n38984 , n38847 );
not ( n38985 , n37512 );
and ( n38986 , n38985 , n38733 );
xor ( n38987 , n38734 , n38823 );
and ( n38988 , n38987 , n37512 );
or ( n38989 , n38986 , n38988 );
and ( n38990 , n38984 , n38989 );
not ( n38991 , n38989 );
and ( n38992 , n38974 , n38975 );
xor ( n38993 , n38991 , n38992 );
and ( n38994 , n38993 , n38847 );
or ( n38995 , n38990 , n38994 );
not ( n38996 , n38995 );
buf ( n38997 , n38996 );
buf ( n38998 , n38997 );
not ( n38999 , n38998 );
or ( n39000 , n38983 , n38999 );
not ( n39001 , n38847 );
not ( n39002 , n37512 );
and ( n39003 , n39002 , n38723 );
xor ( n39004 , n38724 , n38824 );
and ( n39005 , n39004 , n37512 );
or ( n39006 , n39003 , n39005 );
and ( n39007 , n39001 , n39006 );
not ( n39008 , n39006 );
and ( n39009 , n38991 , n38992 );
xor ( n39010 , n39008 , n39009 );
and ( n39011 , n39010 , n38847 );
or ( n39012 , n39007 , n39011 );
not ( n39013 , n39012 );
buf ( n39014 , n39013 );
buf ( n39015 , n39014 );
not ( n39016 , n39015 );
or ( n39017 , n39000 , n39016 );
not ( n39018 , n38847 );
not ( n39019 , n37512 );
and ( n39020 , n39019 , n38713 );
xor ( n39021 , n38714 , n38825 );
and ( n39022 , n39021 , n37512 );
or ( n39023 , n39020 , n39022 );
and ( n39024 , n39018 , n39023 );
not ( n39025 , n39023 );
and ( n39026 , n39008 , n39009 );
xor ( n39027 , n39025 , n39026 );
and ( n39028 , n39027 , n38847 );
or ( n39029 , n39024 , n39028 );
not ( n39030 , n39029 );
buf ( n39031 , n39030 );
buf ( n39032 , n39031 );
not ( n39033 , n39032 );
or ( n39034 , n39017 , n39033 );
not ( n39035 , n38847 );
not ( n39036 , n37512 );
and ( n39037 , n39036 , n38703 );
xor ( n39038 , n38704 , n38826 );
and ( n39039 , n39038 , n37512 );
or ( n39040 , n39037 , n39039 );
and ( n39041 , n39035 , n39040 );
not ( n39042 , n39040 );
and ( n39043 , n39025 , n39026 );
xor ( n39044 , n39042 , n39043 );
and ( n39045 , n39044 , n38847 );
or ( n39046 , n39041 , n39045 );
not ( n39047 , n39046 );
buf ( n39048 , n39047 );
buf ( n39049 , n39048 );
not ( n39050 , n39049 );
or ( n39051 , n39034 , n39050 );
not ( n39052 , n38847 );
not ( n39053 , n37512 );
and ( n39054 , n39053 , n38693 );
xor ( n39055 , n38694 , n38827 );
and ( n39056 , n39055 , n37512 );
or ( n39057 , n39054 , n39056 );
and ( n39058 , n39052 , n39057 );
not ( n39059 , n39057 );
and ( n39060 , n39042 , n39043 );
xor ( n39061 , n39059 , n39060 );
and ( n39062 , n39061 , n38847 );
or ( n39063 , n39058 , n39062 );
not ( n39064 , n39063 );
buf ( n39065 , n39064 );
buf ( n39066 , n39065 );
not ( n39067 , n39066 );
or ( n39068 , n39051 , n39067 );
not ( n39069 , n38847 );
not ( n39070 , n37512 );
and ( n39071 , n39070 , n38683 );
xor ( n39072 , n38684 , n38828 );
and ( n39073 , n39072 , n37512 );
or ( n39074 , n39071 , n39073 );
and ( n39075 , n39069 , n39074 );
not ( n39076 , n39074 );
and ( n39077 , n39059 , n39060 );
xor ( n39078 , n39076 , n39077 );
and ( n39079 , n39078 , n38847 );
or ( n39080 , n39075 , n39079 );
not ( n39081 , n39080 );
buf ( n39082 , n39081 );
buf ( n39083 , n39082 );
not ( n39084 , n39083 );
or ( n39085 , n39068 , n39084 );
not ( n39086 , n38847 );
not ( n39087 , n37512 );
and ( n39088 , n39087 , n38673 );
xor ( n39089 , n38674 , n38829 );
and ( n39090 , n39089 , n37512 );
or ( n39091 , n39088 , n39090 );
and ( n39092 , n39086 , n39091 );
not ( n39093 , n39091 );
and ( n39094 , n39076 , n39077 );
xor ( n39095 , n39093 , n39094 );
and ( n39096 , n39095 , n38847 );
or ( n39097 , n39092 , n39096 );
not ( n39098 , n39097 );
buf ( n39099 , n39098 );
buf ( n39100 , n39099 );
not ( n39101 , n39100 );
or ( n39102 , n39085 , n39101 );
not ( n39103 , n38847 );
not ( n39104 , n37512 );
and ( n39105 , n39104 , n38663 );
xor ( n39106 , n38664 , n38830 );
and ( n39107 , n39106 , n37512 );
or ( n39108 , n39105 , n39107 );
and ( n39109 , n39103 , n39108 );
not ( n39110 , n39108 );
and ( n39111 , n39093 , n39094 );
xor ( n39112 , n39110 , n39111 );
and ( n39113 , n39112 , n38847 );
or ( n39114 , n39109 , n39113 );
not ( n39115 , n39114 );
buf ( n39116 , n39115 );
buf ( n39117 , n39116 );
not ( n39118 , n39117 );
or ( n39119 , n39102 , n39118 );
not ( n39120 , n38847 );
not ( n39121 , n37512 );
and ( n39122 , n39121 , n38653 );
xor ( n39123 , n38654 , n38831 );
and ( n39124 , n39123 , n37512 );
or ( n39125 , n39122 , n39124 );
and ( n39126 , n39120 , n39125 );
not ( n39127 , n39125 );
and ( n39128 , n39110 , n39111 );
xor ( n39129 , n39127 , n39128 );
and ( n39130 , n39129 , n38847 );
or ( n39131 , n39126 , n39130 );
not ( n39132 , n39131 );
buf ( n39133 , n39132 );
buf ( n39134 , n39133 );
not ( n39135 , n39134 );
or ( n39136 , n39119 , n39135 );
not ( n39137 , n38847 );
not ( n39138 , n37512 );
and ( n39139 , n39138 , n38643 );
xor ( n39140 , n38644 , n38832 );
and ( n39141 , n39140 , n37512 );
or ( n39142 , n39139 , n39141 );
and ( n39143 , n39137 , n39142 );
not ( n39144 , n39142 );
and ( n39145 , n39127 , n39128 );
xor ( n39146 , n39144 , n39145 );
and ( n39147 , n39146 , n38847 );
or ( n39148 , n39143 , n39147 );
not ( n39149 , n39148 );
buf ( n39150 , n39149 );
buf ( n39151 , n39150 );
not ( n39152 , n39151 );
or ( n39153 , n39136 , n39152 );
not ( n39154 , n38847 );
not ( n39155 , n37512 );
and ( n39156 , n39155 , n38633 );
xor ( n39157 , n38634 , n38833 );
and ( n39158 , n39157 , n37512 );
or ( n39159 , n39156 , n39158 );
and ( n39160 , n39154 , n39159 );
not ( n39161 , n39159 );
and ( n39162 , n39144 , n39145 );
xor ( n39163 , n39161 , n39162 );
and ( n39164 , n39163 , n38847 );
or ( n39165 , n39160 , n39164 );
not ( n39166 , n39165 );
buf ( n39167 , n39166 );
buf ( n39168 , n39167 );
not ( n39169 , n39168 );
or ( n39170 , n39153 , n39169 );
not ( n39171 , n38847 );
not ( n39172 , n37512 );
and ( n39173 , n39172 , n38623 );
xor ( n39174 , n38624 , n38834 );
and ( n39175 , n39174 , n37512 );
or ( n39176 , n39173 , n39175 );
and ( n39177 , n39171 , n39176 );
not ( n39178 , n39176 );
and ( n39179 , n39161 , n39162 );
xor ( n39180 , n39178 , n39179 );
and ( n39181 , n39180 , n38847 );
or ( n39182 , n39177 , n39181 );
not ( n39183 , n39182 );
buf ( n39184 , n39183 );
buf ( n39185 , n39184 );
not ( n39186 , n39185 );
or ( n39187 , n39170 , n39186 );
not ( n39188 , n38847 );
not ( n39189 , n37512 );
and ( n39190 , n39189 , n38613 );
xor ( n39191 , n38614 , n38835 );
and ( n39192 , n39191 , n37512 );
or ( n39193 , n39190 , n39192 );
and ( n39194 , n39188 , n39193 );
not ( n39195 , n39193 );
and ( n39196 , n39178 , n39179 );
xor ( n39197 , n39195 , n39196 );
and ( n39198 , n39197 , n38847 );
or ( n39199 , n39194 , n39198 );
not ( n39200 , n39199 );
buf ( n39201 , n39200 );
buf ( n39202 , n39201 );
not ( n39203 , n39202 );
or ( n39204 , n39187 , n39203 );
not ( n39205 , n38847 );
not ( n39206 , n37512 );
and ( n39207 , n39206 , n38603 );
xor ( n39208 , n38604 , n38836 );
and ( n39209 , n39208 , n37512 );
or ( n39210 , n39207 , n39209 );
and ( n39211 , n39205 , n39210 );
not ( n39212 , n39210 );
and ( n39213 , n39195 , n39196 );
xor ( n39214 , n39212 , n39213 );
and ( n39215 , n39214 , n38847 );
or ( n39216 , n39211 , n39215 );
not ( n39217 , n39216 );
buf ( n39218 , n39217 );
buf ( n39219 , n39218 );
not ( n39220 , n39219 );
or ( n39221 , n39204 , n39220 );
not ( n39222 , n38847 );
not ( n39223 , n37512 );
and ( n39224 , n39223 , n38593 );
xor ( n39225 , n38594 , n38837 );
and ( n39226 , n39225 , n37512 );
or ( n39227 , n39224 , n39226 );
and ( n39228 , n39222 , n39227 );
not ( n39229 , n39227 );
and ( n39230 , n39212 , n39213 );
xor ( n39231 , n39229 , n39230 );
and ( n39232 , n39231 , n38847 );
or ( n39233 , n39228 , n39232 );
not ( n39234 , n39233 );
buf ( n39235 , n39234 );
buf ( n39236 , n39235 );
not ( n39237 , n39236 );
or ( n39238 , n39221 , n39237 );
not ( n39239 , n38847 );
not ( n39240 , n37512 );
and ( n39241 , n39240 , n38583 );
xor ( n39242 , n38584 , n38838 );
and ( n39243 , n39242 , n37512 );
or ( n39244 , n39241 , n39243 );
and ( n39245 , n39239 , n39244 );
not ( n39246 , n39244 );
and ( n39247 , n39229 , n39230 );
xor ( n39248 , n39246 , n39247 );
and ( n39249 , n39248 , n38847 );
or ( n39250 , n39245 , n39249 );
not ( n39251 , n39250 );
buf ( n39252 , n39251 );
buf ( n39253 , n39252 );
not ( n39254 , n39253 );
or ( n39255 , n39238 , n39254 );
not ( n39256 , n38847 );
not ( n39257 , n37512 );
and ( n39258 , n39257 , n38573 );
xor ( n39259 , n38574 , n38839 );
and ( n39260 , n39259 , n37512 );
or ( n39261 , n39258 , n39260 );
and ( n39262 , n39256 , n39261 );
not ( n39263 , n39261 );
and ( n39264 , n39246 , n39247 );
xor ( n39265 , n39263 , n39264 );
and ( n39266 , n39265 , n38847 );
or ( n39267 , n39262 , n39266 );
not ( n39268 , n39267 );
buf ( n39269 , n39268 );
buf ( n39270 , n39269 );
not ( n39271 , n39270 );
or ( n39272 , n39255 , n39271 );
not ( n39273 , n38847 );
not ( n39274 , n37512 );
and ( n39275 , n39274 , n38563 );
xor ( n39276 , n38564 , n38840 );
and ( n39277 , n39276 , n37512 );
or ( n39278 , n39275 , n39277 );
and ( n39279 , n39273 , n39278 );
not ( n39280 , n39278 );
and ( n39281 , n39263 , n39264 );
xor ( n39282 , n39280 , n39281 );
and ( n39283 , n39282 , n38847 );
or ( n39284 , n39279 , n39283 );
not ( n39285 , n39284 );
buf ( n39286 , n39285 );
buf ( n39287 , n39286 );
not ( n39288 , n39287 );
or ( n39289 , n39272 , n39288 );
not ( n39290 , n38847 );
not ( n39291 , n37512 );
and ( n39292 , n39291 , n38553 );
xor ( n39293 , n38554 , n38841 );
and ( n39294 , n39293 , n37512 );
or ( n39295 , n39292 , n39294 );
and ( n39296 , n39290 , n39295 );
not ( n39297 , n39295 );
and ( n39298 , n39280 , n39281 );
xor ( n39299 , n39297 , n39298 );
and ( n39300 , n39299 , n38847 );
or ( n39301 , n39296 , n39300 );
not ( n39302 , n39301 );
buf ( n39303 , n39302 );
buf ( n39304 , n39303 );
not ( n39305 , n39304 );
or ( n39306 , n39289 , n39305 );
not ( n39307 , n38847 );
not ( n39308 , n37512 );
and ( n39309 , n39308 , n38543 );
xor ( n39310 , n38544 , n38842 );
and ( n39311 , n39310 , n37512 );
or ( n39312 , n39309 , n39311 );
and ( n39313 , n39307 , n39312 );
not ( n39314 , n39312 );
and ( n39315 , n39297 , n39298 );
xor ( n39316 , n39314 , n39315 );
and ( n39317 , n39316 , n38847 );
or ( n39318 , n39313 , n39317 );
not ( n39319 , n39318 );
buf ( n39320 , n39319 );
buf ( n39321 , n39320 );
not ( n39322 , n39321 );
or ( n39323 , n39306 , n39322 );
xor ( n39324 , n38534 , n38843 );
and ( n39325 , n39324 , n37512 );
buf ( n39326 , n39325 );
not ( n39327 , n39326 );
and ( n39328 , n39314 , n39315 );
xor ( n39329 , n39327 , n39328 );
and ( n39330 , n39329 , n38847 );
buf ( n39331 , n39330 );
not ( n39332 , n39331 );
buf ( n39333 , n39332 );
buf ( n39334 , n39333 );
not ( n39335 , n39334 );
or ( n39336 , n39323 , n39335 );
buf ( n39337 , n39336 );
buf ( n39338 , n39337 );
and ( n39339 , n39338 , n38847 );
not ( n39340 , n39339 );
and ( n39341 , n39340 , n38469 );
xor ( n39342 , n38469 , n38847 );
xor ( n39343 , n39342 , n38847 );
and ( n39344 , n39343 , n39339 );
or ( n39345 , n39341 , n39344 );
nor ( n39346 , n35281 , n35283 , n35284 );
and ( n39347 , n39345 , n39346 );
buf ( n39348 , RI15b5d948_1058);
nor ( n39349 , n35286 , n35282 , n35284 );
nor ( n39350 , n35281 , n35282 , n35284 );
or ( n39351 , n39349 , n39350 );
nor ( n39352 , n35286 , n35283 , n35284 );
or ( n39353 , n39351 , n39352 );
and ( n39354 , n35286 , n35283 , n35284 );
or ( n39355 , n39353 , n39354 );
and ( n39356 , n35281 , n35283 , n35284 );
or ( n39357 , n39355 , n39356 );
and ( n39358 , n35281 , n35282 , n35284 );
or ( n39359 , n39357 , n39358 );
and ( n39360 , n39348 , n39359 );
or ( n39361 , n38451 , n39347 , n39360 );
buf ( n39362 , n39361 );
buf ( n39363 , n39362 );
buf ( n39364 , n31655 );
buf ( n39365 , n30987 );
not ( n39366 , n32953 );
buf ( n39367 , RI15b467e8_270);
and ( n39368 , n39366 , n39367 );
buf ( n39369 , RI15b48480_331);
buf ( n39370 , n39369 );
not ( n39371 , n39370 );
buf ( n39372 , n39371 );
not ( n39373 , n39372 );
buf ( n39374 , RI15b49308_362);
not ( n39375 , n39374 );
buf ( n39376 , RI15b484f8_332);
and ( n39377 , n39375 , n39376 );
not ( n39378 , n39376 );
not ( n39379 , n39369 );
xor ( n39380 , n39378 , n39379 );
and ( n39381 , n39380 , n39374 );
or ( n39382 , n39377 , n39381 );
not ( n39383 , n39382 );
buf ( n39384 , n39383 );
buf ( n39385 , n39384 );
not ( n39386 , n39385 );
or ( n39387 , n39373 , n39386 );
not ( n39388 , n39374 );
buf ( n39389 , RI15b48570_333);
and ( n39390 , n39388 , n39389 );
not ( n39391 , n39389 );
and ( n39392 , n39378 , n39379 );
xor ( n39393 , n39391 , n39392 );
and ( n39394 , n39393 , n39374 );
or ( n39395 , n39390 , n39394 );
not ( n39396 , n39395 );
buf ( n39397 , n39396 );
buf ( n39398 , n39397 );
not ( n39399 , n39398 );
or ( n39400 , n39387 , n39399 );
not ( n39401 , n39374 );
buf ( n39402 , RI15b485e8_334);
and ( n39403 , n39401 , n39402 );
not ( n39404 , n39402 );
and ( n39405 , n39391 , n39392 );
xor ( n39406 , n39404 , n39405 );
and ( n39407 , n39406 , n39374 );
or ( n39408 , n39403 , n39407 );
not ( n39409 , n39408 );
buf ( n39410 , n39409 );
buf ( n39411 , n39410 );
not ( n39412 , n39411 );
or ( n39413 , n39400 , n39412 );
not ( n39414 , n39374 );
buf ( n39415 , RI15b48660_335);
and ( n39416 , n39414 , n39415 );
not ( n39417 , n39415 );
and ( n39418 , n39404 , n39405 );
xor ( n39419 , n39417 , n39418 );
and ( n39420 , n39419 , n39374 );
or ( n39421 , n39416 , n39420 );
not ( n39422 , n39421 );
buf ( n39423 , n39422 );
buf ( n39424 , n39423 );
not ( n39425 , n39424 );
or ( n39426 , n39413 , n39425 );
not ( n39427 , n39374 );
buf ( n39428 , RI15b486d8_336);
and ( n39429 , n39427 , n39428 );
not ( n39430 , n39428 );
and ( n39431 , n39417 , n39418 );
xor ( n39432 , n39430 , n39431 );
and ( n39433 , n39432 , n39374 );
or ( n39434 , n39429 , n39433 );
not ( n39435 , n39434 );
buf ( n39436 , n39435 );
buf ( n39437 , n39436 );
not ( n39438 , n39437 );
or ( n39439 , n39426 , n39438 );
not ( n39440 , n39374 );
buf ( n39441 , RI15b48750_337);
and ( n39442 , n39440 , n39441 );
not ( n39443 , n39441 );
and ( n39444 , n39430 , n39431 );
xor ( n39445 , n39443 , n39444 );
and ( n39446 , n39445 , n39374 );
or ( n39447 , n39442 , n39446 );
not ( n39448 , n39447 );
buf ( n39449 , n39448 );
buf ( n39450 , n39449 );
not ( n39451 , n39450 );
or ( n39452 , n39439 , n39451 );
not ( n39453 , n39374 );
buf ( n39454 , RI15b487c8_338);
and ( n39455 , n39453 , n39454 );
not ( n39456 , n39454 );
and ( n39457 , n39443 , n39444 );
xor ( n39458 , n39456 , n39457 );
and ( n39459 , n39458 , n39374 );
or ( n39460 , n39455 , n39459 );
not ( n39461 , n39460 );
buf ( n39462 , n39461 );
buf ( n39463 , n39462 );
not ( n39464 , n39463 );
or ( n39465 , n39452 , n39464 );
not ( n39466 , n39374 );
buf ( n39467 , RI15b48840_339);
and ( n39468 , n39466 , n39467 );
not ( n39469 , n39467 );
and ( n39470 , n39456 , n39457 );
xor ( n39471 , n39469 , n39470 );
and ( n39472 , n39471 , n39374 );
or ( n39473 , n39468 , n39472 );
not ( n39474 , n39473 );
buf ( n39475 , n39474 );
buf ( n39476 , n39475 );
not ( n39477 , n39476 );
or ( n39478 , n39465 , n39477 );
not ( n39479 , n39374 );
buf ( n39480 , RI15b488b8_340);
and ( n39481 , n39479 , n39480 );
not ( n39482 , n39480 );
and ( n39483 , n39469 , n39470 );
xor ( n39484 , n39482 , n39483 );
and ( n39485 , n39484 , n39374 );
or ( n39486 , n39481 , n39485 );
not ( n39487 , n39486 );
buf ( n39488 , n39487 );
buf ( n39489 , n39488 );
not ( n39490 , n39489 );
or ( n39491 , n39478 , n39490 );
not ( n39492 , n39374 );
buf ( n39493 , RI15b48930_341);
and ( n39494 , n39492 , n39493 );
not ( n39495 , n39493 );
and ( n39496 , n39482 , n39483 );
xor ( n39497 , n39495 , n39496 );
and ( n39498 , n39497 , n39374 );
or ( n39499 , n39494 , n39498 );
not ( n39500 , n39499 );
buf ( n39501 , n39500 );
buf ( n39502 , n39501 );
not ( n39503 , n39502 );
or ( n39504 , n39491 , n39503 );
not ( n39505 , n39374 );
buf ( n39506 , RI15b489a8_342);
and ( n39507 , n39505 , n39506 );
not ( n39508 , n39506 );
and ( n39509 , n39495 , n39496 );
xor ( n39510 , n39508 , n39509 );
and ( n39511 , n39510 , n39374 );
or ( n39512 , n39507 , n39511 );
not ( n39513 , n39512 );
buf ( n39514 , n39513 );
buf ( n39515 , n39514 );
not ( n39516 , n39515 );
or ( n39517 , n39504 , n39516 );
not ( n39518 , n39374 );
buf ( n39519 , RI15b48a20_343);
and ( n39520 , n39518 , n39519 );
not ( n39521 , n39519 );
and ( n39522 , n39508 , n39509 );
xor ( n39523 , n39521 , n39522 );
and ( n39524 , n39523 , n39374 );
or ( n39525 , n39520 , n39524 );
not ( n39526 , n39525 );
buf ( n39527 , n39526 );
buf ( n39528 , n39527 );
not ( n39529 , n39528 );
or ( n39530 , n39517 , n39529 );
not ( n39531 , n39374 );
buf ( n39532 , RI15b48a98_344);
and ( n39533 , n39531 , n39532 );
not ( n39534 , n39532 );
and ( n39535 , n39521 , n39522 );
xor ( n39536 , n39534 , n39535 );
and ( n39537 , n39536 , n39374 );
or ( n39538 , n39533 , n39537 );
not ( n39539 , n39538 );
buf ( n39540 , n39539 );
buf ( n39541 , n39540 );
not ( n39542 , n39541 );
or ( n39543 , n39530 , n39542 );
not ( n39544 , n39374 );
buf ( n39545 , RI15b48b10_345);
and ( n39546 , n39544 , n39545 );
not ( n39547 , n39545 );
and ( n39548 , n39534 , n39535 );
xor ( n39549 , n39547 , n39548 );
and ( n39550 , n39549 , n39374 );
or ( n39551 , n39546 , n39550 );
not ( n39552 , n39551 );
buf ( n39553 , n39552 );
buf ( n39554 , n39553 );
not ( n39555 , n39554 );
or ( n39556 , n39543 , n39555 );
not ( n39557 , n39374 );
buf ( n39558 , RI15b48b88_346);
and ( n39559 , n39557 , n39558 );
not ( n39560 , n39558 );
and ( n39561 , n39547 , n39548 );
xor ( n39562 , n39560 , n39561 );
and ( n39563 , n39562 , n39374 );
or ( n39564 , n39559 , n39563 );
not ( n39565 , n39564 );
buf ( n39566 , n39565 );
buf ( n39567 , n39566 );
not ( n39568 , n39567 );
or ( n39569 , n39556 , n39568 );
buf ( n39570 , n39569 );
buf ( n39571 , n39570 );
and ( n39572 , n39571 , n39374 );
not ( n39573 , n39572 );
and ( n39574 , n39573 , n39386 );
xor ( n39575 , n39386 , n39374 );
xor ( n39576 , n39373 , n39374 );
and ( n39577 , n39576 , n39374 );
xor ( n39578 , n39575 , n39577 );
and ( n39579 , n39578 , n39572 );
or ( n39580 , n39574 , n39579 );
and ( n39581 , n39580 , n32953 );
or ( n39582 , n39368 , n39581 );
and ( n39583 , n39582 , n33038 );
or ( n39584 , n32968 , n32967 );
and ( n39585 , n32967 , n39584 );
and ( n39586 , n33067 , n39585 );
not ( n39587 , n39586 );
and ( n39588 , n39587 , n39367 );
buf ( n39589 , n34188 );
not ( n39590 , n39589 );
buf ( n39591 , n39590 );
not ( n39592 , n39591 );
not ( n39593 , n34193 );
and ( n39594 , n39593 , n34195 );
not ( n39595 , n34195 );
not ( n39596 , n34188 );
xor ( n39597 , n39595 , n39596 );
and ( n39598 , n39597 , n34193 );
or ( n39599 , n39594 , n39598 );
not ( n39600 , n39599 );
buf ( n39601 , n39600 );
buf ( n39602 , n39601 );
not ( n39603 , n39602 );
or ( n39604 , n39592 , n39603 );
not ( n39605 , n34193 );
and ( n39606 , n39605 , n34208 );
not ( n39607 , n34208 );
and ( n39608 , n39595 , n39596 );
xor ( n39609 , n39607 , n39608 );
and ( n39610 , n39609 , n34193 );
or ( n39611 , n39606 , n39610 );
not ( n39612 , n39611 );
buf ( n39613 , n39612 );
buf ( n39614 , n39613 );
not ( n39615 , n39614 );
or ( n39616 , n39604 , n39615 );
not ( n39617 , n34193 );
and ( n39618 , n39617 , n34221 );
not ( n39619 , n34221 );
and ( n39620 , n39607 , n39608 );
xor ( n39621 , n39619 , n39620 );
and ( n39622 , n39621 , n34193 );
or ( n39623 , n39618 , n39622 );
not ( n39624 , n39623 );
buf ( n39625 , n39624 );
buf ( n39626 , n39625 );
not ( n39627 , n39626 );
or ( n39628 , n39616 , n39627 );
not ( n39629 , n34193 );
and ( n39630 , n39629 , n34234 );
not ( n39631 , n34234 );
and ( n39632 , n39619 , n39620 );
xor ( n39633 , n39631 , n39632 );
and ( n39634 , n39633 , n34193 );
or ( n39635 , n39630 , n39634 );
not ( n39636 , n39635 );
buf ( n39637 , n39636 );
buf ( n39638 , n39637 );
not ( n39639 , n39638 );
or ( n39640 , n39628 , n39639 );
not ( n39641 , n34193 );
and ( n39642 , n39641 , n34247 );
not ( n39643 , n34247 );
and ( n39644 , n39631 , n39632 );
xor ( n39645 , n39643 , n39644 );
and ( n39646 , n39645 , n34193 );
or ( n39647 , n39642 , n39646 );
not ( n39648 , n39647 );
buf ( n39649 , n39648 );
buf ( n39650 , n39649 );
not ( n39651 , n39650 );
or ( n39652 , n39640 , n39651 );
not ( n39653 , n34193 );
and ( n39654 , n39653 , n34260 );
not ( n39655 , n34260 );
and ( n39656 , n39643 , n39644 );
xor ( n39657 , n39655 , n39656 );
and ( n39658 , n39657 , n34193 );
or ( n39659 , n39654 , n39658 );
not ( n39660 , n39659 );
buf ( n39661 , n39660 );
buf ( n39662 , n39661 );
not ( n39663 , n39662 );
or ( n39664 , n39652 , n39663 );
not ( n39665 , n34193 );
and ( n39666 , n39665 , n34273 );
not ( n39667 , n34273 );
and ( n39668 , n39655 , n39656 );
xor ( n39669 , n39667 , n39668 );
and ( n39670 , n39669 , n34193 );
or ( n39671 , n39666 , n39670 );
not ( n39672 , n39671 );
buf ( n39673 , n39672 );
buf ( n39674 , n39673 );
not ( n39675 , n39674 );
or ( n39676 , n39664 , n39675 );
not ( n39677 , n34193 );
and ( n39678 , n39677 , n34379 );
not ( n39679 , n34379 );
and ( n39680 , n39667 , n39668 );
xor ( n39681 , n39679 , n39680 );
and ( n39682 , n39681 , n34193 );
or ( n39683 , n39678 , n39682 );
not ( n39684 , n39683 );
buf ( n39685 , n39684 );
buf ( n39686 , n39685 );
not ( n39687 , n39686 );
or ( n39688 , n39676 , n39687 );
not ( n39689 , n34193 );
and ( n39690 , n39689 , n34377 );
not ( n39691 , n34377 );
and ( n39692 , n39679 , n39680 );
xor ( n39693 , n39691 , n39692 );
and ( n39694 , n39693 , n34193 );
or ( n39695 , n39690 , n39694 );
not ( n39696 , n39695 );
buf ( n39697 , n39696 );
buf ( n39698 , n39697 );
not ( n39699 , n39698 );
or ( n39700 , n39688 , n39699 );
not ( n39701 , n34193 );
and ( n39702 , n39701 , n34375 );
not ( n39703 , n34375 );
and ( n39704 , n39691 , n39692 );
xor ( n39705 , n39703 , n39704 );
and ( n39706 , n39705 , n34193 );
or ( n39707 , n39702 , n39706 );
not ( n39708 , n39707 );
buf ( n39709 , n39708 );
buf ( n39710 , n39709 );
not ( n39711 , n39710 );
or ( n39712 , n39700 , n39711 );
not ( n39713 , n34193 );
and ( n39714 , n39713 , n34373 );
not ( n39715 , n34373 );
and ( n39716 , n39703 , n39704 );
xor ( n39717 , n39715 , n39716 );
and ( n39718 , n39717 , n34193 );
or ( n39719 , n39714 , n39718 );
not ( n39720 , n39719 );
buf ( n39721 , n39720 );
buf ( n39722 , n39721 );
not ( n39723 , n39722 );
or ( n39724 , n39712 , n39723 );
not ( n39725 , n34193 );
and ( n39726 , n39725 , n34371 );
not ( n39727 , n34371 );
and ( n39728 , n39715 , n39716 );
xor ( n39729 , n39727 , n39728 );
and ( n39730 , n39729 , n34193 );
or ( n39731 , n39726 , n39730 );
not ( n39732 , n39731 );
buf ( n39733 , n39732 );
buf ( n39734 , n39733 );
not ( n39735 , n39734 );
or ( n39736 , n39724 , n39735 );
not ( n39737 , n34193 );
and ( n39738 , n39737 , n34369 );
not ( n39739 , n34369 );
and ( n39740 , n39727 , n39728 );
xor ( n39741 , n39739 , n39740 );
and ( n39742 , n39741 , n34193 );
or ( n39743 , n39738 , n39742 );
not ( n39744 , n39743 );
buf ( n39745 , n39744 );
buf ( n39746 , n39745 );
not ( n39747 , n39746 );
or ( n39748 , n39736 , n39747 );
not ( n39749 , n34193 );
and ( n39750 , n39749 , n34367 );
not ( n39751 , n34367 );
and ( n39752 , n39739 , n39740 );
xor ( n39753 , n39751 , n39752 );
and ( n39754 , n39753 , n34193 );
or ( n39755 , n39750 , n39754 );
not ( n39756 , n39755 );
buf ( n39757 , n39756 );
buf ( n39758 , n39757 );
not ( n39759 , n39758 );
or ( n39760 , n39748 , n39759 );
not ( n39761 , n34193 );
and ( n39762 , n39761 , n34365 );
not ( n39763 , n34365 );
and ( n39764 , n39751 , n39752 );
xor ( n39765 , n39763 , n39764 );
and ( n39766 , n39765 , n34193 );
or ( n39767 , n39762 , n39766 );
not ( n39768 , n39767 );
buf ( n39769 , n39768 );
buf ( n39770 , n39769 );
not ( n39771 , n39770 );
or ( n39772 , n39760 , n39771 );
buf ( n39773 , n39772 );
buf ( n39774 , n39773 );
and ( n39775 , n39774 , n34193 );
not ( n39776 , n39775 );
and ( n39777 , n39776 , n39603 );
xor ( n39778 , n39603 , n34193 );
xor ( n39779 , n39592 , n34193 );
and ( n39780 , n39779 , n34193 );
xor ( n39781 , n39778 , n39780 );
and ( n39782 , n39781 , n39775 );
or ( n39783 , n39777 , n39782 );
and ( n39784 , n39783 , n39586 );
or ( n39785 , n39588 , n39784 );
and ( n39786 , n39785 , n33172 );
or ( n39787 , n33190 , n32924 );
or ( n39788 , n39787 , n32890 );
or ( n39789 , n39788 , n33191 );
or ( n39790 , n39789 , n33193 );
or ( n39791 , n39790 , n33195 );
or ( n39792 , n39791 , n33197 );
or ( n39793 , n39792 , n33199 );
or ( n39794 , n39793 , n33201 );
or ( n39795 , n39794 , n33203 );
and ( n39796 , n39367 , n39795 );
or ( n39797 , n39583 , n39786 , n39796 );
and ( n39798 , n39797 , n33208 );
or ( n39799 , n35057 , n33370 );
or ( n39800 , n39799 , n33373 );
or ( n39801 , n39800 , n33375 );
or ( n39802 , n39801 , n33377 );
or ( n39803 , n39802 , n33379 );
or ( n39804 , n39803 , n33381 );
or ( n39805 , n39804 , n32528 );
and ( n39806 , n39367 , n39805 );
or ( n39807 , C0 , n39798 , n39806 );
buf ( n39808 , n39807 );
buf ( n39809 , n39808 );
buf ( n39810 , n30987 );
buf ( n39811 , n31655 );
buf ( n39812 , n30987 );
and ( n39813 , n31587 , n31007 );
not ( n39814 , n31077 );
and ( n39815 , n39814 , n34011 );
and ( n39816 , n31014 , n31082 );
xor ( n39817 , n31010 , n39816 );
and ( n39818 , n39817 , n31077 );
or ( n39819 , n39815 , n39818 );
and ( n39820 , n39819 , n31373 );
not ( n39821 , n31402 );
and ( n39822 , n39821 , n34011 );
and ( n39823 , n39817 , n31402 );
or ( n39824 , n39822 , n39823 );
and ( n39825 , n39824 , n31408 );
not ( n39826 , n31437 );
and ( n39827 , n39826 , n34011 );
not ( n39828 , n31455 );
and ( n39829 , n39828 , n34062 );
xor ( n39830 , n34011 , n34012 );
and ( n39831 , n39830 , n31455 );
or ( n39832 , n39829 , n39831 );
and ( n39833 , n39832 , n31437 );
or ( n39834 , n39827 , n39833 );
and ( n39835 , n39834 , n31468 );
not ( n39836 , n31497 );
and ( n39837 , n39836 , n34011 );
not ( n39838 , n31454 );
not ( n39839 , n31501 );
and ( n39840 , n39839 , n34062 );
xor ( n39841 , n34063 , n34064 );
and ( n39842 , n39841 , n31501 );
or ( n39843 , n39840 , n39842 );
and ( n39844 , n39838 , n39843 );
and ( n39845 , n39830 , n31454 );
or ( n39846 , n39844 , n39845 );
and ( n39847 , n39846 , n31497 );
or ( n39848 , n39837 , n39847 );
and ( n39849 , n39848 , n31521 );
and ( n39850 , n34011 , n31553 );
or ( n39851 , n39820 , n39825 , n39835 , n39849 , n39850 );
and ( n39852 , n39851 , n31557 );
not ( n39853 , n31452 );
not ( n39854 , n31619 );
and ( n39855 , n39854 , n34119 );
xor ( n39856 , n34120 , n34121 );
and ( n39857 , n39856 , n31619 );
or ( n39858 , n39855 , n39857 );
and ( n39859 , n39853 , n39858 );
and ( n39860 , n34011 , n31452 );
or ( n39861 , n39859 , n39860 );
and ( n39862 , n39861 , n31638 );
buf ( n39863 , n33973 );
and ( n39864 , n34011 , n31650 );
or ( n39865 , C0 , n39813 , n39852 , n39862 , n39863 , n39864 );
buf ( n39866 , n39865 );
buf ( n39867 , n39866 );
buf ( n39868 , n31655 );
buf ( n39869 , n31655 );
and ( n39870 , n31588 , n31007 );
not ( n39871 , n31077 );
and ( n39872 , n39871 , n31459 );
and ( n39873 , n33490 , n31077 );
or ( n39874 , n39872 , n39873 );
and ( n39875 , n39874 , n31373 );
not ( n39876 , n31402 );
and ( n39877 , n39876 , n31459 );
and ( n39878 , n33490 , n31402 );
or ( n39879 , n39877 , n39878 );
and ( n39880 , n39879 , n31408 );
not ( n39881 , n31437 );
and ( n39882 , n39881 , n31459 );
not ( n39883 , n31455 );
and ( n39884 , n39883 , n31505 );
xor ( n39885 , n31459 , n31460 );
and ( n39886 , n39885 , n31455 );
or ( n39887 , n39884 , n39886 );
and ( n39888 , n39887 , n31437 );
or ( n39889 , n39882 , n39888 );
and ( n39890 , n39889 , n31468 );
not ( n39891 , n31497 );
and ( n39892 , n39891 , n31459 );
not ( n39893 , n31454 );
not ( n39894 , n31501 );
and ( n39895 , n39894 , n31505 );
xor ( n39896 , n31506 , n31511 );
and ( n39897 , n39896 , n31501 );
or ( n39898 , n39895 , n39897 );
and ( n39899 , n39893 , n39898 );
and ( n39900 , n39885 , n31454 );
or ( n39901 , n39899 , n39900 );
and ( n39902 , n39901 , n31497 );
or ( n39903 , n39892 , n39902 );
and ( n39904 , n39903 , n31521 );
and ( n39905 , n31459 , n31553 );
or ( n39906 , n39875 , n39880 , n39890 , n39904 , n39905 );
and ( n39907 , n39906 , n31557 );
not ( n39908 , n31452 );
not ( n39909 , n31619 );
and ( n39910 , n39909 , n31624 );
xor ( n39911 , n31625 , n31630 );
and ( n39912 , n39911 , n31619 );
or ( n39913 , n39910 , n39912 );
and ( n39914 , n39908 , n39913 );
and ( n39915 , n31459 , n31452 );
or ( n39916 , n39914 , n39915 );
and ( n39917 , n39916 , n31638 );
and ( n39918 , n31459 , n31650 );
or ( n39919 , C0 , n39870 , n39907 , n39917 , C0 , n39918 );
buf ( n39920 , n39919 );
buf ( n39921 , n39920 );
buf ( n39922 , n30987 );
buf ( n39923 , n30987 );
and ( n39924 , n31507 , n31509 );
and ( n39925 , n31505 , n39924 );
and ( n39926 , n31457 , n39925 );
and ( n39927 , n34062 , n39926 );
and ( n39928 , n34060 , n39927 );
and ( n39929 , n34058 , n39928 );
and ( n39930 , n34056 , n39929 );
and ( n39931 , n34054 , n39930 );
and ( n39932 , n34052 , n39931 );
and ( n39933 , n34050 , n39932 );
and ( n39934 , n34048 , n39933 );
and ( n39935 , n34046 , n39934 );
and ( n39936 , n34044 , n39935 );
and ( n39937 , n34042 , n39936 );
and ( n39938 , n34040 , n39937 );
and ( n39939 , n34038 , n39938 );
and ( n39940 , n33997 , n39939 );
and ( n39941 , n35447 , n39940 );
and ( n39942 , n35445 , n39941 );
and ( n39943 , n35443 , n39942 );
and ( n39944 , n35441 , n39943 );
and ( n39945 , n35439 , n39944 );
and ( n39946 , n35437 , n39945 );
and ( n39947 , n35435 , n39946 );
xor ( n39948 , n35433 , n39947 );
and ( n39949 , n39948 , n31550 );
not ( n39950 , n31041 );
buf ( n39951 , n31041 );
buf ( n39952 , n31041 );
buf ( n39953 , n31041 );
buf ( n39954 , n31041 );
buf ( n39955 , n31041 );
buf ( n39956 , n31041 );
buf ( n39957 , n31041 );
buf ( n39958 , n31041 );
buf ( n39959 , n31041 );
buf ( n39960 , n31041 );
buf ( n39961 , n31041 );
buf ( n39962 , n31041 );
buf ( n39963 , n31041 );
buf ( n39964 , n31041 );
buf ( n39965 , n31041 );
buf ( n39966 , n31041 );
buf ( n39967 , n31041 );
buf ( n39968 , n31041 );
buf ( n39969 , n31041 );
buf ( n39970 , n31041 );
buf ( n39971 , n31041 );
buf ( n39972 , n31041 );
buf ( n39973 , n31041 );
buf ( n39974 , n31041 );
buf ( n39975 , n31041 );
or ( n39976 , n31075 , n33415 );
and ( n39977 , n31044 , n39976 );
or ( n39978 , n31046 , n31048 , n31041 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39977 );
and ( n39979 , n39950 , n39978 );
not ( n39980 , n39979 );
and ( n39981 , n39980 , n35433 );
not ( n39982 , n31026 );
buf ( n39983 , n39982 );
not ( n39984 , n39983 );
not ( n39985 , n39984 );
not ( n39986 , n31022 );
buf ( n39987 , n39986 );
buf ( n39988 , n39987 );
not ( n39989 , n39988 );
not ( n39990 , n39989 );
not ( n39991 , n31018 );
not ( n39992 , n39991 );
buf ( n39993 , n39992 );
buf ( n39994 , n39993 );
not ( n39995 , n39994 );
not ( n39996 , n39995 );
xor ( n39997 , n31014 , n31018 );
not ( n39998 , n39997 );
buf ( n39999 , n39998 );
buf ( n40000 , n39999 );
not ( n40001 , n40000 );
not ( n40002 , n40001 );
nor ( n40003 , n39985 , n39990 , n39996 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40004 , n31173 , n40003 );
nor ( n40005 , n39984 , n39990 , n39996 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40006 , n31175 , n40005 );
nor ( n40007 , n39985 , n39989 , n39996 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40008 , n31177 , n40007 );
nor ( n40009 , n39984 , n39989 , n39996 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40010 , n31179 , n40009 );
nor ( n40011 , n39985 , n39990 , n39995 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40012 , n31181 , n40011 );
nor ( n40013 , n39984 , n39990 , n39995 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40014 , n31183 , n40013 );
nor ( n40015 , n39985 , n39989 , n39995 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40016 , n31185 , n40015 );
nor ( n40017 , n39984 , n39989 , n39995 , n40002 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40018 , n31187 , n40017 );
nor ( n40019 , n39985 , n39990 , n39996 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40020 , n31189 , n40019 );
nor ( n40021 , n39984 , n39990 , n39996 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40022 , n31191 , n40021 );
nor ( n40023 , n39985 , n39989 , n39996 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40024 , n31193 , n40023 );
nor ( n40025 , n39984 , n39989 , n39996 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40026 , n31195 , n40025 );
nor ( n40027 , n39985 , n39990 , n39995 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40028 , n31197 , n40027 );
nor ( n40029 , n39984 , n39990 , n39995 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40030 , n31199 , n40029 );
nor ( n40031 , n39985 , n39989 , n39995 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40032 , n31201 , n40031 );
nor ( n40033 , n39984 , n39989 , n39995 , n40001 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40034 , n31203 , n40033 );
or ( n40035 , n40004 , n40006 , n40008 , n40010 , n40012 , n40014 , n40016 , n40018 , n40020 , n40022 , n40024 , n40026 , n40028 , n40030 , n40032 , n40034 );
and ( n40036 , n31140 , n40003 );
and ( n40037 , n31142 , n40005 );
and ( n40038 , n31144 , n40007 );
and ( n40039 , n31146 , n40009 );
and ( n40040 , n31148 , n40011 );
and ( n40041 , n31150 , n40013 );
and ( n40042 , n31152 , n40015 );
and ( n40043 , n31154 , n40017 );
and ( n40044 , n31156 , n40019 );
and ( n40045 , n31158 , n40021 );
and ( n40046 , n31160 , n40023 );
and ( n40047 , n31162 , n40025 );
and ( n40048 , n31164 , n40027 );
and ( n40049 , n31166 , n40029 );
and ( n40050 , n31168 , n40031 );
and ( n40051 , n31170 , n40033 );
or ( n40052 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 );
and ( n40053 , n31086 , n40003 );
and ( n40054 , n31090 , n40005 );
and ( n40055 , n31094 , n40007 );
and ( n40056 , n31098 , n40009 );
and ( n40057 , n31101 , n40011 );
and ( n40058 , n31105 , n40013 );
and ( n40059 , n31108 , n40015 );
and ( n40060 , n31111 , n40017 );
and ( n40061 , n31114 , n40019 );
and ( n40062 , n31117 , n40021 );
and ( n40063 , n31120 , n40023 );
and ( n40064 , n31123 , n40025 );
and ( n40065 , n31126 , n40027 );
and ( n40066 , n31129 , n40029 );
and ( n40067 , n31132 , n40031 );
and ( n40068 , n31135 , n40033 );
or ( n40069 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 );
not ( n40070 , n31026 );
not ( n40071 , n40070 );
buf ( n40072 , n40071 );
not ( n40073 , n40072 );
not ( n40074 , n40073 );
xnor ( n40075 , n31022 , n31026 );
not ( n40076 , n40075 );
buf ( n40077 , n40076 );
buf ( n40078 , n40077 );
not ( n40079 , n40078 );
not ( n40080 , n40079 );
or ( n40081 , n31022 , n31026 );
xor ( n40082 , n31018 , n40081 );
not ( n40083 , n40082 );
buf ( n40084 , n40083 );
buf ( n40085 , n40084 );
not ( n40086 , n40085 );
not ( n40087 , n40086 );
and ( n40088 , n31018 , n40081 );
xor ( n40089 , n31014 , n40088 );
not ( n40090 , n40089 );
buf ( n40091 , n40090 );
buf ( n40092 , n40091 );
not ( n40093 , n40092 );
not ( n40094 , n40093 );
nor ( n40095 , n40074 , n40080 , n40087 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40096 , n31340 , n40095 );
nor ( n40097 , n40073 , n40080 , n40087 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40098 , n31342 , n40097 );
nor ( n40099 , n40074 , n40079 , n40087 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40100 , n31344 , n40099 );
nor ( n40101 , n40073 , n40079 , n40087 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40102 , n31346 , n40101 );
nor ( n40103 , n40074 , n40080 , n40086 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40104 , n31348 , n40103 );
nor ( n40105 , n40073 , n40080 , n40086 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40106 , n31350 , n40105 );
nor ( n40107 , n40074 , n40079 , n40086 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40108 , n31352 , n40107 );
nor ( n40109 , n40073 , n40079 , n40086 , n40094 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40110 , n31354 , n40109 );
nor ( n40111 , n40074 , n40080 , n40087 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40112 , n31356 , n40111 );
nor ( n40113 , n40073 , n40080 , n40087 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40114 , n31358 , n40113 );
nor ( n40115 , n40074 , n40079 , n40087 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40116 , n31360 , n40115 );
nor ( n40117 , n40073 , n40079 , n40087 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40118 , n31362 , n40117 );
nor ( n40119 , n40074 , n40080 , n40086 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40120 , n31364 , n40119 );
nor ( n40121 , n40073 , n40080 , n40086 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40122 , n31366 , n40121 );
nor ( n40123 , n40074 , n40079 , n40086 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40124 , n31368 , n40123 );
nor ( n40125 , n40073 , n40079 , n40086 , n40093 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n40126 , n31370 , n40125 );
or ( n40127 , n40096 , n40098 , n40100 , n40102 , n40104 , n40106 , n40108 , n40110 , n40112 , n40114 , n40116 , n40118 , n40120 , n40122 , n40124 , n40126 );
and ( n40128 , n40069 , n40127 );
and ( n40129 , n40052 , n40128 );
xor ( n40130 , n40035 , n40129 );
and ( n40131 , n40130 , n39979 );
or ( n40132 , n39981 , n40131 );
and ( n40133 , n40132 , n31538 );
or ( n40134 , n31537 , n31521 );
or ( n40135 , n40134 , n31468 );
or ( n40136 , n40135 , n31408 );
or ( n40137 , n40136 , n31373 );
or ( n40138 , n40137 , n31540 );
or ( n40139 , n40138 , n31542 );
or ( n40140 , n40139 , n31544 );
or ( n40141 , n40140 , n31546 );
or ( n40142 , n40141 , n31548 );
or ( n40143 , n40142 , n31552 );
and ( n40144 , n35433 , n40143 );
or ( n40145 , n39949 , n40133 , n40144 );
and ( n40146 , n40145 , n31557 );
or ( n40147 , n31640 , n33973 );
or ( n40148 , n40147 , n31638 );
or ( n40149 , n40148 , n31641 );
or ( n40150 , n40149 , n31643 );
or ( n40151 , n40150 , n31645 );
or ( n40152 , n40151 , n31647 );
or ( n40153 , n40152 , n31649 );
or ( n40154 , n40153 , n31007 );
and ( n40155 , n35433 , n40154 );
or ( n40156 , C0 , n40146 , n40155 );
buf ( n40157 , n40156 );
buf ( n40158 , n40157 );
buf ( n40159 , RI15b5e5f0_1085);
buf ( n40160 , n40159 );
buf ( n40161 , n31655 );
buf ( n40162 , n30987 );
not ( n40163 , n31658 );
not ( n40164 , n40163 );
and ( n40165 , n40164 , n31820 );
nor ( n40166 , n31673 , n31669 , n31665 , n31661 , n31657 );
not ( n40167 , n40166 );
and ( n40168 , n40167 , n31820 );
and ( n40169 , n32252 , n40166 );
or ( n40170 , n40168 , n40169 );
and ( n40171 , n40170 , n40163 );
or ( n40172 , n40165 , n40171 );
and ( n40173 , n40172 , n32498 );
not ( n40174 , n31673 );
not ( n40175 , n40174 );
buf ( n40176 , n40175 );
not ( n40177 , n40176 );
xor ( n40178 , n31669 , n31673 );
not ( n40179 , n40178 );
buf ( n40180 , n40179 );
buf ( n40181 , n40180 );
not ( n40182 , n40181 );
and ( n40183 , n31669 , n31673 );
xor ( n40184 , n31665 , n40183 );
not ( n40185 , n40184 );
buf ( n40186 , n40185 );
buf ( n40187 , n40186 );
not ( n40188 , n40187 );
and ( n40189 , n31665 , n40183 );
xor ( n40190 , n31661 , n40189 );
not ( n40191 , n40190 );
buf ( n40192 , n40191 );
buf ( n40193 , n40192 );
not ( n40194 , n40193 );
nor ( n40195 , n40177 , n40182 , n40188 , n40194 , C0 );
not ( n40196 , n40195 );
not ( n40197 , n40166 );
and ( n40198 , n40197 , n31820 );
buf ( n40199 , RI15b5e6e0_1087);
buf ( n40200 , RI15b5d9c0_1059);
buf ( n40201 , RI15b5da38_1060);
buf ( n40202 , RI15b5dab0_1061);
buf ( n40203 , RI15b5db28_1062);
buf ( n40204 , RI15b5dba0_1063);
buf ( n40205 , RI15b5dc18_1064);
buf ( n40206 , RI15b5dc90_1065);
buf ( n40207 , RI15b5dd08_1066);
buf ( n40208 , RI15b5dd80_1067);
buf ( n40209 , RI15b5ddf8_1068);
buf ( n40210 , RI15b5de70_1069);
buf ( n40211 , RI15b5dee8_1070);
buf ( n40212 , RI15b5df60_1071);
buf ( n40213 , RI15b5dfd8_1072);
buf ( n40214 , RI15b5e050_1073);
buf ( n40215 , RI15b5e0c8_1074);
buf ( n40216 , RI15b5e140_1075);
buf ( n40217 , RI15b5e1b8_1076);
buf ( n40218 , RI15b5e230_1077);
buf ( n40219 , RI15b5e2a8_1078);
buf ( n40220 , RI15b5e320_1079);
buf ( n40221 , RI15b5e398_1080);
buf ( n40222 , RI15b5e410_1081);
buf ( n40223 , RI15b5e488_1082);
buf ( n40224 , RI15b5e500_1083);
buf ( n40225 , RI15b5e578_1084);
buf ( n40226 , RI15b5e668_1086);
or ( n40227 , n39348 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40159 , n40226 );
and ( n40228 , n40199 , n40227 );
not ( n40229 , n40228 );
buf ( n40230 , RI15b3f948_34);
and ( n40231 , n40229 , n40230 );
buf ( n40232 , RI15b64950_1297);
and ( n40233 , n40232 , n40228 );
or ( n40234 , n40231 , n40233 );
buf ( n40235 , n40234 );
not ( n40236 , n40235 );
buf ( n40237 , n40236 );
not ( n40238 , n40237 );
not ( n40239 , n40228 );
buf ( n40240 , RI15b3eac0_3);
and ( n40241 , n40239 , n40240 );
buf ( n40242 , RI15b657d8_1328);
and ( n40243 , n40242 , n40228 );
or ( n40244 , n40241 , n40243 );
not ( n40245 , n40244 );
not ( n40246 , n40228 );
buf ( n40247 , RI15b3f8d0_33);
and ( n40248 , n40246 , n40247 );
buf ( n40249 , RI15b649c8_1298);
and ( n40250 , n40249 , n40228 );
or ( n40251 , n40248 , n40250 );
and ( n40252 , n40245 , n40251 );
not ( n40253 , n40251 );
not ( n40254 , n40234 );
xor ( n40255 , n40253 , n40254 );
and ( n40256 , n40255 , n40244 );
or ( n40257 , n40252 , n40256 );
not ( n40258 , n40257 );
buf ( n40259 , n40258 );
buf ( n40260 , n40259 );
not ( n40261 , n40260 );
or ( n40262 , n40238 , n40261 );
not ( n40263 , n40244 );
not ( n40264 , n40228 );
buf ( n40265 , RI15b3f858_32);
and ( n40266 , n40264 , n40265 );
buf ( n40267 , RI15b64a40_1299);
and ( n40268 , n40267 , n40228 );
or ( n40269 , n40266 , n40268 );
and ( n40270 , n40263 , n40269 );
not ( n40271 , n40269 );
and ( n40272 , n40253 , n40254 );
xor ( n40273 , n40271 , n40272 );
and ( n40274 , n40273 , n40244 );
or ( n40275 , n40270 , n40274 );
not ( n40276 , n40275 );
buf ( n40277 , n40276 );
buf ( n40278 , n40277 );
not ( n40279 , n40278 );
or ( n40280 , n40262 , n40279 );
not ( n40281 , n40244 );
not ( n40282 , n40228 );
buf ( n40283 , RI15b3f7e0_31);
and ( n40284 , n40282 , n40283 );
buf ( n40285 , RI15b64ab8_1300);
and ( n40286 , n40285 , n40228 );
or ( n40287 , n40284 , n40286 );
and ( n40288 , n40281 , n40287 );
not ( n40289 , n40287 );
and ( n40290 , n40271 , n40272 );
xor ( n40291 , n40289 , n40290 );
and ( n40292 , n40291 , n40244 );
or ( n40293 , n40288 , n40292 );
not ( n40294 , n40293 );
buf ( n40295 , n40294 );
buf ( n40296 , n40295 );
not ( n40297 , n40296 );
or ( n40298 , n40280 , n40297 );
not ( n40299 , n40244 );
not ( n40300 , n40228 );
buf ( n40301 , RI15b3f768_30);
and ( n40302 , n40300 , n40301 );
buf ( n40303 , RI15b64b30_1301);
and ( n40304 , n40303 , n40228 );
or ( n40305 , n40302 , n40304 );
and ( n40306 , n40299 , n40305 );
not ( n40307 , n40305 );
and ( n40308 , n40289 , n40290 );
xor ( n40309 , n40307 , n40308 );
and ( n40310 , n40309 , n40244 );
or ( n40311 , n40306 , n40310 );
not ( n40312 , n40311 );
buf ( n40313 , n40312 );
buf ( n40314 , n40313 );
not ( n40315 , n40314 );
or ( n40316 , n40298 , n40315 );
not ( n40317 , n40244 );
not ( n40318 , n40228 );
buf ( n40319 , RI15b3f6f0_29);
and ( n40320 , n40318 , n40319 );
buf ( n40321 , RI15b64ba8_1302);
and ( n40322 , n40321 , n40228 );
or ( n40323 , n40320 , n40322 );
and ( n40324 , n40317 , n40323 );
not ( n40325 , n40323 );
and ( n40326 , n40307 , n40308 );
xor ( n40327 , n40325 , n40326 );
and ( n40328 , n40327 , n40244 );
or ( n40329 , n40324 , n40328 );
not ( n40330 , n40329 );
buf ( n40331 , n40330 );
buf ( n40332 , n40331 );
not ( n40333 , n40332 );
or ( n40334 , n40316 , n40333 );
not ( n40335 , n40244 );
not ( n40336 , n40228 );
buf ( n40337 , RI15b3f678_28);
and ( n40338 , n40336 , n40337 );
buf ( n40339 , RI15b64c20_1303);
and ( n40340 , n40339 , n40228 );
or ( n40341 , n40338 , n40340 );
and ( n40342 , n40335 , n40341 );
not ( n40343 , n40341 );
and ( n40344 , n40325 , n40326 );
xor ( n40345 , n40343 , n40344 );
and ( n40346 , n40345 , n40244 );
or ( n40347 , n40342 , n40346 );
not ( n40348 , n40347 );
buf ( n40349 , n40348 );
buf ( n40350 , n40349 );
not ( n40351 , n40350 );
or ( n40352 , n40334 , n40351 );
not ( n40353 , n40244 );
not ( n40354 , n40228 );
buf ( n40355 , RI15b3f600_27);
and ( n40356 , n40354 , n40355 );
buf ( n40357 , RI15b64c98_1304);
and ( n40358 , n40357 , n40228 );
or ( n40359 , n40356 , n40358 );
and ( n40360 , n40353 , n40359 );
not ( n40361 , n40359 );
and ( n40362 , n40343 , n40344 );
xor ( n40363 , n40361 , n40362 );
and ( n40364 , n40363 , n40244 );
or ( n40365 , n40360 , n40364 );
not ( n40366 , n40365 );
buf ( n40367 , n40366 );
buf ( n40368 , n40367 );
not ( n40369 , n40368 );
or ( n40370 , n40352 , n40369 );
buf ( n40371 , n40370 );
buf ( n40372 , n40371 );
and ( n40373 , n40372 , n40244 );
not ( n40374 , n40373 );
and ( n40375 , n40374 , n40369 );
xor ( n40376 , n40369 , n40244 );
xor ( n40377 , n40351 , n40244 );
xor ( n40378 , n40333 , n40244 );
xor ( n40379 , n40315 , n40244 );
xor ( n40380 , n40297 , n40244 );
xor ( n40381 , n40279 , n40244 );
xor ( n40382 , n40261 , n40244 );
xor ( n40383 , n40238 , n40244 );
and ( n40384 , n40383 , n40244 );
and ( n40385 , n40382 , n40384 );
and ( n40386 , n40381 , n40385 );
and ( n40387 , n40380 , n40386 );
and ( n40388 , n40379 , n40387 );
and ( n40389 , n40378 , n40388 );
and ( n40390 , n40377 , n40389 );
xor ( n40391 , n40376 , n40390 );
and ( n40392 , n40391 , n40373 );
or ( n40393 , n40375 , n40392 );
and ( n40394 , n40393 , n40166 );
or ( n40395 , n40198 , n40394 );
and ( n40396 , n40196 , n40395 );
and ( n40397 , n40393 , n40195 );
or ( n40398 , n40396 , n40397 );
and ( n40399 , n40398 , n32473 );
not ( n40400 , n32475 );
not ( n40401 , n40195 );
not ( n40402 , n40166 );
and ( n40403 , n40402 , n31820 );
and ( n40404 , n40393 , n40166 );
or ( n40405 , n40403 , n40404 );
and ( n40406 , n40401 , n40405 );
and ( n40407 , n40393 , n40195 );
or ( n40408 , n40406 , n40407 );
and ( n40409 , n40400 , n40408 );
not ( n40410 , n40177 );
not ( n40411 , n40410 );
buf ( n40412 , n40411 );
not ( n40413 , n40412 );
not ( n40414 , n40413 );
not ( n40415 , n40414 );
buf ( n40416 , n40415 );
not ( n40417 , n40416 );
xor ( n40418 , n40182 , n40177 );
not ( n40419 , n40418 );
buf ( n40420 , n40419 );
not ( n40421 , n40420 );
xor ( n40422 , n40421 , n40413 );
not ( n40423 , n40422 );
buf ( n40424 , n40423 );
not ( n40425 , n40424 );
and ( n40426 , n40182 , n40177 );
xor ( n40427 , n40188 , n40426 );
not ( n40428 , n40427 );
buf ( n40429 , n40428 );
not ( n40430 , n40429 );
and ( n40431 , n40421 , n40413 );
xor ( n40432 , n40430 , n40431 );
not ( n40433 , n40432 );
buf ( n40434 , n40433 );
not ( n40435 , n40434 );
and ( n40436 , n40188 , n40426 );
xor ( n40437 , n40194 , n40436 );
not ( n40438 , n40437 );
buf ( n40439 , n40438 );
not ( n40440 , n40439 );
and ( n40441 , n40430 , n40431 );
xor ( n40442 , n40440 , n40441 );
not ( n40443 , n40442 );
buf ( n40444 , n40443 );
not ( n40445 , n40444 );
nor ( n40446 , n40417 , n40425 , n40435 , n40445 , C0 );
not ( n40447 , n40446 );
nor ( n40448 , n40413 , n40421 , n40430 , n40440 , C0 );
not ( n40449 , n40448 );
and ( n40450 , n40449 , n40408 );
not ( n40451 , n40244 );
not ( n40452 , n40228 );
buf ( n40453 , RI15b3f1c8_18);
and ( n40454 , n40452 , n40453 );
buf ( n40455 , RI15b650d0_1313);
and ( n40456 , n40455 , n40228 );
or ( n40457 , n40454 , n40456 );
and ( n40458 , n40451 , n40457 );
not ( n40459 , n40457 );
not ( n40460 , n40228 );
buf ( n40461 , RI15b3f240_19);
and ( n40462 , n40460 , n40461 );
buf ( n40463 , RI15b65058_1312);
and ( n40464 , n40463 , n40228 );
or ( n40465 , n40462 , n40464 );
not ( n40466 , n40465 );
not ( n40467 , n40228 );
buf ( n40468 , RI15b3f2b8_20);
and ( n40469 , n40467 , n40468 );
buf ( n40470 , RI15b64fe0_1311);
and ( n40471 , n40470 , n40228 );
or ( n40472 , n40469 , n40471 );
not ( n40473 , n40472 );
not ( n40474 , n40228 );
buf ( n40475 , RI15b3f330_21);
and ( n40476 , n40474 , n40475 );
buf ( n40477 , RI15b64f68_1310);
and ( n40478 , n40477 , n40228 );
or ( n40479 , n40476 , n40478 );
not ( n40480 , n40479 );
not ( n40481 , n40228 );
buf ( n40482 , RI15b3f3a8_22);
and ( n40483 , n40481 , n40482 );
buf ( n40484 , RI15b64ef0_1309);
and ( n40485 , n40484 , n40228 );
or ( n40486 , n40483 , n40485 );
not ( n40487 , n40486 );
not ( n40488 , n40228 );
buf ( n40489 , RI15b3f420_23);
and ( n40490 , n40488 , n40489 );
buf ( n40491 , RI15b64e78_1308);
and ( n40492 , n40491 , n40228 );
or ( n40493 , n40490 , n40492 );
not ( n40494 , n40493 );
not ( n40495 , n40228 );
buf ( n40496 , RI15b3f498_24);
and ( n40497 , n40495 , n40496 );
buf ( n40498 , RI15b64e00_1307);
and ( n40499 , n40498 , n40228 );
or ( n40500 , n40497 , n40499 );
not ( n40501 , n40500 );
not ( n40502 , n40228 );
buf ( n40503 , RI15b3f510_25);
and ( n40504 , n40502 , n40503 );
buf ( n40505 , RI15b64d88_1306);
and ( n40506 , n40505 , n40228 );
or ( n40507 , n40504 , n40506 );
not ( n40508 , n40507 );
not ( n40509 , n40228 );
buf ( n40510 , RI15b3f588_26);
and ( n40511 , n40509 , n40510 );
buf ( n40512 , RI15b64d10_1305);
and ( n40513 , n40512 , n40228 );
or ( n40514 , n40511 , n40513 );
not ( n40515 , n40514 );
not ( n40516 , n40359 );
not ( n40517 , n40341 );
not ( n40518 , n40323 );
not ( n40519 , n40305 );
not ( n40520 , n40287 );
not ( n40521 , n40269 );
not ( n40522 , n40251 );
not ( n40523 , n40234 );
and ( n40524 , n40522 , n40523 );
and ( n40525 , n40521 , n40524 );
and ( n40526 , n40520 , n40525 );
and ( n40527 , n40519 , n40526 );
and ( n40528 , n40518 , n40527 );
and ( n40529 , n40517 , n40528 );
and ( n40530 , n40516 , n40529 );
and ( n40531 , n40515 , n40530 );
and ( n40532 , n40508 , n40531 );
and ( n40533 , n40501 , n40532 );
and ( n40534 , n40494 , n40533 );
and ( n40535 , n40487 , n40534 );
and ( n40536 , n40480 , n40535 );
and ( n40537 , n40473 , n40536 );
and ( n40538 , n40466 , n40537 );
xor ( n40539 , n40459 , n40538 );
and ( n40540 , n40539 , n40244 );
or ( n40541 , n40458 , n40540 );
not ( n40542 , n40541 );
buf ( n40543 , n40542 );
buf ( n40544 , n40543 );
not ( n40545 , n40544 );
buf ( n40546 , n40545 );
buf ( n40547 , n40546 );
not ( n40548 , n40547 );
buf ( n40549 , n40548 );
not ( n40550 , n40549 );
not ( n40551 , n40244 );
not ( n40552 , n40228 );
buf ( n40553 , RI15b3eb38_4);
and ( n40554 , n40552 , n40553 );
buf ( n40555 , RI15b65760_1327);
and ( n40556 , n40555 , n40228 );
or ( n40557 , n40554 , n40556 );
not ( n40558 , n40557 );
not ( n40559 , n40228 );
buf ( n40560 , RI15b3ebb0_5);
and ( n40561 , n40559 , n40560 );
buf ( n40562 , RI15b656e8_1326);
and ( n40563 , n40562 , n40228 );
or ( n40564 , n40561 , n40563 );
not ( n40565 , n40564 );
not ( n40566 , n40228 );
buf ( n40567 , RI15b3ec28_6);
and ( n40568 , n40566 , n40567 );
buf ( n40569 , RI15b65670_1325);
and ( n40570 , n40569 , n40228 );
or ( n40571 , n40568 , n40570 );
not ( n40572 , n40571 );
not ( n40573 , n40228 );
buf ( n40574 , RI15b3eca0_7);
and ( n40575 , n40573 , n40574 );
buf ( n40576 , RI15b655f8_1324);
and ( n40577 , n40576 , n40228 );
or ( n40578 , n40575 , n40577 );
not ( n40579 , n40578 );
not ( n40580 , n40228 );
buf ( n40581 , RI15b3ed18_8);
and ( n40582 , n40580 , n40581 );
buf ( n40583 , RI15b65580_1323);
and ( n40584 , n40583 , n40228 );
or ( n40585 , n40582 , n40584 );
not ( n40586 , n40585 );
not ( n40587 , n40228 );
buf ( n40588 , RI15b3ed90_9);
and ( n40589 , n40587 , n40588 );
buf ( n40590 , RI15b65508_1322);
and ( n40591 , n40590 , n40228 );
or ( n40592 , n40589 , n40591 );
not ( n40593 , n40592 );
not ( n40594 , n40228 );
buf ( n40595 , RI15b3ee08_10);
and ( n40596 , n40594 , n40595 );
buf ( n40597 , RI15b65490_1321);
and ( n40598 , n40597 , n40228 );
or ( n40599 , n40596 , n40598 );
not ( n40600 , n40599 );
not ( n40601 , n40228 );
buf ( n40602 , RI15b3ee80_11);
and ( n40603 , n40601 , n40602 );
buf ( n40604 , RI15b65418_1320);
and ( n40605 , n40604 , n40228 );
or ( n40606 , n40603 , n40605 );
not ( n40607 , n40606 );
not ( n40608 , n40228 );
buf ( n40609 , RI15b3eef8_12);
and ( n40610 , n40608 , n40609 );
buf ( n40611 , RI15b653a0_1319);
and ( n40612 , n40611 , n40228 );
or ( n40613 , n40610 , n40612 );
not ( n40614 , n40613 );
not ( n40615 , n40228 );
buf ( n40616 , RI15b3ef70_13);
and ( n40617 , n40615 , n40616 );
buf ( n40618 , RI15b65328_1318);
and ( n40619 , n40618 , n40228 );
or ( n40620 , n40617 , n40619 );
not ( n40621 , n40620 );
not ( n40622 , n40228 );
buf ( n40623 , RI15b3efe8_14);
and ( n40624 , n40622 , n40623 );
buf ( n40625 , RI15b652b0_1317);
and ( n40626 , n40625 , n40228 );
or ( n40627 , n40624 , n40626 );
not ( n40628 , n40627 );
not ( n40629 , n40228 );
buf ( n40630 , RI15b3f060_15);
and ( n40631 , n40629 , n40630 );
buf ( n40632 , RI15b65238_1316);
and ( n40633 , n40632 , n40228 );
or ( n40634 , n40631 , n40633 );
not ( n40635 , n40634 );
not ( n40636 , n40228 );
buf ( n40637 , RI15b3f0d8_16);
and ( n40638 , n40636 , n40637 );
buf ( n40639 , RI15b651c0_1315);
and ( n40640 , n40639 , n40228 );
or ( n40641 , n40638 , n40640 );
not ( n40642 , n40641 );
not ( n40643 , n40228 );
buf ( n40644 , RI15b3f150_17);
and ( n40645 , n40643 , n40644 );
buf ( n40646 , RI15b65148_1314);
and ( n40647 , n40646 , n40228 );
or ( n40648 , n40645 , n40647 );
not ( n40649 , n40648 );
and ( n40650 , n40459 , n40538 );
and ( n40651 , n40649 , n40650 );
and ( n40652 , n40642 , n40651 );
and ( n40653 , n40635 , n40652 );
and ( n40654 , n40628 , n40653 );
and ( n40655 , n40621 , n40654 );
and ( n40656 , n40614 , n40655 );
and ( n40657 , n40607 , n40656 );
and ( n40658 , n40600 , n40657 );
and ( n40659 , n40593 , n40658 );
and ( n40660 , n40586 , n40659 );
and ( n40661 , n40579 , n40660 );
and ( n40662 , n40572 , n40661 );
and ( n40663 , n40565 , n40662 );
and ( n40664 , n40558 , n40663 );
xor ( n40665 , n40551 , n40664 );
buf ( n40666 , n40244 );
and ( n40667 , n40665 , n40666 );
buf ( n40668 , n40667 );
not ( n40669 , n40668 );
not ( n40670 , n40669 );
not ( n40671 , n40670 );
not ( n40672 , n40244 );
and ( n40673 , n40672 , n40557 );
xor ( n40674 , n40558 , n40663 );
and ( n40675 , n40674 , n40244 );
or ( n40676 , n40673 , n40675 );
not ( n40677 , n40676 );
buf ( n40678 , n40677 );
buf ( n40679 , n40678 );
not ( n40680 , n40679 );
not ( n40681 , n40680 );
not ( n40682 , n40244 );
and ( n40683 , n40682 , n40564 );
xor ( n40684 , n40565 , n40662 );
and ( n40685 , n40684 , n40244 );
or ( n40686 , n40683 , n40685 );
not ( n40687 , n40686 );
buf ( n40688 , n40687 );
buf ( n40689 , n40688 );
not ( n40690 , n40689 );
not ( n40691 , n40690 );
not ( n40692 , n40244 );
and ( n40693 , n40692 , n40571 );
xor ( n40694 , n40572 , n40661 );
and ( n40695 , n40694 , n40244 );
or ( n40696 , n40693 , n40695 );
not ( n40697 , n40696 );
buf ( n40698 , n40697 );
buf ( n40699 , n40698 );
not ( n40700 , n40699 );
not ( n40701 , n40700 );
not ( n40702 , n40244 );
and ( n40703 , n40702 , n40578 );
xor ( n40704 , n40579 , n40660 );
and ( n40705 , n40704 , n40244 );
or ( n40706 , n40703 , n40705 );
not ( n40707 , n40706 );
buf ( n40708 , n40707 );
buf ( n40709 , n40708 );
not ( n40710 , n40709 );
not ( n40711 , n40710 );
not ( n40712 , n40244 );
and ( n40713 , n40712 , n40585 );
xor ( n40714 , n40586 , n40659 );
and ( n40715 , n40714 , n40244 );
or ( n40716 , n40713 , n40715 );
not ( n40717 , n40716 );
buf ( n40718 , n40717 );
buf ( n40719 , n40718 );
not ( n40720 , n40719 );
not ( n40721 , n40720 );
not ( n40722 , n40244 );
and ( n40723 , n40722 , n40592 );
xor ( n40724 , n40593 , n40658 );
and ( n40725 , n40724 , n40244 );
or ( n40726 , n40723 , n40725 );
not ( n40727 , n40726 );
buf ( n40728 , n40727 );
buf ( n40729 , n40728 );
not ( n40730 , n40729 );
not ( n40731 , n40730 );
not ( n40732 , n40244 );
and ( n40733 , n40732 , n40599 );
xor ( n40734 , n40600 , n40657 );
and ( n40735 , n40734 , n40244 );
or ( n40736 , n40733 , n40735 );
not ( n40737 , n40736 );
buf ( n40738 , n40737 );
buf ( n40739 , n40738 );
not ( n40740 , n40739 );
not ( n40741 , n40740 );
not ( n40742 , n40244 );
and ( n40743 , n40742 , n40606 );
xor ( n40744 , n40607 , n40656 );
and ( n40745 , n40744 , n40244 );
or ( n40746 , n40743 , n40745 );
not ( n40747 , n40746 );
buf ( n40748 , n40747 );
buf ( n40749 , n40748 );
not ( n40750 , n40749 );
not ( n40751 , n40750 );
not ( n40752 , n40244 );
and ( n40753 , n40752 , n40613 );
xor ( n40754 , n40614 , n40655 );
and ( n40755 , n40754 , n40244 );
or ( n40756 , n40753 , n40755 );
not ( n40757 , n40756 );
buf ( n40758 , n40757 );
buf ( n40759 , n40758 );
not ( n40760 , n40759 );
not ( n40761 , n40760 );
not ( n40762 , n40244 );
and ( n40763 , n40762 , n40620 );
xor ( n40764 , n40621 , n40654 );
and ( n40765 , n40764 , n40244 );
or ( n40766 , n40763 , n40765 );
not ( n40767 , n40766 );
buf ( n40768 , n40767 );
buf ( n40769 , n40768 );
not ( n40770 , n40769 );
not ( n40771 , n40770 );
not ( n40772 , n40244 );
and ( n40773 , n40772 , n40627 );
xor ( n40774 , n40628 , n40653 );
and ( n40775 , n40774 , n40244 );
or ( n40776 , n40773 , n40775 );
not ( n40777 , n40776 );
buf ( n40778 , n40777 );
buf ( n40779 , n40778 );
not ( n40780 , n40779 );
not ( n40781 , n40780 );
not ( n40782 , n40244 );
and ( n40783 , n40782 , n40634 );
xor ( n40784 , n40635 , n40652 );
and ( n40785 , n40784 , n40244 );
or ( n40786 , n40783 , n40785 );
not ( n40787 , n40786 );
buf ( n40788 , n40787 );
buf ( n40789 , n40788 );
not ( n40790 , n40789 );
not ( n40791 , n40790 );
not ( n40792 , n40244 );
and ( n40793 , n40792 , n40641 );
xor ( n40794 , n40642 , n40651 );
and ( n40795 , n40794 , n40244 );
or ( n40796 , n40793 , n40795 );
not ( n40797 , n40796 );
buf ( n40798 , n40797 );
buf ( n40799 , n40798 );
not ( n40800 , n40799 );
not ( n40801 , n40800 );
not ( n40802 , n40244 );
and ( n40803 , n40802 , n40648 );
xor ( n40804 , n40649 , n40650 );
and ( n40805 , n40804 , n40244 );
or ( n40806 , n40803 , n40805 );
not ( n40807 , n40806 );
buf ( n40808 , n40807 );
buf ( n40809 , n40808 );
not ( n40810 , n40809 );
not ( n40811 , n40810 );
not ( n40812 , n40545 );
and ( n40813 , n40811 , n40812 );
and ( n40814 , n40801 , n40813 );
and ( n40815 , n40791 , n40814 );
and ( n40816 , n40781 , n40815 );
and ( n40817 , n40771 , n40816 );
and ( n40818 , n40761 , n40817 );
and ( n40819 , n40751 , n40818 );
and ( n40820 , n40741 , n40819 );
and ( n40821 , n40731 , n40820 );
and ( n40822 , n40721 , n40821 );
and ( n40823 , n40711 , n40822 );
and ( n40824 , n40701 , n40823 );
and ( n40825 , n40691 , n40824 );
and ( n40826 , n40681 , n40825 );
and ( n40827 , n40671 , n40826 );
not ( n40828 , n40827 );
and ( n40829 , n40828 , n40244 );
buf ( n40830 , n40829 );
not ( n40831 , n40830 );
not ( n40832 , n40244 );
and ( n40833 , n40832 , n40810 );
xor ( n40834 , n40811 , n40812 );
and ( n40835 , n40834 , n40244 );
or ( n40836 , n40833 , n40835 );
and ( n40837 , n40831 , n40836 );
not ( n40838 , n40836 );
not ( n40839 , n40546 );
xor ( n40840 , n40838 , n40839 );
and ( n40841 , n40840 , n40830 );
or ( n40842 , n40837 , n40841 );
not ( n40843 , n40842 );
buf ( n40844 , n40843 );
buf ( n40845 , n40844 );
not ( n40846 , n40845 );
or ( n40847 , n40550 , n40846 );
not ( n40848 , n40830 );
not ( n40849 , n40244 );
and ( n40850 , n40849 , n40800 );
xor ( n40851 , n40801 , n40813 );
and ( n40852 , n40851 , n40244 );
or ( n40853 , n40850 , n40852 );
and ( n40854 , n40848 , n40853 );
not ( n40855 , n40853 );
and ( n40856 , n40838 , n40839 );
xor ( n40857 , n40855 , n40856 );
and ( n40858 , n40857 , n40830 );
or ( n40859 , n40854 , n40858 );
not ( n40860 , n40859 );
buf ( n40861 , n40860 );
buf ( n40862 , n40861 );
not ( n40863 , n40862 );
or ( n40864 , n40847 , n40863 );
not ( n40865 , n40830 );
not ( n40866 , n40244 );
and ( n40867 , n40866 , n40790 );
xor ( n40868 , n40791 , n40814 );
and ( n40869 , n40868 , n40244 );
or ( n40870 , n40867 , n40869 );
and ( n40871 , n40865 , n40870 );
not ( n40872 , n40870 );
and ( n40873 , n40855 , n40856 );
xor ( n40874 , n40872 , n40873 );
and ( n40875 , n40874 , n40830 );
or ( n40876 , n40871 , n40875 );
not ( n40877 , n40876 );
buf ( n40878 , n40877 );
buf ( n40879 , n40878 );
not ( n40880 , n40879 );
or ( n40881 , n40864 , n40880 );
not ( n40882 , n40830 );
not ( n40883 , n40244 );
and ( n40884 , n40883 , n40780 );
xor ( n40885 , n40781 , n40815 );
and ( n40886 , n40885 , n40244 );
or ( n40887 , n40884 , n40886 );
and ( n40888 , n40882 , n40887 );
not ( n40889 , n40887 );
and ( n40890 , n40872 , n40873 );
xor ( n40891 , n40889 , n40890 );
and ( n40892 , n40891 , n40830 );
or ( n40893 , n40888 , n40892 );
not ( n40894 , n40893 );
buf ( n40895 , n40894 );
buf ( n40896 , n40895 );
not ( n40897 , n40896 );
or ( n40898 , n40881 , n40897 );
not ( n40899 , n40830 );
not ( n40900 , n40244 );
and ( n40901 , n40900 , n40770 );
xor ( n40902 , n40771 , n40816 );
and ( n40903 , n40902 , n40244 );
or ( n40904 , n40901 , n40903 );
and ( n40905 , n40899 , n40904 );
not ( n40906 , n40904 );
and ( n40907 , n40889 , n40890 );
xor ( n40908 , n40906 , n40907 );
and ( n40909 , n40908 , n40830 );
or ( n40910 , n40905 , n40909 );
not ( n40911 , n40910 );
buf ( n40912 , n40911 );
buf ( n40913 , n40912 );
not ( n40914 , n40913 );
or ( n40915 , n40898 , n40914 );
not ( n40916 , n40830 );
not ( n40917 , n40244 );
and ( n40918 , n40917 , n40760 );
xor ( n40919 , n40761 , n40817 );
and ( n40920 , n40919 , n40244 );
or ( n40921 , n40918 , n40920 );
and ( n40922 , n40916 , n40921 );
not ( n40923 , n40921 );
and ( n40924 , n40906 , n40907 );
xor ( n40925 , n40923 , n40924 );
and ( n40926 , n40925 , n40830 );
or ( n40927 , n40922 , n40926 );
not ( n40928 , n40927 );
buf ( n40929 , n40928 );
buf ( n40930 , n40929 );
not ( n40931 , n40930 );
or ( n40932 , n40915 , n40931 );
not ( n40933 , n40830 );
not ( n40934 , n40244 );
and ( n40935 , n40934 , n40750 );
xor ( n40936 , n40751 , n40818 );
and ( n40937 , n40936 , n40244 );
or ( n40938 , n40935 , n40937 );
and ( n40939 , n40933 , n40938 );
not ( n40940 , n40938 );
and ( n40941 , n40923 , n40924 );
xor ( n40942 , n40940 , n40941 );
and ( n40943 , n40942 , n40830 );
or ( n40944 , n40939 , n40943 );
not ( n40945 , n40944 );
buf ( n40946 , n40945 );
buf ( n40947 , n40946 );
not ( n40948 , n40947 );
or ( n40949 , n40932 , n40948 );
buf ( n40950 , n40949 );
buf ( n40951 , n40950 );
and ( n40952 , n40951 , n40830 );
not ( n40953 , n40952 );
and ( n40954 , n40953 , n40948 );
xor ( n40955 , n40948 , n40830 );
xor ( n40956 , n40931 , n40830 );
xor ( n40957 , n40914 , n40830 );
xor ( n40958 , n40897 , n40830 );
xor ( n40959 , n40880 , n40830 );
xor ( n40960 , n40863 , n40830 );
xor ( n40961 , n40846 , n40830 );
xor ( n40962 , n40550 , n40830 );
and ( n40963 , n40962 , n40830 );
and ( n40964 , n40961 , n40963 );
and ( n40965 , n40960 , n40964 );
and ( n40966 , n40959 , n40965 );
and ( n40967 , n40958 , n40966 );
and ( n40968 , n40957 , n40967 );
and ( n40969 , n40956 , n40968 );
xor ( n40970 , n40955 , n40969 );
and ( n40971 , n40970 , n40952 );
or ( n40972 , n40954 , n40971 );
and ( n40973 , n40972 , n40448 );
or ( n40974 , n40450 , n40973 );
and ( n40975 , n40447 , n40974 );
not ( n40976 , n40244 );
and ( n40977 , n40976 , n40599 );
not ( n40978 , n40599 );
not ( n40979 , n40606 );
not ( n40980 , n40613 );
not ( n40981 , n40620 );
not ( n40982 , n40627 );
not ( n40983 , n40634 );
not ( n40984 , n40641 );
not ( n40985 , n40648 );
not ( n40986 , n40457 );
not ( n40987 , n40465 );
not ( n40988 , n40472 );
not ( n40989 , n40479 );
not ( n40990 , n40486 );
not ( n40991 , n40493 );
not ( n40992 , n40500 );
not ( n40993 , n40507 );
not ( n40994 , n40514 );
not ( n40995 , n40359 );
not ( n40996 , n40341 );
not ( n40997 , n40323 );
not ( n40998 , n40305 );
not ( n40999 , n40287 );
not ( n41000 , n40269 );
not ( n41001 , n40251 );
not ( n41002 , n40234 );
and ( n41003 , n41001 , n41002 );
and ( n41004 , n41000 , n41003 );
and ( n41005 , n40999 , n41004 );
and ( n41006 , n40998 , n41005 );
and ( n41007 , n40997 , n41006 );
and ( n41008 , n40996 , n41007 );
and ( n41009 , n40995 , n41008 );
and ( n41010 , n40994 , n41009 );
and ( n41011 , n40993 , n41010 );
and ( n41012 , n40992 , n41011 );
and ( n41013 , n40991 , n41012 );
and ( n41014 , n40990 , n41013 );
and ( n41015 , n40989 , n41014 );
and ( n41016 , n40988 , n41015 );
and ( n41017 , n40987 , n41016 );
and ( n41018 , n40986 , n41017 );
and ( n41019 , n40985 , n41018 );
and ( n41020 , n40984 , n41019 );
and ( n41021 , n40983 , n41020 );
and ( n41022 , n40982 , n41021 );
and ( n41023 , n40981 , n41022 );
and ( n41024 , n40980 , n41023 );
and ( n41025 , n40979 , n41024 );
xor ( n41026 , n40978 , n41025 );
and ( n41027 , n41026 , n40244 );
or ( n41028 , n40977 , n41027 );
not ( n41029 , n41028 );
buf ( n41030 , n41029 );
buf ( n41031 , n41030 );
not ( n41032 , n41031 );
buf ( n41033 , n41032 );
buf ( n41034 , n41033 );
not ( n41035 , n41034 );
buf ( n41036 , n41035 );
not ( n41037 , n41036 );
not ( n41038 , n40244 );
not ( n41039 , n40557 );
not ( n41040 , n40564 );
not ( n41041 , n40571 );
not ( n41042 , n40578 );
not ( n41043 , n40585 );
not ( n41044 , n40592 );
and ( n41045 , n40978 , n41025 );
and ( n41046 , n41044 , n41045 );
and ( n41047 , n41043 , n41046 );
and ( n41048 , n41042 , n41047 );
and ( n41049 , n41041 , n41048 );
and ( n41050 , n41040 , n41049 );
and ( n41051 , n41039 , n41050 );
xor ( n41052 , n41038 , n41051 );
buf ( n41053 , n40244 );
and ( n41054 , n41052 , n41053 );
buf ( n41055 , n41054 );
not ( n41056 , n41055 );
not ( n41057 , n41056 );
not ( n41058 , n41057 );
not ( n41059 , n40244 );
and ( n41060 , n41059 , n40557 );
xor ( n41061 , n41039 , n41050 );
and ( n41062 , n41061 , n40244 );
or ( n41063 , n41060 , n41062 );
not ( n41064 , n41063 );
buf ( n41065 , n41064 );
buf ( n41066 , n41065 );
not ( n41067 , n41066 );
not ( n41068 , n41067 );
not ( n41069 , n40244 );
and ( n41070 , n41069 , n40564 );
xor ( n41071 , n41040 , n41049 );
and ( n41072 , n41071 , n40244 );
or ( n41073 , n41070 , n41072 );
not ( n41074 , n41073 );
buf ( n41075 , n41074 );
buf ( n41076 , n41075 );
not ( n41077 , n41076 );
not ( n41078 , n41077 );
not ( n41079 , n40244 );
and ( n41080 , n41079 , n40571 );
xor ( n41081 , n41041 , n41048 );
and ( n41082 , n41081 , n40244 );
or ( n41083 , n41080 , n41082 );
not ( n41084 , n41083 );
buf ( n41085 , n41084 );
buf ( n41086 , n41085 );
not ( n41087 , n41086 );
not ( n41088 , n41087 );
not ( n41089 , n40244 );
and ( n41090 , n41089 , n40578 );
xor ( n41091 , n41042 , n41047 );
and ( n41092 , n41091 , n40244 );
or ( n41093 , n41090 , n41092 );
not ( n41094 , n41093 );
buf ( n41095 , n41094 );
buf ( n41096 , n41095 );
not ( n41097 , n41096 );
not ( n41098 , n41097 );
not ( n41099 , n40244 );
and ( n41100 , n41099 , n40585 );
xor ( n41101 , n41043 , n41046 );
and ( n41102 , n41101 , n40244 );
or ( n41103 , n41100 , n41102 );
not ( n41104 , n41103 );
buf ( n41105 , n41104 );
buf ( n41106 , n41105 );
not ( n41107 , n41106 );
not ( n41108 , n41107 );
not ( n41109 , n40244 );
and ( n41110 , n41109 , n40592 );
xor ( n41111 , n41044 , n41045 );
and ( n41112 , n41111 , n40244 );
or ( n41113 , n41110 , n41112 );
not ( n41114 , n41113 );
buf ( n41115 , n41114 );
buf ( n41116 , n41115 );
not ( n41117 , n41116 );
not ( n41118 , n41117 );
not ( n41119 , n41032 );
and ( n41120 , n41118 , n41119 );
and ( n41121 , n41108 , n41120 );
and ( n41122 , n41098 , n41121 );
and ( n41123 , n41088 , n41122 );
and ( n41124 , n41078 , n41123 );
and ( n41125 , n41068 , n41124 );
and ( n41126 , n41058 , n41125 );
not ( n41127 , n41126 );
and ( n41128 , n41127 , n40244 );
buf ( n41129 , n41128 );
not ( n41130 , n41129 );
not ( n41131 , n40244 );
and ( n41132 , n41131 , n41117 );
xor ( n41133 , n41118 , n41119 );
and ( n41134 , n41133 , n40244 );
or ( n41135 , n41132 , n41134 );
and ( n41136 , n41130 , n41135 );
not ( n41137 , n41135 );
not ( n41138 , n41033 );
xor ( n41139 , n41137 , n41138 );
and ( n41140 , n41139 , n41129 );
or ( n41141 , n41136 , n41140 );
not ( n41142 , n41141 );
buf ( n41143 , n41142 );
buf ( n41144 , n41143 );
not ( n41145 , n41144 );
or ( n41146 , n41037 , n41145 );
not ( n41147 , n41129 );
not ( n41148 , n40244 );
and ( n41149 , n41148 , n41107 );
xor ( n41150 , n41108 , n41120 );
and ( n41151 , n41150 , n40244 );
or ( n41152 , n41149 , n41151 );
and ( n41153 , n41147 , n41152 );
not ( n41154 , n41152 );
and ( n41155 , n41137 , n41138 );
xor ( n41156 , n41154 , n41155 );
and ( n41157 , n41156 , n41129 );
or ( n41158 , n41153 , n41157 );
not ( n41159 , n41158 );
buf ( n41160 , n41159 );
buf ( n41161 , n41160 );
not ( n41162 , n41161 );
or ( n41163 , n41146 , n41162 );
not ( n41164 , n41129 );
not ( n41165 , n40244 );
and ( n41166 , n41165 , n41097 );
xor ( n41167 , n41098 , n41121 );
and ( n41168 , n41167 , n40244 );
or ( n41169 , n41166 , n41168 );
and ( n41170 , n41164 , n41169 );
not ( n41171 , n41169 );
and ( n41172 , n41154 , n41155 );
xor ( n41173 , n41171 , n41172 );
and ( n41174 , n41173 , n41129 );
or ( n41175 , n41170 , n41174 );
not ( n41176 , n41175 );
buf ( n41177 , n41176 );
buf ( n41178 , n41177 );
not ( n41179 , n41178 );
or ( n41180 , n41163 , n41179 );
not ( n41181 , n41129 );
not ( n41182 , n40244 );
and ( n41183 , n41182 , n41087 );
xor ( n41184 , n41088 , n41122 );
and ( n41185 , n41184 , n40244 );
or ( n41186 , n41183 , n41185 );
and ( n41187 , n41181 , n41186 );
not ( n41188 , n41186 );
and ( n41189 , n41171 , n41172 );
xor ( n41190 , n41188 , n41189 );
and ( n41191 , n41190 , n41129 );
or ( n41192 , n41187 , n41191 );
not ( n41193 , n41192 );
buf ( n41194 , n41193 );
buf ( n41195 , n41194 );
not ( n41196 , n41195 );
or ( n41197 , n41180 , n41196 );
not ( n41198 , n41129 );
not ( n41199 , n40244 );
and ( n41200 , n41199 , n41077 );
xor ( n41201 , n41078 , n41123 );
and ( n41202 , n41201 , n40244 );
or ( n41203 , n41200 , n41202 );
and ( n41204 , n41198 , n41203 );
not ( n41205 , n41203 );
and ( n41206 , n41188 , n41189 );
xor ( n41207 , n41205 , n41206 );
and ( n41208 , n41207 , n41129 );
or ( n41209 , n41204 , n41208 );
not ( n41210 , n41209 );
buf ( n41211 , n41210 );
buf ( n41212 , n41211 );
not ( n41213 , n41212 );
or ( n41214 , n41197 , n41213 );
not ( n41215 , n41129 );
not ( n41216 , n40244 );
and ( n41217 , n41216 , n41067 );
xor ( n41218 , n41068 , n41124 );
and ( n41219 , n41218 , n40244 );
or ( n41220 , n41217 , n41219 );
and ( n41221 , n41215 , n41220 );
not ( n41222 , n41220 );
and ( n41223 , n41205 , n41206 );
xor ( n41224 , n41222 , n41223 );
and ( n41225 , n41224 , n41129 );
or ( n41226 , n41221 , n41225 );
not ( n41227 , n41226 );
buf ( n41228 , n41227 );
buf ( n41229 , n41228 );
not ( n41230 , n41229 );
or ( n41231 , n41214 , n41230 );
xor ( n41232 , n41058 , n41125 );
and ( n41233 , n41232 , n40244 );
buf ( n41234 , n41233 );
not ( n41235 , n41234 );
and ( n41236 , n41222 , n41223 );
xor ( n41237 , n41235 , n41236 );
and ( n41238 , n41237 , n41129 );
buf ( n41239 , n41238 );
not ( n41240 , n41239 );
buf ( n41241 , n41240 );
buf ( n41242 , n41241 );
not ( n41243 , n41242 );
or ( n41244 , n41231 , n41243 );
buf ( n41245 , n41244 );
buf ( n41246 , n41245 );
and ( n41247 , n41246 , n41129 );
not ( n41248 , n41247 );
and ( n41249 , n41248 , n41243 );
xor ( n41250 , n41243 , n41129 );
xor ( n41251 , n41230 , n41129 );
xor ( n41252 , n41213 , n41129 );
xor ( n41253 , n41196 , n41129 );
xor ( n41254 , n41179 , n41129 );
xor ( n41255 , n41162 , n41129 );
xor ( n41256 , n41145 , n41129 );
xor ( n41257 , n41037 , n41129 );
and ( n41258 , n41257 , n41129 );
and ( n41259 , n41256 , n41258 );
and ( n41260 , n41255 , n41259 );
and ( n41261 , n41254 , n41260 );
and ( n41262 , n41253 , n41261 );
and ( n41263 , n41252 , n41262 );
and ( n41264 , n41251 , n41263 );
xor ( n41265 , n41250 , n41264 );
and ( n41266 , n41265 , n41247 );
or ( n41267 , n41249 , n41266 );
and ( n41268 , n41267 , n40446 );
or ( n41269 , n40975 , n41268 );
and ( n41270 , n41269 , n32475 );
or ( n41271 , n40409 , n41270 );
and ( n41272 , n41271 , n32486 );
or ( n41273 , n32491 , n32489 );
or ( n41274 , n41273 , n32492 );
or ( n41275 , n41274 , n32456 );
or ( n41276 , n41275 , n32494 );
or ( n41277 , n41276 , n32496 );
or ( n41278 , n41277 , n32500 );
and ( n41279 , n31820 , n41278 );
or ( n41280 , C0 , n40173 , n40399 , n41272 , n41279 );
buf ( n41281 , n41280 );
buf ( n41282 , n41281 );
not ( n41283 , n31728 );
buf ( n41284 , RI15b62f88_1242);
and ( n41285 , n41283 , n41284 );
buf ( n41286 , RI15b5c7f0_1021);
and ( n41287 , n31732 , n31747 );
xor ( n41288 , n41286 , n41287 );
and ( n41289 , n31748 , n32090 );
xor ( n41290 , n41288 , n41289 );
and ( n41291 , n41290 , n31728 );
or ( n41292 , n41285 , n41291 );
and ( n41293 , n41292 , n32253 );
not ( n41294 , n32283 );
and ( n41295 , n41294 , n41284 );
not ( n41296 , n31823 );
and ( n41297 , n31732 , n32292 );
xor ( n41298 , n41286 , n41297 );
and ( n41299 , n32293 , n32329 );
xor ( n41300 , n41298 , n41299 );
and ( n41301 , n41296 , n41300 );
and ( n41302 , n31732 , n32338 );
xor ( n41303 , n41286 , n41302 );
or ( n41304 , n32339 , n32392 );
xnor ( n41305 , n41303 , n41304 );
and ( n41306 , n41305 , n31823 );
or ( n41307 , n41301 , n41306 );
and ( n41308 , n41307 , n32283 );
or ( n41309 , n41295 , n41308 );
and ( n41310 , n41309 , n32398 );
and ( n41311 , n41284 , n32436 );
or ( n41312 , n41293 , n41310 , n41311 );
and ( n41313 , n41312 , n32456 );
and ( n41314 , n31730 , n32470 );
xor ( n41315 , n41284 , n41314 );
and ( n41316 , n41315 , n32473 );
not ( n41317 , n32475 );
and ( n41318 , n41317 , n41315 );
and ( n41319 , n31730 , n32482 );
xor ( n41320 , n41284 , n41319 );
and ( n41321 , n41320 , n32475 );
or ( n41322 , n41318 , n41321 );
and ( n41323 , n41322 , n32486 );
and ( n41324 , n37573 , n32489 );
and ( n41325 , n41284 , n32501 );
or ( n41326 , C0 , n41313 , n41316 , n41323 , n41324 , n41325 );
buf ( n41327 , n41326 );
buf ( n41328 , n41327 );
buf ( n41329 , n31655 );
buf ( n41330 , n30987 );
and ( n41331 , n33212 , n32528 );
not ( n41332 , n32598 );
and ( n41333 , n41332 , n32975 );
buf ( n41334 , n41333 );
and ( n41335 , n41334 , n32890 );
not ( n41336 , n32919 );
and ( n41337 , n41336 , n32975 );
buf ( n41338 , n41337 );
and ( n41339 , n41338 , n32924 );
not ( n41340 , n32953 );
and ( n41341 , n41340 , n32975 );
not ( n41342 , n32971 );
and ( n41343 , n41342 , n33075 );
xor ( n41344 , n32975 , n33030 );
and ( n41345 , n41344 , n32971 );
or ( n41346 , n41343 , n41345 );
and ( n41347 , n41346 , n32953 );
or ( n41348 , n41341 , n41347 );
and ( n41349 , n41348 , n33038 );
not ( n41350 , n33067 );
and ( n41351 , n41350 , n32975 );
not ( n41352 , n32970 );
not ( n41353 , n33071 );
and ( n41354 , n41353 , n33075 );
xor ( n41355 , n33076 , n33162 );
and ( n41356 , n41355 , n33071 );
or ( n41357 , n41354 , n41356 );
and ( n41358 , n41352 , n41357 );
and ( n41359 , n41344 , n32970 );
or ( n41360 , n41358 , n41359 );
and ( n41361 , n41360 , n33067 );
or ( n41362 , n41351 , n41361 );
and ( n41363 , n41362 , n33172 );
and ( n41364 , n32975 , n33204 );
or ( n41365 , n41335 , n41339 , n41349 , n41363 , n41364 );
and ( n41366 , n41365 , n33208 );
not ( n41367 , n32968 );
not ( n41368 , n33270 );
and ( n41369 , n41368 , n33275 );
xor ( n41370 , n33276 , n33362 );
and ( n41371 , n41370 , n33270 );
or ( n41372 , n41369 , n41371 );
and ( n41373 , n41367 , n41372 );
and ( n41374 , n32975 , n32968 );
or ( n41375 , n41373 , n41374 );
and ( n41376 , n41375 , n33370 );
and ( n41377 , n32975 , n33382 );
or ( n41378 , C0 , n41331 , n41366 , n41376 , C0 , n41377 );
buf ( n41379 , n41378 );
buf ( n41380 , n41379 );
buf ( n41381 , n30987 );
buf ( n41382 , n31655 );
buf ( n41383 , n31655 );
buf ( n41384 , RI15b479b8_308);
buf ( n41385 , n41384 );
buf ( n41386 , n31655 );
not ( n41387 , n34150 );
and ( n41388 , n41387 , n32771 );
not ( n41389 , n32546 );
not ( n41390 , n32538 );
not ( n41391 , n32530 );
and ( n41392 , n41389 , n34153 , n41390 , n32534 , n41391 );
not ( n41393 , n41392 );
and ( n41394 , n41393 , n32771 );
and ( n41395 , n32789 , n41392 );
or ( n41396 , n41394 , n41395 );
and ( n41397 , n41396 , n34150 );
or ( n41398 , n41388 , n41397 );
and ( n41399 , n41398 , n33381 );
not ( n41400 , n34165 );
not ( n41401 , n34177 );
and ( n41402 , n41400 , n34171 , n41401 , n34183 );
not ( n41403 , n41402 );
not ( n41404 , n41392 );
and ( n41405 , n41404 , n32771 );
and ( n41406 , n34301 , n41392 );
or ( n41407 , n41405 , n41406 );
and ( n41408 , n41403 , n41407 );
and ( n41409 , n34301 , n41402 );
or ( n41410 , n41408 , n41409 );
and ( n41411 , n41410 , n33375 );
not ( n41412 , n32968 );
not ( n41413 , n41402 );
not ( n41414 , n41392 );
and ( n41415 , n41414 , n32771 );
and ( n41416 , n34301 , n41392 );
or ( n41417 , n41415 , n41416 );
and ( n41418 , n41413 , n41417 );
and ( n41419 , n34301 , n41402 );
or ( n41420 , n41418 , n41419 );
and ( n41421 , n41412 , n41420 );
not ( n41422 , n34325 );
not ( n41423 , n34344 );
and ( n41424 , n41422 , n34334 , n41423 , n34354 );
not ( n41425 , n41424 );
not ( n41426 , n34321 );
not ( n41427 , n34339 );
and ( n41428 , n41426 , n34357 , n41427 , n34349 );
not ( n41429 , n41428 );
and ( n41430 , n41429 , n41420 );
and ( n41431 , n34761 , n41428 );
or ( n41432 , n41430 , n41431 );
and ( n41433 , n41425 , n41432 );
and ( n41434 , n35050 , n41424 );
or ( n41435 , n41433 , n41434 );
and ( n41436 , n41435 , n32968 );
or ( n41437 , n41421 , n41436 );
and ( n41438 , n41437 , n33370 );
and ( n41439 , n32771 , n35062 );
or ( n41440 , C0 , n41399 , n41411 , n41438 , n41439 );
buf ( n41441 , n41440 );
buf ( n41442 , n41441 );
buf ( n41443 , n30987 );
buf ( n41444 , n30987 );
buf ( n41445 , n31655 );
not ( n41446 , n34150 );
and ( n41447 , n41446 , n32805 );
not ( n41448 , n41392 );
and ( n41449 , n41448 , n32805 );
and ( n41450 , n32823 , n41392 );
or ( n41451 , n41449 , n41450 );
and ( n41452 , n41451 , n34150 );
or ( n41453 , n41447 , n41452 );
and ( n41454 , n41453 , n33381 );
not ( n41455 , n41402 );
not ( n41456 , n41392 );
and ( n41457 , n41456 , n32805 );
not ( n41458 , n34287 );
and ( n41459 , n41458 , n34257 );
xor ( n41460 , n34257 , n34193 );
and ( n41461 , n34290 , n34298 );
xor ( n41462 , n41460 , n41461 );
and ( n41463 , n41462 , n34287 );
or ( n41464 , n41459 , n41463 );
and ( n41465 , n41464 , n41392 );
or ( n41466 , n41457 , n41465 );
and ( n41467 , n41455 , n41466 );
and ( n41468 , n41464 , n41402 );
or ( n41469 , n41467 , n41468 );
and ( n41470 , n41469 , n33375 );
not ( n41471 , n32968 );
not ( n41472 , n41402 );
not ( n41473 , n41392 );
and ( n41474 , n41473 , n32805 );
and ( n41475 , n41464 , n41392 );
or ( n41476 , n41474 , n41475 );
and ( n41477 , n41472 , n41476 );
and ( n41478 , n41464 , n41402 );
or ( n41479 , n41477 , n41478 );
and ( n41480 , n41471 , n41479 );
not ( n41481 , n41424 );
not ( n41482 , n41428 );
and ( n41483 , n41482 , n41479 );
not ( n41484 , n34747 );
and ( n41485 , n41484 , n34709 );
xor ( n41486 , n34709 , n34625 );
and ( n41487 , n34750 , n34758 );
xor ( n41488 , n41486 , n41487 );
and ( n41489 , n41488 , n34747 );
or ( n41490 , n41485 , n41489 );
and ( n41491 , n41490 , n41428 );
or ( n41492 , n41483 , n41491 );
and ( n41493 , n41481 , n41492 );
not ( n41494 , n35036 );
and ( n41495 , n41494 , n35002 );
xor ( n41496 , n35002 , n34918 );
and ( n41497 , n35039 , n35047 );
xor ( n41498 , n41496 , n41497 );
and ( n41499 , n41498 , n35036 );
or ( n41500 , n41495 , n41499 );
and ( n41501 , n41500 , n41424 );
or ( n41502 , n41493 , n41501 );
and ( n41503 , n41502 , n32968 );
or ( n41504 , n41480 , n41503 );
and ( n41505 , n41504 , n33370 );
and ( n41506 , n32805 , n35062 );
or ( n41507 , C0 , n41454 , n41470 , n41505 , n41506 );
buf ( n41508 , n41507 );
buf ( n41509 , n41508 );
buf ( n41510 , RI15b47b98_312);
buf ( n41511 , n41510 );
buf ( n41512 , n31655 );
buf ( n41513 , n30987 );
buf ( n41514 , n30987 );
buf ( n41515 , RI15b52278_668);
not ( n41516 , n41515 );
buf ( n41517 , RI15b52458_672);
not ( n41518 , n41517 );
and ( n41519 , n41516 , n41518 );
buf ( n41520 , RI15b523e0_671);
and ( n41521 , n41519 , n41520 );
buf ( n41522 , RI15b52368_670);
not ( n41523 , n41522 );
and ( n41524 , n41521 , n41523 );
buf ( n41525 , RI15b522f0_669);
and ( n41526 , n41524 , n41525 );
buf ( n41527 , RI15b51300_635);
buf ( n41528 , RI15b51378_636);
buf ( n41529 , RI15b513f0_637);
buf ( n41530 , RI15b51468_638);
nor ( n41531 , n41527 , n41528 , n41529 , n41530 );
and ( n41532 , n41526 , n41531 );
not ( n41533 , n41532 );
and ( n41534 , n41533 , n34221 );
buf ( n41535 , RI15b534c0_707);
and ( n41536 , n41535 , n41532 );
or ( n41537 , n41534 , n41536 );
buf ( n41538 , n41537 );
buf ( n41539 , n41538 );
buf ( n41540 , n31655 );
buf ( n41541 , n30987 );
and ( n41542 , n33131 , n33133 );
and ( n41543 , n33129 , n41542 );
xor ( n41544 , n33127 , n41543 );
and ( n41545 , n41544 , n33201 );
not ( n41546 , n32562 );
buf ( n41547 , n32562 );
buf ( n41548 , n32562 );
buf ( n41549 , n32562 );
buf ( n41550 , n32562 );
buf ( n41551 , n32562 );
buf ( n41552 , n32562 );
buf ( n41553 , n32562 );
buf ( n41554 , n32562 );
buf ( n41555 , n32562 );
buf ( n41556 , n32562 );
buf ( n41557 , n32562 );
buf ( n41558 , n32562 );
buf ( n41559 , n32562 );
buf ( n41560 , n32562 );
buf ( n41561 , n32562 );
buf ( n41562 , n32562 );
buf ( n41563 , n32562 );
buf ( n41564 , n32562 );
buf ( n41565 , n32562 );
buf ( n41566 , n32562 );
buf ( n41567 , n32562 );
buf ( n41568 , n32562 );
buf ( n41569 , n32562 );
buf ( n41570 , n32562 );
buf ( n41571 , n32562 );
xor ( n41572 , n32546 , n32547 );
or ( n41573 , n32596 , n41572 );
and ( n41574 , n32565 , n41573 );
or ( n41575 , n32567 , n32569 , n32562 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41574 );
and ( n41576 , n41546 , n41575 );
not ( n41577 , n41576 );
and ( n41578 , n41577 , n33127 );
buf ( n41579 , n32753 );
and ( n41580 , n41579 , n41576 );
or ( n41581 , n41578 , n41580 );
and ( n41582 , n41581 , n33189 );
or ( n41583 , n33188 , n33172 );
or ( n41584 , n41583 , n33038 );
or ( n41585 , n41584 , n32924 );
or ( n41586 , n41585 , n32890 );
or ( n41587 , n41586 , n33191 );
or ( n41588 , n41587 , n33193 );
or ( n41589 , n41588 , n33195 );
or ( n41590 , n41589 , n33197 );
or ( n41591 , n41590 , n33199 );
or ( n41592 , n41591 , n33203 );
and ( n41593 , n33127 , n41592 );
or ( n41594 , n41545 , n41582 , n41593 );
and ( n41595 , n41594 , n33208 );
and ( n41596 , n33127 , n39805 );
or ( n41597 , C0 , n41595 , n41596 );
buf ( n41598 , n41597 );
buf ( n41599 , n41598 );
buf ( n41600 , n30987 );
buf ( n41601 , n31655 );
buf ( n41602 , n31655 );
not ( n41603 , n31437 );
buf ( n41604 , RI15b52f98_696);
and ( n41605 , n41603 , n41604 );
buf ( n41606 , RI15b548e8_750);
buf ( n41607 , n41606 );
not ( n41608 , n41607 );
buf ( n41609 , n41608 );
not ( n41610 , n41609 );
buf ( n41611 , RI15b55770_781);
not ( n41612 , n41611 );
buf ( n41613 , RI15b54960_751);
and ( n41614 , n41612 , n41613 );
not ( n41615 , n41613 );
not ( n41616 , n41606 );
xor ( n41617 , n41615 , n41616 );
and ( n41618 , n41617 , n41611 );
or ( n41619 , n41614 , n41618 );
not ( n41620 , n41619 );
buf ( n41621 , n41620 );
buf ( n41622 , n41621 );
not ( n41623 , n41622 );
or ( n41624 , n41610 , n41623 );
not ( n41625 , n41611 );
buf ( n41626 , RI15b549d8_752);
and ( n41627 , n41625 , n41626 );
not ( n41628 , n41626 );
and ( n41629 , n41615 , n41616 );
xor ( n41630 , n41628 , n41629 );
and ( n41631 , n41630 , n41611 );
or ( n41632 , n41627 , n41631 );
not ( n41633 , n41632 );
buf ( n41634 , n41633 );
buf ( n41635 , n41634 );
not ( n41636 , n41635 );
or ( n41637 , n41624 , n41636 );
not ( n41638 , n41611 );
buf ( n41639 , RI15b54a50_753);
and ( n41640 , n41638 , n41639 );
not ( n41641 , n41639 );
and ( n41642 , n41628 , n41629 );
xor ( n41643 , n41641 , n41642 );
and ( n41644 , n41643 , n41611 );
or ( n41645 , n41640 , n41644 );
not ( n41646 , n41645 );
buf ( n41647 , n41646 );
buf ( n41648 , n41647 );
not ( n41649 , n41648 );
or ( n41650 , n41637 , n41649 );
not ( n41651 , n41611 );
buf ( n41652 , RI15b54ac8_754);
and ( n41653 , n41651 , n41652 );
not ( n41654 , n41652 );
and ( n41655 , n41641 , n41642 );
xor ( n41656 , n41654 , n41655 );
and ( n41657 , n41656 , n41611 );
or ( n41658 , n41653 , n41657 );
not ( n41659 , n41658 );
buf ( n41660 , n41659 );
buf ( n41661 , n41660 );
not ( n41662 , n41661 );
or ( n41663 , n41650 , n41662 );
not ( n41664 , n41611 );
buf ( n41665 , RI15b54b40_755);
and ( n41666 , n41664 , n41665 );
not ( n41667 , n41665 );
and ( n41668 , n41654 , n41655 );
xor ( n41669 , n41667 , n41668 );
and ( n41670 , n41669 , n41611 );
or ( n41671 , n41666 , n41670 );
not ( n41672 , n41671 );
buf ( n41673 , n41672 );
buf ( n41674 , n41673 );
not ( n41675 , n41674 );
or ( n41676 , n41663 , n41675 );
not ( n41677 , n41611 );
buf ( n41678 , RI15b54bb8_756);
and ( n41679 , n41677 , n41678 );
not ( n41680 , n41678 );
and ( n41681 , n41667 , n41668 );
xor ( n41682 , n41680 , n41681 );
and ( n41683 , n41682 , n41611 );
or ( n41684 , n41679 , n41683 );
not ( n41685 , n41684 );
buf ( n41686 , n41685 );
buf ( n41687 , n41686 );
not ( n41688 , n41687 );
or ( n41689 , n41676 , n41688 );
not ( n41690 , n41611 );
buf ( n41691 , RI15b54c30_757);
and ( n41692 , n41690 , n41691 );
not ( n41693 , n41691 );
and ( n41694 , n41680 , n41681 );
xor ( n41695 , n41693 , n41694 );
and ( n41696 , n41695 , n41611 );
or ( n41697 , n41692 , n41696 );
not ( n41698 , n41697 );
buf ( n41699 , n41698 );
buf ( n41700 , n41699 );
not ( n41701 , n41700 );
or ( n41702 , n41689 , n41701 );
not ( n41703 , n41611 );
buf ( n41704 , RI15b54ca8_758);
and ( n41705 , n41703 , n41704 );
not ( n41706 , n41704 );
and ( n41707 , n41693 , n41694 );
xor ( n41708 , n41706 , n41707 );
and ( n41709 , n41708 , n41611 );
or ( n41710 , n41705 , n41709 );
not ( n41711 , n41710 );
buf ( n41712 , n41711 );
buf ( n41713 , n41712 );
not ( n41714 , n41713 );
or ( n41715 , n41702 , n41714 );
not ( n41716 , n41611 );
buf ( n41717 , RI15b54d20_759);
and ( n41718 , n41716 , n41717 );
not ( n41719 , n41717 );
and ( n41720 , n41706 , n41707 );
xor ( n41721 , n41719 , n41720 );
and ( n41722 , n41721 , n41611 );
or ( n41723 , n41718 , n41722 );
not ( n41724 , n41723 );
buf ( n41725 , n41724 );
buf ( n41726 , n41725 );
not ( n41727 , n41726 );
or ( n41728 , n41715 , n41727 );
not ( n41729 , n41611 );
buf ( n41730 , RI15b54d98_760);
and ( n41731 , n41729 , n41730 );
not ( n41732 , n41730 );
and ( n41733 , n41719 , n41720 );
xor ( n41734 , n41732 , n41733 );
and ( n41735 , n41734 , n41611 );
or ( n41736 , n41731 , n41735 );
not ( n41737 , n41736 );
buf ( n41738 , n41737 );
buf ( n41739 , n41738 );
not ( n41740 , n41739 );
or ( n41741 , n41728 , n41740 );
not ( n41742 , n41611 );
buf ( n41743 , RI15b54e10_761);
and ( n41744 , n41742 , n41743 );
not ( n41745 , n41743 );
and ( n41746 , n41732 , n41733 );
xor ( n41747 , n41745 , n41746 );
and ( n41748 , n41747 , n41611 );
or ( n41749 , n41744 , n41748 );
not ( n41750 , n41749 );
buf ( n41751 , n41750 );
buf ( n41752 , n41751 );
not ( n41753 , n41752 );
or ( n41754 , n41741 , n41753 );
not ( n41755 , n41611 );
buf ( n41756 , RI15b54e88_762);
and ( n41757 , n41755 , n41756 );
not ( n41758 , n41756 );
and ( n41759 , n41745 , n41746 );
xor ( n41760 , n41758 , n41759 );
and ( n41761 , n41760 , n41611 );
or ( n41762 , n41757 , n41761 );
not ( n41763 , n41762 );
buf ( n41764 , n41763 );
buf ( n41765 , n41764 );
not ( n41766 , n41765 );
or ( n41767 , n41754 , n41766 );
not ( n41768 , n41611 );
buf ( n41769 , RI15b54f00_763);
and ( n41770 , n41768 , n41769 );
not ( n41771 , n41769 );
and ( n41772 , n41758 , n41759 );
xor ( n41773 , n41771 , n41772 );
and ( n41774 , n41773 , n41611 );
or ( n41775 , n41770 , n41774 );
not ( n41776 , n41775 );
buf ( n41777 , n41776 );
buf ( n41778 , n41777 );
not ( n41779 , n41778 );
or ( n41780 , n41767 , n41779 );
not ( n41781 , n41611 );
buf ( n41782 , RI15b54f78_764);
and ( n41783 , n41781 , n41782 );
not ( n41784 , n41782 );
and ( n41785 , n41771 , n41772 );
xor ( n41786 , n41784 , n41785 );
and ( n41787 , n41786 , n41611 );
or ( n41788 , n41783 , n41787 );
not ( n41789 , n41788 );
buf ( n41790 , n41789 );
buf ( n41791 , n41790 );
not ( n41792 , n41791 );
or ( n41793 , n41780 , n41792 );
not ( n41794 , n41611 );
buf ( n41795 , RI15b54ff0_765);
and ( n41796 , n41794 , n41795 );
not ( n41797 , n41795 );
and ( n41798 , n41784 , n41785 );
xor ( n41799 , n41797 , n41798 );
and ( n41800 , n41799 , n41611 );
or ( n41801 , n41796 , n41800 );
not ( n41802 , n41801 );
buf ( n41803 , n41802 );
buf ( n41804 , n41803 );
not ( n41805 , n41804 );
or ( n41806 , n41793 , n41805 );
buf ( n41807 , n41806 );
buf ( n41808 , n41807 );
and ( n41809 , n41808 , n41611 );
not ( n41810 , n41809 );
and ( n41811 , n41810 , n41714 );
xor ( n41812 , n41714 , n41611 );
xor ( n41813 , n41701 , n41611 );
xor ( n41814 , n41688 , n41611 );
xor ( n41815 , n41675 , n41611 );
xor ( n41816 , n41662 , n41611 );
xor ( n41817 , n41649 , n41611 );
xor ( n41818 , n41636 , n41611 );
xor ( n41819 , n41623 , n41611 );
xor ( n41820 , n41610 , n41611 );
and ( n41821 , n41820 , n41611 );
and ( n41822 , n41819 , n41821 );
and ( n41823 , n41818 , n41822 );
and ( n41824 , n41817 , n41823 );
and ( n41825 , n41816 , n41824 );
and ( n41826 , n41815 , n41825 );
and ( n41827 , n41814 , n41826 );
and ( n41828 , n41813 , n41827 );
xor ( n41829 , n41812 , n41828 );
and ( n41830 , n41829 , n41809 );
or ( n41831 , n41811 , n41830 );
and ( n41832 , n41831 , n31437 );
or ( n41833 , n41605 , n41832 );
and ( n41834 , n41833 , n31468 );
or ( n41835 , n31452 , n31451 );
and ( n41836 , n31451 , n41835 );
and ( n41837 , n31497 , n41836 );
not ( n41838 , n41837 );
and ( n41839 , n41838 , n41604 );
buf ( n41840 , RI15b514e0_639);
buf ( n41841 , RI15b515d0_641);
buf ( n41842 , RI15b51648_642);
buf ( n41843 , RI15b516c0_643);
buf ( n41844 , RI15b51738_644);
buf ( n41845 , RI15b517b0_645);
buf ( n41846 , RI15b51828_646);
buf ( n41847 , RI15b518a0_647);
buf ( n41848 , RI15b51918_648);
buf ( n41849 , RI15b51990_649);
buf ( n41850 , RI15b51a08_650);
buf ( n41851 , RI15b51a80_651);
buf ( n41852 , RI15b51af8_652);
buf ( n41853 , RI15b51b70_653);
buf ( n41854 , RI15b51be8_654);
buf ( n41855 , RI15b51c60_655);
buf ( n41856 , RI15b51cd8_656);
buf ( n41857 , RI15b51d50_657);
buf ( n41858 , RI15b51dc8_658);
buf ( n41859 , RI15b51e40_659);
buf ( n41860 , RI15b51eb8_660);
buf ( n41861 , RI15b51f30_661);
buf ( n41862 , RI15b51fa8_662);
buf ( n41863 , RI15b52020_663);
buf ( n41864 , RI15b52098_664);
buf ( n41865 , RI15b52110_665);
buf ( n41866 , RI15b52188_666);
buf ( n41867 , RI15b52200_667);
or ( n41868 , n41840 , n35544 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 );
and ( n41869 , n41515 , n41868 );
not ( n41870 , n41869 );
and ( n41871 , n41870 , n34188 );
and ( n41872 , n40232 , n41869 );
or ( n41873 , n41871 , n41872 );
buf ( n41874 , n41873 );
not ( n41875 , n41874 );
buf ( n41876 , n41875 );
not ( n41877 , n41876 );
not ( n41878 , n41869 );
and ( n41879 , n41878 , n34193 );
and ( n41880 , n40242 , n41869 );
or ( n41881 , n41879 , n41880 );
not ( n41882 , n41881 );
not ( n41883 , n41869 );
and ( n41884 , n41883 , n34195 );
and ( n41885 , n40249 , n41869 );
or ( n41886 , n41884 , n41885 );
and ( n41887 , n41882 , n41886 );
not ( n41888 , n41886 );
not ( n41889 , n41873 );
xor ( n41890 , n41888 , n41889 );
and ( n41891 , n41890 , n41881 );
or ( n41892 , n41887 , n41891 );
not ( n41893 , n41892 );
buf ( n41894 , n41893 );
buf ( n41895 , n41894 );
not ( n41896 , n41895 );
or ( n41897 , n41877 , n41896 );
not ( n41898 , n41881 );
not ( n41899 , n41869 );
and ( n41900 , n41899 , n34208 );
and ( n41901 , n40267 , n41869 );
or ( n41902 , n41900 , n41901 );
and ( n41903 , n41898 , n41902 );
not ( n41904 , n41902 );
and ( n41905 , n41888 , n41889 );
xor ( n41906 , n41904 , n41905 );
and ( n41907 , n41906 , n41881 );
or ( n41908 , n41903 , n41907 );
not ( n41909 , n41908 );
buf ( n41910 , n41909 );
buf ( n41911 , n41910 );
not ( n41912 , n41911 );
or ( n41913 , n41897 , n41912 );
not ( n41914 , n41881 );
not ( n41915 , n41869 );
and ( n41916 , n41915 , n34221 );
and ( n41917 , n40285 , n41869 );
or ( n41918 , n41916 , n41917 );
and ( n41919 , n41914 , n41918 );
not ( n41920 , n41918 );
and ( n41921 , n41904 , n41905 );
xor ( n41922 , n41920 , n41921 );
and ( n41923 , n41922 , n41881 );
or ( n41924 , n41919 , n41923 );
not ( n41925 , n41924 );
buf ( n41926 , n41925 );
buf ( n41927 , n41926 );
not ( n41928 , n41927 );
or ( n41929 , n41913 , n41928 );
not ( n41930 , n41881 );
not ( n41931 , n41869 );
and ( n41932 , n41931 , n34234 );
and ( n41933 , n40303 , n41869 );
or ( n41934 , n41932 , n41933 );
and ( n41935 , n41930 , n41934 );
not ( n41936 , n41934 );
and ( n41937 , n41920 , n41921 );
xor ( n41938 , n41936 , n41937 );
and ( n41939 , n41938 , n41881 );
or ( n41940 , n41935 , n41939 );
not ( n41941 , n41940 );
buf ( n41942 , n41941 );
buf ( n41943 , n41942 );
not ( n41944 , n41943 );
or ( n41945 , n41929 , n41944 );
not ( n41946 , n41881 );
not ( n41947 , n41869 );
and ( n41948 , n41947 , n34247 );
and ( n41949 , n40321 , n41869 );
or ( n41950 , n41948 , n41949 );
and ( n41951 , n41946 , n41950 );
not ( n41952 , n41950 );
and ( n41953 , n41936 , n41937 );
xor ( n41954 , n41952 , n41953 );
and ( n41955 , n41954 , n41881 );
or ( n41956 , n41951 , n41955 );
not ( n41957 , n41956 );
buf ( n41958 , n41957 );
buf ( n41959 , n41958 );
not ( n41960 , n41959 );
or ( n41961 , n41945 , n41960 );
not ( n41962 , n41881 );
not ( n41963 , n41869 );
and ( n41964 , n41963 , n34260 );
and ( n41965 , n40339 , n41869 );
or ( n41966 , n41964 , n41965 );
and ( n41967 , n41962 , n41966 );
not ( n41968 , n41966 );
and ( n41969 , n41952 , n41953 );
xor ( n41970 , n41968 , n41969 );
and ( n41971 , n41970 , n41881 );
or ( n41972 , n41967 , n41971 );
not ( n41973 , n41972 );
buf ( n41974 , n41973 );
buf ( n41975 , n41974 );
not ( n41976 , n41975 );
or ( n41977 , n41961 , n41976 );
not ( n41978 , n41881 );
not ( n41979 , n41869 );
and ( n41980 , n41979 , n34273 );
and ( n41981 , n40357 , n41869 );
or ( n41982 , n41980 , n41981 );
and ( n41983 , n41978 , n41982 );
not ( n41984 , n41982 );
and ( n41985 , n41968 , n41969 );
xor ( n41986 , n41984 , n41985 );
and ( n41987 , n41986 , n41881 );
or ( n41988 , n41983 , n41987 );
not ( n41989 , n41988 );
buf ( n41990 , n41989 );
buf ( n41991 , n41990 );
not ( n41992 , n41991 );
or ( n41993 , n41977 , n41992 );
not ( n41994 , n41881 );
not ( n41995 , n41869 );
and ( n41996 , n41995 , n34379 );
and ( n41997 , n40512 , n41869 );
or ( n41998 , n41996 , n41997 );
and ( n41999 , n41994 , n41998 );
not ( n42000 , n41998 );
and ( n42001 , n41984 , n41985 );
xor ( n42002 , n42000 , n42001 );
and ( n42003 , n42002 , n41881 );
or ( n42004 , n41999 , n42003 );
not ( n42005 , n42004 );
buf ( n42006 , n42005 );
buf ( n42007 , n42006 );
not ( n42008 , n42007 );
or ( n42009 , n41993 , n42008 );
not ( n42010 , n41881 );
not ( n42011 , n41869 );
and ( n42012 , n42011 , n34377 );
and ( n42013 , n40505 , n41869 );
or ( n42014 , n42012 , n42013 );
and ( n42015 , n42010 , n42014 );
not ( n42016 , n42014 );
and ( n42017 , n42000 , n42001 );
xor ( n42018 , n42016 , n42017 );
and ( n42019 , n42018 , n41881 );
or ( n42020 , n42015 , n42019 );
not ( n42021 , n42020 );
buf ( n42022 , n42021 );
buf ( n42023 , n42022 );
not ( n42024 , n42023 );
or ( n42025 , n42009 , n42024 );
not ( n42026 , n41881 );
not ( n42027 , n41869 );
and ( n42028 , n42027 , n34375 );
and ( n42029 , n40498 , n41869 );
or ( n42030 , n42028 , n42029 );
and ( n42031 , n42026 , n42030 );
not ( n42032 , n42030 );
and ( n42033 , n42016 , n42017 );
xor ( n42034 , n42032 , n42033 );
and ( n42035 , n42034 , n41881 );
or ( n42036 , n42031 , n42035 );
not ( n42037 , n42036 );
buf ( n42038 , n42037 );
buf ( n42039 , n42038 );
not ( n42040 , n42039 );
or ( n42041 , n42025 , n42040 );
not ( n42042 , n41881 );
not ( n42043 , n41869 );
and ( n42044 , n42043 , n34373 );
and ( n42045 , n40491 , n41869 );
or ( n42046 , n42044 , n42045 );
and ( n42047 , n42042 , n42046 );
not ( n42048 , n42046 );
and ( n42049 , n42032 , n42033 );
xor ( n42050 , n42048 , n42049 );
and ( n42051 , n42050 , n41881 );
or ( n42052 , n42047 , n42051 );
not ( n42053 , n42052 );
buf ( n42054 , n42053 );
buf ( n42055 , n42054 );
not ( n42056 , n42055 );
or ( n42057 , n42041 , n42056 );
not ( n42058 , n41881 );
not ( n42059 , n41869 );
and ( n42060 , n42059 , n34371 );
and ( n42061 , n40484 , n41869 );
or ( n42062 , n42060 , n42061 );
and ( n42063 , n42058 , n42062 );
not ( n42064 , n42062 );
and ( n42065 , n42048 , n42049 );
xor ( n42066 , n42064 , n42065 );
and ( n42067 , n42066 , n41881 );
or ( n42068 , n42063 , n42067 );
not ( n42069 , n42068 );
buf ( n42070 , n42069 );
buf ( n42071 , n42070 );
not ( n42072 , n42071 );
or ( n42073 , n42057 , n42072 );
not ( n42074 , n41881 );
not ( n42075 , n41869 );
and ( n42076 , n42075 , n34369 );
and ( n42077 , n40477 , n41869 );
or ( n42078 , n42076 , n42077 );
and ( n42079 , n42074 , n42078 );
not ( n42080 , n42078 );
and ( n42081 , n42064 , n42065 );
xor ( n42082 , n42080 , n42081 );
and ( n42083 , n42082 , n41881 );
or ( n42084 , n42079 , n42083 );
not ( n42085 , n42084 );
buf ( n42086 , n42085 );
buf ( n42087 , n42086 );
not ( n42088 , n42087 );
or ( n42089 , n42073 , n42088 );
not ( n42090 , n41881 );
not ( n42091 , n41869 );
and ( n42092 , n42091 , n34367 );
and ( n42093 , n40470 , n41869 );
or ( n42094 , n42092 , n42093 );
and ( n42095 , n42090 , n42094 );
not ( n42096 , n42094 );
and ( n42097 , n42080 , n42081 );
xor ( n42098 , n42096 , n42097 );
and ( n42099 , n42098 , n41881 );
or ( n42100 , n42095 , n42099 );
not ( n42101 , n42100 );
buf ( n42102 , n42101 );
buf ( n42103 , n42102 );
not ( n42104 , n42103 );
or ( n42105 , n42089 , n42104 );
not ( n42106 , n41881 );
not ( n42107 , n41869 );
and ( n42108 , n42107 , n34365 );
and ( n42109 , n40463 , n41869 );
or ( n42110 , n42108 , n42109 );
and ( n42111 , n42106 , n42110 );
not ( n42112 , n42110 );
and ( n42113 , n42096 , n42097 );
xor ( n42114 , n42112 , n42113 );
and ( n42115 , n42114 , n41881 );
or ( n42116 , n42111 , n42115 );
not ( n42117 , n42116 );
buf ( n42118 , n42117 );
buf ( n42119 , n42118 );
not ( n42120 , n42119 );
or ( n42121 , n42105 , n42120 );
buf ( n42122 , n42121 );
buf ( n42123 , n42122 );
and ( n42124 , n42123 , n41881 );
not ( n42125 , n42124 );
and ( n42126 , n42125 , n42008 );
xor ( n42127 , n42008 , n41881 );
xor ( n42128 , n41992 , n41881 );
xor ( n42129 , n41976 , n41881 );
xor ( n42130 , n41960 , n41881 );
xor ( n42131 , n41944 , n41881 );
xor ( n42132 , n41928 , n41881 );
xor ( n42133 , n41912 , n41881 );
xor ( n42134 , n41896 , n41881 );
xor ( n42135 , n41877 , n41881 );
and ( n42136 , n42135 , n41881 );
and ( n42137 , n42134 , n42136 );
and ( n42138 , n42133 , n42137 );
and ( n42139 , n42132 , n42138 );
and ( n42140 , n42131 , n42139 );
and ( n42141 , n42130 , n42140 );
and ( n42142 , n42129 , n42141 );
and ( n42143 , n42128 , n42142 );
xor ( n42144 , n42127 , n42143 );
and ( n42145 , n42144 , n42124 );
or ( n42146 , n42126 , n42145 );
and ( n42147 , n42146 , n41837 );
or ( n42148 , n41839 , n42147 );
and ( n42149 , n42148 , n31521 );
or ( n42150 , n31539 , n31408 );
or ( n42151 , n42150 , n31373 );
or ( n42152 , n42151 , n31540 );
or ( n42153 , n42152 , n31542 );
or ( n42154 , n42153 , n31544 );
or ( n42155 , n42154 , n31546 );
or ( n42156 , n42155 , n31548 );
or ( n42157 , n42156 , n31550 );
or ( n42158 , n42157 , n31552 );
and ( n42159 , n41604 , n42158 );
or ( n42160 , n41834 , n42149 , n42159 );
and ( n42161 , n42160 , n31557 );
and ( n42162 , n41604 , n40154 );
or ( n42163 , C0 , n42161 , n42162 );
buf ( n42164 , n42163 );
buf ( n42165 , n42164 );
buf ( n42166 , n30987 );
not ( n42167 , n40163 );
and ( n42168 , n42167 , n31828 );
not ( n42169 , n31673 );
not ( n42170 , n31657 );
and ( n42171 , n42169 , n31669 , n31665 , n31661 , n42170 );
not ( n42172 , n42171 );
and ( n42173 , n42172 , n31828 );
and ( n42174 , n32235 , n42171 );
or ( n42175 , n42173 , n42174 );
and ( n42176 , n42175 , n40163 );
or ( n42177 , n42168 , n42176 );
and ( n42178 , n42177 , n32498 );
not ( n42179 , n40177 );
and ( n42180 , n42179 , n40182 , n40188 , n40194 , C1 );
not ( n42181 , n42180 );
not ( n42182 , n42171 );
and ( n42183 , n42182 , n31828 );
not ( n42184 , n40373 );
and ( n42185 , n42184 , n40351 );
xor ( n42186 , n40377 , n40389 );
and ( n42187 , n42186 , n40373 );
or ( n42188 , n42185 , n42187 );
and ( n42189 , n42188 , n42171 );
or ( n42190 , n42183 , n42189 );
and ( n42191 , n42181 , n42190 );
and ( n42192 , n42188 , n42180 );
or ( n42193 , n42191 , n42192 );
and ( n42194 , n42193 , n32473 );
not ( n42195 , n32475 );
not ( n42196 , n42180 );
not ( n42197 , n42171 );
and ( n42198 , n42197 , n31828 );
and ( n42199 , n42188 , n42171 );
or ( n42200 , n42198 , n42199 );
and ( n42201 , n42196 , n42200 );
and ( n42202 , n42188 , n42180 );
or ( n42203 , n42201 , n42202 );
and ( n42204 , n42195 , n42203 );
not ( n42205 , n40417 );
and ( n42206 , n42205 , n40425 , n40435 , n40445 , C1 );
not ( n42207 , n42206 );
not ( n42208 , n40413 );
and ( n42209 , n42208 , n40421 , n40430 , n40440 , C1 );
not ( n42210 , n42209 );
and ( n42211 , n42210 , n42203 );
not ( n42212 , n40952 );
and ( n42213 , n42212 , n40931 );
xor ( n42214 , n40956 , n40968 );
and ( n42215 , n42214 , n40952 );
or ( n42216 , n42213 , n42215 );
and ( n42217 , n42216 , n42209 );
or ( n42218 , n42211 , n42217 );
and ( n42219 , n42207 , n42218 );
not ( n42220 , n41247 );
and ( n42221 , n42220 , n41230 );
xor ( n42222 , n41251 , n41263 );
and ( n42223 , n42222 , n41247 );
or ( n42224 , n42221 , n42223 );
and ( n42225 , n42224 , n42206 );
or ( n42226 , n42219 , n42225 );
and ( n42227 , n42226 , n32475 );
or ( n42228 , n42204 , n42227 );
and ( n42229 , n42228 , n32486 );
and ( n42230 , n31828 , n41278 );
or ( n42231 , C0 , n42178 , n42194 , n42229 , n42230 );
buf ( n42232 , n42231 );
buf ( n42233 , n42232 );
buf ( n42234 , n30987 );
not ( n42235 , n40163 );
and ( n42236 , n42235 , n31887 );
not ( n42237 , n31669 );
nor ( n42238 , n31673 , n42237 , n31665 , n31661 , n31657 );
not ( n42239 , n42238 );
and ( n42240 , n42239 , n31887 );
and ( n42241 , n32218 , n42238 );
or ( n42242 , n42240 , n42241 );
and ( n42243 , n42242 , n40163 );
or ( n42244 , n42236 , n42243 );
and ( n42245 , n42244 , n32498 );
not ( n42246 , n40182 );
nor ( n42247 , n40177 , n42246 , n40188 , n40194 , C0 );
not ( n42248 , n42247 );
not ( n42249 , n42238 );
and ( n42250 , n42249 , n31887 );
not ( n42251 , n40373 );
and ( n42252 , n42251 , n40333 );
xor ( n42253 , n40378 , n40388 );
and ( n42254 , n42253 , n40373 );
or ( n42255 , n42252 , n42254 );
and ( n42256 , n42255 , n42238 );
or ( n42257 , n42250 , n42256 );
and ( n42258 , n42248 , n42257 );
and ( n42259 , n42255 , n42247 );
or ( n42260 , n42258 , n42259 );
and ( n42261 , n42260 , n32473 );
not ( n42262 , n32475 );
not ( n42263 , n42247 );
not ( n42264 , n42238 );
and ( n42265 , n42264 , n31887 );
and ( n42266 , n42255 , n42238 );
or ( n42267 , n42265 , n42266 );
and ( n42268 , n42263 , n42267 );
and ( n42269 , n42255 , n42247 );
or ( n42270 , n42268 , n42269 );
and ( n42271 , n42262 , n42270 );
not ( n42272 , n40425 );
nor ( n42273 , n40417 , n42272 , n40435 , n40445 , C0 );
not ( n42274 , n42273 );
not ( n42275 , n40421 );
nor ( n42276 , n40413 , n42275 , n40430 , n40440 , C0 );
not ( n42277 , n42276 );
and ( n42278 , n42277 , n42270 );
not ( n42279 , n40952 );
and ( n42280 , n42279 , n40914 );
xor ( n42281 , n40957 , n40967 );
and ( n42282 , n42281 , n40952 );
or ( n42283 , n42280 , n42282 );
and ( n42284 , n42283 , n42276 );
or ( n42285 , n42278 , n42284 );
and ( n42286 , n42274 , n42285 );
not ( n42287 , n41247 );
and ( n42288 , n42287 , n41213 );
xor ( n42289 , n41252 , n41262 );
and ( n42290 , n42289 , n41247 );
or ( n42291 , n42288 , n42290 );
and ( n42292 , n42291 , n42273 );
or ( n42293 , n42286 , n42292 );
and ( n42294 , n42293 , n32475 );
or ( n42295 , n42271 , n42294 );
and ( n42296 , n42295 , n32486 );
and ( n42297 , n31887 , n41278 );
or ( n42298 , C0 , n42245 , n42261 , n42296 , n42297 );
buf ( n42299 , n42298 );
buf ( n42300 , n42299 );
buf ( n42301 , n31655 );
buf ( n42302 , n30987 );
xor ( n42303 , n34048 , n39933 );
and ( n42304 , n42303 , n31550 );
not ( n42305 , n39979 );
and ( n42306 , n42305 , n34048 );
not ( n42307 , n31026 );
buf ( n42308 , n42307 );
not ( n42309 , n42308 );
not ( n42310 , n42309 );
not ( n42311 , n31022 );
not ( n42312 , n42311 );
buf ( n42313 , n42312 );
buf ( n42314 , n42313 );
not ( n42315 , n42314 );
not ( n42316 , n42315 );
xor ( n42317 , n31018 , n31022 );
not ( n42318 , n42317 );
buf ( n42319 , n42318 );
buf ( n42320 , n42319 );
not ( n42321 , n42320 );
not ( n42322 , n42321 );
and ( n42323 , n31018 , n31022 );
xor ( n42324 , n31014 , n42323 );
not ( n42325 , n42324 );
buf ( n42326 , n42325 );
buf ( n42327 , n42326 );
not ( n42328 , n42327 );
not ( n42329 , n42328 );
nor ( n42330 , n42310 , n42316 , n42322 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42331 , n31206 , n42330 );
nor ( n42332 , n42309 , n42316 , n42322 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42333 , n31208 , n42332 );
nor ( n42334 , n42310 , n42315 , n42322 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42335 , n31210 , n42334 );
nor ( n42336 , n42309 , n42315 , n42322 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42337 , n31212 , n42336 );
nor ( n42338 , n42310 , n42316 , n42321 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42339 , n31214 , n42338 );
nor ( n42340 , n42309 , n42316 , n42321 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42341 , n31216 , n42340 );
nor ( n42342 , n42310 , n42315 , n42321 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42343 , n31218 , n42342 );
nor ( n42344 , n42309 , n42315 , n42321 , n42329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42345 , n31220 , n42344 );
nor ( n42346 , n42310 , n42316 , n42322 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42347 , n31222 , n42346 );
nor ( n42348 , n42309 , n42316 , n42322 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42349 , n31224 , n42348 );
nor ( n42350 , n42310 , n42315 , n42322 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42351 , n31226 , n42350 );
nor ( n42352 , n42309 , n42315 , n42322 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42353 , n31228 , n42352 );
nor ( n42354 , n42310 , n42316 , n42321 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42355 , n31230 , n42354 );
nor ( n42356 , n42309 , n42316 , n42321 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42357 , n31232 , n42356 );
nor ( n42358 , n42310 , n42315 , n42321 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42359 , n31234 , n42358 );
nor ( n42360 , n42309 , n42315 , n42321 , n42328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n42361 , n31236 , n42360 );
or ( n42362 , n42331 , n42333 , n42335 , n42337 , n42339 , n42341 , n42343 , n42345 , n42347 , n42349 , n42351 , n42353 , n42355 , n42357 , n42359 , n42361 );
and ( n42363 , n42362 , n39979 );
or ( n42364 , n42306 , n42363 );
and ( n42365 , n42364 , n31538 );
and ( n42366 , n34048 , n40143 );
or ( n42367 , n42304 , n42365 , n42366 );
and ( n42368 , n42367 , n31557 );
and ( n42369 , n34048 , n40154 );
or ( n42370 , C0 , n42368 , n42369 );
buf ( n42371 , n42370 );
buf ( n42372 , n42371 );
buf ( n42373 , n31655 );
not ( n42374 , n33419 );
and ( n42375 , n42374 , n31566 );
buf ( n42376 , RI15b50b08_618);
buf ( n42377 , RI15b50a90_617);
buf ( n42378 , RI15b50a18_616);
buf ( n42379 , RI15b509a0_615);
and ( n42380 , n33422 , n33463 );
and ( n42381 , n42379 , n42380 );
and ( n42382 , n42378 , n42381 );
and ( n42383 , n42377 , n42382 );
xor ( n42384 , n42376 , n42383 );
xor ( n42385 , n42377 , n42382 );
xor ( n42386 , n42378 , n42381 );
xor ( n42387 , n42379 , n42380 );
and ( n42388 , n33464 , n33701 );
and ( n42389 , n42387 , n42388 );
and ( n42390 , n42386 , n42389 );
and ( n42391 , n42385 , n42390 );
xor ( n42392 , n42384 , n42391 );
and ( n42393 , n42392 , n33419 );
or ( n42394 , n42375 , n42393 );
and ( n42395 , n42394 , n31529 );
not ( n42396 , n33734 );
and ( n42397 , n42396 , n31566 );
not ( n42398 , n33533 );
and ( n42399 , n33422 , n33756 );
and ( n42400 , n42379 , n42399 );
and ( n42401 , n42378 , n42400 );
and ( n42402 , n42377 , n42401 );
xor ( n42403 , n42376 , n42402 );
xor ( n42404 , n42377 , n42401 );
xor ( n42405 , n42378 , n42400 );
xor ( n42406 , n42379 , n42399 );
and ( n42407 , n33757 , n33819 );
and ( n42408 , n42406 , n42407 );
and ( n42409 , n42405 , n42408 );
and ( n42410 , n42404 , n42409 );
xor ( n42411 , n42403 , n42410 );
and ( n42412 , n42398 , n42411 );
and ( n42413 , n33422 , n33841 );
and ( n42414 , n42379 , n42413 );
and ( n42415 , n42378 , n42414 );
and ( n42416 , n42377 , n42415 );
xor ( n42417 , n42376 , n42416 );
xor ( n42418 , n42377 , n42415 );
xor ( n42419 , n42378 , n42414 );
xor ( n42420 , n42379 , n42413 );
or ( n42421 , n33842 , n33921 );
or ( n42422 , n42420 , n42421 );
or ( n42423 , n42419 , n42422 );
or ( n42424 , n42418 , n42423 );
xnor ( n42425 , n42417 , n42424 );
and ( n42426 , n42425 , n33533 );
or ( n42427 , n42412 , n42426 );
and ( n42428 , n42427 , n33734 );
or ( n42429 , n42397 , n42428 );
and ( n42430 , n42429 , n31527 );
and ( n42431 , n31566 , n33942 );
or ( n42432 , n42395 , n42430 , n42431 );
and ( n42433 , n42432 , n31557 );
and ( n42434 , n35488 , n31643 );
not ( n42435 , n31452 );
and ( n42436 , n42435 , n35488 );
and ( n42437 , n31570 , n33967 );
and ( n42438 , n31569 , n42437 );
and ( n42439 , n31568 , n42438 );
and ( n42440 , n31567 , n42439 );
xor ( n42441 , n31566 , n42440 );
and ( n42442 , n42441 , n31452 );
or ( n42443 , n42436 , n42442 );
and ( n42444 , n42443 , n31638 );
and ( n42445 , n35392 , n33973 );
and ( n42446 , n31566 , n33978 );
or ( n42447 , C0 , n42433 , n42434 , n42444 , n42445 , n42446 );
buf ( n42448 , n42447 );
buf ( n42449 , n42448 );
buf ( n42450 , n30987 );
buf ( n42451 , n30987 );
and ( n42452 , n31578 , n31007 );
not ( n42453 , n31077 );
and ( n42454 , n42453 , n34002 );
buf ( n42455 , n42454 );
and ( n42456 , n42455 , n31373 );
not ( n42457 , n31402 );
and ( n42458 , n42457 , n34002 );
buf ( n42459 , n42458 );
and ( n42460 , n42459 , n31408 );
not ( n42461 , n31437 );
and ( n42462 , n42461 , n34002 );
not ( n42463 , n31455 );
and ( n42464 , n42463 , n34044 );
xor ( n42465 , n34002 , n34021 );
and ( n42466 , n42465 , n31455 );
or ( n42467 , n42464 , n42466 );
and ( n42468 , n42467 , n31437 );
or ( n42469 , n42462 , n42468 );
and ( n42470 , n42469 , n31468 );
not ( n42471 , n31497 );
and ( n42472 , n42471 , n34002 );
not ( n42473 , n31454 );
not ( n42474 , n31501 );
and ( n42475 , n42474 , n34044 );
xor ( n42476 , n34045 , n34073 );
and ( n42477 , n42476 , n31501 );
or ( n42478 , n42475 , n42477 );
and ( n42479 , n42473 , n42478 );
and ( n42480 , n42465 , n31454 );
or ( n42481 , n42479 , n42480 );
and ( n42482 , n42481 , n31497 );
or ( n42483 , n42472 , n42482 );
and ( n42484 , n42483 , n31521 );
and ( n42485 , n34002 , n31553 );
or ( n42486 , n42456 , n42460 , n42470 , n42484 , n42485 );
and ( n42487 , n42486 , n31557 );
not ( n42488 , n31452 );
not ( n42489 , n31619 );
and ( n42490 , n42489 , n34101 );
xor ( n42491 , n34102 , n34130 );
and ( n42492 , n42491 , n31619 );
or ( n42493 , n42490 , n42492 );
and ( n42494 , n42488 , n42493 );
and ( n42495 , n34002 , n31452 );
or ( n42496 , n42494 , n42495 );
and ( n42497 , n42496 , n31638 );
buf ( n42498 , n33973 );
and ( n42499 , n34002 , n31650 );
or ( n42500 , C0 , n42452 , n42487 , n42497 , n42498 , n42499 );
buf ( n42501 , n42500 );
buf ( n42502 , n42501 );
buf ( n42503 , n31655 );
buf ( n42504 , n31655 );
buf ( n42505 , n30987 );
not ( n42506 , n34150 );
and ( n42507 , n42506 , n32817 );
not ( n42508 , n34154 );
and ( n42509 , n42508 , n32817 );
and ( n42510 , n32823 , n34154 );
or ( n42511 , n42509 , n42510 );
and ( n42512 , n42511 , n34150 );
or ( n42513 , n42507 , n42512 );
and ( n42514 , n42513 , n33381 );
not ( n42515 , n34184 );
not ( n42516 , n34154 );
and ( n42517 , n42516 , n32817 );
and ( n42518 , n41464 , n34154 );
or ( n42519 , n42517 , n42518 );
and ( n42520 , n42515 , n42519 );
and ( n42521 , n41464 , n34184 );
or ( n42522 , n42520 , n42521 );
and ( n42523 , n42522 , n33375 );
not ( n42524 , n32968 );
not ( n42525 , n34184 );
not ( n42526 , n34154 );
and ( n42527 , n42526 , n32817 );
and ( n42528 , n41464 , n34154 );
or ( n42529 , n42527 , n42528 );
and ( n42530 , n42525 , n42529 );
and ( n42531 , n41464 , n34184 );
or ( n42532 , n42530 , n42531 );
and ( n42533 , n42524 , n42532 );
not ( n42534 , n34355 );
not ( n42535 , n34358 );
and ( n42536 , n42535 , n42532 );
and ( n42537 , n41490 , n34358 );
or ( n42538 , n42536 , n42537 );
and ( n42539 , n42534 , n42538 );
and ( n42540 , n41500 , n34355 );
or ( n42541 , n42539 , n42540 );
and ( n42542 , n42541 , n32968 );
or ( n42543 , n42533 , n42542 );
and ( n42544 , n42543 , n33370 );
and ( n42545 , n32817 , n35062 );
or ( n42546 , C0 , n42514 , n42523 , n42544 , n42545 );
buf ( n42547 , n42546 );
buf ( n42548 , n42547 );
not ( n42549 , n34150 );
and ( n42550 , n42549 , n32716 );
not ( n42551 , n34154 );
and ( n42552 , n42551 , n32716 );
and ( n42553 , n32722 , n34154 );
or ( n42554 , n42552 , n42553 );
and ( n42555 , n42554 , n34150 );
or ( n42556 , n42550 , n42555 );
and ( n42557 , n42556 , n33381 );
not ( n42558 , n34184 );
not ( n42559 , n34154 );
and ( n42560 , n42559 , n32716 );
not ( n42561 , n34287 );
and ( n42562 , n42561 , n34218 );
xor ( n42563 , n34292 , n34296 );
and ( n42564 , n42563 , n34287 );
or ( n42565 , n42562 , n42564 );
and ( n42566 , n42565 , n34154 );
or ( n42567 , n42560 , n42566 );
and ( n42568 , n42558 , n42567 );
and ( n42569 , n42565 , n34184 );
or ( n42570 , n42568 , n42569 );
and ( n42571 , n42570 , n33375 );
not ( n42572 , n32968 );
not ( n42573 , n34184 );
not ( n42574 , n34154 );
and ( n42575 , n42574 , n32716 );
and ( n42576 , n42565 , n34154 );
or ( n42577 , n42575 , n42576 );
and ( n42578 , n42573 , n42577 );
and ( n42579 , n42565 , n34184 );
or ( n42580 , n42578 , n42579 );
and ( n42581 , n42572 , n42580 );
not ( n42582 , n34355 );
not ( n42583 , n34358 );
and ( n42584 , n42583 , n42580 );
not ( n42585 , n34747 );
and ( n42586 , n42585 , n34658 );
xor ( n42587 , n34752 , n34756 );
and ( n42588 , n42587 , n34747 );
or ( n42589 , n42586 , n42588 );
and ( n42590 , n42589 , n34358 );
or ( n42591 , n42584 , n42590 );
and ( n42592 , n42582 , n42591 );
not ( n42593 , n35036 );
and ( n42594 , n42593 , n34951 );
xor ( n42595 , n35041 , n35045 );
and ( n42596 , n42595 , n35036 );
or ( n42597 , n42594 , n42596 );
and ( n42598 , n42597 , n34355 );
or ( n42599 , n42592 , n42598 );
and ( n42600 , n42599 , n32968 );
or ( n42601 , n42581 , n42600 );
and ( n42602 , n42601 , n33370 );
and ( n42603 , n32716 , n35062 );
or ( n42604 , C0 , n42557 , n42571 , n42602 , n42603 );
buf ( n42605 , n42604 );
buf ( n42606 , n42605 );
buf ( n42607 , n30987 );
buf ( n42608 , n31655 );
not ( n42609 , n32953 );
buf ( n42610 , RI15b46e00_283);
and ( n42611 , n42609 , n42610 );
not ( n42612 , n39572 );
and ( n42613 , n42612 , n39555 );
xor ( n42614 , n39555 , n39374 );
xor ( n42615 , n39542 , n39374 );
xor ( n42616 , n39529 , n39374 );
xor ( n42617 , n39516 , n39374 );
xor ( n42618 , n39503 , n39374 );
xor ( n42619 , n39490 , n39374 );
xor ( n42620 , n39477 , n39374 );
xor ( n42621 , n39464 , n39374 );
xor ( n42622 , n39451 , n39374 );
xor ( n42623 , n39438 , n39374 );
xor ( n42624 , n39425 , n39374 );
xor ( n42625 , n39412 , n39374 );
xor ( n42626 , n39399 , n39374 );
and ( n42627 , n39575 , n39577 );
and ( n42628 , n42626 , n42627 );
and ( n42629 , n42625 , n42628 );
and ( n42630 , n42624 , n42629 );
and ( n42631 , n42623 , n42630 );
and ( n42632 , n42622 , n42631 );
and ( n42633 , n42621 , n42632 );
and ( n42634 , n42620 , n42633 );
and ( n42635 , n42619 , n42634 );
and ( n42636 , n42618 , n42635 );
and ( n42637 , n42617 , n42636 );
and ( n42638 , n42616 , n42637 );
and ( n42639 , n42615 , n42638 );
xor ( n42640 , n42614 , n42639 );
and ( n42641 , n42640 , n39572 );
or ( n42642 , n42613 , n42641 );
and ( n42643 , n42642 , n32953 );
or ( n42644 , n42611 , n42643 );
and ( n42645 , n42644 , n33038 );
not ( n42646 , n39586 );
and ( n42647 , n42646 , n42610 );
not ( n42648 , n39775 );
and ( n42649 , n42648 , n39759 );
xor ( n42650 , n39759 , n34193 );
xor ( n42651 , n39747 , n34193 );
xor ( n42652 , n39735 , n34193 );
xor ( n42653 , n39723 , n34193 );
xor ( n42654 , n39711 , n34193 );
xor ( n42655 , n39699 , n34193 );
xor ( n42656 , n39687 , n34193 );
xor ( n42657 , n39675 , n34193 );
xor ( n42658 , n39663 , n34193 );
xor ( n42659 , n39651 , n34193 );
xor ( n42660 , n39639 , n34193 );
xor ( n42661 , n39627 , n34193 );
xor ( n42662 , n39615 , n34193 );
and ( n42663 , n39778 , n39780 );
and ( n42664 , n42662 , n42663 );
and ( n42665 , n42661 , n42664 );
and ( n42666 , n42660 , n42665 );
and ( n42667 , n42659 , n42666 );
and ( n42668 , n42658 , n42667 );
and ( n42669 , n42657 , n42668 );
and ( n42670 , n42656 , n42669 );
and ( n42671 , n42655 , n42670 );
and ( n42672 , n42654 , n42671 );
and ( n42673 , n42653 , n42672 );
and ( n42674 , n42652 , n42673 );
and ( n42675 , n42651 , n42674 );
xor ( n42676 , n42650 , n42675 );
and ( n42677 , n42676 , n39775 );
or ( n42678 , n42649 , n42677 );
and ( n42679 , n42678 , n39586 );
or ( n42680 , n42647 , n42679 );
and ( n42681 , n42680 , n33172 );
and ( n42682 , n42610 , n39795 );
or ( n42683 , n42645 , n42681 , n42682 );
and ( n42684 , n42683 , n33208 );
and ( n42685 , n42610 , n39805 );
or ( n42686 , C0 , n42684 , n42685 );
buf ( n42687 , n42686 );
buf ( n42688 , n42687 );
buf ( n42689 , n31655 );
buf ( n42690 , n30987 );
buf ( n42691 , n30987 );
buf ( n42692 , n31655 );
buf ( n42693 , n31655 );
buf ( n42694 , n30987 );
buf ( n42695 , RI15b4b180_427);
buf ( n42696 , n42695 );
not ( n42697 , n42696 );
buf ( n42698 , n42697 );
not ( n42699 , n42698 );
not ( n42700 , n35592 );
and ( n42701 , n42700 , n33003 );
not ( n42702 , n33003 );
not ( n42703 , n42695 );
xor ( n42704 , n42702 , n42703 );
and ( n42705 , n42704 , n35592 );
or ( n42706 , n42701 , n42705 );
not ( n42707 , n42706 );
buf ( n42708 , n42707 );
buf ( n42709 , n42708 );
not ( n42710 , n42709 );
or ( n42711 , n42699 , n42710 );
buf ( n42712 , n42711 );
buf ( n42713 , n42712 );
and ( n42714 , n42713 , n35592 );
not ( n42715 , n42714 );
and ( n42716 , n42715 , n42699 );
xor ( n42717 , n42699 , n35592 );
xor ( n42718 , n42717 , n35592 );
and ( n42719 , n42718 , n42714 );
or ( n42720 , n42716 , n42719 );
not ( n42721 , n42720 );
not ( n42722 , n42714 );
and ( n42723 , n42722 , n42710 );
xor ( n42724 , n42710 , n35592 );
and ( n42725 , n42717 , n35592 );
xor ( n42726 , n42724 , n42725 );
and ( n42727 , n42726 , n42714 );
or ( n42728 , n42723 , n42727 );
not ( n42729 , n42728 );
and ( n42730 , n42724 , n42725 );
buf ( n42731 , n42730 );
and ( n42732 , n42731 , n42714 );
buf ( n42733 , n42732 );
nor ( n42734 , n42721 , n42729 , n42733 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n42735 , n42734 );
nor ( n42736 , n42720 , n42729 , n42733 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n42737 , n42736 );
or ( n42738 , n42735 , n42737 , C0 , C0 );
buf ( n42739 , RI15b48228_326);
not ( n42740 , n32968 );
buf ( n42741 , RI15b482a0_327);
buf ( n42742 , n42741 );
buf ( n42743 , n42741 );
buf ( n42744 , n42741 );
buf ( n42745 , n42741 );
buf ( n42746 , n42741 );
buf ( n42747 , n42741 );
buf ( n42748 , n42741 );
buf ( n42749 , n42741 );
buf ( n42750 , n42741 );
buf ( n42751 , n42741 );
buf ( n42752 , n42741 );
buf ( n42753 , n42741 );
buf ( n42754 , n42741 );
buf ( n42755 , n42741 );
buf ( n42756 , n42741 );
buf ( n42757 , n42741 );
buf ( n42758 , n42741 );
buf ( n42759 , n42741 );
buf ( n42760 , n42741 );
buf ( n42761 , n42741 );
buf ( n42762 , n42741 );
buf ( n42763 , n42741 );
buf ( n42764 , n42741 );
buf ( n42765 , n42741 );
buf ( n42766 , n42741 );
buf ( n42767 , n42741 );
buf ( n42768 , n42741 );
buf ( n42769 , n42741 );
buf ( n42770 , n42741 );
nor ( n42771 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 );
and ( n42772 , n42738 , n42771 );
buf ( n42773 , n42734 );
buf ( n42774 , n42736 );
or ( n42775 , C0 , n42773 , n42774 , C0 , C0 );
not ( n42776 , n42739 );
buf ( n42777 , n42741 );
buf ( n42778 , n42741 );
buf ( n42779 , n42741 );
buf ( n42780 , n42741 );
buf ( n42781 , n42741 );
buf ( n42782 , n42741 );
buf ( n42783 , n42741 );
buf ( n42784 , n42741 );
buf ( n42785 , n42741 );
buf ( n42786 , n42741 );
buf ( n42787 , n42741 );
buf ( n42788 , n42741 );
buf ( n42789 , n42741 );
buf ( n42790 , n42741 );
buf ( n42791 , n42741 );
buf ( n42792 , n42741 );
buf ( n42793 , n42741 );
buf ( n42794 , n42741 );
buf ( n42795 , n42741 );
buf ( n42796 , n42741 );
buf ( n42797 , n42741 );
buf ( n42798 , n42741 );
buf ( n42799 , n42741 );
buf ( n42800 , n42741 );
buf ( n42801 , n42741 );
buf ( n42802 , n42741 );
buf ( n42803 , n42741 );
buf ( n42804 , n42741 );
buf ( n42805 , n42741 );
nor ( n42806 , n42776 , n32968 , n42741 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 );
and ( n42807 , n42775 , n42806 );
buf ( n42808 , n42734 );
buf ( n42809 , n42736 );
nor ( n42810 , n42720 , n42728 , n42733 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n42811 , n42810 );
or ( n42812 , C0 , n42808 , n42809 , C0 , n42811 );
buf ( n42813 , n42741 );
buf ( n42814 , n42741 );
buf ( n42815 , n42741 );
buf ( n42816 , n42741 );
buf ( n42817 , n42741 );
buf ( n42818 , n42741 );
buf ( n42819 , n42741 );
buf ( n42820 , n42741 );
buf ( n42821 , n42741 );
buf ( n42822 , n42741 );
buf ( n42823 , n42741 );
buf ( n42824 , n42741 );
buf ( n42825 , n42741 );
buf ( n42826 , n42741 );
buf ( n42827 , n42741 );
buf ( n42828 , n42741 );
buf ( n42829 , n42741 );
buf ( n42830 , n42741 );
buf ( n42831 , n42741 );
buf ( n42832 , n42741 );
buf ( n42833 , n42741 );
buf ( n42834 , n42741 );
buf ( n42835 , n42741 );
buf ( n42836 , n42741 );
buf ( n42837 , n42741 );
buf ( n42838 , n42741 );
buf ( n42839 , n42741 );
buf ( n42840 , n42741 );
buf ( n42841 , n42741 );
nor ( n42842 , n42739 , n32968 , n42741 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 );
and ( n42843 , n42812 , n42842 );
or ( n42844 , C0 , n42772 , n42807 , n42843 );
buf ( n42845 , n42844 );
buf ( n42846 , n42845 );
buf ( n42847 , n30987 );
buf ( n42848 , n31655 );
buf ( n42849 , n30987 );
buf ( n42850 , n31655 );
buf ( n42851 , n31655 );
buf ( n42852 , n30987 );
not ( n42853 , n35592 );
and ( n42854 , n42853 , n33003 );
not ( n42855 , n33003 );
not ( n42856 , n42695 );
xor ( n42857 , n42855 , n42856 );
and ( n42858 , n42857 , n35592 );
or ( n42859 , n42854 , n42858 );
not ( n42860 , n42859 );
buf ( n42861 , n42860 );
buf ( n42862 , n42861 );
not ( n42863 , n42862 );
buf ( n42864 , n42863 );
buf ( n42865 , n42864 );
not ( n42866 , n42865 );
buf ( n42867 , n42866 );
not ( n42868 , n42867 );
not ( n42869 , n35592 );
not ( n42870 , n32600 );
not ( n42871 , n32975 );
not ( n42872 , n32976 );
not ( n42873 , n32977 );
not ( n42874 , n32978 );
not ( n42875 , n32979 );
not ( n42876 , n32980 );
not ( n42877 , n32981 );
not ( n42878 , n32982 );
not ( n42879 , n32983 );
not ( n42880 , n32984 );
not ( n42881 , n32985 );
not ( n42882 , n32986 );
not ( n42883 , n32987 );
not ( n42884 , n32988 );
not ( n42885 , n32989 );
not ( n42886 , n32990 );
not ( n42887 , n32991 );
not ( n42888 , n32992 );
not ( n42889 , n32993 );
not ( n42890 , n32994 );
not ( n42891 , n32995 );
not ( n42892 , n32996 );
not ( n42893 , n32997 );
not ( n42894 , n32998 );
not ( n42895 , n32999 );
not ( n42896 , n33000 );
not ( n42897 , n33001 );
not ( n42898 , n33002 );
and ( n42899 , n42855 , n42856 );
and ( n42900 , n42898 , n42899 );
and ( n42901 , n42897 , n42900 );
and ( n42902 , n42896 , n42901 );
and ( n42903 , n42895 , n42902 );
and ( n42904 , n42894 , n42903 );
and ( n42905 , n42893 , n42904 );
and ( n42906 , n42892 , n42905 );
and ( n42907 , n42891 , n42906 );
and ( n42908 , n42890 , n42907 );
and ( n42909 , n42889 , n42908 );
and ( n42910 , n42888 , n42909 );
and ( n42911 , n42887 , n42910 );
and ( n42912 , n42886 , n42911 );
and ( n42913 , n42885 , n42912 );
and ( n42914 , n42884 , n42913 );
and ( n42915 , n42883 , n42914 );
and ( n42916 , n42882 , n42915 );
and ( n42917 , n42881 , n42916 );
and ( n42918 , n42880 , n42917 );
and ( n42919 , n42879 , n42918 );
and ( n42920 , n42878 , n42919 );
and ( n42921 , n42877 , n42920 );
and ( n42922 , n42876 , n42921 );
and ( n42923 , n42875 , n42922 );
and ( n42924 , n42874 , n42923 );
and ( n42925 , n42873 , n42924 );
and ( n42926 , n42872 , n42925 );
and ( n42927 , n42871 , n42926 );
and ( n42928 , n42870 , n42927 );
xor ( n42929 , n42869 , n42928 );
buf ( n42930 , n35592 );
and ( n42931 , n42929 , n42930 );
buf ( n42932 , n42931 );
not ( n42933 , n42932 );
not ( n42934 , n42933 );
not ( n42935 , n42934 );
not ( n42936 , n35592 );
and ( n42937 , n42936 , n32600 );
xor ( n42938 , n42870 , n42927 );
and ( n42939 , n42938 , n35592 );
or ( n42940 , n42937 , n42939 );
not ( n42941 , n42940 );
buf ( n42942 , n42941 );
buf ( n42943 , n42942 );
not ( n42944 , n42943 );
not ( n42945 , n42944 );
not ( n42946 , n35592 );
and ( n42947 , n42946 , n32975 );
xor ( n42948 , n42871 , n42926 );
and ( n42949 , n42948 , n35592 );
or ( n42950 , n42947 , n42949 );
not ( n42951 , n42950 );
buf ( n42952 , n42951 );
buf ( n42953 , n42952 );
not ( n42954 , n42953 );
not ( n42955 , n42954 );
not ( n42956 , n35592 );
and ( n42957 , n42956 , n32976 );
xor ( n42958 , n42872 , n42925 );
and ( n42959 , n42958 , n35592 );
or ( n42960 , n42957 , n42959 );
not ( n42961 , n42960 );
buf ( n42962 , n42961 );
buf ( n42963 , n42962 );
not ( n42964 , n42963 );
not ( n42965 , n42964 );
not ( n42966 , n35592 );
and ( n42967 , n42966 , n32977 );
xor ( n42968 , n42873 , n42924 );
and ( n42969 , n42968 , n35592 );
or ( n42970 , n42967 , n42969 );
not ( n42971 , n42970 );
buf ( n42972 , n42971 );
buf ( n42973 , n42972 );
not ( n42974 , n42973 );
not ( n42975 , n42974 );
not ( n42976 , n35592 );
and ( n42977 , n42976 , n32978 );
xor ( n42978 , n42874 , n42923 );
and ( n42979 , n42978 , n35592 );
or ( n42980 , n42977 , n42979 );
not ( n42981 , n42980 );
buf ( n42982 , n42981 );
buf ( n42983 , n42982 );
not ( n42984 , n42983 );
not ( n42985 , n42984 );
not ( n42986 , n35592 );
and ( n42987 , n42986 , n32979 );
xor ( n42988 , n42875 , n42922 );
and ( n42989 , n42988 , n35592 );
or ( n42990 , n42987 , n42989 );
not ( n42991 , n42990 );
buf ( n42992 , n42991 );
buf ( n42993 , n42992 );
not ( n42994 , n42993 );
not ( n42995 , n42994 );
not ( n42996 , n35592 );
and ( n42997 , n42996 , n32980 );
xor ( n42998 , n42876 , n42921 );
and ( n42999 , n42998 , n35592 );
or ( n43000 , n42997 , n42999 );
not ( n43001 , n43000 );
buf ( n43002 , n43001 );
buf ( n43003 , n43002 );
not ( n43004 , n43003 );
not ( n43005 , n43004 );
not ( n43006 , n35592 );
and ( n43007 , n43006 , n32981 );
xor ( n43008 , n42877 , n42920 );
and ( n43009 , n43008 , n35592 );
or ( n43010 , n43007 , n43009 );
not ( n43011 , n43010 );
buf ( n43012 , n43011 );
buf ( n43013 , n43012 );
not ( n43014 , n43013 );
not ( n43015 , n43014 );
not ( n43016 , n35592 );
and ( n43017 , n43016 , n32982 );
xor ( n43018 , n42878 , n42919 );
and ( n43019 , n43018 , n35592 );
or ( n43020 , n43017 , n43019 );
not ( n43021 , n43020 );
buf ( n43022 , n43021 );
buf ( n43023 , n43022 );
not ( n43024 , n43023 );
not ( n43025 , n43024 );
not ( n43026 , n35592 );
and ( n43027 , n43026 , n32983 );
xor ( n43028 , n42879 , n42918 );
and ( n43029 , n43028 , n35592 );
or ( n43030 , n43027 , n43029 );
not ( n43031 , n43030 );
buf ( n43032 , n43031 );
buf ( n43033 , n43032 );
not ( n43034 , n43033 );
not ( n43035 , n43034 );
not ( n43036 , n35592 );
and ( n43037 , n43036 , n32984 );
xor ( n43038 , n42880 , n42917 );
and ( n43039 , n43038 , n35592 );
or ( n43040 , n43037 , n43039 );
not ( n43041 , n43040 );
buf ( n43042 , n43041 );
buf ( n43043 , n43042 );
not ( n43044 , n43043 );
not ( n43045 , n43044 );
not ( n43046 , n35592 );
and ( n43047 , n43046 , n32985 );
xor ( n43048 , n42881 , n42916 );
and ( n43049 , n43048 , n35592 );
or ( n43050 , n43047 , n43049 );
not ( n43051 , n43050 );
buf ( n43052 , n43051 );
buf ( n43053 , n43052 );
not ( n43054 , n43053 );
not ( n43055 , n43054 );
not ( n43056 , n35592 );
and ( n43057 , n43056 , n32986 );
xor ( n43058 , n42882 , n42915 );
and ( n43059 , n43058 , n35592 );
or ( n43060 , n43057 , n43059 );
not ( n43061 , n43060 );
buf ( n43062 , n43061 );
buf ( n43063 , n43062 );
not ( n43064 , n43063 );
not ( n43065 , n43064 );
not ( n43066 , n35592 );
and ( n43067 , n43066 , n32987 );
xor ( n43068 , n42883 , n42914 );
and ( n43069 , n43068 , n35592 );
or ( n43070 , n43067 , n43069 );
not ( n43071 , n43070 );
buf ( n43072 , n43071 );
buf ( n43073 , n43072 );
not ( n43074 , n43073 );
not ( n43075 , n43074 );
not ( n43076 , n35592 );
and ( n43077 , n43076 , n32988 );
xor ( n43078 , n42884 , n42913 );
and ( n43079 , n43078 , n35592 );
or ( n43080 , n43077 , n43079 );
not ( n43081 , n43080 );
buf ( n43082 , n43081 );
buf ( n43083 , n43082 );
not ( n43084 , n43083 );
not ( n43085 , n43084 );
not ( n43086 , n35592 );
and ( n43087 , n43086 , n32989 );
xor ( n43088 , n42885 , n42912 );
and ( n43089 , n43088 , n35592 );
or ( n43090 , n43087 , n43089 );
not ( n43091 , n43090 );
buf ( n43092 , n43091 );
buf ( n43093 , n43092 );
not ( n43094 , n43093 );
not ( n43095 , n43094 );
not ( n43096 , n35592 );
and ( n43097 , n43096 , n32990 );
xor ( n43098 , n42886 , n42911 );
and ( n43099 , n43098 , n35592 );
or ( n43100 , n43097 , n43099 );
not ( n43101 , n43100 );
buf ( n43102 , n43101 );
buf ( n43103 , n43102 );
not ( n43104 , n43103 );
not ( n43105 , n43104 );
not ( n43106 , n35592 );
and ( n43107 , n43106 , n32991 );
xor ( n43108 , n42887 , n42910 );
and ( n43109 , n43108 , n35592 );
or ( n43110 , n43107 , n43109 );
not ( n43111 , n43110 );
buf ( n43112 , n43111 );
buf ( n43113 , n43112 );
not ( n43114 , n43113 );
not ( n43115 , n43114 );
not ( n43116 , n35592 );
and ( n43117 , n43116 , n32992 );
xor ( n43118 , n42888 , n42909 );
and ( n43119 , n43118 , n35592 );
or ( n43120 , n43117 , n43119 );
not ( n43121 , n43120 );
buf ( n43122 , n43121 );
buf ( n43123 , n43122 );
not ( n43124 , n43123 );
not ( n43125 , n43124 );
not ( n43126 , n35592 );
and ( n43127 , n43126 , n32993 );
xor ( n43128 , n42889 , n42908 );
and ( n43129 , n43128 , n35592 );
or ( n43130 , n43127 , n43129 );
not ( n43131 , n43130 );
buf ( n43132 , n43131 );
buf ( n43133 , n43132 );
not ( n43134 , n43133 );
not ( n43135 , n43134 );
not ( n43136 , n35592 );
and ( n43137 , n43136 , n32994 );
xor ( n43138 , n42890 , n42907 );
and ( n43139 , n43138 , n35592 );
or ( n43140 , n43137 , n43139 );
not ( n43141 , n43140 );
buf ( n43142 , n43141 );
buf ( n43143 , n43142 );
not ( n43144 , n43143 );
not ( n43145 , n43144 );
not ( n43146 , n35592 );
and ( n43147 , n43146 , n32995 );
xor ( n43148 , n42891 , n42906 );
and ( n43149 , n43148 , n35592 );
or ( n43150 , n43147 , n43149 );
not ( n43151 , n43150 );
buf ( n43152 , n43151 );
buf ( n43153 , n43152 );
not ( n43154 , n43153 );
not ( n43155 , n43154 );
not ( n43156 , n35592 );
and ( n43157 , n43156 , n32996 );
xor ( n43158 , n42892 , n42905 );
and ( n43159 , n43158 , n35592 );
or ( n43160 , n43157 , n43159 );
not ( n43161 , n43160 );
buf ( n43162 , n43161 );
buf ( n43163 , n43162 );
not ( n43164 , n43163 );
not ( n43165 , n43164 );
not ( n43166 , n35592 );
and ( n43167 , n43166 , n32997 );
xor ( n43168 , n42893 , n42904 );
and ( n43169 , n43168 , n35592 );
or ( n43170 , n43167 , n43169 );
not ( n43171 , n43170 );
buf ( n43172 , n43171 );
buf ( n43173 , n43172 );
not ( n43174 , n43173 );
not ( n43175 , n43174 );
not ( n43176 , n35592 );
and ( n43177 , n43176 , n32998 );
xor ( n43178 , n42894 , n42903 );
and ( n43179 , n43178 , n35592 );
or ( n43180 , n43177 , n43179 );
not ( n43181 , n43180 );
buf ( n43182 , n43181 );
buf ( n43183 , n43182 );
not ( n43184 , n43183 );
not ( n43185 , n43184 );
not ( n43186 , n35592 );
and ( n43187 , n43186 , n32999 );
xor ( n43188 , n42895 , n42902 );
and ( n43189 , n43188 , n35592 );
or ( n43190 , n43187 , n43189 );
not ( n43191 , n43190 );
buf ( n43192 , n43191 );
buf ( n43193 , n43192 );
not ( n43194 , n43193 );
not ( n43195 , n43194 );
not ( n43196 , n35592 );
and ( n43197 , n43196 , n33000 );
xor ( n43198 , n42896 , n42901 );
and ( n43199 , n43198 , n35592 );
or ( n43200 , n43197 , n43199 );
not ( n43201 , n43200 );
buf ( n43202 , n43201 );
buf ( n43203 , n43202 );
not ( n43204 , n43203 );
not ( n43205 , n43204 );
not ( n43206 , n35592 );
and ( n43207 , n43206 , n33001 );
xor ( n43208 , n42897 , n42900 );
and ( n43209 , n43208 , n35592 );
or ( n43210 , n43207 , n43209 );
not ( n43211 , n43210 );
buf ( n43212 , n43211 );
buf ( n43213 , n43212 );
not ( n43214 , n43213 );
not ( n43215 , n43214 );
not ( n43216 , n35592 );
and ( n43217 , n43216 , n33002 );
xor ( n43218 , n42898 , n42899 );
and ( n43219 , n43218 , n35592 );
or ( n43220 , n43217 , n43219 );
not ( n43221 , n43220 );
buf ( n43222 , n43221 );
buf ( n43223 , n43222 );
not ( n43224 , n43223 );
not ( n43225 , n43224 );
not ( n43226 , n42863 );
and ( n43227 , n43225 , n43226 );
and ( n43228 , n43215 , n43227 );
and ( n43229 , n43205 , n43228 );
and ( n43230 , n43195 , n43229 );
and ( n43231 , n43185 , n43230 );
and ( n43232 , n43175 , n43231 );
and ( n43233 , n43165 , n43232 );
and ( n43234 , n43155 , n43233 );
and ( n43235 , n43145 , n43234 );
and ( n43236 , n43135 , n43235 );
and ( n43237 , n43125 , n43236 );
and ( n43238 , n43115 , n43237 );
and ( n43239 , n43105 , n43238 );
and ( n43240 , n43095 , n43239 );
and ( n43241 , n43085 , n43240 );
and ( n43242 , n43075 , n43241 );
and ( n43243 , n43065 , n43242 );
and ( n43244 , n43055 , n43243 );
and ( n43245 , n43045 , n43244 );
and ( n43246 , n43035 , n43245 );
and ( n43247 , n43025 , n43246 );
and ( n43248 , n43015 , n43247 );
and ( n43249 , n43005 , n43248 );
and ( n43250 , n42995 , n43249 );
and ( n43251 , n42985 , n43250 );
and ( n43252 , n42975 , n43251 );
and ( n43253 , n42965 , n43252 );
and ( n43254 , n42955 , n43253 );
and ( n43255 , n42945 , n43254 );
and ( n43256 , n42935 , n43255 );
not ( n43257 , n43256 );
and ( n43258 , n43257 , n35592 );
buf ( n43259 , n43258 );
not ( n43260 , n43259 );
not ( n43261 , n35592 );
and ( n43262 , n43261 , n43224 );
xor ( n43263 , n43225 , n43226 );
and ( n43264 , n43263 , n35592 );
or ( n43265 , n43262 , n43264 );
and ( n43266 , n43260 , n43265 );
not ( n43267 , n43265 );
not ( n43268 , n42864 );
xor ( n43269 , n43267 , n43268 );
and ( n43270 , n43269 , n43259 );
or ( n43271 , n43266 , n43270 );
not ( n43272 , n43271 );
buf ( n43273 , n43272 );
buf ( n43274 , n43273 );
not ( n43275 , n43274 );
or ( n43276 , n42868 , n43275 );
not ( n43277 , n43259 );
not ( n43278 , n35592 );
and ( n43279 , n43278 , n43214 );
xor ( n43280 , n43215 , n43227 );
and ( n43281 , n43280 , n35592 );
or ( n43282 , n43279 , n43281 );
and ( n43283 , n43277 , n43282 );
not ( n43284 , n43282 );
and ( n43285 , n43267 , n43268 );
xor ( n43286 , n43284 , n43285 );
and ( n43287 , n43286 , n43259 );
or ( n43288 , n43283 , n43287 );
not ( n43289 , n43288 );
buf ( n43290 , n43289 );
buf ( n43291 , n43290 );
not ( n43292 , n43291 );
or ( n43293 , n43276 , n43292 );
not ( n43294 , n43259 );
not ( n43295 , n35592 );
and ( n43296 , n43295 , n43204 );
xor ( n43297 , n43205 , n43228 );
and ( n43298 , n43297 , n35592 );
or ( n43299 , n43296 , n43298 );
and ( n43300 , n43294 , n43299 );
not ( n43301 , n43299 );
and ( n43302 , n43284 , n43285 );
xor ( n43303 , n43301 , n43302 );
and ( n43304 , n43303 , n43259 );
or ( n43305 , n43300 , n43304 );
not ( n43306 , n43305 );
buf ( n43307 , n43306 );
buf ( n43308 , n43307 );
not ( n43309 , n43308 );
or ( n43310 , n43293 , n43309 );
not ( n43311 , n43259 );
not ( n43312 , n35592 );
and ( n43313 , n43312 , n43194 );
xor ( n43314 , n43195 , n43229 );
and ( n43315 , n43314 , n35592 );
or ( n43316 , n43313 , n43315 );
and ( n43317 , n43311 , n43316 );
not ( n43318 , n43316 );
and ( n43319 , n43301 , n43302 );
xor ( n43320 , n43318 , n43319 );
and ( n43321 , n43320 , n43259 );
or ( n43322 , n43317 , n43321 );
not ( n43323 , n43322 );
buf ( n43324 , n43323 );
buf ( n43325 , n43324 );
not ( n43326 , n43325 );
or ( n43327 , n43310 , n43326 );
not ( n43328 , n43259 );
not ( n43329 , n35592 );
and ( n43330 , n43329 , n43184 );
xor ( n43331 , n43185 , n43230 );
and ( n43332 , n43331 , n35592 );
or ( n43333 , n43330 , n43332 );
and ( n43334 , n43328 , n43333 );
not ( n43335 , n43333 );
and ( n43336 , n43318 , n43319 );
xor ( n43337 , n43335 , n43336 );
and ( n43338 , n43337 , n43259 );
or ( n43339 , n43334 , n43338 );
not ( n43340 , n43339 );
buf ( n43341 , n43340 );
buf ( n43342 , n43341 );
not ( n43343 , n43342 );
or ( n43344 , n43327 , n43343 );
not ( n43345 , n43259 );
not ( n43346 , n35592 );
and ( n43347 , n43346 , n43174 );
xor ( n43348 , n43175 , n43231 );
and ( n43349 , n43348 , n35592 );
or ( n43350 , n43347 , n43349 );
and ( n43351 , n43345 , n43350 );
not ( n43352 , n43350 );
and ( n43353 , n43335 , n43336 );
xor ( n43354 , n43352 , n43353 );
and ( n43355 , n43354 , n43259 );
or ( n43356 , n43351 , n43355 );
not ( n43357 , n43356 );
buf ( n43358 , n43357 );
buf ( n43359 , n43358 );
not ( n43360 , n43359 );
or ( n43361 , n43344 , n43360 );
not ( n43362 , n43259 );
not ( n43363 , n35592 );
and ( n43364 , n43363 , n43164 );
xor ( n43365 , n43165 , n43232 );
and ( n43366 , n43365 , n35592 );
or ( n43367 , n43364 , n43366 );
and ( n43368 , n43362 , n43367 );
not ( n43369 , n43367 );
and ( n43370 , n43352 , n43353 );
xor ( n43371 , n43369 , n43370 );
and ( n43372 , n43371 , n43259 );
or ( n43373 , n43368 , n43372 );
not ( n43374 , n43373 );
buf ( n43375 , n43374 );
buf ( n43376 , n43375 );
not ( n43377 , n43376 );
or ( n43378 , n43361 , n43377 );
not ( n43379 , n43259 );
not ( n43380 , n35592 );
and ( n43381 , n43380 , n43154 );
xor ( n43382 , n43155 , n43233 );
and ( n43383 , n43382 , n35592 );
or ( n43384 , n43381 , n43383 );
and ( n43385 , n43379 , n43384 );
not ( n43386 , n43384 );
and ( n43387 , n43369 , n43370 );
xor ( n43388 , n43386 , n43387 );
and ( n43389 , n43388 , n43259 );
or ( n43390 , n43385 , n43389 );
not ( n43391 , n43390 );
buf ( n43392 , n43391 );
buf ( n43393 , n43392 );
not ( n43394 , n43393 );
or ( n43395 , n43378 , n43394 );
not ( n43396 , n43259 );
not ( n43397 , n35592 );
and ( n43398 , n43397 , n43144 );
xor ( n43399 , n43145 , n43234 );
and ( n43400 , n43399 , n35592 );
or ( n43401 , n43398 , n43400 );
and ( n43402 , n43396 , n43401 );
not ( n43403 , n43401 );
and ( n43404 , n43386 , n43387 );
xor ( n43405 , n43403 , n43404 );
and ( n43406 , n43405 , n43259 );
or ( n43407 , n43402 , n43406 );
not ( n43408 , n43407 );
buf ( n43409 , n43408 );
buf ( n43410 , n43409 );
not ( n43411 , n43410 );
or ( n43412 , n43395 , n43411 );
not ( n43413 , n43259 );
not ( n43414 , n35592 );
and ( n43415 , n43414 , n43134 );
xor ( n43416 , n43135 , n43235 );
and ( n43417 , n43416 , n35592 );
or ( n43418 , n43415 , n43417 );
and ( n43419 , n43413 , n43418 );
not ( n43420 , n43418 );
and ( n43421 , n43403 , n43404 );
xor ( n43422 , n43420 , n43421 );
and ( n43423 , n43422 , n43259 );
or ( n43424 , n43419 , n43423 );
not ( n43425 , n43424 );
buf ( n43426 , n43425 );
buf ( n43427 , n43426 );
not ( n43428 , n43427 );
or ( n43429 , n43412 , n43428 );
not ( n43430 , n43259 );
not ( n43431 , n35592 );
and ( n43432 , n43431 , n43124 );
xor ( n43433 , n43125 , n43236 );
and ( n43434 , n43433 , n35592 );
or ( n43435 , n43432 , n43434 );
and ( n43436 , n43430 , n43435 );
not ( n43437 , n43435 );
and ( n43438 , n43420 , n43421 );
xor ( n43439 , n43437 , n43438 );
and ( n43440 , n43439 , n43259 );
or ( n43441 , n43436 , n43440 );
not ( n43442 , n43441 );
buf ( n43443 , n43442 );
buf ( n43444 , n43443 );
not ( n43445 , n43444 );
or ( n43446 , n43429 , n43445 );
not ( n43447 , n43259 );
not ( n43448 , n35592 );
and ( n43449 , n43448 , n43114 );
xor ( n43450 , n43115 , n43237 );
and ( n43451 , n43450 , n35592 );
or ( n43452 , n43449 , n43451 );
and ( n43453 , n43447 , n43452 );
not ( n43454 , n43452 );
and ( n43455 , n43437 , n43438 );
xor ( n43456 , n43454 , n43455 );
and ( n43457 , n43456 , n43259 );
or ( n43458 , n43453 , n43457 );
not ( n43459 , n43458 );
buf ( n43460 , n43459 );
buf ( n43461 , n43460 );
not ( n43462 , n43461 );
or ( n43463 , n43446 , n43462 );
not ( n43464 , n43259 );
not ( n43465 , n35592 );
and ( n43466 , n43465 , n43104 );
xor ( n43467 , n43105 , n43238 );
and ( n43468 , n43467 , n35592 );
or ( n43469 , n43466 , n43468 );
and ( n43470 , n43464 , n43469 );
not ( n43471 , n43469 );
and ( n43472 , n43454 , n43455 );
xor ( n43473 , n43471 , n43472 );
and ( n43474 , n43473 , n43259 );
or ( n43475 , n43470 , n43474 );
not ( n43476 , n43475 );
buf ( n43477 , n43476 );
buf ( n43478 , n43477 );
not ( n43479 , n43478 );
or ( n43480 , n43463 , n43479 );
not ( n43481 , n43259 );
not ( n43482 , n35592 );
and ( n43483 , n43482 , n43094 );
xor ( n43484 , n43095 , n43239 );
and ( n43485 , n43484 , n35592 );
or ( n43486 , n43483 , n43485 );
and ( n43487 , n43481 , n43486 );
not ( n43488 , n43486 );
and ( n43489 , n43471 , n43472 );
xor ( n43490 , n43488 , n43489 );
and ( n43491 , n43490 , n43259 );
or ( n43492 , n43487 , n43491 );
not ( n43493 , n43492 );
buf ( n43494 , n43493 );
buf ( n43495 , n43494 );
not ( n43496 , n43495 );
or ( n43497 , n43480 , n43496 );
not ( n43498 , n43259 );
not ( n43499 , n35592 );
and ( n43500 , n43499 , n43084 );
xor ( n43501 , n43085 , n43240 );
and ( n43502 , n43501 , n35592 );
or ( n43503 , n43500 , n43502 );
and ( n43504 , n43498 , n43503 );
not ( n43505 , n43503 );
and ( n43506 , n43488 , n43489 );
xor ( n43507 , n43505 , n43506 );
and ( n43508 , n43507 , n43259 );
or ( n43509 , n43504 , n43508 );
not ( n43510 , n43509 );
buf ( n43511 , n43510 );
buf ( n43512 , n43511 );
not ( n43513 , n43512 );
or ( n43514 , n43497 , n43513 );
not ( n43515 , n43259 );
not ( n43516 , n35592 );
and ( n43517 , n43516 , n43074 );
xor ( n43518 , n43075 , n43241 );
and ( n43519 , n43518 , n35592 );
or ( n43520 , n43517 , n43519 );
and ( n43521 , n43515 , n43520 );
not ( n43522 , n43520 );
and ( n43523 , n43505 , n43506 );
xor ( n43524 , n43522 , n43523 );
and ( n43525 , n43524 , n43259 );
or ( n43526 , n43521 , n43525 );
not ( n43527 , n43526 );
buf ( n43528 , n43527 );
buf ( n43529 , n43528 );
not ( n43530 , n43529 );
or ( n43531 , n43514 , n43530 );
not ( n43532 , n43259 );
not ( n43533 , n35592 );
and ( n43534 , n43533 , n43064 );
xor ( n43535 , n43065 , n43242 );
and ( n43536 , n43535 , n35592 );
or ( n43537 , n43534 , n43536 );
and ( n43538 , n43532 , n43537 );
not ( n43539 , n43537 );
and ( n43540 , n43522 , n43523 );
xor ( n43541 , n43539 , n43540 );
and ( n43542 , n43541 , n43259 );
or ( n43543 , n43538 , n43542 );
not ( n43544 , n43543 );
buf ( n43545 , n43544 );
buf ( n43546 , n43545 );
not ( n43547 , n43546 );
or ( n43548 , n43531 , n43547 );
not ( n43549 , n43259 );
not ( n43550 , n35592 );
and ( n43551 , n43550 , n43054 );
xor ( n43552 , n43055 , n43243 );
and ( n43553 , n43552 , n35592 );
or ( n43554 , n43551 , n43553 );
and ( n43555 , n43549 , n43554 );
not ( n43556 , n43554 );
and ( n43557 , n43539 , n43540 );
xor ( n43558 , n43556 , n43557 );
and ( n43559 , n43558 , n43259 );
or ( n43560 , n43555 , n43559 );
not ( n43561 , n43560 );
buf ( n43562 , n43561 );
buf ( n43563 , n43562 );
not ( n43564 , n43563 );
or ( n43565 , n43548 , n43564 );
not ( n43566 , n43259 );
not ( n43567 , n35592 );
and ( n43568 , n43567 , n43044 );
xor ( n43569 , n43045 , n43244 );
and ( n43570 , n43569 , n35592 );
or ( n43571 , n43568 , n43570 );
and ( n43572 , n43566 , n43571 );
not ( n43573 , n43571 );
and ( n43574 , n43556 , n43557 );
xor ( n43575 , n43573 , n43574 );
and ( n43576 , n43575 , n43259 );
or ( n43577 , n43572 , n43576 );
not ( n43578 , n43577 );
buf ( n43579 , n43578 );
buf ( n43580 , n43579 );
not ( n43581 , n43580 );
or ( n43582 , n43565 , n43581 );
not ( n43583 , n43259 );
not ( n43584 , n35592 );
and ( n43585 , n43584 , n43034 );
xor ( n43586 , n43035 , n43245 );
and ( n43587 , n43586 , n35592 );
or ( n43588 , n43585 , n43587 );
and ( n43589 , n43583 , n43588 );
not ( n43590 , n43588 );
and ( n43591 , n43573 , n43574 );
xor ( n43592 , n43590 , n43591 );
and ( n43593 , n43592 , n43259 );
or ( n43594 , n43589 , n43593 );
not ( n43595 , n43594 );
buf ( n43596 , n43595 );
buf ( n43597 , n43596 );
not ( n43598 , n43597 );
or ( n43599 , n43582 , n43598 );
not ( n43600 , n43259 );
not ( n43601 , n35592 );
and ( n43602 , n43601 , n43024 );
xor ( n43603 , n43025 , n43246 );
and ( n43604 , n43603 , n35592 );
or ( n43605 , n43602 , n43604 );
and ( n43606 , n43600 , n43605 );
not ( n43607 , n43605 );
and ( n43608 , n43590 , n43591 );
xor ( n43609 , n43607 , n43608 );
and ( n43610 , n43609 , n43259 );
or ( n43611 , n43606 , n43610 );
not ( n43612 , n43611 );
buf ( n43613 , n43612 );
buf ( n43614 , n43613 );
not ( n43615 , n43614 );
or ( n43616 , n43599 , n43615 );
not ( n43617 , n43259 );
not ( n43618 , n35592 );
and ( n43619 , n43618 , n43014 );
xor ( n43620 , n43015 , n43247 );
and ( n43621 , n43620 , n35592 );
or ( n43622 , n43619 , n43621 );
and ( n43623 , n43617 , n43622 );
not ( n43624 , n43622 );
and ( n43625 , n43607 , n43608 );
xor ( n43626 , n43624 , n43625 );
and ( n43627 , n43626 , n43259 );
or ( n43628 , n43623 , n43627 );
not ( n43629 , n43628 );
buf ( n43630 , n43629 );
buf ( n43631 , n43630 );
not ( n43632 , n43631 );
or ( n43633 , n43616 , n43632 );
not ( n43634 , n43259 );
not ( n43635 , n35592 );
and ( n43636 , n43635 , n43004 );
xor ( n43637 , n43005 , n43248 );
and ( n43638 , n43637 , n35592 );
or ( n43639 , n43636 , n43638 );
and ( n43640 , n43634 , n43639 );
not ( n43641 , n43639 );
and ( n43642 , n43624 , n43625 );
xor ( n43643 , n43641 , n43642 );
and ( n43644 , n43643 , n43259 );
or ( n43645 , n43640 , n43644 );
not ( n43646 , n43645 );
buf ( n43647 , n43646 );
buf ( n43648 , n43647 );
not ( n43649 , n43648 );
or ( n43650 , n43633 , n43649 );
not ( n43651 , n43259 );
not ( n43652 , n35592 );
and ( n43653 , n43652 , n42994 );
xor ( n43654 , n42995 , n43249 );
and ( n43655 , n43654 , n35592 );
or ( n43656 , n43653 , n43655 );
and ( n43657 , n43651 , n43656 );
not ( n43658 , n43656 );
and ( n43659 , n43641 , n43642 );
xor ( n43660 , n43658 , n43659 );
and ( n43661 , n43660 , n43259 );
or ( n43662 , n43657 , n43661 );
not ( n43663 , n43662 );
buf ( n43664 , n43663 );
buf ( n43665 , n43664 );
not ( n43666 , n43665 );
or ( n43667 , n43650 , n43666 );
not ( n43668 , n43259 );
not ( n43669 , n35592 );
and ( n43670 , n43669 , n42984 );
xor ( n43671 , n42985 , n43250 );
and ( n43672 , n43671 , n35592 );
or ( n43673 , n43670 , n43672 );
and ( n43674 , n43668 , n43673 );
not ( n43675 , n43673 );
and ( n43676 , n43658 , n43659 );
xor ( n43677 , n43675 , n43676 );
and ( n43678 , n43677 , n43259 );
or ( n43679 , n43674 , n43678 );
not ( n43680 , n43679 );
buf ( n43681 , n43680 );
buf ( n43682 , n43681 );
not ( n43683 , n43682 );
or ( n43684 , n43667 , n43683 );
not ( n43685 , n43259 );
not ( n43686 , n35592 );
and ( n43687 , n43686 , n42974 );
xor ( n43688 , n42975 , n43251 );
and ( n43689 , n43688 , n35592 );
or ( n43690 , n43687 , n43689 );
and ( n43691 , n43685 , n43690 );
not ( n43692 , n43690 );
and ( n43693 , n43675 , n43676 );
xor ( n43694 , n43692 , n43693 );
and ( n43695 , n43694 , n43259 );
or ( n43696 , n43691 , n43695 );
not ( n43697 , n43696 );
buf ( n43698 , n43697 );
buf ( n43699 , n43698 );
not ( n43700 , n43699 );
or ( n43701 , n43684 , n43700 );
not ( n43702 , n43259 );
not ( n43703 , n35592 );
and ( n43704 , n43703 , n42964 );
xor ( n43705 , n42965 , n43252 );
and ( n43706 , n43705 , n35592 );
or ( n43707 , n43704 , n43706 );
and ( n43708 , n43702 , n43707 );
not ( n43709 , n43707 );
and ( n43710 , n43692 , n43693 );
xor ( n43711 , n43709 , n43710 );
and ( n43712 , n43711 , n43259 );
or ( n43713 , n43708 , n43712 );
not ( n43714 , n43713 );
buf ( n43715 , n43714 );
buf ( n43716 , n43715 );
not ( n43717 , n43716 );
or ( n43718 , n43701 , n43717 );
not ( n43719 , n43259 );
not ( n43720 , n35592 );
and ( n43721 , n43720 , n42954 );
xor ( n43722 , n42955 , n43253 );
and ( n43723 , n43722 , n35592 );
or ( n43724 , n43721 , n43723 );
and ( n43725 , n43719 , n43724 );
not ( n43726 , n43724 );
and ( n43727 , n43709 , n43710 );
xor ( n43728 , n43726 , n43727 );
and ( n43729 , n43728 , n43259 );
or ( n43730 , n43725 , n43729 );
not ( n43731 , n43730 );
buf ( n43732 , n43731 );
buf ( n43733 , n43732 );
not ( n43734 , n43733 );
or ( n43735 , n43718 , n43734 );
not ( n43736 , n43259 );
not ( n43737 , n35592 );
and ( n43738 , n43737 , n42944 );
xor ( n43739 , n42945 , n43254 );
and ( n43740 , n43739 , n35592 );
or ( n43741 , n43738 , n43740 );
and ( n43742 , n43736 , n43741 );
not ( n43743 , n43741 );
and ( n43744 , n43726 , n43727 );
xor ( n43745 , n43743 , n43744 );
and ( n43746 , n43745 , n43259 );
or ( n43747 , n43742 , n43746 );
not ( n43748 , n43747 );
buf ( n43749 , n43748 );
buf ( n43750 , n43749 );
not ( n43751 , n43750 );
or ( n43752 , n43735 , n43751 );
buf ( n43753 , n43752 );
buf ( n43754 , n43753 );
and ( n43755 , n43754 , n43259 );
not ( n43756 , n43755 );
and ( n43757 , n43756 , n43360 );
xor ( n43758 , n43360 , n43259 );
xor ( n43759 , n43343 , n43259 );
xor ( n43760 , n43326 , n43259 );
xor ( n43761 , n43309 , n43259 );
xor ( n43762 , n43292 , n43259 );
xor ( n43763 , n43275 , n43259 );
xor ( n43764 , n42868 , n43259 );
and ( n43765 , n43764 , n43259 );
and ( n43766 , n43763 , n43765 );
and ( n43767 , n43762 , n43766 );
and ( n43768 , n43761 , n43767 );
and ( n43769 , n43760 , n43768 );
and ( n43770 , n43759 , n43769 );
xor ( n43771 , n43758 , n43770 );
and ( n43772 , n43771 , n43755 );
or ( n43773 , n43757 , n43772 );
and ( n43774 , n32961 , n32957 , n32959 );
and ( n43775 , n43773 , n43774 );
not ( n43776 , n35592 );
and ( n43777 , n43776 , n33002 );
not ( n43778 , n33002 );
not ( n43779 , n33003 );
not ( n43780 , n42695 );
and ( n43781 , n43779 , n43780 );
xor ( n43782 , n43778 , n43781 );
and ( n43783 , n43782 , n35592 );
or ( n43784 , n43777 , n43783 );
not ( n43785 , n43784 );
buf ( n43786 , n43785 );
buf ( n43787 , n43786 );
not ( n43788 , n43787 );
buf ( n43789 , n43788 );
buf ( n43790 , n43789 );
not ( n43791 , n43790 );
buf ( n43792 , n43791 );
not ( n43793 , n43792 );
not ( n43794 , n35592 );
not ( n43795 , n32600 );
not ( n43796 , n32975 );
not ( n43797 , n32976 );
not ( n43798 , n32977 );
not ( n43799 , n32978 );
not ( n43800 , n32979 );
not ( n43801 , n32980 );
not ( n43802 , n32981 );
not ( n43803 , n32982 );
not ( n43804 , n32983 );
not ( n43805 , n32984 );
not ( n43806 , n32985 );
not ( n43807 , n32986 );
not ( n43808 , n32987 );
not ( n43809 , n32988 );
not ( n43810 , n32989 );
not ( n43811 , n32990 );
not ( n43812 , n32991 );
not ( n43813 , n32992 );
not ( n43814 , n32993 );
not ( n43815 , n32994 );
not ( n43816 , n32995 );
not ( n43817 , n32996 );
not ( n43818 , n32997 );
not ( n43819 , n32998 );
not ( n43820 , n32999 );
not ( n43821 , n33000 );
not ( n43822 , n33001 );
and ( n43823 , n43778 , n43781 );
and ( n43824 , n43822 , n43823 );
and ( n43825 , n43821 , n43824 );
and ( n43826 , n43820 , n43825 );
and ( n43827 , n43819 , n43826 );
and ( n43828 , n43818 , n43827 );
and ( n43829 , n43817 , n43828 );
and ( n43830 , n43816 , n43829 );
and ( n43831 , n43815 , n43830 );
and ( n43832 , n43814 , n43831 );
and ( n43833 , n43813 , n43832 );
and ( n43834 , n43812 , n43833 );
and ( n43835 , n43811 , n43834 );
and ( n43836 , n43810 , n43835 );
and ( n43837 , n43809 , n43836 );
and ( n43838 , n43808 , n43837 );
and ( n43839 , n43807 , n43838 );
and ( n43840 , n43806 , n43839 );
and ( n43841 , n43805 , n43840 );
and ( n43842 , n43804 , n43841 );
and ( n43843 , n43803 , n43842 );
and ( n43844 , n43802 , n43843 );
and ( n43845 , n43801 , n43844 );
and ( n43846 , n43800 , n43845 );
and ( n43847 , n43799 , n43846 );
and ( n43848 , n43798 , n43847 );
and ( n43849 , n43797 , n43848 );
and ( n43850 , n43796 , n43849 );
and ( n43851 , n43795 , n43850 );
xor ( n43852 , n43794 , n43851 );
buf ( n43853 , n35592 );
and ( n43854 , n43852 , n43853 );
buf ( n43855 , n43854 );
not ( n43856 , n43855 );
not ( n43857 , n43856 );
not ( n43858 , n43857 );
not ( n43859 , n35592 );
and ( n43860 , n43859 , n32600 );
xor ( n43861 , n43795 , n43850 );
and ( n43862 , n43861 , n35592 );
or ( n43863 , n43860 , n43862 );
not ( n43864 , n43863 );
buf ( n43865 , n43864 );
buf ( n43866 , n43865 );
not ( n43867 , n43866 );
not ( n43868 , n43867 );
not ( n43869 , n35592 );
and ( n43870 , n43869 , n32975 );
xor ( n43871 , n43796 , n43849 );
and ( n43872 , n43871 , n35592 );
or ( n43873 , n43870 , n43872 );
not ( n43874 , n43873 );
buf ( n43875 , n43874 );
buf ( n43876 , n43875 );
not ( n43877 , n43876 );
not ( n43878 , n43877 );
not ( n43879 , n35592 );
and ( n43880 , n43879 , n32976 );
xor ( n43881 , n43797 , n43848 );
and ( n43882 , n43881 , n35592 );
or ( n43883 , n43880 , n43882 );
not ( n43884 , n43883 );
buf ( n43885 , n43884 );
buf ( n43886 , n43885 );
not ( n43887 , n43886 );
not ( n43888 , n43887 );
not ( n43889 , n35592 );
and ( n43890 , n43889 , n32977 );
xor ( n43891 , n43798 , n43847 );
and ( n43892 , n43891 , n35592 );
or ( n43893 , n43890 , n43892 );
not ( n43894 , n43893 );
buf ( n43895 , n43894 );
buf ( n43896 , n43895 );
not ( n43897 , n43896 );
not ( n43898 , n43897 );
not ( n43899 , n35592 );
and ( n43900 , n43899 , n32978 );
xor ( n43901 , n43799 , n43846 );
and ( n43902 , n43901 , n35592 );
or ( n43903 , n43900 , n43902 );
not ( n43904 , n43903 );
buf ( n43905 , n43904 );
buf ( n43906 , n43905 );
not ( n43907 , n43906 );
not ( n43908 , n43907 );
not ( n43909 , n35592 );
and ( n43910 , n43909 , n32979 );
xor ( n43911 , n43800 , n43845 );
and ( n43912 , n43911 , n35592 );
or ( n43913 , n43910 , n43912 );
not ( n43914 , n43913 );
buf ( n43915 , n43914 );
buf ( n43916 , n43915 );
not ( n43917 , n43916 );
not ( n43918 , n43917 );
not ( n43919 , n35592 );
and ( n43920 , n43919 , n32980 );
xor ( n43921 , n43801 , n43844 );
and ( n43922 , n43921 , n35592 );
or ( n43923 , n43920 , n43922 );
not ( n43924 , n43923 );
buf ( n43925 , n43924 );
buf ( n43926 , n43925 );
not ( n43927 , n43926 );
not ( n43928 , n43927 );
not ( n43929 , n35592 );
and ( n43930 , n43929 , n32981 );
xor ( n43931 , n43802 , n43843 );
and ( n43932 , n43931 , n35592 );
or ( n43933 , n43930 , n43932 );
not ( n43934 , n43933 );
buf ( n43935 , n43934 );
buf ( n43936 , n43935 );
not ( n43937 , n43936 );
not ( n43938 , n43937 );
not ( n43939 , n35592 );
and ( n43940 , n43939 , n32982 );
xor ( n43941 , n43803 , n43842 );
and ( n43942 , n43941 , n35592 );
or ( n43943 , n43940 , n43942 );
not ( n43944 , n43943 );
buf ( n43945 , n43944 );
buf ( n43946 , n43945 );
not ( n43947 , n43946 );
not ( n43948 , n43947 );
not ( n43949 , n35592 );
and ( n43950 , n43949 , n32983 );
xor ( n43951 , n43804 , n43841 );
and ( n43952 , n43951 , n35592 );
or ( n43953 , n43950 , n43952 );
not ( n43954 , n43953 );
buf ( n43955 , n43954 );
buf ( n43956 , n43955 );
not ( n43957 , n43956 );
not ( n43958 , n43957 );
not ( n43959 , n35592 );
and ( n43960 , n43959 , n32984 );
xor ( n43961 , n43805 , n43840 );
and ( n43962 , n43961 , n35592 );
or ( n43963 , n43960 , n43962 );
not ( n43964 , n43963 );
buf ( n43965 , n43964 );
buf ( n43966 , n43965 );
not ( n43967 , n43966 );
not ( n43968 , n43967 );
not ( n43969 , n35592 );
and ( n43970 , n43969 , n32985 );
xor ( n43971 , n43806 , n43839 );
and ( n43972 , n43971 , n35592 );
or ( n43973 , n43970 , n43972 );
not ( n43974 , n43973 );
buf ( n43975 , n43974 );
buf ( n43976 , n43975 );
not ( n43977 , n43976 );
not ( n43978 , n43977 );
not ( n43979 , n35592 );
and ( n43980 , n43979 , n32986 );
xor ( n43981 , n43807 , n43838 );
and ( n43982 , n43981 , n35592 );
or ( n43983 , n43980 , n43982 );
not ( n43984 , n43983 );
buf ( n43985 , n43984 );
buf ( n43986 , n43985 );
not ( n43987 , n43986 );
not ( n43988 , n43987 );
not ( n43989 , n35592 );
and ( n43990 , n43989 , n32987 );
xor ( n43991 , n43808 , n43837 );
and ( n43992 , n43991 , n35592 );
or ( n43993 , n43990 , n43992 );
not ( n43994 , n43993 );
buf ( n43995 , n43994 );
buf ( n43996 , n43995 );
not ( n43997 , n43996 );
not ( n43998 , n43997 );
not ( n43999 , n35592 );
and ( n44000 , n43999 , n32988 );
xor ( n44001 , n43809 , n43836 );
and ( n44002 , n44001 , n35592 );
or ( n44003 , n44000 , n44002 );
not ( n44004 , n44003 );
buf ( n44005 , n44004 );
buf ( n44006 , n44005 );
not ( n44007 , n44006 );
not ( n44008 , n44007 );
not ( n44009 , n35592 );
and ( n44010 , n44009 , n32989 );
xor ( n44011 , n43810 , n43835 );
and ( n44012 , n44011 , n35592 );
or ( n44013 , n44010 , n44012 );
not ( n44014 , n44013 );
buf ( n44015 , n44014 );
buf ( n44016 , n44015 );
not ( n44017 , n44016 );
not ( n44018 , n44017 );
not ( n44019 , n35592 );
and ( n44020 , n44019 , n32990 );
xor ( n44021 , n43811 , n43834 );
and ( n44022 , n44021 , n35592 );
or ( n44023 , n44020 , n44022 );
not ( n44024 , n44023 );
buf ( n44025 , n44024 );
buf ( n44026 , n44025 );
not ( n44027 , n44026 );
not ( n44028 , n44027 );
not ( n44029 , n35592 );
and ( n44030 , n44029 , n32991 );
xor ( n44031 , n43812 , n43833 );
and ( n44032 , n44031 , n35592 );
or ( n44033 , n44030 , n44032 );
not ( n44034 , n44033 );
buf ( n44035 , n44034 );
buf ( n44036 , n44035 );
not ( n44037 , n44036 );
not ( n44038 , n44037 );
not ( n44039 , n35592 );
and ( n44040 , n44039 , n32992 );
xor ( n44041 , n43813 , n43832 );
and ( n44042 , n44041 , n35592 );
or ( n44043 , n44040 , n44042 );
not ( n44044 , n44043 );
buf ( n44045 , n44044 );
buf ( n44046 , n44045 );
not ( n44047 , n44046 );
not ( n44048 , n44047 );
not ( n44049 , n35592 );
and ( n44050 , n44049 , n32993 );
xor ( n44051 , n43814 , n43831 );
and ( n44052 , n44051 , n35592 );
or ( n44053 , n44050 , n44052 );
not ( n44054 , n44053 );
buf ( n44055 , n44054 );
buf ( n44056 , n44055 );
not ( n44057 , n44056 );
not ( n44058 , n44057 );
not ( n44059 , n35592 );
and ( n44060 , n44059 , n32994 );
xor ( n44061 , n43815 , n43830 );
and ( n44062 , n44061 , n35592 );
or ( n44063 , n44060 , n44062 );
not ( n44064 , n44063 );
buf ( n44065 , n44064 );
buf ( n44066 , n44065 );
not ( n44067 , n44066 );
not ( n44068 , n44067 );
not ( n44069 , n35592 );
and ( n44070 , n44069 , n32995 );
xor ( n44071 , n43816 , n43829 );
and ( n44072 , n44071 , n35592 );
or ( n44073 , n44070 , n44072 );
not ( n44074 , n44073 );
buf ( n44075 , n44074 );
buf ( n44076 , n44075 );
not ( n44077 , n44076 );
not ( n44078 , n44077 );
not ( n44079 , n35592 );
and ( n44080 , n44079 , n32996 );
xor ( n44081 , n43817 , n43828 );
and ( n44082 , n44081 , n35592 );
or ( n44083 , n44080 , n44082 );
not ( n44084 , n44083 );
buf ( n44085 , n44084 );
buf ( n44086 , n44085 );
not ( n44087 , n44086 );
not ( n44088 , n44087 );
not ( n44089 , n35592 );
and ( n44090 , n44089 , n32997 );
xor ( n44091 , n43818 , n43827 );
and ( n44092 , n44091 , n35592 );
or ( n44093 , n44090 , n44092 );
not ( n44094 , n44093 );
buf ( n44095 , n44094 );
buf ( n44096 , n44095 );
not ( n44097 , n44096 );
not ( n44098 , n44097 );
not ( n44099 , n35592 );
and ( n44100 , n44099 , n32998 );
xor ( n44101 , n43819 , n43826 );
and ( n44102 , n44101 , n35592 );
or ( n44103 , n44100 , n44102 );
not ( n44104 , n44103 );
buf ( n44105 , n44104 );
buf ( n44106 , n44105 );
not ( n44107 , n44106 );
not ( n44108 , n44107 );
not ( n44109 , n35592 );
and ( n44110 , n44109 , n32999 );
xor ( n44111 , n43820 , n43825 );
and ( n44112 , n44111 , n35592 );
or ( n44113 , n44110 , n44112 );
not ( n44114 , n44113 );
buf ( n44115 , n44114 );
buf ( n44116 , n44115 );
not ( n44117 , n44116 );
not ( n44118 , n44117 );
not ( n44119 , n35592 );
and ( n44120 , n44119 , n33000 );
xor ( n44121 , n43821 , n43824 );
and ( n44122 , n44121 , n35592 );
or ( n44123 , n44120 , n44122 );
not ( n44124 , n44123 );
buf ( n44125 , n44124 );
buf ( n44126 , n44125 );
not ( n44127 , n44126 );
not ( n44128 , n44127 );
not ( n44129 , n35592 );
and ( n44130 , n44129 , n33001 );
xor ( n44131 , n43822 , n43823 );
and ( n44132 , n44131 , n35592 );
or ( n44133 , n44130 , n44132 );
not ( n44134 , n44133 );
buf ( n44135 , n44134 );
buf ( n44136 , n44135 );
not ( n44137 , n44136 );
not ( n44138 , n44137 );
not ( n44139 , n43788 );
and ( n44140 , n44138 , n44139 );
and ( n44141 , n44128 , n44140 );
and ( n44142 , n44118 , n44141 );
and ( n44143 , n44108 , n44142 );
and ( n44144 , n44098 , n44143 );
and ( n44145 , n44088 , n44144 );
and ( n44146 , n44078 , n44145 );
and ( n44147 , n44068 , n44146 );
and ( n44148 , n44058 , n44147 );
and ( n44149 , n44048 , n44148 );
and ( n44150 , n44038 , n44149 );
and ( n44151 , n44028 , n44150 );
and ( n44152 , n44018 , n44151 );
and ( n44153 , n44008 , n44152 );
and ( n44154 , n43998 , n44153 );
and ( n44155 , n43988 , n44154 );
and ( n44156 , n43978 , n44155 );
and ( n44157 , n43968 , n44156 );
and ( n44158 , n43958 , n44157 );
and ( n44159 , n43948 , n44158 );
and ( n44160 , n43938 , n44159 );
and ( n44161 , n43928 , n44160 );
and ( n44162 , n43918 , n44161 );
and ( n44163 , n43908 , n44162 );
and ( n44164 , n43898 , n44163 );
and ( n44165 , n43888 , n44164 );
and ( n44166 , n43878 , n44165 );
and ( n44167 , n43868 , n44166 );
and ( n44168 , n43858 , n44167 );
not ( n44169 , n44168 );
and ( n44170 , n44169 , n35592 );
buf ( n44171 , n44170 );
not ( n44172 , n44171 );
not ( n44173 , n35592 );
and ( n44174 , n44173 , n44137 );
xor ( n44175 , n44138 , n44139 );
and ( n44176 , n44175 , n35592 );
or ( n44177 , n44174 , n44176 );
and ( n44178 , n44172 , n44177 );
not ( n44179 , n44177 );
not ( n44180 , n43789 );
xor ( n44181 , n44179 , n44180 );
and ( n44182 , n44181 , n44171 );
or ( n44183 , n44178 , n44182 );
not ( n44184 , n44183 );
buf ( n44185 , n44184 );
buf ( n44186 , n44185 );
not ( n44187 , n44186 );
or ( n44188 , n43793 , n44187 );
not ( n44189 , n44171 );
not ( n44190 , n35592 );
and ( n44191 , n44190 , n44127 );
xor ( n44192 , n44128 , n44140 );
and ( n44193 , n44192 , n35592 );
or ( n44194 , n44191 , n44193 );
and ( n44195 , n44189 , n44194 );
not ( n44196 , n44194 );
and ( n44197 , n44179 , n44180 );
xor ( n44198 , n44196 , n44197 );
and ( n44199 , n44198 , n44171 );
or ( n44200 , n44195 , n44199 );
not ( n44201 , n44200 );
buf ( n44202 , n44201 );
buf ( n44203 , n44202 );
not ( n44204 , n44203 );
or ( n44205 , n44188 , n44204 );
not ( n44206 , n44171 );
not ( n44207 , n35592 );
and ( n44208 , n44207 , n44117 );
xor ( n44209 , n44118 , n44141 );
and ( n44210 , n44209 , n35592 );
or ( n44211 , n44208 , n44210 );
and ( n44212 , n44206 , n44211 );
not ( n44213 , n44211 );
and ( n44214 , n44196 , n44197 );
xor ( n44215 , n44213 , n44214 );
and ( n44216 , n44215 , n44171 );
or ( n44217 , n44212 , n44216 );
not ( n44218 , n44217 );
buf ( n44219 , n44218 );
buf ( n44220 , n44219 );
not ( n44221 , n44220 );
or ( n44222 , n44205 , n44221 );
not ( n44223 , n44171 );
not ( n44224 , n35592 );
and ( n44225 , n44224 , n44107 );
xor ( n44226 , n44108 , n44142 );
and ( n44227 , n44226 , n35592 );
or ( n44228 , n44225 , n44227 );
and ( n44229 , n44223 , n44228 );
not ( n44230 , n44228 );
and ( n44231 , n44213 , n44214 );
xor ( n44232 , n44230 , n44231 );
and ( n44233 , n44232 , n44171 );
or ( n44234 , n44229 , n44233 );
not ( n44235 , n44234 );
buf ( n44236 , n44235 );
buf ( n44237 , n44236 );
not ( n44238 , n44237 );
or ( n44239 , n44222 , n44238 );
not ( n44240 , n44171 );
not ( n44241 , n35592 );
and ( n44242 , n44241 , n44097 );
xor ( n44243 , n44098 , n44143 );
and ( n44244 , n44243 , n35592 );
or ( n44245 , n44242 , n44244 );
and ( n44246 , n44240 , n44245 );
not ( n44247 , n44245 );
and ( n44248 , n44230 , n44231 );
xor ( n44249 , n44247 , n44248 );
and ( n44250 , n44249 , n44171 );
or ( n44251 , n44246 , n44250 );
not ( n44252 , n44251 );
buf ( n44253 , n44252 );
buf ( n44254 , n44253 );
not ( n44255 , n44254 );
or ( n44256 , n44239 , n44255 );
not ( n44257 , n44171 );
not ( n44258 , n35592 );
and ( n44259 , n44258 , n44087 );
xor ( n44260 , n44088 , n44144 );
and ( n44261 , n44260 , n35592 );
or ( n44262 , n44259 , n44261 );
and ( n44263 , n44257 , n44262 );
not ( n44264 , n44262 );
and ( n44265 , n44247 , n44248 );
xor ( n44266 , n44264 , n44265 );
and ( n44267 , n44266 , n44171 );
or ( n44268 , n44263 , n44267 );
not ( n44269 , n44268 );
buf ( n44270 , n44269 );
buf ( n44271 , n44270 );
not ( n44272 , n44271 );
or ( n44273 , n44256 , n44272 );
not ( n44274 , n44171 );
not ( n44275 , n35592 );
and ( n44276 , n44275 , n44077 );
xor ( n44277 , n44078 , n44145 );
and ( n44278 , n44277 , n35592 );
or ( n44279 , n44276 , n44278 );
and ( n44280 , n44274 , n44279 );
not ( n44281 , n44279 );
and ( n44282 , n44264 , n44265 );
xor ( n44283 , n44281 , n44282 );
and ( n44284 , n44283 , n44171 );
or ( n44285 , n44280 , n44284 );
not ( n44286 , n44285 );
buf ( n44287 , n44286 );
buf ( n44288 , n44287 );
not ( n44289 , n44288 );
or ( n44290 , n44273 , n44289 );
not ( n44291 , n44171 );
not ( n44292 , n35592 );
and ( n44293 , n44292 , n44067 );
xor ( n44294 , n44068 , n44146 );
and ( n44295 , n44294 , n35592 );
or ( n44296 , n44293 , n44295 );
and ( n44297 , n44291 , n44296 );
not ( n44298 , n44296 );
and ( n44299 , n44281 , n44282 );
xor ( n44300 , n44298 , n44299 );
and ( n44301 , n44300 , n44171 );
or ( n44302 , n44297 , n44301 );
not ( n44303 , n44302 );
buf ( n44304 , n44303 );
buf ( n44305 , n44304 );
not ( n44306 , n44305 );
or ( n44307 , n44290 , n44306 );
not ( n44308 , n44171 );
not ( n44309 , n35592 );
and ( n44310 , n44309 , n44057 );
xor ( n44311 , n44058 , n44147 );
and ( n44312 , n44311 , n35592 );
or ( n44313 , n44310 , n44312 );
and ( n44314 , n44308 , n44313 );
not ( n44315 , n44313 );
and ( n44316 , n44298 , n44299 );
xor ( n44317 , n44315 , n44316 );
and ( n44318 , n44317 , n44171 );
or ( n44319 , n44314 , n44318 );
not ( n44320 , n44319 );
buf ( n44321 , n44320 );
buf ( n44322 , n44321 );
not ( n44323 , n44322 );
or ( n44324 , n44307 , n44323 );
not ( n44325 , n44171 );
not ( n44326 , n35592 );
and ( n44327 , n44326 , n44047 );
xor ( n44328 , n44048 , n44148 );
and ( n44329 , n44328 , n35592 );
or ( n44330 , n44327 , n44329 );
and ( n44331 , n44325 , n44330 );
not ( n44332 , n44330 );
and ( n44333 , n44315 , n44316 );
xor ( n44334 , n44332 , n44333 );
and ( n44335 , n44334 , n44171 );
or ( n44336 , n44331 , n44335 );
not ( n44337 , n44336 );
buf ( n44338 , n44337 );
buf ( n44339 , n44338 );
not ( n44340 , n44339 );
or ( n44341 , n44324 , n44340 );
not ( n44342 , n44171 );
not ( n44343 , n35592 );
and ( n44344 , n44343 , n44037 );
xor ( n44345 , n44038 , n44149 );
and ( n44346 , n44345 , n35592 );
or ( n44347 , n44344 , n44346 );
and ( n44348 , n44342 , n44347 );
not ( n44349 , n44347 );
and ( n44350 , n44332 , n44333 );
xor ( n44351 , n44349 , n44350 );
and ( n44352 , n44351 , n44171 );
or ( n44353 , n44348 , n44352 );
not ( n44354 , n44353 );
buf ( n44355 , n44354 );
buf ( n44356 , n44355 );
not ( n44357 , n44356 );
or ( n44358 , n44341 , n44357 );
not ( n44359 , n44171 );
not ( n44360 , n35592 );
and ( n44361 , n44360 , n44027 );
xor ( n44362 , n44028 , n44150 );
and ( n44363 , n44362 , n35592 );
or ( n44364 , n44361 , n44363 );
and ( n44365 , n44359 , n44364 );
not ( n44366 , n44364 );
and ( n44367 , n44349 , n44350 );
xor ( n44368 , n44366 , n44367 );
and ( n44369 , n44368 , n44171 );
or ( n44370 , n44365 , n44369 );
not ( n44371 , n44370 );
buf ( n44372 , n44371 );
buf ( n44373 , n44372 );
not ( n44374 , n44373 );
or ( n44375 , n44358 , n44374 );
not ( n44376 , n44171 );
not ( n44377 , n35592 );
and ( n44378 , n44377 , n44017 );
xor ( n44379 , n44018 , n44151 );
and ( n44380 , n44379 , n35592 );
or ( n44381 , n44378 , n44380 );
and ( n44382 , n44376 , n44381 );
not ( n44383 , n44381 );
and ( n44384 , n44366 , n44367 );
xor ( n44385 , n44383 , n44384 );
and ( n44386 , n44385 , n44171 );
or ( n44387 , n44382 , n44386 );
not ( n44388 , n44387 );
buf ( n44389 , n44388 );
buf ( n44390 , n44389 );
not ( n44391 , n44390 );
or ( n44392 , n44375 , n44391 );
not ( n44393 , n44171 );
not ( n44394 , n35592 );
and ( n44395 , n44394 , n44007 );
xor ( n44396 , n44008 , n44152 );
and ( n44397 , n44396 , n35592 );
or ( n44398 , n44395 , n44397 );
and ( n44399 , n44393 , n44398 );
not ( n44400 , n44398 );
and ( n44401 , n44383 , n44384 );
xor ( n44402 , n44400 , n44401 );
and ( n44403 , n44402 , n44171 );
or ( n44404 , n44399 , n44403 );
not ( n44405 , n44404 );
buf ( n44406 , n44405 );
buf ( n44407 , n44406 );
not ( n44408 , n44407 );
or ( n44409 , n44392 , n44408 );
not ( n44410 , n44171 );
not ( n44411 , n35592 );
and ( n44412 , n44411 , n43997 );
xor ( n44413 , n43998 , n44153 );
and ( n44414 , n44413 , n35592 );
or ( n44415 , n44412 , n44414 );
and ( n44416 , n44410 , n44415 );
not ( n44417 , n44415 );
and ( n44418 , n44400 , n44401 );
xor ( n44419 , n44417 , n44418 );
and ( n44420 , n44419 , n44171 );
or ( n44421 , n44416 , n44420 );
not ( n44422 , n44421 );
buf ( n44423 , n44422 );
buf ( n44424 , n44423 );
not ( n44425 , n44424 );
or ( n44426 , n44409 , n44425 );
not ( n44427 , n44171 );
not ( n44428 , n35592 );
and ( n44429 , n44428 , n43987 );
xor ( n44430 , n43988 , n44154 );
and ( n44431 , n44430 , n35592 );
or ( n44432 , n44429 , n44431 );
and ( n44433 , n44427 , n44432 );
not ( n44434 , n44432 );
and ( n44435 , n44417 , n44418 );
xor ( n44436 , n44434 , n44435 );
and ( n44437 , n44436 , n44171 );
or ( n44438 , n44433 , n44437 );
not ( n44439 , n44438 );
buf ( n44440 , n44439 );
buf ( n44441 , n44440 );
not ( n44442 , n44441 );
or ( n44443 , n44426 , n44442 );
not ( n44444 , n44171 );
not ( n44445 , n35592 );
and ( n44446 , n44445 , n43977 );
xor ( n44447 , n43978 , n44155 );
and ( n44448 , n44447 , n35592 );
or ( n44449 , n44446 , n44448 );
and ( n44450 , n44444 , n44449 );
not ( n44451 , n44449 );
and ( n44452 , n44434 , n44435 );
xor ( n44453 , n44451 , n44452 );
and ( n44454 , n44453 , n44171 );
or ( n44455 , n44450 , n44454 );
not ( n44456 , n44455 );
buf ( n44457 , n44456 );
buf ( n44458 , n44457 );
not ( n44459 , n44458 );
or ( n44460 , n44443 , n44459 );
not ( n44461 , n44171 );
not ( n44462 , n35592 );
and ( n44463 , n44462 , n43967 );
xor ( n44464 , n43968 , n44156 );
and ( n44465 , n44464 , n35592 );
or ( n44466 , n44463 , n44465 );
and ( n44467 , n44461 , n44466 );
not ( n44468 , n44466 );
and ( n44469 , n44451 , n44452 );
xor ( n44470 , n44468 , n44469 );
and ( n44471 , n44470 , n44171 );
or ( n44472 , n44467 , n44471 );
not ( n44473 , n44472 );
buf ( n44474 , n44473 );
buf ( n44475 , n44474 );
not ( n44476 , n44475 );
or ( n44477 , n44460 , n44476 );
not ( n44478 , n44171 );
not ( n44479 , n35592 );
and ( n44480 , n44479 , n43957 );
xor ( n44481 , n43958 , n44157 );
and ( n44482 , n44481 , n35592 );
or ( n44483 , n44480 , n44482 );
and ( n44484 , n44478 , n44483 );
not ( n44485 , n44483 );
and ( n44486 , n44468 , n44469 );
xor ( n44487 , n44485 , n44486 );
and ( n44488 , n44487 , n44171 );
or ( n44489 , n44484 , n44488 );
not ( n44490 , n44489 );
buf ( n44491 , n44490 );
buf ( n44492 , n44491 );
not ( n44493 , n44492 );
or ( n44494 , n44477 , n44493 );
not ( n44495 , n44171 );
not ( n44496 , n35592 );
and ( n44497 , n44496 , n43947 );
xor ( n44498 , n43948 , n44158 );
and ( n44499 , n44498 , n35592 );
or ( n44500 , n44497 , n44499 );
and ( n44501 , n44495 , n44500 );
not ( n44502 , n44500 );
and ( n44503 , n44485 , n44486 );
xor ( n44504 , n44502 , n44503 );
and ( n44505 , n44504 , n44171 );
or ( n44506 , n44501 , n44505 );
not ( n44507 , n44506 );
buf ( n44508 , n44507 );
buf ( n44509 , n44508 );
not ( n44510 , n44509 );
or ( n44511 , n44494 , n44510 );
not ( n44512 , n44171 );
not ( n44513 , n35592 );
and ( n44514 , n44513 , n43937 );
xor ( n44515 , n43938 , n44159 );
and ( n44516 , n44515 , n35592 );
or ( n44517 , n44514 , n44516 );
and ( n44518 , n44512 , n44517 );
not ( n44519 , n44517 );
and ( n44520 , n44502 , n44503 );
xor ( n44521 , n44519 , n44520 );
and ( n44522 , n44521 , n44171 );
or ( n44523 , n44518 , n44522 );
not ( n44524 , n44523 );
buf ( n44525 , n44524 );
buf ( n44526 , n44525 );
not ( n44527 , n44526 );
or ( n44528 , n44511 , n44527 );
not ( n44529 , n44171 );
not ( n44530 , n35592 );
and ( n44531 , n44530 , n43927 );
xor ( n44532 , n43928 , n44160 );
and ( n44533 , n44532 , n35592 );
or ( n44534 , n44531 , n44533 );
and ( n44535 , n44529 , n44534 );
not ( n44536 , n44534 );
and ( n44537 , n44519 , n44520 );
xor ( n44538 , n44536 , n44537 );
and ( n44539 , n44538 , n44171 );
or ( n44540 , n44535 , n44539 );
not ( n44541 , n44540 );
buf ( n44542 , n44541 );
buf ( n44543 , n44542 );
not ( n44544 , n44543 );
or ( n44545 , n44528 , n44544 );
not ( n44546 , n44171 );
not ( n44547 , n35592 );
and ( n44548 , n44547 , n43917 );
xor ( n44549 , n43918 , n44161 );
and ( n44550 , n44549 , n35592 );
or ( n44551 , n44548 , n44550 );
and ( n44552 , n44546 , n44551 );
not ( n44553 , n44551 );
and ( n44554 , n44536 , n44537 );
xor ( n44555 , n44553 , n44554 );
and ( n44556 , n44555 , n44171 );
or ( n44557 , n44552 , n44556 );
not ( n44558 , n44557 );
buf ( n44559 , n44558 );
buf ( n44560 , n44559 );
not ( n44561 , n44560 );
or ( n44562 , n44545 , n44561 );
not ( n44563 , n44171 );
not ( n44564 , n35592 );
and ( n44565 , n44564 , n43907 );
xor ( n44566 , n43908 , n44162 );
and ( n44567 , n44566 , n35592 );
or ( n44568 , n44565 , n44567 );
and ( n44569 , n44563 , n44568 );
not ( n44570 , n44568 );
and ( n44571 , n44553 , n44554 );
xor ( n44572 , n44570 , n44571 );
and ( n44573 , n44572 , n44171 );
or ( n44574 , n44569 , n44573 );
not ( n44575 , n44574 );
buf ( n44576 , n44575 );
buf ( n44577 , n44576 );
not ( n44578 , n44577 );
or ( n44579 , n44562 , n44578 );
not ( n44580 , n44171 );
not ( n44581 , n35592 );
and ( n44582 , n44581 , n43897 );
xor ( n44583 , n43898 , n44163 );
and ( n44584 , n44583 , n35592 );
or ( n44585 , n44582 , n44584 );
and ( n44586 , n44580 , n44585 );
not ( n44587 , n44585 );
and ( n44588 , n44570 , n44571 );
xor ( n44589 , n44587 , n44588 );
and ( n44590 , n44589 , n44171 );
or ( n44591 , n44586 , n44590 );
not ( n44592 , n44591 );
buf ( n44593 , n44592 );
buf ( n44594 , n44593 );
not ( n44595 , n44594 );
or ( n44596 , n44579 , n44595 );
not ( n44597 , n44171 );
not ( n44598 , n35592 );
and ( n44599 , n44598 , n43887 );
xor ( n44600 , n43888 , n44164 );
and ( n44601 , n44600 , n35592 );
or ( n44602 , n44599 , n44601 );
and ( n44603 , n44597 , n44602 );
not ( n44604 , n44602 );
and ( n44605 , n44587 , n44588 );
xor ( n44606 , n44604 , n44605 );
and ( n44607 , n44606 , n44171 );
or ( n44608 , n44603 , n44607 );
not ( n44609 , n44608 );
buf ( n44610 , n44609 );
buf ( n44611 , n44610 );
not ( n44612 , n44611 );
or ( n44613 , n44596 , n44612 );
not ( n44614 , n44171 );
not ( n44615 , n35592 );
and ( n44616 , n44615 , n43877 );
xor ( n44617 , n43878 , n44165 );
and ( n44618 , n44617 , n35592 );
or ( n44619 , n44616 , n44618 );
and ( n44620 , n44614 , n44619 );
not ( n44621 , n44619 );
and ( n44622 , n44604 , n44605 );
xor ( n44623 , n44621 , n44622 );
and ( n44624 , n44623 , n44171 );
or ( n44625 , n44620 , n44624 );
not ( n44626 , n44625 );
buf ( n44627 , n44626 );
buf ( n44628 , n44627 );
not ( n44629 , n44628 );
or ( n44630 , n44613 , n44629 );
not ( n44631 , n44171 );
not ( n44632 , n35592 );
and ( n44633 , n44632 , n43867 );
xor ( n44634 , n43868 , n44166 );
and ( n44635 , n44634 , n35592 );
or ( n44636 , n44633 , n44635 );
and ( n44637 , n44631 , n44636 );
not ( n44638 , n44636 );
and ( n44639 , n44621 , n44622 );
xor ( n44640 , n44638 , n44639 );
and ( n44641 , n44640 , n44171 );
or ( n44642 , n44637 , n44641 );
not ( n44643 , n44642 );
buf ( n44644 , n44643 );
buf ( n44645 , n44644 );
not ( n44646 , n44645 );
or ( n44647 , n44630 , n44646 );
xor ( n44648 , n43858 , n44167 );
and ( n44649 , n44648 , n35592 );
buf ( n44650 , n44649 );
not ( n44651 , n44650 );
and ( n44652 , n44638 , n44639 );
xor ( n44653 , n44651 , n44652 );
and ( n44654 , n44653 , n44171 );
buf ( n44655 , n44654 );
not ( n44656 , n44655 );
buf ( n44657 , n44656 );
buf ( n44658 , n44657 );
not ( n44659 , n44658 );
or ( n44660 , n44647 , n44659 );
buf ( n44661 , n44660 );
buf ( n44662 , n44661 );
and ( n44663 , n44662 , n44171 );
not ( n44664 , n44663 );
and ( n44665 , n44664 , n44272 );
xor ( n44666 , n44272 , n44171 );
xor ( n44667 , n44255 , n44171 );
xor ( n44668 , n44238 , n44171 );
xor ( n44669 , n44221 , n44171 );
xor ( n44670 , n44204 , n44171 );
xor ( n44671 , n44187 , n44171 );
xor ( n44672 , n43793 , n44171 );
and ( n44673 , n44672 , n44171 );
and ( n44674 , n44671 , n44673 );
and ( n44675 , n44670 , n44674 );
and ( n44676 , n44669 , n44675 );
and ( n44677 , n44668 , n44676 );
and ( n44678 , n44667 , n44677 );
xor ( n44679 , n44666 , n44678 );
and ( n44680 , n44679 , n44663 );
or ( n44681 , n44665 , n44680 );
nor ( n44682 , n32956 , n32958 , n32959 );
and ( n44683 , n44681 , n44682 );
buf ( n44684 , RI15b45348_226);
nor ( n44685 , n32961 , n32957 , n32959 );
nor ( n44686 , n32956 , n32957 , n32959 );
or ( n44687 , n44685 , n44686 );
nor ( n44688 , n32961 , n32958 , n32959 );
or ( n44689 , n44687 , n44688 );
and ( n44690 , n32961 , n32958 , n32959 );
or ( n44691 , n44689 , n44690 );
and ( n44692 , n32956 , n32958 , n32959 );
or ( n44693 , n44691 , n44692 );
and ( n44694 , n32956 , n32957 , n32959 );
or ( n44695 , n44693 , n44694 );
and ( n44696 , n44684 , n44695 );
or ( n44697 , n43775 , n44683 , n44696 );
buf ( n44698 , n44697 );
buf ( n44699 , n44698 );
buf ( n44700 , n31655 );
buf ( n44701 , n30987 );
buf ( n44702 , RI15b4c080_459);
and ( n44703 , n31447 , n31451 );
not ( n44704 , n44703 );
and ( n44705 , n31077 , n44704 );
and ( n44706 , n44702 , n44705 );
and ( n44707 , n44706 , n31373 );
and ( n44708 , n31402 , n31450 );
and ( n44709 , n44702 , n44708 );
and ( n44710 , n44709 , n31408 );
and ( n44711 , n31437 , n44704 );
and ( n44712 , n44702 , n44711 );
and ( n44713 , n44712 , n31468 );
and ( n44714 , n31497 , n31450 );
and ( n44715 , n44702 , n44714 );
and ( n44716 , n44715 , n31521 );
and ( n44717 , n33419 , n31529 );
and ( n44718 , n33734 , n31527 );
or ( n44719 , n44707 , n44710 , n44713 , n44716 , n44717 , n44718 , C0 );
and ( n44720 , n44719 , n31557 );
and ( n44721 , n44702 , n40154 );
or ( n44722 , C0 , n44720 , n44721 );
buf ( n44723 , n44722 );
buf ( n44724 , n44723 );
buf ( n44725 , n30987 );
buf ( n44726 , n31655 );
not ( n44727 , n31728 );
and ( n44728 , n44727 , n32459 );
xor ( n44729 , n31825 , n31858 );
xor ( n44730 , n44729 , n32084 );
and ( n44731 , n44730 , n31728 );
or ( n44732 , n44728 , n44731 );
and ( n44733 , n44732 , n32253 );
not ( n44734 , n32283 );
and ( n44735 , n44734 , n32459 );
not ( n44736 , n31823 );
xor ( n44737 , n32296 , n31858 );
xor ( n44738 , n44737 , n32323 );
and ( n44739 , n44736 , n44738 );
xor ( n44740 , n32344 , n32346 );
xor ( n44741 , n44740 , n32386 );
and ( n44742 , n44741 , n31823 );
or ( n44743 , n44739 , n44742 );
and ( n44744 , n44743 , n32283 );
or ( n44745 , n44735 , n44744 );
and ( n44746 , n44745 , n32398 );
and ( n44747 , n32459 , n32436 );
or ( n44748 , n44733 , n44746 , n44747 );
and ( n44749 , n44748 , n32456 );
xor ( n44750 , n32459 , n32468 );
and ( n44751 , n44750 , n32473 );
not ( n44752 , n32475 );
and ( n44753 , n44752 , n44750 );
xor ( n44754 , n32459 , n32480 );
and ( n44755 , n44754 , n32475 );
or ( n44756 , n44753 , n44755 );
and ( n44757 , n44756 , n32486 );
and ( n44758 , n37577 , n32489 );
and ( n44759 , n32459 , n32501 );
or ( n44760 , C0 , n44749 , n44751 , n44757 , n44758 , n44759 );
buf ( n44761 , n44760 );
buf ( n44762 , n44761 );
buf ( n44763 , RI15b55680_779);
buf ( n44764 , RI15b55608_778);
buf ( n44765 , RI15b55590_777);
buf ( n44766 , RI15b55518_776);
buf ( n44767 , RI15b554a0_775);
buf ( n44768 , RI15b55428_774);
buf ( n44769 , RI15b553b0_773);
buf ( n44770 , RI15b55338_772);
buf ( n44771 , RI15b552c0_771);
buf ( n44772 , RI15b55248_770);
buf ( n44773 , RI15b551d0_769);
buf ( n44774 , RI15b55158_768);
buf ( n44775 , RI15b550e0_767);
buf ( n44776 , RI15b55068_766);
and ( n44777 , n41613 , n41606 );
and ( n44778 , n41626 , n44777 );
and ( n44779 , n41639 , n44778 );
and ( n44780 , n41652 , n44779 );
and ( n44781 , n41665 , n44780 );
and ( n44782 , n41678 , n44781 );
and ( n44783 , n41691 , n44782 );
and ( n44784 , n41704 , n44783 );
and ( n44785 , n41717 , n44784 );
and ( n44786 , n41730 , n44785 );
and ( n44787 , n41743 , n44786 );
and ( n44788 , n41756 , n44787 );
and ( n44789 , n41769 , n44788 );
and ( n44790 , n41782 , n44789 );
and ( n44791 , n41795 , n44790 );
and ( n44792 , n44776 , n44791 );
and ( n44793 , n44775 , n44792 );
and ( n44794 , n44774 , n44793 );
and ( n44795 , n44773 , n44794 );
and ( n44796 , n44772 , n44795 );
and ( n44797 , n44771 , n44796 );
and ( n44798 , n44770 , n44797 );
and ( n44799 , n44769 , n44798 );
and ( n44800 , n44768 , n44799 );
and ( n44801 , n44767 , n44800 );
and ( n44802 , n44766 , n44801 );
and ( n44803 , n44765 , n44802 );
and ( n44804 , n44764 , n44803 );
xor ( n44805 , n44763 , n44804 );
and ( n44806 , n44805 , n31548 );
and ( n44807 , n31402 , n31451 );
not ( n44808 , n44807 );
and ( n44809 , n44808 , n44763 );
not ( n44810 , n41869 );
and ( n44811 , n44810 , n34419 );
and ( n44812 , n40562 , n41869 );
or ( n44813 , n44811 , n44812 );
and ( n44814 , n44813 , n44807 );
or ( n44815 , n44809 , n44814 );
and ( n44816 , n44815 , n31408 );
and ( n44817 , n31497 , n31451 );
not ( n44818 , n44817 );
and ( n44819 , n44818 , n44763 );
buf ( n44820 , n41873 );
not ( n44821 , n44820 );
buf ( n44822 , n44821 );
not ( n44823 , n44822 );
not ( n44824 , n41881 );
and ( n44825 , n44824 , n41886 );
not ( n44826 , n41886 );
not ( n44827 , n41873 );
xor ( n44828 , n44826 , n44827 );
and ( n44829 , n44828 , n41881 );
or ( n44830 , n44825 , n44829 );
not ( n44831 , n44830 );
buf ( n44832 , n44831 );
buf ( n44833 , n44832 );
not ( n44834 , n44833 );
or ( n44835 , n44823 , n44834 );
not ( n44836 , n41881 );
and ( n44837 , n44836 , n41902 );
not ( n44838 , n41902 );
and ( n44839 , n44826 , n44827 );
xor ( n44840 , n44838 , n44839 );
and ( n44841 , n44840 , n41881 );
or ( n44842 , n44837 , n44841 );
not ( n44843 , n44842 );
buf ( n44844 , n44843 );
buf ( n44845 , n44844 );
not ( n44846 , n44845 );
or ( n44847 , n44835 , n44846 );
not ( n44848 , n41881 );
and ( n44849 , n44848 , n41918 );
not ( n44850 , n41918 );
and ( n44851 , n44838 , n44839 );
xor ( n44852 , n44850 , n44851 );
and ( n44853 , n44852 , n41881 );
or ( n44854 , n44849 , n44853 );
not ( n44855 , n44854 );
buf ( n44856 , n44855 );
buf ( n44857 , n44856 );
not ( n44858 , n44857 );
or ( n44859 , n44847 , n44858 );
not ( n44860 , n41881 );
and ( n44861 , n44860 , n41934 );
not ( n44862 , n41934 );
and ( n44863 , n44850 , n44851 );
xor ( n44864 , n44862 , n44863 );
and ( n44865 , n44864 , n41881 );
or ( n44866 , n44861 , n44865 );
not ( n44867 , n44866 );
buf ( n44868 , n44867 );
buf ( n44869 , n44868 );
not ( n44870 , n44869 );
or ( n44871 , n44859 , n44870 );
not ( n44872 , n41881 );
and ( n44873 , n44872 , n41950 );
not ( n44874 , n41950 );
and ( n44875 , n44862 , n44863 );
xor ( n44876 , n44874 , n44875 );
and ( n44877 , n44876 , n41881 );
or ( n44878 , n44873 , n44877 );
not ( n44879 , n44878 );
buf ( n44880 , n44879 );
buf ( n44881 , n44880 );
not ( n44882 , n44881 );
or ( n44883 , n44871 , n44882 );
not ( n44884 , n41881 );
and ( n44885 , n44884 , n41966 );
not ( n44886 , n41966 );
and ( n44887 , n44874 , n44875 );
xor ( n44888 , n44886 , n44887 );
and ( n44889 , n44888 , n41881 );
or ( n44890 , n44885 , n44889 );
not ( n44891 , n44890 );
buf ( n44892 , n44891 );
buf ( n44893 , n44892 );
not ( n44894 , n44893 );
or ( n44895 , n44883 , n44894 );
not ( n44896 , n41881 );
and ( n44897 , n44896 , n41982 );
not ( n44898 , n41982 );
and ( n44899 , n44886 , n44887 );
xor ( n44900 , n44898 , n44899 );
and ( n44901 , n44900 , n41881 );
or ( n44902 , n44897 , n44901 );
not ( n44903 , n44902 );
buf ( n44904 , n44903 );
buf ( n44905 , n44904 );
not ( n44906 , n44905 );
or ( n44907 , n44895 , n44906 );
not ( n44908 , n41881 );
and ( n44909 , n44908 , n41998 );
not ( n44910 , n41998 );
and ( n44911 , n44898 , n44899 );
xor ( n44912 , n44910 , n44911 );
and ( n44913 , n44912 , n41881 );
or ( n44914 , n44909 , n44913 );
not ( n44915 , n44914 );
buf ( n44916 , n44915 );
buf ( n44917 , n44916 );
not ( n44918 , n44917 );
or ( n44919 , n44907 , n44918 );
not ( n44920 , n41881 );
and ( n44921 , n44920 , n42014 );
not ( n44922 , n42014 );
and ( n44923 , n44910 , n44911 );
xor ( n44924 , n44922 , n44923 );
and ( n44925 , n44924 , n41881 );
or ( n44926 , n44921 , n44925 );
not ( n44927 , n44926 );
buf ( n44928 , n44927 );
buf ( n44929 , n44928 );
not ( n44930 , n44929 );
or ( n44931 , n44919 , n44930 );
not ( n44932 , n41881 );
and ( n44933 , n44932 , n42030 );
not ( n44934 , n42030 );
and ( n44935 , n44922 , n44923 );
xor ( n44936 , n44934 , n44935 );
and ( n44937 , n44936 , n41881 );
or ( n44938 , n44933 , n44937 );
not ( n44939 , n44938 );
buf ( n44940 , n44939 );
buf ( n44941 , n44940 );
not ( n44942 , n44941 );
or ( n44943 , n44931 , n44942 );
not ( n44944 , n41881 );
and ( n44945 , n44944 , n42046 );
not ( n44946 , n42046 );
and ( n44947 , n44934 , n44935 );
xor ( n44948 , n44946 , n44947 );
and ( n44949 , n44948 , n41881 );
or ( n44950 , n44945 , n44949 );
not ( n44951 , n44950 );
buf ( n44952 , n44951 );
buf ( n44953 , n44952 );
not ( n44954 , n44953 );
or ( n44955 , n44943 , n44954 );
not ( n44956 , n41881 );
and ( n44957 , n44956 , n42062 );
not ( n44958 , n42062 );
and ( n44959 , n44946 , n44947 );
xor ( n44960 , n44958 , n44959 );
and ( n44961 , n44960 , n41881 );
or ( n44962 , n44957 , n44961 );
not ( n44963 , n44962 );
buf ( n44964 , n44963 );
buf ( n44965 , n44964 );
not ( n44966 , n44965 );
or ( n44967 , n44955 , n44966 );
not ( n44968 , n41881 );
and ( n44969 , n44968 , n42078 );
not ( n44970 , n42078 );
and ( n44971 , n44958 , n44959 );
xor ( n44972 , n44970 , n44971 );
and ( n44973 , n44972 , n41881 );
or ( n44974 , n44969 , n44973 );
not ( n44975 , n44974 );
buf ( n44976 , n44975 );
buf ( n44977 , n44976 );
not ( n44978 , n44977 );
or ( n44979 , n44967 , n44978 );
not ( n44980 , n41881 );
and ( n44981 , n44980 , n42094 );
not ( n44982 , n42094 );
and ( n44983 , n44970 , n44971 );
xor ( n44984 , n44982 , n44983 );
and ( n44985 , n44984 , n41881 );
or ( n44986 , n44981 , n44985 );
not ( n44987 , n44986 );
buf ( n44988 , n44987 );
buf ( n44989 , n44988 );
not ( n44990 , n44989 );
or ( n44991 , n44979 , n44990 );
buf ( n44992 , n44991 );
buf ( n44993 , n44992 );
and ( n44994 , n44993 , n41881 );
not ( n44995 , n44994 );
and ( n44996 , n44995 , n44978 );
xor ( n44997 , n44978 , n41881 );
xor ( n44998 , n44966 , n41881 );
xor ( n44999 , n44954 , n41881 );
xor ( n45000 , n44942 , n41881 );
xor ( n45001 , n44930 , n41881 );
xor ( n45002 , n44918 , n41881 );
xor ( n45003 , n44906 , n41881 );
xor ( n45004 , n44894 , n41881 );
xor ( n45005 , n44882 , n41881 );
xor ( n45006 , n44870 , n41881 );
xor ( n45007 , n44858 , n41881 );
xor ( n45008 , n44846 , n41881 );
xor ( n45009 , n44834 , n41881 );
xor ( n45010 , n44823 , n41881 );
and ( n45011 , n45010 , n41881 );
and ( n45012 , n45009 , n45011 );
and ( n45013 , n45008 , n45012 );
and ( n45014 , n45007 , n45013 );
and ( n45015 , n45006 , n45014 );
and ( n45016 , n45005 , n45015 );
and ( n45017 , n45004 , n45016 );
and ( n45018 , n45003 , n45017 );
and ( n45019 , n45002 , n45018 );
and ( n45020 , n45001 , n45019 );
and ( n45021 , n45000 , n45020 );
and ( n45022 , n44999 , n45021 );
and ( n45023 , n44998 , n45022 );
xor ( n45024 , n44997 , n45023 );
and ( n45025 , n45024 , n44994 );
or ( n45026 , n44996 , n45025 );
and ( n45027 , n45026 , n44817 );
or ( n45028 , n44819 , n45027 );
and ( n45029 , n45028 , n31521 );
not ( n45030 , n31041 );
buf ( n45031 , n31041 );
buf ( n45032 , n31041 );
buf ( n45033 , n31041 );
buf ( n45034 , n31041 );
buf ( n45035 , n31041 );
buf ( n45036 , n31041 );
buf ( n45037 , n31041 );
buf ( n45038 , n31041 );
buf ( n45039 , n31041 );
buf ( n45040 , n31041 );
buf ( n45041 , n31041 );
buf ( n45042 , n31041 );
buf ( n45043 , n31041 );
buf ( n45044 , n31041 );
buf ( n45045 , n31041 );
buf ( n45046 , n31041 );
buf ( n45047 , n31041 );
buf ( n45048 , n31041 );
buf ( n45049 , n31041 );
buf ( n45050 , n31041 );
buf ( n45051 , n31041 );
buf ( n45052 , n31041 );
buf ( n45053 , n31041 );
buf ( n45054 , n31041 );
buf ( n45055 , n31041 );
or ( n45056 , n31075 , n33415 );
and ( n45057 , n31044 , n45056 );
or ( n45058 , n31046 , n31048 , n31041 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45057 );
and ( n45059 , n45030 , n45058 );
not ( n45060 , n45059 );
and ( n45061 , n45060 , n44763 );
and ( n45062 , n31307 , n40003 );
and ( n45063 , n31309 , n40005 );
and ( n45064 , n31311 , n40007 );
and ( n45065 , n31313 , n40009 );
and ( n45066 , n31315 , n40011 );
and ( n45067 , n31317 , n40013 );
and ( n45068 , n31319 , n40015 );
and ( n45069 , n31321 , n40017 );
and ( n45070 , n31323 , n40019 );
and ( n45071 , n31325 , n40021 );
and ( n45072 , n31327 , n40023 );
and ( n45073 , n31329 , n40025 );
and ( n45074 , n31331 , n40027 );
and ( n45075 , n31333 , n40029 );
and ( n45076 , n31335 , n40031 );
and ( n45077 , n31337 , n40033 );
or ( n45078 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 );
and ( n45079 , n31274 , n40003 );
and ( n45080 , n31276 , n40005 );
and ( n45081 , n31278 , n40007 );
and ( n45082 , n31280 , n40009 );
and ( n45083 , n31282 , n40011 );
and ( n45084 , n31284 , n40013 );
and ( n45085 , n31286 , n40015 );
and ( n45086 , n31288 , n40017 );
and ( n45087 , n31290 , n40019 );
and ( n45088 , n31292 , n40021 );
and ( n45089 , n31294 , n40023 );
and ( n45090 , n31296 , n40025 );
and ( n45091 , n31298 , n40027 );
and ( n45092 , n31300 , n40029 );
and ( n45093 , n31302 , n40031 );
and ( n45094 , n31304 , n40033 );
or ( n45095 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 );
and ( n45096 , n31240 , n40003 );
and ( n45097 , n31242 , n40005 );
and ( n45098 , n31244 , n40007 );
and ( n45099 , n31246 , n40009 );
and ( n45100 , n31248 , n40011 );
and ( n45101 , n31250 , n40013 );
and ( n45102 , n31252 , n40015 );
and ( n45103 , n31254 , n40017 );
and ( n45104 , n31256 , n40019 );
and ( n45105 , n31258 , n40021 );
and ( n45106 , n31260 , n40023 );
and ( n45107 , n31262 , n40025 );
and ( n45108 , n31264 , n40027 );
and ( n45109 , n31266 , n40029 );
and ( n45110 , n31268 , n40031 );
and ( n45111 , n31270 , n40033 );
or ( n45112 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 );
and ( n45113 , n31206 , n40003 );
and ( n45114 , n31208 , n40005 );
and ( n45115 , n31210 , n40007 );
and ( n45116 , n31212 , n40009 );
and ( n45117 , n31214 , n40011 );
and ( n45118 , n31216 , n40013 );
and ( n45119 , n31218 , n40015 );
and ( n45120 , n31220 , n40017 );
and ( n45121 , n31222 , n40019 );
and ( n45122 , n31224 , n40021 );
and ( n45123 , n31226 , n40023 );
and ( n45124 , n31228 , n40025 );
and ( n45125 , n31230 , n40027 );
and ( n45126 , n31232 , n40029 );
and ( n45127 , n31234 , n40031 );
and ( n45128 , n31236 , n40033 );
or ( n45129 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 );
and ( n45130 , n40069 , n40127 );
and ( n45131 , n40052 , n45130 );
and ( n45132 , n40035 , n45131 );
and ( n45133 , n45129 , n45132 );
and ( n45134 , n45112 , n45133 );
and ( n45135 , n45095 , n45134 );
xor ( n45136 , n45078 , n45135 );
and ( n45137 , n45136 , n45059 );
or ( n45138 , n45061 , n45137 );
and ( n45139 , n45138 , n31536 );
or ( n45140 , n31535 , n31538 );
or ( n45141 , n45140 , n31468 );
or ( n45142 , n45141 , n31373 );
or ( n45143 , n45142 , n31540 );
or ( n45144 , n45143 , n31542 );
or ( n45145 , n45144 , n31544 );
or ( n45146 , n45145 , n31546 );
or ( n45147 , n45146 , n31550 );
or ( n45148 , n45147 , n31552 );
and ( n45149 , n44763 , n45148 );
or ( n45150 , n44806 , n44816 , n45029 , n45139 , n45149 );
and ( n45151 , n45150 , n31557 );
and ( n45152 , n44763 , n40154 );
or ( n45153 , C0 , n45151 , n45152 );
buf ( n45154 , n45153 );
buf ( n45155 , n45154 );
buf ( n45156 , n31655 );
buf ( n45157 , n30987 );
not ( n45158 , n40163 );
and ( n45159 , n45158 , n31953 );
not ( n45160 , n31665 );
nor ( n45161 , n31673 , n31669 , n45160 , n31661 , n31657 );
not ( n45162 , n45161 );
and ( n45163 , n45162 , n31953 );
and ( n45164 , n32183 , n45161 );
or ( n45165 , n45163 , n45164 );
and ( n45166 , n45165 , n40163 );
or ( n45167 , n45159 , n45166 );
and ( n45168 , n45167 , n32498 );
not ( n45169 , n40188 );
nor ( n45170 , n40177 , n40182 , n45169 , n40194 , C0 );
not ( n45171 , n45170 );
not ( n45172 , n45161 );
and ( n45173 , n45172 , n31953 );
not ( n45174 , n40373 );
and ( n45175 , n45174 , n40297 );
xor ( n45176 , n40380 , n40386 );
and ( n45177 , n45176 , n40373 );
or ( n45178 , n45175 , n45177 );
and ( n45179 , n45178 , n45161 );
or ( n45180 , n45173 , n45179 );
and ( n45181 , n45171 , n45180 );
and ( n45182 , n45178 , n45170 );
or ( n45183 , n45181 , n45182 );
and ( n45184 , n45183 , n32473 );
not ( n45185 , n32475 );
not ( n45186 , n45170 );
not ( n45187 , n45161 );
and ( n45188 , n45187 , n31953 );
and ( n45189 , n45178 , n45161 );
or ( n45190 , n45188 , n45189 );
and ( n45191 , n45186 , n45190 );
and ( n45192 , n45178 , n45170 );
or ( n45193 , n45191 , n45192 );
and ( n45194 , n45185 , n45193 );
not ( n45195 , n40435 );
nor ( n45196 , n40417 , n40425 , n45195 , n40445 , C0 );
not ( n45197 , n45196 );
not ( n45198 , n40430 );
nor ( n45199 , n40413 , n40421 , n45198 , n40440 , C0 );
not ( n45200 , n45199 );
and ( n45201 , n45200 , n45193 );
not ( n45202 , n40952 );
and ( n45203 , n45202 , n40880 );
xor ( n45204 , n40959 , n40965 );
and ( n45205 , n45204 , n40952 );
or ( n45206 , n45203 , n45205 );
and ( n45207 , n45206 , n45199 );
or ( n45208 , n45201 , n45207 );
and ( n45209 , n45197 , n45208 );
not ( n45210 , n41247 );
and ( n45211 , n45210 , n41179 );
xor ( n45212 , n41254 , n41260 );
and ( n45213 , n45212 , n41247 );
or ( n45214 , n45211 , n45213 );
and ( n45215 , n45214 , n45196 );
or ( n45216 , n45209 , n45215 );
and ( n45217 , n45216 , n32475 );
or ( n45218 , n45194 , n45217 );
and ( n45219 , n45218 , n32486 );
and ( n45220 , n31953 , n41278 );
or ( n45221 , C0 , n45168 , n45184 , n45219 , n45220 );
buf ( n45222 , n45221 );
buf ( n45223 , n45222 );
buf ( n45224 , n30987 );
not ( n45225 , n40163 );
and ( n45226 , n45225 , n31871 );
and ( n45227 , n42169 , n31669 , n45160 , n31661 , n42170 );
not ( n45228 , n45227 );
and ( n45229 , n45228 , n31871 );
and ( n45230 , n32218 , n45227 );
or ( n45231 , n45229 , n45230 );
and ( n45232 , n45231 , n40163 );
or ( n45233 , n45226 , n45232 );
and ( n45234 , n45233 , n32498 );
and ( n45235 , n42179 , n40182 , n45169 , n40194 , C1 );
not ( n45236 , n45235 );
not ( n45237 , n45227 );
and ( n45238 , n45237 , n31871 );
and ( n45239 , n42255 , n45227 );
or ( n45240 , n45238 , n45239 );
and ( n45241 , n45236 , n45240 );
and ( n45242 , n42255 , n45235 );
or ( n45243 , n45241 , n45242 );
and ( n45244 , n45243 , n32473 );
not ( n45245 , n32475 );
not ( n45246 , n45235 );
not ( n45247 , n45227 );
and ( n45248 , n45247 , n31871 );
and ( n45249 , n42255 , n45227 );
or ( n45250 , n45248 , n45249 );
and ( n45251 , n45246 , n45250 );
and ( n45252 , n42255 , n45235 );
or ( n45253 , n45251 , n45252 );
and ( n45254 , n45245 , n45253 );
and ( n45255 , n42205 , n40425 , n45195 , n40445 , C1 );
not ( n45256 , n45255 );
and ( n45257 , n42208 , n40421 , n45198 , n40440 , C1 );
not ( n45258 , n45257 );
and ( n45259 , n45258 , n45253 );
and ( n45260 , n42283 , n45257 );
or ( n45261 , n45259 , n45260 );
and ( n45262 , n45256 , n45261 );
and ( n45263 , n42291 , n45255 );
or ( n45264 , n45262 , n45263 );
and ( n45265 , n45264 , n32475 );
or ( n45266 , n45254 , n45265 );
and ( n45267 , n45266 , n32486 );
and ( n45268 , n31871 , n41278 );
or ( n45269 , C0 , n45234 , n45244 , n45267 , n45268 );
buf ( n45270 , n45269 );
buf ( n45271 , n45270 );
buf ( n45272 , RI15b52908_682);
and ( n45273 , n45272 , n31645 );
and ( n45274 , n31077 , n31447 );
not ( n45275 , n45274 );
buf ( n45276 , RI15b53f10_729);
and ( n45277 , n45275 , n45276 );
buf ( n45278 , n45277 );
and ( n45279 , n45278 , n31373 );
and ( n45280 , n31437 , n31447 );
not ( n45281 , n45280 );
and ( n45282 , n45281 , n45276 );
not ( n45283 , n41611 );
and ( n45284 , n45283 , n44776 );
not ( n45285 , n44776 );
not ( n45286 , n41795 );
not ( n45287 , n41782 );
not ( n45288 , n41769 );
not ( n45289 , n41756 );
not ( n45290 , n41743 );
not ( n45291 , n41730 );
not ( n45292 , n41717 );
not ( n45293 , n41704 );
not ( n45294 , n41691 );
not ( n45295 , n41678 );
not ( n45296 , n41665 );
not ( n45297 , n41652 );
not ( n45298 , n41639 );
not ( n45299 , n41626 );
not ( n45300 , n41613 );
not ( n45301 , n41606 );
and ( n45302 , n45300 , n45301 );
and ( n45303 , n45299 , n45302 );
and ( n45304 , n45298 , n45303 );
and ( n45305 , n45297 , n45304 );
and ( n45306 , n45296 , n45305 );
and ( n45307 , n45295 , n45306 );
and ( n45308 , n45294 , n45307 );
and ( n45309 , n45293 , n45308 );
and ( n45310 , n45292 , n45309 );
and ( n45311 , n45291 , n45310 );
and ( n45312 , n45290 , n45311 );
and ( n45313 , n45289 , n45312 );
and ( n45314 , n45288 , n45313 );
and ( n45315 , n45287 , n45314 );
and ( n45316 , n45286 , n45315 );
xor ( n45317 , n45285 , n45316 );
and ( n45318 , n45317 , n41611 );
or ( n45319 , n45284 , n45318 );
not ( n45320 , n45319 );
buf ( n45321 , n45320 );
buf ( n45322 , n45321 );
not ( n45323 , n45322 );
buf ( n45324 , n45323 );
buf ( n45325 , n45324 );
not ( n45326 , n45325 );
buf ( n45327 , n45326 );
not ( n45328 , n45327 );
not ( n45329 , n41611 );
buf ( n45330 , RI15b556f8_780);
not ( n45331 , n45330 );
not ( n45332 , n44763 );
not ( n45333 , n44764 );
not ( n45334 , n44765 );
not ( n45335 , n44766 );
not ( n45336 , n44767 );
not ( n45337 , n44768 );
not ( n45338 , n44769 );
not ( n45339 , n44770 );
not ( n45340 , n44771 );
not ( n45341 , n44772 );
not ( n45342 , n44773 );
not ( n45343 , n44774 );
not ( n45344 , n44775 );
and ( n45345 , n45285 , n45316 );
and ( n45346 , n45344 , n45345 );
and ( n45347 , n45343 , n45346 );
and ( n45348 , n45342 , n45347 );
and ( n45349 , n45341 , n45348 );
and ( n45350 , n45340 , n45349 );
and ( n45351 , n45339 , n45350 );
and ( n45352 , n45338 , n45351 );
and ( n45353 , n45337 , n45352 );
and ( n45354 , n45336 , n45353 );
and ( n45355 , n45335 , n45354 );
and ( n45356 , n45334 , n45355 );
and ( n45357 , n45333 , n45356 );
and ( n45358 , n45332 , n45357 );
and ( n45359 , n45331 , n45358 );
xor ( n45360 , n45329 , n45359 );
buf ( n45361 , n41611 );
and ( n45362 , n45360 , n45361 );
buf ( n45363 , n45362 );
not ( n45364 , n45363 );
not ( n45365 , n45364 );
not ( n45366 , n45365 );
not ( n45367 , n41611 );
and ( n45368 , n45367 , n45330 );
xor ( n45369 , n45331 , n45358 );
and ( n45370 , n45369 , n41611 );
or ( n45371 , n45368 , n45370 );
not ( n45372 , n45371 );
buf ( n45373 , n45372 );
buf ( n45374 , n45373 );
not ( n45375 , n45374 );
not ( n45376 , n45375 );
not ( n45377 , n41611 );
and ( n45378 , n45377 , n44763 );
xor ( n45379 , n45332 , n45357 );
and ( n45380 , n45379 , n41611 );
or ( n45381 , n45378 , n45380 );
not ( n45382 , n45381 );
buf ( n45383 , n45382 );
buf ( n45384 , n45383 );
not ( n45385 , n45384 );
not ( n45386 , n45385 );
not ( n45387 , n41611 );
and ( n45388 , n45387 , n44764 );
xor ( n45389 , n45333 , n45356 );
and ( n45390 , n45389 , n41611 );
or ( n45391 , n45388 , n45390 );
not ( n45392 , n45391 );
buf ( n45393 , n45392 );
buf ( n45394 , n45393 );
not ( n45395 , n45394 );
not ( n45396 , n45395 );
not ( n45397 , n41611 );
and ( n45398 , n45397 , n44765 );
xor ( n45399 , n45334 , n45355 );
and ( n45400 , n45399 , n41611 );
or ( n45401 , n45398 , n45400 );
not ( n45402 , n45401 );
buf ( n45403 , n45402 );
buf ( n45404 , n45403 );
not ( n45405 , n45404 );
not ( n45406 , n45405 );
not ( n45407 , n41611 );
and ( n45408 , n45407 , n44766 );
xor ( n45409 , n45335 , n45354 );
and ( n45410 , n45409 , n41611 );
or ( n45411 , n45408 , n45410 );
not ( n45412 , n45411 );
buf ( n45413 , n45412 );
buf ( n45414 , n45413 );
not ( n45415 , n45414 );
not ( n45416 , n45415 );
not ( n45417 , n41611 );
and ( n45418 , n45417 , n44767 );
xor ( n45419 , n45336 , n45353 );
and ( n45420 , n45419 , n41611 );
or ( n45421 , n45418 , n45420 );
not ( n45422 , n45421 );
buf ( n45423 , n45422 );
buf ( n45424 , n45423 );
not ( n45425 , n45424 );
not ( n45426 , n45425 );
not ( n45427 , n41611 );
and ( n45428 , n45427 , n44768 );
xor ( n45429 , n45337 , n45352 );
and ( n45430 , n45429 , n41611 );
or ( n45431 , n45428 , n45430 );
not ( n45432 , n45431 );
buf ( n45433 , n45432 );
buf ( n45434 , n45433 );
not ( n45435 , n45434 );
not ( n45436 , n45435 );
not ( n45437 , n41611 );
and ( n45438 , n45437 , n44769 );
xor ( n45439 , n45338 , n45351 );
and ( n45440 , n45439 , n41611 );
or ( n45441 , n45438 , n45440 );
not ( n45442 , n45441 );
buf ( n45443 , n45442 );
buf ( n45444 , n45443 );
not ( n45445 , n45444 );
not ( n45446 , n45445 );
not ( n45447 , n41611 );
and ( n45448 , n45447 , n44770 );
xor ( n45449 , n45339 , n45350 );
and ( n45450 , n45449 , n41611 );
or ( n45451 , n45448 , n45450 );
not ( n45452 , n45451 );
buf ( n45453 , n45452 );
buf ( n45454 , n45453 );
not ( n45455 , n45454 );
not ( n45456 , n45455 );
not ( n45457 , n41611 );
and ( n45458 , n45457 , n44771 );
xor ( n45459 , n45340 , n45349 );
and ( n45460 , n45459 , n41611 );
or ( n45461 , n45458 , n45460 );
not ( n45462 , n45461 );
buf ( n45463 , n45462 );
buf ( n45464 , n45463 );
not ( n45465 , n45464 );
not ( n45466 , n45465 );
not ( n45467 , n41611 );
and ( n45468 , n45467 , n44772 );
xor ( n45469 , n45341 , n45348 );
and ( n45470 , n45469 , n41611 );
or ( n45471 , n45468 , n45470 );
not ( n45472 , n45471 );
buf ( n45473 , n45472 );
buf ( n45474 , n45473 );
not ( n45475 , n45474 );
not ( n45476 , n45475 );
not ( n45477 , n41611 );
and ( n45478 , n45477 , n44773 );
xor ( n45479 , n45342 , n45347 );
and ( n45480 , n45479 , n41611 );
or ( n45481 , n45478 , n45480 );
not ( n45482 , n45481 );
buf ( n45483 , n45482 );
buf ( n45484 , n45483 );
not ( n45485 , n45484 );
not ( n45486 , n45485 );
not ( n45487 , n41611 );
and ( n45488 , n45487 , n44774 );
xor ( n45489 , n45343 , n45346 );
and ( n45490 , n45489 , n41611 );
or ( n45491 , n45488 , n45490 );
not ( n45492 , n45491 );
buf ( n45493 , n45492 );
buf ( n45494 , n45493 );
not ( n45495 , n45494 );
not ( n45496 , n45495 );
not ( n45497 , n41611 );
and ( n45498 , n45497 , n44775 );
xor ( n45499 , n45344 , n45345 );
and ( n45500 , n45499 , n41611 );
or ( n45501 , n45498 , n45500 );
not ( n45502 , n45501 );
buf ( n45503 , n45502 );
buf ( n45504 , n45503 );
not ( n45505 , n45504 );
not ( n45506 , n45505 );
not ( n45507 , n45323 );
and ( n45508 , n45506 , n45507 );
and ( n45509 , n45496 , n45508 );
and ( n45510 , n45486 , n45509 );
and ( n45511 , n45476 , n45510 );
and ( n45512 , n45466 , n45511 );
and ( n45513 , n45456 , n45512 );
and ( n45514 , n45446 , n45513 );
and ( n45515 , n45436 , n45514 );
and ( n45516 , n45426 , n45515 );
and ( n45517 , n45416 , n45516 );
and ( n45518 , n45406 , n45517 );
and ( n45519 , n45396 , n45518 );
and ( n45520 , n45386 , n45519 );
and ( n45521 , n45376 , n45520 );
and ( n45522 , n45366 , n45521 );
not ( n45523 , n45522 );
and ( n45524 , n45523 , n41611 );
buf ( n45525 , n45524 );
not ( n45526 , n45525 );
not ( n45527 , n41611 );
and ( n45528 , n45527 , n45505 );
xor ( n45529 , n45506 , n45507 );
and ( n45530 , n45529 , n41611 );
or ( n45531 , n45528 , n45530 );
and ( n45532 , n45526 , n45531 );
not ( n45533 , n45531 );
not ( n45534 , n45324 );
xor ( n45535 , n45533 , n45534 );
and ( n45536 , n45535 , n45525 );
or ( n45537 , n45532 , n45536 );
not ( n45538 , n45537 );
buf ( n45539 , n45538 );
buf ( n45540 , n45539 );
not ( n45541 , n45540 );
or ( n45542 , n45328 , n45541 );
not ( n45543 , n45525 );
not ( n45544 , n41611 );
and ( n45545 , n45544 , n45495 );
xor ( n45546 , n45496 , n45508 );
and ( n45547 , n45546 , n41611 );
or ( n45548 , n45545 , n45547 );
and ( n45549 , n45543 , n45548 );
not ( n45550 , n45548 );
and ( n45551 , n45533 , n45534 );
xor ( n45552 , n45550 , n45551 );
and ( n45553 , n45552 , n45525 );
or ( n45554 , n45549 , n45553 );
not ( n45555 , n45554 );
buf ( n45556 , n45555 );
buf ( n45557 , n45556 );
not ( n45558 , n45557 );
or ( n45559 , n45542 , n45558 );
not ( n45560 , n45525 );
not ( n45561 , n41611 );
and ( n45562 , n45561 , n45485 );
xor ( n45563 , n45486 , n45509 );
and ( n45564 , n45563 , n41611 );
or ( n45565 , n45562 , n45564 );
and ( n45566 , n45560 , n45565 );
not ( n45567 , n45565 );
and ( n45568 , n45550 , n45551 );
xor ( n45569 , n45567 , n45568 );
and ( n45570 , n45569 , n45525 );
or ( n45571 , n45566 , n45570 );
not ( n45572 , n45571 );
buf ( n45573 , n45572 );
buf ( n45574 , n45573 );
not ( n45575 , n45574 );
or ( n45576 , n45559 , n45575 );
not ( n45577 , n45525 );
not ( n45578 , n41611 );
and ( n45579 , n45578 , n45475 );
xor ( n45580 , n45476 , n45510 );
and ( n45581 , n45580 , n41611 );
or ( n45582 , n45579 , n45581 );
and ( n45583 , n45577 , n45582 );
not ( n45584 , n45582 );
and ( n45585 , n45567 , n45568 );
xor ( n45586 , n45584 , n45585 );
and ( n45587 , n45586 , n45525 );
or ( n45588 , n45583 , n45587 );
not ( n45589 , n45588 );
buf ( n45590 , n45589 );
buf ( n45591 , n45590 );
not ( n45592 , n45591 );
or ( n45593 , n45576 , n45592 );
not ( n45594 , n45525 );
not ( n45595 , n41611 );
and ( n45596 , n45595 , n45465 );
xor ( n45597 , n45466 , n45511 );
and ( n45598 , n45597 , n41611 );
or ( n45599 , n45596 , n45598 );
and ( n45600 , n45594 , n45599 );
not ( n45601 , n45599 );
and ( n45602 , n45584 , n45585 );
xor ( n45603 , n45601 , n45602 );
and ( n45604 , n45603 , n45525 );
or ( n45605 , n45600 , n45604 );
not ( n45606 , n45605 );
buf ( n45607 , n45606 );
buf ( n45608 , n45607 );
not ( n45609 , n45608 );
or ( n45610 , n45593 , n45609 );
not ( n45611 , n45525 );
not ( n45612 , n41611 );
and ( n45613 , n45612 , n45455 );
xor ( n45614 , n45456 , n45512 );
and ( n45615 , n45614 , n41611 );
or ( n45616 , n45613 , n45615 );
and ( n45617 , n45611 , n45616 );
not ( n45618 , n45616 );
and ( n45619 , n45601 , n45602 );
xor ( n45620 , n45618 , n45619 );
and ( n45621 , n45620 , n45525 );
or ( n45622 , n45617 , n45621 );
not ( n45623 , n45622 );
buf ( n45624 , n45623 );
buf ( n45625 , n45624 );
not ( n45626 , n45625 );
or ( n45627 , n45610 , n45626 );
not ( n45628 , n45525 );
not ( n45629 , n41611 );
and ( n45630 , n45629 , n45445 );
xor ( n45631 , n45446 , n45513 );
and ( n45632 , n45631 , n41611 );
or ( n45633 , n45630 , n45632 );
and ( n45634 , n45628 , n45633 );
not ( n45635 , n45633 );
and ( n45636 , n45618 , n45619 );
xor ( n45637 , n45635 , n45636 );
and ( n45638 , n45637 , n45525 );
or ( n45639 , n45634 , n45638 );
not ( n45640 , n45639 );
buf ( n45641 , n45640 );
buf ( n45642 , n45641 );
not ( n45643 , n45642 );
or ( n45644 , n45627 , n45643 );
not ( n45645 , n45525 );
not ( n45646 , n41611 );
and ( n45647 , n45646 , n45435 );
xor ( n45648 , n45436 , n45514 );
and ( n45649 , n45648 , n41611 );
or ( n45650 , n45647 , n45649 );
and ( n45651 , n45645 , n45650 );
not ( n45652 , n45650 );
and ( n45653 , n45635 , n45636 );
xor ( n45654 , n45652 , n45653 );
and ( n45655 , n45654 , n45525 );
or ( n45656 , n45651 , n45655 );
not ( n45657 , n45656 );
buf ( n45658 , n45657 );
buf ( n45659 , n45658 );
not ( n45660 , n45659 );
or ( n45661 , n45644 , n45660 );
not ( n45662 , n45525 );
not ( n45663 , n41611 );
and ( n45664 , n45663 , n45425 );
xor ( n45665 , n45426 , n45515 );
and ( n45666 , n45665 , n41611 );
or ( n45667 , n45664 , n45666 );
and ( n45668 , n45662 , n45667 );
not ( n45669 , n45667 );
and ( n45670 , n45652 , n45653 );
xor ( n45671 , n45669 , n45670 );
and ( n45672 , n45671 , n45525 );
or ( n45673 , n45668 , n45672 );
not ( n45674 , n45673 );
buf ( n45675 , n45674 );
buf ( n45676 , n45675 );
not ( n45677 , n45676 );
or ( n45678 , n45661 , n45677 );
not ( n45679 , n45525 );
not ( n45680 , n41611 );
and ( n45681 , n45680 , n45415 );
xor ( n45682 , n45416 , n45516 );
and ( n45683 , n45682 , n41611 );
or ( n45684 , n45681 , n45683 );
and ( n45685 , n45679 , n45684 );
not ( n45686 , n45684 );
and ( n45687 , n45669 , n45670 );
xor ( n45688 , n45686 , n45687 );
and ( n45689 , n45688 , n45525 );
or ( n45690 , n45685 , n45689 );
not ( n45691 , n45690 );
buf ( n45692 , n45691 );
buf ( n45693 , n45692 );
not ( n45694 , n45693 );
or ( n45695 , n45678 , n45694 );
not ( n45696 , n45525 );
not ( n45697 , n41611 );
and ( n45698 , n45697 , n45405 );
xor ( n45699 , n45406 , n45517 );
and ( n45700 , n45699 , n41611 );
or ( n45701 , n45698 , n45700 );
and ( n45702 , n45696 , n45701 );
not ( n45703 , n45701 );
and ( n45704 , n45686 , n45687 );
xor ( n45705 , n45703 , n45704 );
and ( n45706 , n45705 , n45525 );
or ( n45707 , n45702 , n45706 );
not ( n45708 , n45707 );
buf ( n45709 , n45708 );
buf ( n45710 , n45709 );
not ( n45711 , n45710 );
or ( n45712 , n45695 , n45711 );
not ( n45713 , n45525 );
not ( n45714 , n41611 );
and ( n45715 , n45714 , n45395 );
xor ( n45716 , n45396 , n45518 );
and ( n45717 , n45716 , n41611 );
or ( n45718 , n45715 , n45717 );
and ( n45719 , n45713 , n45718 );
not ( n45720 , n45718 );
and ( n45721 , n45703 , n45704 );
xor ( n45722 , n45720 , n45721 );
and ( n45723 , n45722 , n45525 );
or ( n45724 , n45719 , n45723 );
not ( n45725 , n45724 );
buf ( n45726 , n45725 );
buf ( n45727 , n45726 );
not ( n45728 , n45727 );
or ( n45729 , n45712 , n45728 );
not ( n45730 , n45525 );
not ( n45731 , n41611 );
and ( n45732 , n45731 , n45385 );
xor ( n45733 , n45386 , n45519 );
and ( n45734 , n45733 , n41611 );
or ( n45735 , n45732 , n45734 );
and ( n45736 , n45730 , n45735 );
not ( n45737 , n45735 );
and ( n45738 , n45720 , n45721 );
xor ( n45739 , n45737 , n45738 );
and ( n45740 , n45739 , n45525 );
or ( n45741 , n45736 , n45740 );
not ( n45742 , n45741 );
buf ( n45743 , n45742 );
buf ( n45744 , n45743 );
not ( n45745 , n45744 );
or ( n45746 , n45729 , n45745 );
not ( n45747 , n45525 );
not ( n45748 , n41611 );
and ( n45749 , n45748 , n45375 );
xor ( n45750 , n45376 , n45520 );
and ( n45751 , n45750 , n41611 );
or ( n45752 , n45749 , n45751 );
and ( n45753 , n45747 , n45752 );
not ( n45754 , n45752 );
and ( n45755 , n45737 , n45738 );
xor ( n45756 , n45754 , n45755 );
and ( n45757 , n45756 , n45525 );
or ( n45758 , n45753 , n45757 );
not ( n45759 , n45758 );
buf ( n45760 , n45759 );
buf ( n45761 , n45760 );
not ( n45762 , n45761 );
or ( n45763 , n45746 , n45762 );
buf ( n45764 , n45763 );
buf ( n45765 , n45764 );
and ( n45766 , n45765 , n45525 );
not ( n45767 , n45766 );
and ( n45768 , n45767 , n45677 );
xor ( n45769 , n45677 , n45525 );
xor ( n45770 , n45660 , n45525 );
xor ( n45771 , n45643 , n45525 );
xor ( n45772 , n45626 , n45525 );
xor ( n45773 , n45609 , n45525 );
xor ( n45774 , n45592 , n45525 );
xor ( n45775 , n45575 , n45525 );
xor ( n45776 , n45558 , n45525 );
xor ( n45777 , n45541 , n45525 );
xor ( n45778 , n45328 , n45525 );
and ( n45779 , n45778 , n45525 );
and ( n45780 , n45777 , n45779 );
and ( n45781 , n45776 , n45780 );
and ( n45782 , n45775 , n45781 );
and ( n45783 , n45774 , n45782 );
and ( n45784 , n45773 , n45783 );
and ( n45785 , n45772 , n45784 );
and ( n45786 , n45771 , n45785 );
and ( n45787 , n45770 , n45786 );
xor ( n45788 , n45769 , n45787 );
and ( n45789 , n45788 , n45766 );
or ( n45790 , n45768 , n45789 );
and ( n45791 , n45790 , n45280 );
or ( n45792 , n45282 , n45791 );
and ( n45793 , n45792 , n31468 );
or ( n45794 , n31539 , n31521 );
or ( n45795 , n45794 , n31408 );
or ( n45796 , n45795 , n31540 );
or ( n45797 , n45796 , n31542 );
or ( n45798 , n45797 , n31544 );
or ( n45799 , n45798 , n31546 );
or ( n45800 , n45799 , n31548 );
or ( n45801 , n45800 , n31550 );
or ( n45802 , n45801 , n31552 );
and ( n45803 , n45276 , n45802 );
or ( n45804 , n45279 , n45793 , n45803 );
and ( n45805 , n45804 , n31557 );
or ( n45806 , n40150 , n31647 );
or ( n45807 , n45806 , n31649 );
or ( n45808 , n45807 , n31007 );
and ( n45809 , n45276 , n45808 );
or ( n45810 , C0 , n45273 , n45805 , n45809 );
buf ( n45811 , n45810 );
buf ( n45812 , n45811 );
buf ( n45813 , n31655 );
buf ( n45814 , n30987 );
buf ( n45815 , n30987 );
buf ( n45816 , n30987 );
not ( n45817 , n40163 );
and ( n45818 , n45817 , n32046 );
not ( n45819 , n45227 );
and ( n45820 , n45819 , n32046 );
and ( n45821 , n32130 , n45227 );
or ( n45822 , n45820 , n45821 );
and ( n45823 , n45822 , n40163 );
or ( n45824 , n45818 , n45823 );
and ( n45825 , n45824 , n32498 );
not ( n45826 , n45235 );
not ( n45827 , n45227 );
and ( n45828 , n45827 , n32046 );
not ( n45829 , n40373 );
and ( n45830 , n45829 , n40238 );
xor ( n45831 , n40383 , n40244 );
and ( n45832 , n45831 , n40373 );
or ( n45833 , n45830 , n45832 );
and ( n45834 , n45833 , n45227 );
or ( n45835 , n45828 , n45834 );
and ( n45836 , n45826 , n45835 );
and ( n45837 , n45833 , n45235 );
or ( n45838 , n45836 , n45837 );
and ( n45839 , n45838 , n32473 );
not ( n45840 , n32475 );
not ( n45841 , n45235 );
not ( n45842 , n45227 );
and ( n45843 , n45842 , n32046 );
and ( n45844 , n45833 , n45227 );
or ( n45845 , n45843 , n45844 );
and ( n45846 , n45841 , n45845 );
and ( n45847 , n45833 , n45235 );
or ( n45848 , n45846 , n45847 );
and ( n45849 , n45840 , n45848 );
not ( n45850 , n45255 );
not ( n45851 , n45257 );
and ( n45852 , n45851 , n45848 );
not ( n45853 , n40952 );
and ( n45854 , n45853 , n40550 );
xor ( n45855 , n40962 , n40830 );
and ( n45856 , n45855 , n40952 );
or ( n45857 , n45854 , n45856 );
and ( n45858 , n45857 , n45257 );
or ( n45859 , n45852 , n45858 );
and ( n45860 , n45850 , n45859 );
not ( n45861 , n41247 );
and ( n45862 , n45861 , n41037 );
xor ( n45863 , n41257 , n41129 );
and ( n45864 , n45863 , n41247 );
or ( n45865 , n45862 , n45864 );
and ( n45866 , n45865 , n45255 );
or ( n45867 , n45860 , n45866 );
and ( n45868 , n45867 , n32475 );
or ( n45869 , n45849 , n45868 );
and ( n45870 , n45869 , n32486 );
and ( n45871 , n32046 , n41278 );
or ( n45872 , C0 , n45825 , n45839 , n45870 , n45871 );
buf ( n45873 , n45872 );
buf ( n45874 , n45873 );
buf ( n45875 , RI15b52b60_687);
and ( n45876 , n45875 , n31645 );
not ( n45877 , n45274 );
and ( n45878 , n45877 , n35533 );
buf ( n45879 , n45878 );
and ( n45880 , n45879 , n31373 );
not ( n45881 , n45280 );
and ( n45882 , n45881 , n35533 );
not ( n45883 , n45766 );
and ( n45884 , n45883 , n45762 );
xor ( n45885 , n45762 , n45525 );
xor ( n45886 , n45745 , n45525 );
xor ( n45887 , n45728 , n45525 );
xor ( n45888 , n45711 , n45525 );
xor ( n45889 , n45694 , n45525 );
and ( n45890 , n45769 , n45787 );
and ( n45891 , n45889 , n45890 );
and ( n45892 , n45888 , n45891 );
and ( n45893 , n45887 , n45892 );
and ( n45894 , n45886 , n45893 );
xor ( n45895 , n45885 , n45894 );
and ( n45896 , n45895 , n45766 );
or ( n45897 , n45884 , n45896 );
and ( n45898 , n45897 , n45280 );
or ( n45899 , n45882 , n45898 );
and ( n45900 , n45899 , n31468 );
and ( n45901 , n35533 , n45802 );
or ( n45902 , n45880 , n45900 , n45901 );
and ( n45903 , n45902 , n31557 );
and ( n45904 , n35533 , n45808 );
or ( n45905 , C0 , n45876 , n45903 , n45904 );
buf ( n45906 , n45905 );
buf ( n45907 , n45906 );
buf ( n45908 , n30987 );
buf ( n45909 , n31655 );
buf ( n45910 , n31655 );
and ( n45911 , n33237 , n32528 );
not ( n45912 , n32598 );
and ( n45913 , n45912 , n33000 );
and ( n45914 , n32543 , n32547 );
and ( n45915 , n32539 , n45914 );
and ( n45916 , n32535 , n45915 );
xor ( n45917 , n32531 , n45916 );
and ( n45918 , n45917 , n32598 );
or ( n45919 , n45913 , n45918 );
and ( n45920 , n45919 , n32890 );
not ( n45921 , n32919 );
and ( n45922 , n45921 , n33000 );
and ( n45923 , n45917 , n32919 );
or ( n45924 , n45922 , n45923 );
and ( n45925 , n45924 , n32924 );
not ( n45926 , n32953 );
and ( n45927 , n45926 , n33000 );
not ( n45928 , n32971 );
and ( n45929 , n45928 , n33125 );
xor ( n45930 , n33000 , n33005 );
and ( n45931 , n45930 , n32971 );
or ( n45932 , n45929 , n45931 );
and ( n45933 , n45932 , n32953 );
or ( n45934 , n45927 , n45933 );
and ( n45935 , n45934 , n33038 );
not ( n45936 , n33067 );
and ( n45937 , n45936 , n33000 );
not ( n45938 , n32970 );
not ( n45939 , n33071 );
and ( n45940 , n45939 , n33125 );
xor ( n45941 , n33126 , n33137 );
and ( n45942 , n45941 , n33071 );
or ( n45943 , n45940 , n45942 );
and ( n45944 , n45938 , n45943 );
and ( n45945 , n45930 , n32970 );
or ( n45946 , n45944 , n45945 );
and ( n45947 , n45946 , n33067 );
or ( n45948 , n45937 , n45947 );
and ( n45949 , n45948 , n33172 );
and ( n45950 , n33000 , n33204 );
or ( n45951 , n45920 , n45925 , n45935 , n45949 , n45950 );
and ( n45952 , n45951 , n33208 );
not ( n45953 , n32968 );
not ( n45954 , n33270 );
and ( n45955 , n45954 , n33325 );
xor ( n45956 , n33326 , n33337 );
and ( n45957 , n45956 , n33270 );
or ( n45958 , n45955 , n45957 );
and ( n45959 , n45953 , n45958 );
and ( n45960 , n33000 , n32968 );
or ( n45961 , n45959 , n45960 );
and ( n45962 , n45961 , n33370 );
buf ( n45963 , n35056 );
and ( n45964 , n33000 , n33382 );
or ( n45965 , C0 , n45911 , n45952 , n45962 , n45963 , n45964 );
buf ( n45966 , n45965 );
buf ( n45967 , n45966 );
buf ( n45968 , n30987 );
buf ( n45969 , n30987 );
and ( n45970 , n32463 , n32500 );
not ( n45971 , n35211 );
and ( n45972 , n45971 , n37585 );
and ( n45973 , n31763 , n35211 );
or ( n45974 , n45972 , n45973 );
and ( n45975 , n45974 , n32421 );
not ( n45976 , n35245 );
and ( n45977 , n45976 , n37585 );
and ( n45978 , n31763 , n35245 );
or ( n45979 , n45977 , n45978 );
and ( n45980 , n45979 , n32419 );
not ( n45981 , n35278 );
and ( n45982 , n45981 , n37585 );
not ( n45983 , n35295 );
buf ( n45984 , RI15b61d40_1203);
and ( n45985 , n45983 , n45984 );
xor ( n45986 , n37585 , n37514 );
and ( n45987 , n45986 , n35295 );
or ( n45988 , n45985 , n45987 );
and ( n45989 , n45988 , n35278 );
or ( n45990 , n45982 , n45989 );
and ( n45991 , n45990 , n32417 );
not ( n45992 , n35331 );
and ( n45993 , n45992 , n37585 );
not ( n45994 , n35294 );
buf ( n45995 , RI15b62ad8_1232);
not ( n45996 , n45995 );
and ( n45997 , n45996 , n45984 );
not ( n45998 , n45984 );
buf ( n45999 , RI15b61cc8_1202);
not ( n46000 , n45999 );
not ( n46001 , n35297 );
and ( n46002 , n46000 , n46001 );
xor ( n46003 , n45998 , n46002 );
and ( n46004 , n46003 , n45995 );
or ( n46005 , n45997 , n46004 );
and ( n46006 , n45994 , n46005 );
and ( n46007 , n45986 , n35294 );
or ( n46008 , n46006 , n46007 );
and ( n46009 , n46008 , n35331 );
or ( n46010 , n45993 , n46009 );
and ( n46011 , n46010 , n32415 );
and ( n46012 , n37585 , n35354 );
or ( n46013 , n45975 , n45980 , n45991 , n46011 , n46012 );
and ( n46014 , n46013 , n32456 );
not ( n46015 , n32475 );
buf ( n46016 , RI15b639d8_1264);
buf ( n46017 , RI15b63960_1263);
buf ( n46018 , RI15b638e8_1262);
buf ( n46019 , RI15b63870_1261);
buf ( n46020 , RI15b637f8_1260);
buf ( n46021 , RI15b63780_1259);
buf ( n46022 , RI15b63708_1258);
buf ( n46023 , RI15b63690_1257);
buf ( n46024 , RI15b63618_1256);
buf ( n46025 , RI15b635a0_1255);
buf ( n46026 , RI15b63528_1254);
buf ( n46027 , RI15b634b0_1253);
buf ( n46028 , RI15b63438_1252);
buf ( n46029 , RI15b633c0_1251);
buf ( n46030 , RI15b63348_1250);
buf ( n46031 , RI15b632d0_1249);
buf ( n46032 , RI15b63258_1248);
buf ( n46033 , RI15b631e0_1247);
buf ( n46034 , RI15b63168_1246);
buf ( n46035 , RI15b630f0_1245);
buf ( n46036 , RI15b63078_1244);
buf ( n46037 , RI15b63000_1243);
and ( n46038 , n41284 , n41314 );
and ( n46039 , n46037 , n46038 );
and ( n46040 , n46036 , n46039 );
and ( n46041 , n46035 , n46040 );
and ( n46042 , n46034 , n46041 );
and ( n46043 , n46033 , n46042 );
and ( n46044 , n46032 , n46043 );
and ( n46045 , n46031 , n46044 );
and ( n46046 , n46030 , n46045 );
and ( n46047 , n46029 , n46046 );
and ( n46048 , n46028 , n46047 );
and ( n46049 , n46027 , n46048 );
and ( n46050 , n46026 , n46049 );
and ( n46051 , n46025 , n46050 );
and ( n46052 , n46024 , n46051 );
and ( n46053 , n46023 , n46052 );
and ( n46054 , n46022 , n46053 );
and ( n46055 , n46021 , n46054 );
and ( n46056 , n46020 , n46055 );
and ( n46057 , n46019 , n46056 );
and ( n46058 , n46018 , n46057 );
and ( n46059 , n46017 , n46058 );
xor ( n46060 , n46016 , n46059 );
not ( n46061 , n46060 );
xor ( n46062 , n32463 , n32464 );
and ( n46063 , n46061 , n46062 );
not ( n46064 , n46062 );
not ( n46065 , n32464 );
not ( n46066 , n46065 );
not ( n46067 , n35182 );
and ( n46068 , n46066 , n46067 );
xor ( n46069 , n46064 , n46068 );
and ( n46070 , n46069 , n46060 );
or ( n46071 , n46063 , n46070 );
and ( n46072 , n46015 , n46071 );
and ( n46073 , n37585 , n32475 );
or ( n46074 , n46072 , n46073 );
and ( n46075 , n46074 , n32486 );
and ( n46076 , n37585 , n35367 );
or ( n46077 , C0 , n45970 , n46014 , n46075 , C0 , n46076 );
buf ( n46078 , n46077 );
buf ( n46079 , n46078 );
buf ( n46080 , n31655 );
buf ( n46081 , RI15b5f658_1120);
and ( n46082 , n46081 , n32494 );
and ( n46083 , n35211 , n35288 );
not ( n46084 , n46083 );
buf ( n46085 , RI15b5fdd8_1136);
and ( n46086 , n46084 , n46085 );
buf ( n46087 , RI15b60d50_1169);
buf ( n46088 , n46087 );
not ( n46089 , n46088 );
buf ( n46090 , n46089 );
not ( n46091 , n46090 );
buf ( n46092 , RI15b61bd8_1200);
not ( n46093 , n46092 );
buf ( n46094 , RI15b60dc8_1170);
and ( n46095 , n46093 , n46094 );
not ( n46096 , n46094 );
not ( n46097 , n46087 );
xor ( n46098 , n46096 , n46097 );
and ( n46099 , n46098 , n46092 );
or ( n46100 , n46095 , n46099 );
not ( n46101 , n46100 );
buf ( n46102 , n46101 );
buf ( n46103 , n46102 );
not ( n46104 , n46103 );
or ( n46105 , n46091 , n46104 );
not ( n46106 , n46092 );
buf ( n46107 , RI15b60e40_1171);
and ( n46108 , n46106 , n46107 );
not ( n46109 , n46107 );
and ( n46110 , n46096 , n46097 );
xor ( n46111 , n46109 , n46110 );
and ( n46112 , n46111 , n46092 );
or ( n46113 , n46108 , n46112 );
not ( n46114 , n46113 );
buf ( n46115 , n46114 );
buf ( n46116 , n46115 );
not ( n46117 , n46116 );
or ( n46118 , n46105 , n46117 );
not ( n46119 , n46092 );
buf ( n46120 , RI15b60eb8_1172);
and ( n46121 , n46119 , n46120 );
not ( n46122 , n46120 );
and ( n46123 , n46109 , n46110 );
xor ( n46124 , n46122 , n46123 );
and ( n46125 , n46124 , n46092 );
or ( n46126 , n46121 , n46125 );
not ( n46127 , n46126 );
buf ( n46128 , n46127 );
buf ( n46129 , n46128 );
not ( n46130 , n46129 );
or ( n46131 , n46118 , n46130 );
not ( n46132 , n46092 );
buf ( n46133 , RI15b60f30_1173);
and ( n46134 , n46132 , n46133 );
not ( n46135 , n46133 );
and ( n46136 , n46122 , n46123 );
xor ( n46137 , n46135 , n46136 );
and ( n46138 , n46137 , n46092 );
or ( n46139 , n46134 , n46138 );
not ( n46140 , n46139 );
buf ( n46141 , n46140 );
buf ( n46142 , n46141 );
not ( n46143 , n46142 );
or ( n46144 , n46131 , n46143 );
not ( n46145 , n46092 );
buf ( n46146 , RI15b60fa8_1174);
and ( n46147 , n46145 , n46146 );
not ( n46148 , n46146 );
and ( n46149 , n46135 , n46136 );
xor ( n46150 , n46148 , n46149 );
and ( n46151 , n46150 , n46092 );
or ( n46152 , n46147 , n46151 );
not ( n46153 , n46152 );
buf ( n46154 , n46153 );
buf ( n46155 , n46154 );
not ( n46156 , n46155 );
or ( n46157 , n46144 , n46156 );
not ( n46158 , n46092 );
buf ( n46159 , RI15b61020_1175);
and ( n46160 , n46158 , n46159 );
not ( n46161 , n46159 );
and ( n46162 , n46148 , n46149 );
xor ( n46163 , n46161 , n46162 );
and ( n46164 , n46163 , n46092 );
or ( n46165 , n46160 , n46164 );
not ( n46166 , n46165 );
buf ( n46167 , n46166 );
buf ( n46168 , n46167 );
not ( n46169 , n46168 );
or ( n46170 , n46157 , n46169 );
not ( n46171 , n46092 );
buf ( n46172 , RI15b61098_1176);
and ( n46173 , n46171 , n46172 );
not ( n46174 , n46172 );
and ( n46175 , n46161 , n46162 );
xor ( n46176 , n46174 , n46175 );
and ( n46177 , n46176 , n46092 );
or ( n46178 , n46173 , n46177 );
not ( n46179 , n46178 );
buf ( n46180 , n46179 );
buf ( n46181 , n46180 );
not ( n46182 , n46181 );
or ( n46183 , n46170 , n46182 );
not ( n46184 , n46092 );
buf ( n46185 , RI15b61110_1177);
and ( n46186 , n46184 , n46185 );
not ( n46187 , n46185 );
and ( n46188 , n46174 , n46175 );
xor ( n46189 , n46187 , n46188 );
and ( n46190 , n46189 , n46092 );
or ( n46191 , n46186 , n46190 );
not ( n46192 , n46191 );
buf ( n46193 , n46192 );
buf ( n46194 , n46193 );
not ( n46195 , n46194 );
or ( n46196 , n46183 , n46195 );
not ( n46197 , n46092 );
buf ( n46198 , RI15b61188_1178);
and ( n46199 , n46197 , n46198 );
not ( n46200 , n46198 );
and ( n46201 , n46187 , n46188 );
xor ( n46202 , n46200 , n46201 );
and ( n46203 , n46202 , n46092 );
or ( n46204 , n46199 , n46203 );
not ( n46205 , n46204 );
buf ( n46206 , n46205 );
buf ( n46207 , n46206 );
not ( n46208 , n46207 );
or ( n46209 , n46196 , n46208 );
not ( n46210 , n46092 );
buf ( n46211 , RI15b61200_1179);
and ( n46212 , n46210 , n46211 );
not ( n46213 , n46211 );
and ( n46214 , n46200 , n46201 );
xor ( n46215 , n46213 , n46214 );
and ( n46216 , n46215 , n46092 );
or ( n46217 , n46212 , n46216 );
not ( n46218 , n46217 );
buf ( n46219 , n46218 );
buf ( n46220 , n46219 );
not ( n46221 , n46220 );
or ( n46222 , n46209 , n46221 );
not ( n46223 , n46092 );
buf ( n46224 , RI15b61278_1180);
and ( n46225 , n46223 , n46224 );
not ( n46226 , n46224 );
and ( n46227 , n46213 , n46214 );
xor ( n46228 , n46226 , n46227 );
and ( n46229 , n46228 , n46092 );
or ( n46230 , n46225 , n46229 );
not ( n46231 , n46230 );
buf ( n46232 , n46231 );
buf ( n46233 , n46232 );
not ( n46234 , n46233 );
or ( n46235 , n46222 , n46234 );
not ( n46236 , n46092 );
buf ( n46237 , RI15b612f0_1181);
and ( n46238 , n46236 , n46237 );
not ( n46239 , n46237 );
and ( n46240 , n46226 , n46227 );
xor ( n46241 , n46239 , n46240 );
and ( n46242 , n46241 , n46092 );
or ( n46243 , n46238 , n46242 );
not ( n46244 , n46243 );
buf ( n46245 , n46244 );
buf ( n46246 , n46245 );
not ( n46247 , n46246 );
or ( n46248 , n46235 , n46247 );
not ( n46249 , n46092 );
buf ( n46250 , RI15b61368_1182);
and ( n46251 , n46249 , n46250 );
not ( n46252 , n46250 );
and ( n46253 , n46239 , n46240 );
xor ( n46254 , n46252 , n46253 );
and ( n46255 , n46254 , n46092 );
or ( n46256 , n46251 , n46255 );
not ( n46257 , n46256 );
buf ( n46258 , n46257 );
buf ( n46259 , n46258 );
not ( n46260 , n46259 );
or ( n46261 , n46248 , n46260 );
not ( n46262 , n46092 );
buf ( n46263 , RI15b613e0_1183);
and ( n46264 , n46262 , n46263 );
not ( n46265 , n46263 );
and ( n46266 , n46252 , n46253 );
xor ( n46267 , n46265 , n46266 );
and ( n46268 , n46267 , n46092 );
or ( n46269 , n46264 , n46268 );
not ( n46270 , n46269 );
buf ( n46271 , n46270 );
buf ( n46272 , n46271 );
not ( n46273 , n46272 );
or ( n46274 , n46261 , n46273 );
not ( n46275 , n46092 );
buf ( n46276 , RI15b61458_1184);
and ( n46277 , n46275 , n46276 );
not ( n46278 , n46276 );
and ( n46279 , n46265 , n46266 );
xor ( n46280 , n46278 , n46279 );
and ( n46281 , n46280 , n46092 );
or ( n46282 , n46277 , n46281 );
not ( n46283 , n46282 );
buf ( n46284 , n46283 );
buf ( n46285 , n46284 );
not ( n46286 , n46285 );
or ( n46287 , n46274 , n46286 );
buf ( n46288 , n46287 );
buf ( n46289 , n46288 );
and ( n46290 , n46289 , n46092 );
not ( n46291 , n46290 );
and ( n46292 , n46291 , n46260 );
xor ( n46293 , n46260 , n46092 );
xor ( n46294 , n46247 , n46092 );
xor ( n46295 , n46234 , n46092 );
xor ( n46296 , n46221 , n46092 );
xor ( n46297 , n46208 , n46092 );
xor ( n46298 , n46195 , n46092 );
xor ( n46299 , n46182 , n46092 );
xor ( n46300 , n46169 , n46092 );
xor ( n46301 , n46156 , n46092 );
xor ( n46302 , n46143 , n46092 );
xor ( n46303 , n46130 , n46092 );
xor ( n46304 , n46117 , n46092 );
xor ( n46305 , n46104 , n46092 );
xor ( n46306 , n46091 , n46092 );
and ( n46307 , n46306 , n46092 );
and ( n46308 , n46305 , n46307 );
and ( n46309 , n46304 , n46308 );
and ( n46310 , n46303 , n46309 );
and ( n46311 , n46302 , n46310 );
and ( n46312 , n46301 , n46311 );
and ( n46313 , n46300 , n46312 );
and ( n46314 , n46299 , n46313 );
and ( n46315 , n46298 , n46314 );
and ( n46316 , n46297 , n46315 );
and ( n46317 , n46296 , n46316 );
and ( n46318 , n46295 , n46317 );
and ( n46319 , n46294 , n46318 );
xor ( n46320 , n46293 , n46319 );
and ( n46321 , n46320 , n46290 );
or ( n46322 , n46292 , n46321 );
and ( n46323 , n46322 , n46083 );
or ( n46324 , n46086 , n46323 );
and ( n46325 , n46324 , n32421 );
and ( n46326 , n35278 , n35288 );
not ( n46327 , n46326 );
and ( n46328 , n46327 , n46085 );
and ( n46329 , n46322 , n46326 );
or ( n46330 , n46328 , n46329 );
and ( n46331 , n46330 , n32417 );
or ( n46332 , n35347 , n32415 );
or ( n46333 , n46332 , n32419 );
or ( n46334 , n46333 , n32423 );
or ( n46335 , n46334 , n32425 );
or ( n46336 , n46335 , n32427 );
or ( n46337 , n46336 , n32429 );
or ( n46338 , n46337 , n32431 );
or ( n46339 , n46338 , n32433 );
or ( n46340 , n46339 , n32435 );
and ( n46341 , n46085 , n46340 );
or ( n46342 , n46325 , n46331 , n46341 );
and ( n46343 , n46342 , n32456 );
or ( n46344 , n41273 , n32486 );
or ( n46345 , n46344 , n32492 );
or ( n46346 , n46345 , n32473 );
or ( n46347 , n46346 , n32496 );
or ( n46348 , n46347 , n32498 );
or ( n46349 , n46348 , n32500 );
and ( n46350 , n46085 , n46349 );
or ( n46351 , C0 , n46082 , n46343 , n46350 );
buf ( n46352 , n46351 );
buf ( n46353 , n46352 );
buf ( n46354 , n31655 );
buf ( n46355 , n30987 );
not ( n46356 , n31010 );
not ( n46357 , n46356 );
and ( n46358 , n46357 , n31146 );
not ( n46359 , n31025 );
not ( n46360 , n31021 );
not ( n46361 , n31009 );
and ( n46362 , n46359 , n46360 , n31017 , n31013 , n46361 );
not ( n46363 , n46362 );
and ( n46364 , n46363 , n31146 );
and ( n46365 , n31172 , n46362 );
or ( n46366 , n46364 , n46365 );
and ( n46367 , n46366 , n46356 );
or ( n46368 , n46358 , n46367 );
and ( n46369 , n46368 , n31649 );
not ( n46370 , n31025 );
not ( n46371 , n46370 );
buf ( n46372 , n46371 );
not ( n46373 , n46372 );
not ( n46374 , n46373 );
xor ( n46375 , n31021 , n31025 );
not ( n46376 , n46375 );
buf ( n46377 , n46376 );
buf ( n46378 , n46377 );
not ( n46379 , n46378 );
not ( n46380 , n46379 );
and ( n46381 , n31021 , n31025 );
xor ( n46382 , n31017 , n46381 );
not ( n46383 , n46382 );
buf ( n46384 , n46383 );
buf ( n46385 , n46384 );
not ( n46386 , n46385 );
and ( n46387 , n31017 , n46381 );
xor ( n46388 , n31013 , n46387 );
not ( n46389 , n46388 );
buf ( n46390 , n46389 );
buf ( n46391 , n46390 );
not ( n46392 , n46391 );
and ( n46393 , n46374 , n46380 , n46386 , n46392 , C1 );
not ( n46394 , n46393 );
not ( n46395 , n46362 );
and ( n46396 , n46395 , n31146 );
buf ( n46397 , n41873 );
not ( n46398 , n46397 );
buf ( n46399 , n46398 );
not ( n46400 , n46399 );
not ( n46401 , n41881 );
and ( n46402 , n46401 , n41886 );
not ( n46403 , n41886 );
not ( n46404 , n41873 );
xor ( n46405 , n46403 , n46404 );
and ( n46406 , n46405 , n41881 );
or ( n46407 , n46402 , n46406 );
not ( n46408 , n46407 );
buf ( n46409 , n46408 );
buf ( n46410 , n46409 );
not ( n46411 , n46410 );
or ( n46412 , n46400 , n46411 );
not ( n46413 , n41881 );
and ( n46414 , n46413 , n41902 );
not ( n46415 , n41902 );
and ( n46416 , n46403 , n46404 );
xor ( n46417 , n46415 , n46416 );
and ( n46418 , n46417 , n41881 );
or ( n46419 , n46414 , n46418 );
not ( n46420 , n46419 );
buf ( n46421 , n46420 );
buf ( n46422 , n46421 );
not ( n46423 , n46422 );
or ( n46424 , n46412 , n46423 );
not ( n46425 , n41881 );
and ( n46426 , n46425 , n41918 );
not ( n46427 , n41918 );
and ( n46428 , n46415 , n46416 );
xor ( n46429 , n46427 , n46428 );
and ( n46430 , n46429 , n41881 );
or ( n46431 , n46426 , n46430 );
not ( n46432 , n46431 );
buf ( n46433 , n46432 );
buf ( n46434 , n46433 );
not ( n46435 , n46434 );
or ( n46436 , n46424 , n46435 );
not ( n46437 , n41881 );
and ( n46438 , n46437 , n41934 );
not ( n46439 , n41934 );
and ( n46440 , n46427 , n46428 );
xor ( n46441 , n46439 , n46440 );
and ( n46442 , n46441 , n41881 );
or ( n46443 , n46438 , n46442 );
not ( n46444 , n46443 );
buf ( n46445 , n46444 );
buf ( n46446 , n46445 );
not ( n46447 , n46446 );
or ( n46448 , n46436 , n46447 );
not ( n46449 , n41881 );
and ( n46450 , n46449 , n41950 );
not ( n46451 , n41950 );
and ( n46452 , n46439 , n46440 );
xor ( n46453 , n46451 , n46452 );
and ( n46454 , n46453 , n41881 );
or ( n46455 , n46450 , n46454 );
not ( n46456 , n46455 );
buf ( n46457 , n46456 );
buf ( n46458 , n46457 );
not ( n46459 , n46458 );
or ( n46460 , n46448 , n46459 );
not ( n46461 , n41881 );
and ( n46462 , n46461 , n41966 );
not ( n46463 , n41966 );
and ( n46464 , n46451 , n46452 );
xor ( n46465 , n46463 , n46464 );
and ( n46466 , n46465 , n41881 );
or ( n46467 , n46462 , n46466 );
not ( n46468 , n46467 );
buf ( n46469 , n46468 );
buf ( n46470 , n46469 );
not ( n46471 , n46470 );
or ( n46472 , n46460 , n46471 );
not ( n46473 , n41881 );
and ( n46474 , n46473 , n41982 );
not ( n46475 , n41982 );
and ( n46476 , n46463 , n46464 );
xor ( n46477 , n46475 , n46476 );
and ( n46478 , n46477 , n41881 );
or ( n46479 , n46474 , n46478 );
not ( n46480 , n46479 );
buf ( n46481 , n46480 );
buf ( n46482 , n46481 );
not ( n46483 , n46482 );
or ( n46484 , n46472 , n46483 );
buf ( n46485 , n46484 );
buf ( n46486 , n46485 );
and ( n46487 , n46486 , n41881 );
not ( n46488 , n46487 );
and ( n46489 , n46488 , n46411 );
xor ( n46490 , n46411 , n41881 );
xor ( n46491 , n46400 , n41881 );
and ( n46492 , n46491 , n41881 );
xor ( n46493 , n46490 , n46492 );
and ( n46494 , n46493 , n46487 );
or ( n46495 , n46489 , n46494 );
and ( n46496 , n46495 , n46362 );
or ( n46497 , n46396 , n46496 );
and ( n46498 , n46394 , n46497 );
and ( n46499 , n46495 , n46393 );
or ( n46500 , n46498 , n46499 );
and ( n46501 , n46500 , n31643 );
not ( n46502 , n31452 );
not ( n46503 , n46393 );
not ( n46504 , n46362 );
and ( n46505 , n46504 , n31146 );
and ( n46506 , n46495 , n46362 );
or ( n46507 , n46505 , n46506 );
and ( n46508 , n46503 , n46507 );
and ( n46509 , n46495 , n46393 );
or ( n46510 , n46508 , n46509 );
and ( n46511 , n46502 , n46510 );
not ( n46512 , n46373 );
not ( n46513 , n46512 );
buf ( n46514 , n46513 );
not ( n46515 , n46514 );
not ( n46516 , n46515 );
not ( n46517 , n46516 );
buf ( n46518 , n46517 );
not ( n46519 , n46518 );
not ( n46520 , n46519 );
xor ( n46521 , n46379 , n46373 );
not ( n46522 , n46521 );
buf ( n46523 , n46522 );
not ( n46524 , n46523 );
xor ( n46525 , n46524 , n46515 );
not ( n46526 , n46525 );
buf ( n46527 , n46526 );
not ( n46528 , n46527 );
not ( n46529 , n46528 );
and ( n46530 , n46379 , n46373 );
xor ( n46531 , n46386 , n46530 );
not ( n46532 , n46531 );
buf ( n46533 , n46532 );
not ( n46534 , n46533 );
and ( n46535 , n46524 , n46515 );
xor ( n46536 , n46534 , n46535 );
not ( n46537 , n46536 );
buf ( n46538 , n46537 );
not ( n46539 , n46538 );
and ( n46540 , n46386 , n46530 );
xor ( n46541 , n46392 , n46540 );
not ( n46542 , n46541 );
buf ( n46543 , n46542 );
not ( n46544 , n46543 );
and ( n46545 , n46534 , n46535 );
xor ( n46546 , n46544 , n46545 );
not ( n46547 , n46546 );
buf ( n46548 , n46547 );
not ( n46549 , n46548 );
and ( n46550 , n46520 , n46529 , n46539 , n46549 , C1 );
not ( n46551 , n46550 );
not ( n46552 , n46515 );
not ( n46553 , n46524 );
and ( n46554 , n46552 , n46553 , n46534 , n46544 , C1 );
not ( n46555 , n46554 );
and ( n46556 , n46555 , n46510 );
not ( n46557 , n41881 );
not ( n46558 , n41869 );
and ( n46559 , n46558 , n34362 );
and ( n46560 , n40455 , n41869 );
or ( n46561 , n46559 , n46560 );
and ( n46562 , n46557 , n46561 );
not ( n46563 , n46561 );
not ( n46564 , n42110 );
not ( n46565 , n42094 );
not ( n46566 , n42078 );
not ( n46567 , n42062 );
not ( n46568 , n42046 );
not ( n46569 , n42030 );
not ( n46570 , n42014 );
not ( n46571 , n41998 );
not ( n46572 , n41982 );
not ( n46573 , n41966 );
not ( n46574 , n41950 );
not ( n46575 , n41934 );
not ( n46576 , n41918 );
not ( n46577 , n41902 );
not ( n46578 , n41886 );
not ( n46579 , n41873 );
and ( n46580 , n46578 , n46579 );
and ( n46581 , n46577 , n46580 );
and ( n46582 , n46576 , n46581 );
and ( n46583 , n46575 , n46582 );
and ( n46584 , n46574 , n46583 );
and ( n46585 , n46573 , n46584 );
and ( n46586 , n46572 , n46585 );
and ( n46587 , n46571 , n46586 );
and ( n46588 , n46570 , n46587 );
and ( n46589 , n46569 , n46588 );
and ( n46590 , n46568 , n46589 );
and ( n46591 , n46567 , n46590 );
and ( n46592 , n46566 , n46591 );
and ( n46593 , n46565 , n46592 );
and ( n46594 , n46564 , n46593 );
xor ( n46595 , n46563 , n46594 );
and ( n46596 , n46595 , n41881 );
or ( n46597 , n46562 , n46596 );
not ( n46598 , n46597 );
buf ( n46599 , n46598 );
buf ( n46600 , n46599 );
not ( n46601 , n46600 );
buf ( n46602 , n46601 );
buf ( n46603 , n46602 );
not ( n46604 , n46603 );
buf ( n46605 , n46604 );
not ( n46606 , n46605 );
not ( n46607 , n41881 );
not ( n46608 , n41869 );
and ( n46609 , n46608 , n34417 );
and ( n46610 , n40555 , n41869 );
or ( n46611 , n46609 , n46610 );
not ( n46612 , n46611 );
not ( n46613 , n44813 );
not ( n46614 , n41869 );
and ( n46615 , n46614 , n34421 );
and ( n46616 , n40569 , n41869 );
or ( n46617 , n46615 , n46616 );
not ( n46618 , n46617 );
not ( n46619 , n41869 );
and ( n46620 , n46619 , n34423 );
and ( n46621 , n40576 , n41869 );
or ( n46622 , n46620 , n46621 );
not ( n46623 , n46622 );
not ( n46624 , n41869 );
and ( n46625 , n46624 , n34425 );
and ( n46626 , n40583 , n41869 );
or ( n46627 , n46625 , n46626 );
not ( n46628 , n46627 );
not ( n46629 , n41869 );
and ( n46630 , n46629 , n34427 );
and ( n46631 , n40590 , n41869 );
or ( n46632 , n46630 , n46631 );
not ( n46633 , n46632 );
not ( n46634 , n41869 );
and ( n46635 , n46634 , n34429 );
and ( n46636 , n40597 , n41869 );
or ( n46637 , n46635 , n46636 );
not ( n46638 , n46637 );
not ( n46639 , n41869 );
and ( n46640 , n46639 , n34431 );
and ( n46641 , n40604 , n41869 );
or ( n46642 , n46640 , n46641 );
not ( n46643 , n46642 );
not ( n46644 , n41869 );
and ( n46645 , n46644 , n34433 );
and ( n46646 , n40611 , n41869 );
or ( n46647 , n46645 , n46646 );
not ( n46648 , n46647 );
not ( n46649 , n41869 );
and ( n46650 , n46649 , n34435 );
and ( n46651 , n40618 , n41869 );
or ( n46652 , n46650 , n46651 );
not ( n46653 , n46652 );
not ( n46654 , n41869 );
and ( n46655 , n46654 , n34437 );
and ( n46656 , n40625 , n41869 );
or ( n46657 , n46655 , n46656 );
not ( n46658 , n46657 );
not ( n46659 , n41869 );
and ( n46660 , n46659 , n34439 );
and ( n46661 , n40632 , n41869 );
or ( n46662 , n46660 , n46661 );
not ( n46663 , n46662 );
not ( n46664 , n41869 );
and ( n46665 , n46664 , n34441 );
and ( n46666 , n40639 , n41869 );
or ( n46667 , n46665 , n46666 );
not ( n46668 , n46667 );
not ( n46669 , n41869 );
and ( n46670 , n46669 , n34443 );
and ( n46671 , n40646 , n41869 );
or ( n46672 , n46670 , n46671 );
not ( n46673 , n46672 );
and ( n46674 , n46563 , n46594 );
and ( n46675 , n46673 , n46674 );
and ( n46676 , n46668 , n46675 );
and ( n46677 , n46663 , n46676 );
and ( n46678 , n46658 , n46677 );
and ( n46679 , n46653 , n46678 );
and ( n46680 , n46648 , n46679 );
and ( n46681 , n46643 , n46680 );
and ( n46682 , n46638 , n46681 );
and ( n46683 , n46633 , n46682 );
and ( n46684 , n46628 , n46683 );
and ( n46685 , n46623 , n46684 );
and ( n46686 , n46618 , n46685 );
and ( n46687 , n46613 , n46686 );
and ( n46688 , n46612 , n46687 );
xor ( n46689 , n46607 , n46688 );
buf ( n46690 , n41881 );
and ( n46691 , n46689 , n46690 );
buf ( n46692 , n46691 );
not ( n46693 , n46692 );
not ( n46694 , n46693 );
not ( n46695 , n46694 );
not ( n46696 , n41881 );
and ( n46697 , n46696 , n46611 );
xor ( n46698 , n46612 , n46687 );
and ( n46699 , n46698 , n41881 );
or ( n46700 , n46697 , n46699 );
not ( n46701 , n46700 );
buf ( n46702 , n46701 );
buf ( n46703 , n46702 );
not ( n46704 , n46703 );
not ( n46705 , n46704 );
not ( n46706 , n41881 );
and ( n46707 , n46706 , n44813 );
xor ( n46708 , n46613 , n46686 );
and ( n46709 , n46708 , n41881 );
or ( n46710 , n46707 , n46709 );
not ( n46711 , n46710 );
buf ( n46712 , n46711 );
buf ( n46713 , n46712 );
not ( n46714 , n46713 );
not ( n46715 , n46714 );
not ( n46716 , n41881 );
and ( n46717 , n46716 , n46617 );
xor ( n46718 , n46618 , n46685 );
and ( n46719 , n46718 , n41881 );
or ( n46720 , n46717 , n46719 );
not ( n46721 , n46720 );
buf ( n46722 , n46721 );
buf ( n46723 , n46722 );
not ( n46724 , n46723 );
not ( n46725 , n46724 );
not ( n46726 , n41881 );
and ( n46727 , n46726 , n46622 );
xor ( n46728 , n46623 , n46684 );
and ( n46729 , n46728 , n41881 );
or ( n46730 , n46727 , n46729 );
not ( n46731 , n46730 );
buf ( n46732 , n46731 );
buf ( n46733 , n46732 );
not ( n46734 , n46733 );
not ( n46735 , n46734 );
not ( n46736 , n41881 );
and ( n46737 , n46736 , n46627 );
xor ( n46738 , n46628 , n46683 );
and ( n46739 , n46738 , n41881 );
or ( n46740 , n46737 , n46739 );
not ( n46741 , n46740 );
buf ( n46742 , n46741 );
buf ( n46743 , n46742 );
not ( n46744 , n46743 );
not ( n46745 , n46744 );
not ( n46746 , n41881 );
and ( n46747 , n46746 , n46632 );
xor ( n46748 , n46633 , n46682 );
and ( n46749 , n46748 , n41881 );
or ( n46750 , n46747 , n46749 );
not ( n46751 , n46750 );
buf ( n46752 , n46751 );
buf ( n46753 , n46752 );
not ( n46754 , n46753 );
not ( n46755 , n46754 );
not ( n46756 , n41881 );
and ( n46757 , n46756 , n46637 );
xor ( n46758 , n46638 , n46681 );
and ( n46759 , n46758 , n41881 );
or ( n46760 , n46757 , n46759 );
not ( n46761 , n46760 );
buf ( n46762 , n46761 );
buf ( n46763 , n46762 );
not ( n46764 , n46763 );
not ( n46765 , n46764 );
not ( n46766 , n41881 );
and ( n46767 , n46766 , n46642 );
xor ( n46768 , n46643 , n46680 );
and ( n46769 , n46768 , n41881 );
or ( n46770 , n46767 , n46769 );
not ( n46771 , n46770 );
buf ( n46772 , n46771 );
buf ( n46773 , n46772 );
not ( n46774 , n46773 );
not ( n46775 , n46774 );
not ( n46776 , n41881 );
and ( n46777 , n46776 , n46647 );
xor ( n46778 , n46648 , n46679 );
and ( n46779 , n46778 , n41881 );
or ( n46780 , n46777 , n46779 );
not ( n46781 , n46780 );
buf ( n46782 , n46781 );
buf ( n46783 , n46782 );
not ( n46784 , n46783 );
not ( n46785 , n46784 );
not ( n46786 , n41881 );
and ( n46787 , n46786 , n46652 );
xor ( n46788 , n46653 , n46678 );
and ( n46789 , n46788 , n41881 );
or ( n46790 , n46787 , n46789 );
not ( n46791 , n46790 );
buf ( n46792 , n46791 );
buf ( n46793 , n46792 );
not ( n46794 , n46793 );
not ( n46795 , n46794 );
not ( n46796 , n41881 );
and ( n46797 , n46796 , n46657 );
xor ( n46798 , n46658 , n46677 );
and ( n46799 , n46798 , n41881 );
or ( n46800 , n46797 , n46799 );
not ( n46801 , n46800 );
buf ( n46802 , n46801 );
buf ( n46803 , n46802 );
not ( n46804 , n46803 );
not ( n46805 , n46804 );
not ( n46806 , n41881 );
and ( n46807 , n46806 , n46662 );
xor ( n46808 , n46663 , n46676 );
and ( n46809 , n46808 , n41881 );
or ( n46810 , n46807 , n46809 );
not ( n46811 , n46810 );
buf ( n46812 , n46811 );
buf ( n46813 , n46812 );
not ( n46814 , n46813 );
not ( n46815 , n46814 );
not ( n46816 , n41881 );
and ( n46817 , n46816 , n46667 );
xor ( n46818 , n46668 , n46675 );
and ( n46819 , n46818 , n41881 );
or ( n46820 , n46817 , n46819 );
not ( n46821 , n46820 );
buf ( n46822 , n46821 );
buf ( n46823 , n46822 );
not ( n46824 , n46823 );
not ( n46825 , n46824 );
not ( n46826 , n41881 );
and ( n46827 , n46826 , n46672 );
xor ( n46828 , n46673 , n46674 );
and ( n46829 , n46828 , n41881 );
or ( n46830 , n46827 , n46829 );
not ( n46831 , n46830 );
buf ( n46832 , n46831 );
buf ( n46833 , n46832 );
not ( n46834 , n46833 );
not ( n46835 , n46834 );
not ( n46836 , n46601 );
and ( n46837 , n46835 , n46836 );
and ( n46838 , n46825 , n46837 );
and ( n46839 , n46815 , n46838 );
and ( n46840 , n46805 , n46839 );
and ( n46841 , n46795 , n46840 );
and ( n46842 , n46785 , n46841 );
and ( n46843 , n46775 , n46842 );
and ( n46844 , n46765 , n46843 );
and ( n46845 , n46755 , n46844 );
and ( n46846 , n46745 , n46845 );
and ( n46847 , n46735 , n46846 );
and ( n46848 , n46725 , n46847 );
and ( n46849 , n46715 , n46848 );
and ( n46850 , n46705 , n46849 );
and ( n46851 , n46695 , n46850 );
not ( n46852 , n46851 );
and ( n46853 , n46852 , n41881 );
buf ( n46854 , n46853 );
not ( n46855 , n46854 );
not ( n46856 , n41881 );
and ( n46857 , n46856 , n46834 );
xor ( n46858 , n46835 , n46836 );
and ( n46859 , n46858 , n41881 );
or ( n46860 , n46857 , n46859 );
and ( n46861 , n46855 , n46860 );
not ( n46862 , n46860 );
not ( n46863 , n46602 );
xor ( n46864 , n46862 , n46863 );
and ( n46865 , n46864 , n46854 );
or ( n46866 , n46861 , n46865 );
not ( n46867 , n46866 );
buf ( n46868 , n46867 );
buf ( n46869 , n46868 );
not ( n46870 , n46869 );
or ( n46871 , n46606 , n46870 );
not ( n46872 , n46854 );
not ( n46873 , n41881 );
and ( n46874 , n46873 , n46824 );
xor ( n46875 , n46825 , n46837 );
and ( n46876 , n46875 , n41881 );
or ( n46877 , n46874 , n46876 );
and ( n46878 , n46872 , n46877 );
not ( n46879 , n46877 );
and ( n46880 , n46862 , n46863 );
xor ( n46881 , n46879 , n46880 );
and ( n46882 , n46881 , n46854 );
or ( n46883 , n46878 , n46882 );
not ( n46884 , n46883 );
buf ( n46885 , n46884 );
buf ( n46886 , n46885 );
not ( n46887 , n46886 );
or ( n46888 , n46871 , n46887 );
not ( n46889 , n46854 );
not ( n46890 , n41881 );
and ( n46891 , n46890 , n46814 );
xor ( n46892 , n46815 , n46838 );
and ( n46893 , n46892 , n41881 );
or ( n46894 , n46891 , n46893 );
and ( n46895 , n46889 , n46894 );
not ( n46896 , n46894 );
and ( n46897 , n46879 , n46880 );
xor ( n46898 , n46896 , n46897 );
and ( n46899 , n46898 , n46854 );
or ( n46900 , n46895 , n46899 );
not ( n46901 , n46900 );
buf ( n46902 , n46901 );
buf ( n46903 , n46902 );
not ( n46904 , n46903 );
or ( n46905 , n46888 , n46904 );
not ( n46906 , n46854 );
not ( n46907 , n41881 );
and ( n46908 , n46907 , n46804 );
xor ( n46909 , n46805 , n46839 );
and ( n46910 , n46909 , n41881 );
or ( n46911 , n46908 , n46910 );
and ( n46912 , n46906 , n46911 );
not ( n46913 , n46911 );
and ( n46914 , n46896 , n46897 );
xor ( n46915 , n46913 , n46914 );
and ( n46916 , n46915 , n46854 );
or ( n46917 , n46912 , n46916 );
not ( n46918 , n46917 );
buf ( n46919 , n46918 );
buf ( n46920 , n46919 );
not ( n46921 , n46920 );
or ( n46922 , n46905 , n46921 );
not ( n46923 , n46854 );
not ( n46924 , n41881 );
and ( n46925 , n46924 , n46794 );
xor ( n46926 , n46795 , n46840 );
and ( n46927 , n46926 , n41881 );
or ( n46928 , n46925 , n46927 );
and ( n46929 , n46923 , n46928 );
not ( n46930 , n46928 );
and ( n46931 , n46913 , n46914 );
xor ( n46932 , n46930 , n46931 );
and ( n46933 , n46932 , n46854 );
or ( n46934 , n46929 , n46933 );
not ( n46935 , n46934 );
buf ( n46936 , n46935 );
buf ( n46937 , n46936 );
not ( n46938 , n46937 );
or ( n46939 , n46922 , n46938 );
not ( n46940 , n46854 );
not ( n46941 , n41881 );
and ( n46942 , n46941 , n46784 );
xor ( n46943 , n46785 , n46841 );
and ( n46944 , n46943 , n41881 );
or ( n46945 , n46942 , n46944 );
and ( n46946 , n46940 , n46945 );
not ( n46947 , n46945 );
and ( n46948 , n46930 , n46931 );
xor ( n46949 , n46947 , n46948 );
and ( n46950 , n46949 , n46854 );
or ( n46951 , n46946 , n46950 );
not ( n46952 , n46951 );
buf ( n46953 , n46952 );
buf ( n46954 , n46953 );
not ( n46955 , n46954 );
or ( n46956 , n46939 , n46955 );
not ( n46957 , n46854 );
not ( n46958 , n41881 );
and ( n46959 , n46958 , n46774 );
xor ( n46960 , n46775 , n46842 );
and ( n46961 , n46960 , n41881 );
or ( n46962 , n46959 , n46961 );
and ( n46963 , n46957 , n46962 );
not ( n46964 , n46962 );
and ( n46965 , n46947 , n46948 );
xor ( n46966 , n46964 , n46965 );
and ( n46967 , n46966 , n46854 );
or ( n46968 , n46963 , n46967 );
not ( n46969 , n46968 );
buf ( n46970 , n46969 );
buf ( n46971 , n46970 );
not ( n46972 , n46971 );
or ( n46973 , n46956 , n46972 );
buf ( n46974 , n46973 );
buf ( n46975 , n46974 );
and ( n46976 , n46975 , n46854 );
not ( n46977 , n46976 );
and ( n46978 , n46977 , n46870 );
xor ( n46979 , n46870 , n46854 );
xor ( n46980 , n46606 , n46854 );
and ( n46981 , n46980 , n46854 );
xor ( n46982 , n46979 , n46981 );
and ( n46983 , n46982 , n46976 );
or ( n46984 , n46978 , n46983 );
and ( n46985 , n46984 , n46554 );
or ( n46986 , n46556 , n46985 );
and ( n46987 , n46551 , n46986 );
not ( n46988 , n41881 );
and ( n46989 , n46988 , n46637 );
not ( n46990 , n46637 );
not ( n46991 , n46642 );
not ( n46992 , n46647 );
not ( n46993 , n46652 );
not ( n46994 , n46657 );
not ( n46995 , n46662 );
not ( n46996 , n46667 );
not ( n46997 , n46672 );
not ( n46998 , n46561 );
not ( n46999 , n42110 );
not ( n47000 , n42094 );
not ( n47001 , n42078 );
not ( n47002 , n42062 );
not ( n47003 , n42046 );
not ( n47004 , n42030 );
not ( n47005 , n42014 );
not ( n47006 , n41998 );
not ( n47007 , n41982 );
not ( n47008 , n41966 );
not ( n47009 , n41950 );
not ( n47010 , n41934 );
not ( n47011 , n41918 );
not ( n47012 , n41902 );
not ( n47013 , n41886 );
not ( n47014 , n41873 );
and ( n47015 , n47013 , n47014 );
and ( n47016 , n47012 , n47015 );
and ( n47017 , n47011 , n47016 );
and ( n47018 , n47010 , n47017 );
and ( n47019 , n47009 , n47018 );
and ( n47020 , n47008 , n47019 );
and ( n47021 , n47007 , n47020 );
and ( n47022 , n47006 , n47021 );
and ( n47023 , n47005 , n47022 );
and ( n47024 , n47004 , n47023 );
and ( n47025 , n47003 , n47024 );
and ( n47026 , n47002 , n47025 );
and ( n47027 , n47001 , n47026 );
and ( n47028 , n47000 , n47027 );
and ( n47029 , n46999 , n47028 );
and ( n47030 , n46998 , n47029 );
and ( n47031 , n46997 , n47030 );
and ( n47032 , n46996 , n47031 );
and ( n47033 , n46995 , n47032 );
and ( n47034 , n46994 , n47033 );
and ( n47035 , n46993 , n47034 );
and ( n47036 , n46992 , n47035 );
and ( n47037 , n46991 , n47036 );
xor ( n47038 , n46990 , n47037 );
and ( n47039 , n47038 , n41881 );
or ( n47040 , n46989 , n47039 );
not ( n47041 , n47040 );
buf ( n47042 , n47041 );
buf ( n47043 , n47042 );
not ( n47044 , n47043 );
buf ( n47045 , n47044 );
buf ( n47046 , n47045 );
not ( n47047 , n47046 );
buf ( n47048 , n47047 );
not ( n47049 , n47048 );
not ( n47050 , n41881 );
not ( n47051 , n46611 );
not ( n47052 , n44813 );
not ( n47053 , n46617 );
not ( n47054 , n46622 );
not ( n47055 , n46627 );
not ( n47056 , n46632 );
and ( n47057 , n46990 , n47037 );
and ( n47058 , n47056 , n47057 );
and ( n47059 , n47055 , n47058 );
and ( n47060 , n47054 , n47059 );
and ( n47061 , n47053 , n47060 );
and ( n47062 , n47052 , n47061 );
and ( n47063 , n47051 , n47062 );
xor ( n47064 , n47050 , n47063 );
buf ( n47065 , n41881 );
and ( n47066 , n47064 , n47065 );
buf ( n47067 , n47066 );
not ( n47068 , n47067 );
not ( n47069 , n47068 );
not ( n47070 , n47069 );
not ( n47071 , n41881 );
and ( n47072 , n47071 , n46611 );
xor ( n47073 , n47051 , n47062 );
and ( n47074 , n47073 , n41881 );
or ( n47075 , n47072 , n47074 );
not ( n47076 , n47075 );
buf ( n47077 , n47076 );
buf ( n47078 , n47077 );
not ( n47079 , n47078 );
not ( n47080 , n47079 );
not ( n47081 , n41881 );
and ( n47082 , n47081 , n44813 );
xor ( n47083 , n47052 , n47061 );
and ( n47084 , n47083 , n41881 );
or ( n47085 , n47082 , n47084 );
not ( n47086 , n47085 );
buf ( n47087 , n47086 );
buf ( n47088 , n47087 );
not ( n47089 , n47088 );
not ( n47090 , n47089 );
not ( n47091 , n41881 );
and ( n47092 , n47091 , n46617 );
xor ( n47093 , n47053 , n47060 );
and ( n47094 , n47093 , n41881 );
or ( n47095 , n47092 , n47094 );
not ( n47096 , n47095 );
buf ( n47097 , n47096 );
buf ( n47098 , n47097 );
not ( n47099 , n47098 );
not ( n47100 , n47099 );
not ( n47101 , n41881 );
and ( n47102 , n47101 , n46622 );
xor ( n47103 , n47054 , n47059 );
and ( n47104 , n47103 , n41881 );
or ( n47105 , n47102 , n47104 );
not ( n47106 , n47105 );
buf ( n47107 , n47106 );
buf ( n47108 , n47107 );
not ( n47109 , n47108 );
not ( n47110 , n47109 );
not ( n47111 , n41881 );
and ( n47112 , n47111 , n46627 );
xor ( n47113 , n47055 , n47058 );
and ( n47114 , n47113 , n41881 );
or ( n47115 , n47112 , n47114 );
not ( n47116 , n47115 );
buf ( n47117 , n47116 );
buf ( n47118 , n47117 );
not ( n47119 , n47118 );
not ( n47120 , n47119 );
not ( n47121 , n41881 );
and ( n47122 , n47121 , n46632 );
xor ( n47123 , n47056 , n47057 );
and ( n47124 , n47123 , n41881 );
or ( n47125 , n47122 , n47124 );
not ( n47126 , n47125 );
buf ( n47127 , n47126 );
buf ( n47128 , n47127 );
not ( n47129 , n47128 );
not ( n47130 , n47129 );
not ( n47131 , n47044 );
and ( n47132 , n47130 , n47131 );
and ( n47133 , n47120 , n47132 );
and ( n47134 , n47110 , n47133 );
and ( n47135 , n47100 , n47134 );
and ( n47136 , n47090 , n47135 );
and ( n47137 , n47080 , n47136 );
and ( n47138 , n47070 , n47137 );
not ( n47139 , n47138 );
and ( n47140 , n47139 , n41881 );
buf ( n47141 , n47140 );
not ( n47142 , n47141 );
not ( n47143 , n41881 );
and ( n47144 , n47143 , n47129 );
xor ( n47145 , n47130 , n47131 );
and ( n47146 , n47145 , n41881 );
or ( n47147 , n47144 , n47146 );
and ( n47148 , n47142 , n47147 );
not ( n47149 , n47147 );
not ( n47150 , n47045 );
xor ( n47151 , n47149 , n47150 );
and ( n47152 , n47151 , n47141 );
or ( n47153 , n47148 , n47152 );
not ( n47154 , n47153 );
buf ( n47155 , n47154 );
buf ( n47156 , n47155 );
not ( n47157 , n47156 );
or ( n47158 , n47049 , n47157 );
not ( n47159 , n47141 );
not ( n47160 , n41881 );
and ( n47161 , n47160 , n47119 );
xor ( n47162 , n47120 , n47132 );
and ( n47163 , n47162 , n41881 );
or ( n47164 , n47161 , n47163 );
and ( n47165 , n47159 , n47164 );
not ( n47166 , n47164 );
and ( n47167 , n47149 , n47150 );
xor ( n47168 , n47166 , n47167 );
and ( n47169 , n47168 , n47141 );
or ( n47170 , n47165 , n47169 );
not ( n47171 , n47170 );
buf ( n47172 , n47171 );
buf ( n47173 , n47172 );
not ( n47174 , n47173 );
or ( n47175 , n47158 , n47174 );
not ( n47176 , n47141 );
not ( n47177 , n41881 );
and ( n47178 , n47177 , n47109 );
xor ( n47179 , n47110 , n47133 );
and ( n47180 , n47179 , n41881 );
or ( n47181 , n47178 , n47180 );
and ( n47182 , n47176 , n47181 );
not ( n47183 , n47181 );
and ( n47184 , n47166 , n47167 );
xor ( n47185 , n47183 , n47184 );
and ( n47186 , n47185 , n47141 );
or ( n47187 , n47182 , n47186 );
not ( n47188 , n47187 );
buf ( n47189 , n47188 );
buf ( n47190 , n47189 );
not ( n47191 , n47190 );
or ( n47192 , n47175 , n47191 );
not ( n47193 , n47141 );
not ( n47194 , n41881 );
and ( n47195 , n47194 , n47099 );
xor ( n47196 , n47100 , n47134 );
and ( n47197 , n47196 , n41881 );
or ( n47198 , n47195 , n47197 );
and ( n47199 , n47193 , n47198 );
not ( n47200 , n47198 );
and ( n47201 , n47183 , n47184 );
xor ( n47202 , n47200 , n47201 );
and ( n47203 , n47202 , n47141 );
or ( n47204 , n47199 , n47203 );
not ( n47205 , n47204 );
buf ( n47206 , n47205 );
buf ( n47207 , n47206 );
not ( n47208 , n47207 );
or ( n47209 , n47192 , n47208 );
not ( n47210 , n47141 );
not ( n47211 , n41881 );
and ( n47212 , n47211 , n47089 );
xor ( n47213 , n47090 , n47135 );
and ( n47214 , n47213 , n41881 );
or ( n47215 , n47212 , n47214 );
and ( n47216 , n47210 , n47215 );
not ( n47217 , n47215 );
and ( n47218 , n47200 , n47201 );
xor ( n47219 , n47217 , n47218 );
and ( n47220 , n47219 , n47141 );
or ( n47221 , n47216 , n47220 );
not ( n47222 , n47221 );
buf ( n47223 , n47222 );
buf ( n47224 , n47223 );
not ( n47225 , n47224 );
or ( n47226 , n47209 , n47225 );
not ( n47227 , n47141 );
not ( n47228 , n41881 );
and ( n47229 , n47228 , n47079 );
xor ( n47230 , n47080 , n47136 );
and ( n47231 , n47230 , n41881 );
or ( n47232 , n47229 , n47231 );
and ( n47233 , n47227 , n47232 );
not ( n47234 , n47232 );
and ( n47235 , n47217 , n47218 );
xor ( n47236 , n47234 , n47235 );
and ( n47237 , n47236 , n47141 );
or ( n47238 , n47233 , n47237 );
not ( n47239 , n47238 );
buf ( n47240 , n47239 );
buf ( n47241 , n47240 );
not ( n47242 , n47241 );
or ( n47243 , n47226 , n47242 );
xor ( n47244 , n47070 , n47137 );
and ( n47245 , n47244 , n41881 );
buf ( n47246 , n47245 );
not ( n47247 , n47246 );
and ( n47248 , n47234 , n47235 );
xor ( n47249 , n47247 , n47248 );
and ( n47250 , n47249 , n47141 );
buf ( n47251 , n47250 );
not ( n47252 , n47251 );
buf ( n47253 , n47252 );
buf ( n47254 , n47253 );
not ( n47255 , n47254 );
or ( n47256 , n47243 , n47255 );
buf ( n47257 , n47256 );
buf ( n47258 , n47257 );
and ( n47259 , n47258 , n47141 );
not ( n47260 , n47259 );
and ( n47261 , n47260 , n47157 );
xor ( n47262 , n47157 , n47141 );
xor ( n47263 , n47049 , n47141 );
and ( n47264 , n47263 , n47141 );
xor ( n47265 , n47262 , n47264 );
and ( n47266 , n47265 , n47259 );
or ( n47267 , n47261 , n47266 );
and ( n47268 , n47267 , n46550 );
or ( n47269 , n46987 , n47268 );
and ( n47270 , n47269 , n31452 );
or ( n47271 , n46511 , n47270 );
and ( n47272 , n47271 , n31638 );
or ( n47273 , n40147 , n31641 );
or ( n47274 , n47273 , n31557 );
or ( n47275 , n47274 , n31645 );
or ( n47276 , n47275 , n31647 );
or ( n47277 , n47276 , n31007 );
and ( n47278 , n31146 , n47277 );
or ( n47279 , C0 , n46369 , n46501 , n47272 , n47278 );
buf ( n47280 , n47279 );
buf ( n47281 , n47280 );
buf ( n47282 , n31655 );
buf ( n47283 , RI15b62100_1211);
buf ( n47284 , RI15b62088_1210);
buf ( n47285 , RI15b62010_1209);
buf ( n47286 , RI15b61f98_1208);
buf ( n47287 , RI15b61f20_1207);
buf ( n47288 , RI15b61ea8_1206);
buf ( n47289 , RI15b61e30_1205);
buf ( n47290 , RI15b61db8_1204);
and ( n47291 , n45999 , n35297 );
and ( n47292 , n45984 , n47291 );
and ( n47293 , n47290 , n47292 );
and ( n47294 , n47289 , n47293 );
and ( n47295 , n47288 , n47294 );
and ( n47296 , n47287 , n47295 );
and ( n47297 , n47286 , n47296 );
and ( n47298 , n47285 , n47297 );
and ( n47299 , n47284 , n47298 );
xor ( n47300 , n47283 , n47299 );
and ( n47301 , n47300 , n32433 );
not ( n47302 , n31689 );
buf ( n47303 , n31689 );
buf ( n47304 , n31689 );
buf ( n47305 , n31689 );
buf ( n47306 , n31689 );
buf ( n47307 , n31689 );
buf ( n47308 , n31689 );
buf ( n47309 , n31689 );
buf ( n47310 , n31689 );
buf ( n47311 , n31689 );
buf ( n47312 , n31689 );
buf ( n47313 , n31689 );
buf ( n47314 , n31689 );
buf ( n47315 , n31689 );
buf ( n47316 , n31689 );
buf ( n47317 , n31689 );
buf ( n47318 , n31689 );
buf ( n47319 , n31689 );
buf ( n47320 , n31689 );
buf ( n47321 , n31689 );
buf ( n47322 , n31689 );
buf ( n47323 , n31689 );
buf ( n47324 , n31689 );
buf ( n47325 , n31689 );
buf ( n47326 , n31689 );
buf ( n47327 , n31689 );
or ( n47328 , n31723 , n31724 );
and ( n47329 , n31721 , n47328 );
or ( n47330 , n31692 , n31694 , n31689 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47329 );
and ( n47331 , n47302 , n47330 );
not ( n47332 , n47331 );
and ( n47333 , n47332 , n47283 );
not ( n47334 , n31674 );
buf ( n47335 , n47334 );
not ( n47336 , n47335 );
not ( n47337 , n47336 );
not ( n47338 , n31670 );
not ( n47339 , n47338 );
buf ( n47340 , n47339 );
buf ( n47341 , n47340 );
not ( n47342 , n47341 );
not ( n47343 , n47342 );
xor ( n47344 , n31666 , n31670 );
not ( n47345 , n47344 );
buf ( n47346 , n47345 );
buf ( n47347 , n47346 );
not ( n47348 , n47347 );
not ( n47349 , n47348 );
and ( n47350 , n31666 , n31670 );
xor ( n47351 , n31662 , n47350 );
not ( n47352 , n47351 );
buf ( n47353 , n47352 );
buf ( n47354 , n47353 );
not ( n47355 , n47354 );
not ( n47356 , n47355 );
nor ( n47357 , n47337 , n47343 , n47349 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47358 , n31966 , n47357 );
nor ( n47359 , n47336 , n47343 , n47349 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47360 , n31968 , n47359 );
nor ( n47361 , n47337 , n47342 , n47349 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47362 , n31970 , n47361 );
nor ( n47363 , n47336 , n47342 , n47349 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47364 , n31972 , n47363 );
nor ( n47365 , n47337 , n47343 , n47348 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47366 , n31974 , n47365 );
nor ( n47367 , n47336 , n47343 , n47348 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47368 , n31976 , n47367 );
nor ( n47369 , n47337 , n47342 , n47348 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47370 , n31978 , n47369 );
nor ( n47371 , n47336 , n47342 , n47348 , n47356 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47372 , n31980 , n47371 );
nor ( n47373 , n47337 , n47343 , n47349 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47374 , n31982 , n47373 );
nor ( n47375 , n47336 , n47343 , n47349 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47376 , n31984 , n47375 );
nor ( n47377 , n47337 , n47342 , n47349 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47378 , n31986 , n47377 );
nor ( n47379 , n47336 , n47342 , n47349 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47380 , n31988 , n47379 );
nor ( n47381 , n47337 , n47343 , n47348 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47382 , n31990 , n47381 );
nor ( n47383 , n47336 , n47343 , n47348 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47384 , n31992 , n47383 );
nor ( n47385 , n47337 , n47342 , n47348 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47386 , n31994 , n47385 );
nor ( n47387 , n47336 , n47342 , n47348 , n47355 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n47388 , n31996 , n47387 );
or ( n47389 , n47358 , n47360 , n47362 , n47364 , n47366 , n47368 , n47370 , n47372 , n47374 , n47376 , n47378 , n47380 , n47382 , n47384 , n47386 , n47388 );
and ( n47390 , n47389 , n47331 );
or ( n47391 , n47333 , n47390 );
and ( n47392 , n47391 , n32413 );
or ( n47393 , n35346 , n32415 );
or ( n47394 , n47393 , n32417 );
or ( n47395 , n47394 , n32419 );
or ( n47396 , n47395 , n32421 );
or ( n47397 , n47396 , n32423 );
or ( n47398 , n47397 , n32425 );
or ( n47399 , n47398 , n32427 );
or ( n47400 , n47399 , n32429 );
or ( n47401 , n47400 , n32431 );
or ( n47402 , n47401 , n32435 );
and ( n47403 , n47283 , n47402 );
or ( n47404 , n47301 , n47392 , n47403 );
and ( n47405 , n47404 , n32456 );
or ( n47406 , n46346 , n32494 );
or ( n47407 , n47406 , n32496 );
or ( n47408 , n47407 , n32498 );
or ( n47409 , n47408 , n32500 );
and ( n47410 , n47283 , n47409 );
or ( n47411 , C0 , n47405 , n47410 );
buf ( n47412 , n47411 );
buf ( n47413 , n47412 );
not ( n47414 , n35542 );
and ( n47415 , n47414 , n41847 );
buf ( n47416 , RI15b45438_228);
and ( n47417 , n47416 , n35542 );
or ( n47418 , n47415 , n47417 );
buf ( n47419 , n47418 );
buf ( n47420 , n47419 );
not ( n47421 , n46356 );
and ( n47422 , n47421 , n31333 );
nor ( n47423 , n31025 , n46360 , n31017 , n31013 , n31009 );
not ( n47424 , n47423 );
and ( n47425 , n47424 , n31333 );
and ( n47426 , n31339 , n47423 );
or ( n47427 , n47425 , n47426 );
and ( n47428 , n47427 , n46356 );
or ( n47429 , n47422 , n47428 );
and ( n47430 , n47429 , n31649 );
nor ( n47431 , n46373 , n46380 , n46386 , n46392 , C0 );
not ( n47432 , n47431 );
not ( n47433 , n47423 );
and ( n47434 , n47433 , n31333 );
not ( n47435 , n46487 );
and ( n47436 , n47435 , n46471 );
xor ( n47437 , n46471 , n41881 );
xor ( n47438 , n46459 , n41881 );
xor ( n47439 , n46447 , n41881 );
xor ( n47440 , n46435 , n41881 );
xor ( n47441 , n46423 , n41881 );
and ( n47442 , n46490 , n46492 );
and ( n47443 , n47441 , n47442 );
and ( n47444 , n47440 , n47443 );
and ( n47445 , n47439 , n47444 );
and ( n47446 , n47438 , n47445 );
xor ( n47447 , n47437 , n47446 );
and ( n47448 , n47447 , n46487 );
or ( n47449 , n47436 , n47448 );
and ( n47450 , n47449 , n47423 );
or ( n47451 , n47434 , n47450 );
and ( n47452 , n47432 , n47451 );
and ( n47453 , n47449 , n47431 );
or ( n47454 , n47452 , n47453 );
and ( n47455 , n47454 , n31643 );
not ( n47456 , n31452 );
not ( n47457 , n47431 );
not ( n47458 , n47423 );
and ( n47459 , n47458 , n31333 );
and ( n47460 , n47449 , n47423 );
or ( n47461 , n47459 , n47460 );
and ( n47462 , n47457 , n47461 );
and ( n47463 , n47449 , n47431 );
or ( n47464 , n47462 , n47463 );
and ( n47465 , n47456 , n47464 );
nor ( n47466 , n46519 , n46529 , n46539 , n46549 , C0 );
not ( n47467 , n47466 );
nor ( n47468 , n46515 , n46553 , n46534 , n46544 , C0 );
not ( n47469 , n47468 );
and ( n47470 , n47469 , n47464 );
not ( n47471 , n46976 );
and ( n47472 , n47471 , n46955 );
xor ( n47473 , n46955 , n46854 );
xor ( n47474 , n46938 , n46854 );
xor ( n47475 , n46921 , n46854 );
xor ( n47476 , n46904 , n46854 );
xor ( n47477 , n46887 , n46854 );
and ( n47478 , n46979 , n46981 );
and ( n47479 , n47477 , n47478 );
and ( n47480 , n47476 , n47479 );
and ( n47481 , n47475 , n47480 );
and ( n47482 , n47474 , n47481 );
xor ( n47483 , n47473 , n47482 );
and ( n47484 , n47483 , n46976 );
or ( n47485 , n47472 , n47484 );
and ( n47486 , n47485 , n47468 );
or ( n47487 , n47470 , n47486 );
and ( n47488 , n47467 , n47487 );
not ( n47489 , n47259 );
and ( n47490 , n47489 , n47242 );
xor ( n47491 , n47242 , n47141 );
xor ( n47492 , n47225 , n47141 );
xor ( n47493 , n47208 , n47141 );
xor ( n47494 , n47191 , n47141 );
xor ( n47495 , n47174 , n47141 );
and ( n47496 , n47262 , n47264 );
and ( n47497 , n47495 , n47496 );
and ( n47498 , n47494 , n47497 );
and ( n47499 , n47493 , n47498 );
and ( n47500 , n47492 , n47499 );
xor ( n47501 , n47491 , n47500 );
and ( n47502 , n47501 , n47259 );
or ( n47503 , n47490 , n47502 );
and ( n47504 , n47503 , n47466 );
or ( n47505 , n47488 , n47504 );
and ( n47506 , n47505 , n31452 );
or ( n47507 , n47465 , n47506 );
and ( n47508 , n47507 , n31638 );
and ( n47509 , n31333 , n47277 );
or ( n47510 , C0 , n47430 , n47455 , n47508 , n47509 );
buf ( n47511 , n47510 );
buf ( n47512 , n47511 );
buf ( n47513 , n31655 );
buf ( n47514 , n31655 );
buf ( n47515 , n30987 );
buf ( n47516 , n31655 );
buf ( n47517 , RI15b477d8_304);
buf ( n47518 , n47517 );
not ( n47519 , n34150 );
and ( n47520 , n47519 , n32737 );
not ( n47521 , n41392 );
and ( n47522 , n47521 , n32737 );
and ( n47523 , n32755 , n41392 );
or ( n47524 , n47522 , n47523 );
and ( n47525 , n47524 , n34150 );
or ( n47526 , n47520 , n47525 );
and ( n47527 , n47526 , n33381 );
not ( n47528 , n41402 );
not ( n47529 , n41392 );
and ( n47530 , n47529 , n32737 );
and ( n47531 , n35083 , n41392 );
or ( n47532 , n47530 , n47531 );
and ( n47533 , n47528 , n47532 );
and ( n47534 , n35083 , n41402 );
or ( n47535 , n47533 , n47534 );
and ( n47536 , n47535 , n33375 );
not ( n47537 , n32968 );
not ( n47538 , n41402 );
not ( n47539 , n41392 );
and ( n47540 , n47539 , n32737 );
and ( n47541 , n35083 , n41392 );
or ( n47542 , n47540 , n47541 );
and ( n47543 , n47538 , n47542 );
and ( n47544 , n35083 , n41402 );
or ( n47545 , n47543 , n47544 );
and ( n47546 , n47537 , n47545 );
not ( n47547 , n41424 );
not ( n47548 , n41428 );
and ( n47549 , n47548 , n47545 );
and ( n47550 , n35107 , n41428 );
or ( n47551 , n47549 , n47550 );
and ( n47552 , n47547 , n47551 );
and ( n47553 , n35115 , n41424 );
or ( n47554 , n47552 , n47553 );
and ( n47555 , n47554 , n32968 );
or ( n47556 , n47546 , n47555 );
and ( n47557 , n47556 , n33370 );
and ( n47558 , n32737 , n35062 );
or ( n47559 , C0 , n47527 , n47536 , n47557 , n47558 );
buf ( n47560 , n47559 );
buf ( n47561 , n47560 );
buf ( n47562 , n31655 );
buf ( n47563 , n30987 );
buf ( n47564 , n30987 );
not ( n47565 , n31728 );
and ( n47566 , n47565 , n46022 );
buf ( n47567 , RI15b5cf70_1037);
buf ( n47568 , RI15b5cef8_1036);
buf ( n47569 , RI15b5ce80_1035);
buf ( n47570 , RI15b5ce08_1034);
buf ( n47571 , RI15b5cd90_1033);
buf ( n47572 , RI15b5cd18_1032);
buf ( n47573 , RI15b5cca0_1031);
buf ( n47574 , RI15b5cc28_1030);
buf ( n47575 , RI15b5cbb0_1029);
buf ( n47576 , RI15b5cb38_1028);
buf ( n47577 , RI15b5cac0_1027);
buf ( n47578 , RI15b5ca48_1026);
buf ( n47579 , RI15b5c9d0_1025);
buf ( n47580 , RI15b5c958_1024);
buf ( n47581 , RI15b5c8e0_1023);
buf ( n47582 , RI15b5c868_1022);
and ( n47583 , n41286 , n41287 );
and ( n47584 , n47582 , n47583 );
and ( n47585 , n47581 , n47584 );
and ( n47586 , n47580 , n47585 );
and ( n47587 , n47579 , n47586 );
and ( n47588 , n47578 , n47587 );
and ( n47589 , n47577 , n47588 );
and ( n47590 , n47576 , n47589 );
and ( n47591 , n47575 , n47590 );
and ( n47592 , n47574 , n47591 );
and ( n47593 , n47573 , n47592 );
and ( n47594 , n47572 , n47593 );
and ( n47595 , n47571 , n47594 );
and ( n47596 , n47570 , n47595 );
and ( n47597 , n47569 , n47596 );
and ( n47598 , n47568 , n47597 );
xor ( n47599 , n47567 , n47598 );
xor ( n47600 , n47568 , n47597 );
xor ( n47601 , n47569 , n47596 );
xor ( n47602 , n47570 , n47595 );
xor ( n47603 , n47571 , n47594 );
xor ( n47604 , n47572 , n47593 );
xor ( n47605 , n47573 , n47592 );
xor ( n47606 , n47574 , n47591 );
xor ( n47607 , n47575 , n47590 );
xor ( n47608 , n47576 , n47589 );
xor ( n47609 , n47577 , n47588 );
xor ( n47610 , n47578 , n47587 );
xor ( n47611 , n47579 , n47586 );
xor ( n47612 , n47580 , n47585 );
xor ( n47613 , n47581 , n47584 );
xor ( n47614 , n47582 , n47583 );
and ( n47615 , n41288 , n41289 );
and ( n47616 , n47614 , n47615 );
and ( n47617 , n47613 , n47616 );
and ( n47618 , n47612 , n47617 );
and ( n47619 , n47611 , n47618 );
and ( n47620 , n47610 , n47619 );
and ( n47621 , n47609 , n47620 );
and ( n47622 , n47608 , n47621 );
and ( n47623 , n47607 , n47622 );
and ( n47624 , n47606 , n47623 );
and ( n47625 , n47605 , n47624 );
and ( n47626 , n47604 , n47625 );
and ( n47627 , n47603 , n47626 );
and ( n47628 , n47602 , n47627 );
and ( n47629 , n47601 , n47628 );
and ( n47630 , n47600 , n47629 );
xor ( n47631 , n47599 , n47630 );
and ( n47632 , n47631 , n31728 );
or ( n47633 , n47566 , n47632 );
and ( n47634 , n47633 , n32253 );
not ( n47635 , n32283 );
and ( n47636 , n47635 , n46022 );
not ( n47637 , n31823 );
and ( n47638 , n41286 , n41297 );
and ( n47639 , n47582 , n47638 );
and ( n47640 , n47581 , n47639 );
and ( n47641 , n47580 , n47640 );
and ( n47642 , n47579 , n47641 );
and ( n47643 , n47578 , n47642 );
and ( n47644 , n47577 , n47643 );
and ( n47645 , n47576 , n47644 );
and ( n47646 , n47575 , n47645 );
and ( n47647 , n47574 , n47646 );
and ( n47648 , n47573 , n47647 );
and ( n47649 , n47572 , n47648 );
and ( n47650 , n47571 , n47649 );
and ( n47651 , n47570 , n47650 );
and ( n47652 , n47569 , n47651 );
and ( n47653 , n47568 , n47652 );
xor ( n47654 , n47567 , n47653 );
xor ( n47655 , n47568 , n47652 );
xor ( n47656 , n47569 , n47651 );
xor ( n47657 , n47570 , n47650 );
xor ( n47658 , n47571 , n47649 );
xor ( n47659 , n47572 , n47648 );
xor ( n47660 , n47573 , n47647 );
xor ( n47661 , n47574 , n47646 );
xor ( n47662 , n47575 , n47645 );
xor ( n47663 , n47576 , n47644 );
xor ( n47664 , n47577 , n47643 );
xor ( n47665 , n47578 , n47642 );
xor ( n47666 , n47579 , n47641 );
xor ( n47667 , n47580 , n47640 );
xor ( n47668 , n47581 , n47639 );
xor ( n47669 , n47582 , n47638 );
and ( n47670 , n41298 , n41299 );
and ( n47671 , n47669 , n47670 );
and ( n47672 , n47668 , n47671 );
and ( n47673 , n47667 , n47672 );
and ( n47674 , n47666 , n47673 );
and ( n47675 , n47665 , n47674 );
and ( n47676 , n47664 , n47675 );
and ( n47677 , n47663 , n47676 );
and ( n47678 , n47662 , n47677 );
and ( n47679 , n47661 , n47678 );
and ( n47680 , n47660 , n47679 );
and ( n47681 , n47659 , n47680 );
and ( n47682 , n47658 , n47681 );
and ( n47683 , n47657 , n47682 );
and ( n47684 , n47656 , n47683 );
and ( n47685 , n47655 , n47684 );
xor ( n47686 , n47654 , n47685 );
and ( n47687 , n47637 , n47686 );
and ( n47688 , n41286 , n41302 );
and ( n47689 , n47582 , n47688 );
and ( n47690 , n47581 , n47689 );
and ( n47691 , n47580 , n47690 );
and ( n47692 , n47579 , n47691 );
and ( n47693 , n47578 , n47692 );
and ( n47694 , n47577 , n47693 );
and ( n47695 , n47576 , n47694 );
and ( n47696 , n47575 , n47695 );
and ( n47697 , n47574 , n47696 );
and ( n47698 , n47573 , n47697 );
and ( n47699 , n47572 , n47698 );
and ( n47700 , n47571 , n47699 );
and ( n47701 , n47570 , n47700 );
and ( n47702 , n47569 , n47701 );
and ( n47703 , n47568 , n47702 );
xor ( n47704 , n47567 , n47703 );
xor ( n47705 , n47568 , n47702 );
xor ( n47706 , n47569 , n47701 );
xor ( n47707 , n47570 , n47700 );
xor ( n47708 , n47571 , n47699 );
xor ( n47709 , n47572 , n47698 );
xor ( n47710 , n47573 , n47697 );
xor ( n47711 , n47574 , n47696 );
xor ( n47712 , n47575 , n47695 );
xor ( n47713 , n47576 , n47694 );
xor ( n47714 , n47577 , n47693 );
xor ( n47715 , n47578 , n47692 );
xor ( n47716 , n47579 , n47691 );
xor ( n47717 , n47580 , n47690 );
xor ( n47718 , n47581 , n47689 );
xor ( n47719 , n47582 , n47688 );
or ( n47720 , n41303 , n41304 );
or ( n47721 , n47719 , n47720 );
or ( n47722 , n47718 , n47721 );
or ( n47723 , n47717 , n47722 );
or ( n47724 , n47716 , n47723 );
or ( n47725 , n47715 , n47724 );
or ( n47726 , n47714 , n47725 );
or ( n47727 , n47713 , n47726 );
or ( n47728 , n47712 , n47727 );
or ( n47729 , n47711 , n47728 );
or ( n47730 , n47710 , n47729 );
or ( n47731 , n47709 , n47730 );
or ( n47732 , n47708 , n47731 );
or ( n47733 , n47707 , n47732 );
or ( n47734 , n47706 , n47733 );
or ( n47735 , n47705 , n47734 );
xnor ( n47736 , n47704 , n47735 );
and ( n47737 , n47736 , n31823 );
or ( n47738 , n47687 , n47737 );
and ( n47739 , n47738 , n32283 );
or ( n47740 , n47636 , n47739 );
and ( n47741 , n47740 , n32398 );
and ( n47742 , n46022 , n32436 );
or ( n47743 , n47634 , n47741 , n47742 );
and ( n47744 , n47743 , n32456 );
xor ( n47745 , n46022 , n46053 );
and ( n47746 , n47745 , n32473 );
not ( n47747 , n32475 );
and ( n47748 , n47747 , n47745 );
and ( n47749 , n41284 , n41319 );
and ( n47750 , n46037 , n47749 );
and ( n47751 , n46036 , n47750 );
and ( n47752 , n46035 , n47751 );
and ( n47753 , n46034 , n47752 );
and ( n47754 , n46033 , n47753 );
and ( n47755 , n46032 , n47754 );
and ( n47756 , n46031 , n47755 );
and ( n47757 , n46030 , n47756 );
and ( n47758 , n46029 , n47757 );
and ( n47759 , n46028 , n47758 );
and ( n47760 , n46027 , n47759 );
and ( n47761 , n46026 , n47760 );
and ( n47762 , n46025 , n47761 );
and ( n47763 , n46024 , n47762 );
and ( n47764 , n46023 , n47763 );
xor ( n47765 , n46022 , n47764 );
and ( n47766 , n47765 , n32475 );
or ( n47767 , n47748 , n47766 );
and ( n47768 , n47767 , n32486 );
and ( n47769 , n37541 , n32489 );
and ( n47770 , n46022 , n32501 );
or ( n47771 , C0 , n47744 , n47746 , n47768 , n47769 , n47770 );
buf ( n47772 , n47771 );
buf ( n47773 , n47772 );
and ( n47774 , n33228 , n32528 );
not ( n47775 , n32598 );
and ( n47776 , n47775 , n32991 );
buf ( n47777 , n47776 );
and ( n47778 , n47777 , n32890 );
not ( n47779 , n32919 );
and ( n47780 , n47779 , n32991 );
buf ( n47781 , n47780 );
and ( n47782 , n47781 , n32924 );
not ( n47783 , n32953 );
and ( n47784 , n47783 , n32991 );
not ( n47785 , n32971 );
and ( n47786 , n47785 , n33107 );
xor ( n47787 , n32991 , n33014 );
and ( n47788 , n47787 , n32971 );
or ( n47789 , n47786 , n47788 );
and ( n47790 , n47789 , n32953 );
or ( n47791 , n47784 , n47790 );
and ( n47792 , n47791 , n33038 );
not ( n47793 , n33067 );
and ( n47794 , n47793 , n32991 );
not ( n47795 , n32970 );
not ( n47796 , n33071 );
and ( n47797 , n47796 , n33107 );
xor ( n47798 , n33108 , n33146 );
and ( n47799 , n47798 , n33071 );
or ( n47800 , n47797 , n47799 );
and ( n47801 , n47795 , n47800 );
and ( n47802 , n47787 , n32970 );
or ( n47803 , n47801 , n47802 );
and ( n47804 , n47803 , n33067 );
or ( n47805 , n47794 , n47804 );
and ( n47806 , n47805 , n33172 );
and ( n47807 , n32991 , n33204 );
or ( n47808 , n47778 , n47782 , n47792 , n47806 , n47807 );
and ( n47809 , n47808 , n33208 );
not ( n47810 , n32968 );
not ( n47811 , n33270 );
and ( n47812 , n47811 , n33307 );
xor ( n47813 , n33308 , n33346 );
and ( n47814 , n47813 , n33270 );
or ( n47815 , n47812 , n47814 );
and ( n47816 , n47810 , n47815 );
and ( n47817 , n32991 , n32968 );
or ( n47818 , n47816 , n47817 );
and ( n47819 , n47818 , n33370 );
buf ( n47820 , n35056 );
and ( n47821 , n32991 , n33382 );
or ( n47822 , C0 , n47774 , n47809 , n47819 , n47820 , n47821 );
buf ( n47823 , n47822 );
buf ( n47824 , n47823 );
buf ( n47825 , n30987 );
buf ( n47826 , n31655 );
buf ( n47827 , n31655 );
buf ( n47828 , n30987 );
not ( n47829 , n46356 );
and ( n47830 , n47829 , n31342 );
and ( n47831 , n46359 , n31021 , n31017 , n31013 , n46361 );
not ( n47832 , n47831 );
and ( n47833 , n47832 , n31342 );
and ( n47834 , n31372 , n47831 );
or ( n47835 , n47833 , n47834 );
and ( n47836 , n47835 , n46356 );
or ( n47837 , n47830 , n47836 );
and ( n47838 , n47837 , n31649 );
and ( n47839 , n46374 , n46379 , n46386 , n46392 , C1 );
not ( n47840 , n47839 );
not ( n47841 , n47831 );
and ( n47842 , n47841 , n31342 );
not ( n47843 , n46487 );
and ( n47844 , n47843 , n46483 );
xor ( n47845 , n46483 , n41881 );
and ( n47846 , n47437 , n47446 );
xor ( n47847 , n47845 , n47846 );
and ( n47848 , n47847 , n46487 );
or ( n47849 , n47844 , n47848 );
and ( n47850 , n47849 , n47831 );
or ( n47851 , n47842 , n47850 );
and ( n47852 , n47840 , n47851 );
and ( n47853 , n47849 , n47839 );
or ( n47854 , n47852 , n47853 );
and ( n47855 , n47854 , n31643 );
not ( n47856 , n31452 );
not ( n47857 , n47839 );
not ( n47858 , n47831 );
and ( n47859 , n47858 , n31342 );
and ( n47860 , n47849 , n47831 );
or ( n47861 , n47859 , n47860 );
and ( n47862 , n47857 , n47861 );
and ( n47863 , n47849 , n47839 );
or ( n47864 , n47862 , n47863 );
and ( n47865 , n47856 , n47864 );
and ( n47866 , n46520 , n46528 , n46539 , n46549 , C1 );
not ( n47867 , n47866 );
and ( n47868 , n46552 , n46524 , n46534 , n46544 , C1 );
not ( n47869 , n47868 );
and ( n47870 , n47869 , n47864 );
not ( n47871 , n46976 );
and ( n47872 , n47871 , n46972 );
xor ( n47873 , n46972 , n46854 );
and ( n47874 , n47473 , n47482 );
xor ( n47875 , n47873 , n47874 );
and ( n47876 , n47875 , n46976 );
or ( n47877 , n47872 , n47876 );
and ( n47878 , n47877 , n47868 );
or ( n47879 , n47870 , n47878 );
and ( n47880 , n47867 , n47879 );
not ( n47881 , n47259 );
and ( n47882 , n47881 , n47255 );
xor ( n47883 , n47255 , n47141 );
and ( n47884 , n47491 , n47500 );
xor ( n47885 , n47883 , n47884 );
and ( n47886 , n47885 , n47259 );
or ( n47887 , n47882 , n47886 );
and ( n47888 , n47887 , n47866 );
or ( n47889 , n47880 , n47888 );
and ( n47890 , n47889 , n31452 );
or ( n47891 , n47865 , n47890 );
and ( n47892 , n47891 , n31638 );
and ( n47893 , n31342 , n47277 );
or ( n47894 , C0 , n47838 , n47855 , n47892 , n47893 );
buf ( n47895 , n47894 );
buf ( n47896 , n47895 );
buf ( n47897 , n31655 );
buf ( n47898 , n30987 );
not ( n47899 , n35278 );
buf ( n47900 , RI15b5f388_1114);
and ( n47901 , n47899 , n47900 );
not ( n47902 , n46290 );
and ( n47903 , n47902 , n46182 );
xor ( n47904 , n46299 , n46313 );
and ( n47905 , n47904 , n46290 );
or ( n47906 , n47903 , n47905 );
and ( n47907 , n47906 , n35278 );
or ( n47908 , n47901 , n47907 );
and ( n47909 , n47908 , n32417 );
or ( n47910 , n32475 , n35292 );
and ( n47911 , n35292 , n47910 );
and ( n47912 , n35331 , n47911 );
not ( n47913 , n47912 );
and ( n47914 , n47913 , n47900 );
buf ( n47915 , n40234 );
not ( n47916 , n47915 );
buf ( n47917 , n47916 );
not ( n47918 , n47917 );
not ( n47919 , n40244 );
and ( n47920 , n47919 , n40251 );
not ( n47921 , n40251 );
not ( n47922 , n40234 );
xor ( n47923 , n47921 , n47922 );
and ( n47924 , n47923 , n40244 );
or ( n47925 , n47920 , n47924 );
not ( n47926 , n47925 );
buf ( n47927 , n47926 );
buf ( n47928 , n47927 );
not ( n47929 , n47928 );
or ( n47930 , n47918 , n47929 );
not ( n47931 , n40244 );
and ( n47932 , n47931 , n40269 );
not ( n47933 , n40269 );
and ( n47934 , n47921 , n47922 );
xor ( n47935 , n47933 , n47934 );
and ( n47936 , n47935 , n40244 );
or ( n47937 , n47932 , n47936 );
not ( n47938 , n47937 );
buf ( n47939 , n47938 );
buf ( n47940 , n47939 );
not ( n47941 , n47940 );
or ( n47942 , n47930 , n47941 );
not ( n47943 , n40244 );
and ( n47944 , n47943 , n40287 );
not ( n47945 , n40287 );
and ( n47946 , n47933 , n47934 );
xor ( n47947 , n47945 , n47946 );
and ( n47948 , n47947 , n40244 );
or ( n47949 , n47944 , n47948 );
not ( n47950 , n47949 );
buf ( n47951 , n47950 );
buf ( n47952 , n47951 );
not ( n47953 , n47952 );
or ( n47954 , n47942 , n47953 );
not ( n47955 , n40244 );
and ( n47956 , n47955 , n40305 );
not ( n47957 , n40305 );
and ( n47958 , n47945 , n47946 );
xor ( n47959 , n47957 , n47958 );
and ( n47960 , n47959 , n40244 );
or ( n47961 , n47956 , n47960 );
not ( n47962 , n47961 );
buf ( n47963 , n47962 );
buf ( n47964 , n47963 );
not ( n47965 , n47964 );
or ( n47966 , n47954 , n47965 );
not ( n47967 , n40244 );
and ( n47968 , n47967 , n40323 );
not ( n47969 , n40323 );
and ( n47970 , n47957 , n47958 );
xor ( n47971 , n47969 , n47970 );
and ( n47972 , n47971 , n40244 );
or ( n47973 , n47968 , n47972 );
not ( n47974 , n47973 );
buf ( n47975 , n47974 );
buf ( n47976 , n47975 );
not ( n47977 , n47976 );
or ( n47978 , n47966 , n47977 );
not ( n47979 , n40244 );
and ( n47980 , n47979 , n40341 );
not ( n47981 , n40341 );
and ( n47982 , n47969 , n47970 );
xor ( n47983 , n47981 , n47982 );
and ( n47984 , n47983 , n40244 );
or ( n47985 , n47980 , n47984 );
not ( n47986 , n47985 );
buf ( n47987 , n47986 );
buf ( n47988 , n47987 );
not ( n47989 , n47988 );
or ( n47990 , n47978 , n47989 );
not ( n47991 , n40244 );
and ( n47992 , n47991 , n40359 );
not ( n47993 , n40359 );
and ( n47994 , n47981 , n47982 );
xor ( n47995 , n47993 , n47994 );
and ( n47996 , n47995 , n40244 );
or ( n47997 , n47992 , n47996 );
not ( n47998 , n47997 );
buf ( n47999 , n47998 );
buf ( n48000 , n47999 );
not ( n48001 , n48000 );
or ( n48002 , n47990 , n48001 );
not ( n48003 , n40244 );
and ( n48004 , n48003 , n40514 );
not ( n48005 , n40514 );
and ( n48006 , n47993 , n47994 );
xor ( n48007 , n48005 , n48006 );
and ( n48008 , n48007 , n40244 );
or ( n48009 , n48004 , n48008 );
not ( n48010 , n48009 );
buf ( n48011 , n48010 );
buf ( n48012 , n48011 );
not ( n48013 , n48012 );
or ( n48014 , n48002 , n48013 );
not ( n48015 , n40244 );
and ( n48016 , n48015 , n40507 );
not ( n48017 , n40507 );
and ( n48018 , n48005 , n48006 );
xor ( n48019 , n48017 , n48018 );
and ( n48020 , n48019 , n40244 );
or ( n48021 , n48016 , n48020 );
not ( n48022 , n48021 );
buf ( n48023 , n48022 );
buf ( n48024 , n48023 );
not ( n48025 , n48024 );
or ( n48026 , n48014 , n48025 );
not ( n48027 , n40244 );
and ( n48028 , n48027 , n40500 );
not ( n48029 , n40500 );
and ( n48030 , n48017 , n48018 );
xor ( n48031 , n48029 , n48030 );
and ( n48032 , n48031 , n40244 );
or ( n48033 , n48028 , n48032 );
not ( n48034 , n48033 );
buf ( n48035 , n48034 );
buf ( n48036 , n48035 );
not ( n48037 , n48036 );
or ( n48038 , n48026 , n48037 );
not ( n48039 , n40244 );
and ( n48040 , n48039 , n40493 );
not ( n48041 , n40493 );
and ( n48042 , n48029 , n48030 );
xor ( n48043 , n48041 , n48042 );
and ( n48044 , n48043 , n40244 );
or ( n48045 , n48040 , n48044 );
not ( n48046 , n48045 );
buf ( n48047 , n48046 );
buf ( n48048 , n48047 );
not ( n48049 , n48048 );
or ( n48050 , n48038 , n48049 );
not ( n48051 , n40244 );
and ( n48052 , n48051 , n40486 );
not ( n48053 , n40486 );
and ( n48054 , n48041 , n48042 );
xor ( n48055 , n48053 , n48054 );
and ( n48056 , n48055 , n40244 );
or ( n48057 , n48052 , n48056 );
not ( n48058 , n48057 );
buf ( n48059 , n48058 );
buf ( n48060 , n48059 );
not ( n48061 , n48060 );
or ( n48062 , n48050 , n48061 );
not ( n48063 , n40244 );
and ( n48064 , n48063 , n40479 );
not ( n48065 , n40479 );
and ( n48066 , n48053 , n48054 );
xor ( n48067 , n48065 , n48066 );
and ( n48068 , n48067 , n40244 );
or ( n48069 , n48064 , n48068 );
not ( n48070 , n48069 );
buf ( n48071 , n48070 );
buf ( n48072 , n48071 );
not ( n48073 , n48072 );
or ( n48074 , n48062 , n48073 );
not ( n48075 , n40244 );
and ( n48076 , n48075 , n40472 );
not ( n48077 , n40472 );
and ( n48078 , n48065 , n48066 );
xor ( n48079 , n48077 , n48078 );
and ( n48080 , n48079 , n40244 );
or ( n48081 , n48076 , n48080 );
not ( n48082 , n48081 );
buf ( n48083 , n48082 );
buf ( n48084 , n48083 );
not ( n48085 , n48084 );
or ( n48086 , n48074 , n48085 );
not ( n48087 , n40244 );
and ( n48088 , n48087 , n40465 );
not ( n48089 , n40465 );
and ( n48090 , n48077 , n48078 );
xor ( n48091 , n48089 , n48090 );
and ( n48092 , n48091 , n40244 );
or ( n48093 , n48088 , n48092 );
not ( n48094 , n48093 );
buf ( n48095 , n48094 );
buf ( n48096 , n48095 );
not ( n48097 , n48096 );
or ( n48098 , n48086 , n48097 );
buf ( n48099 , n48098 );
buf ( n48100 , n48099 );
and ( n48101 , n48100 , n40244 );
not ( n48102 , n48101 );
and ( n48103 , n48102 , n48001 );
xor ( n48104 , n48001 , n40244 );
xor ( n48105 , n47989 , n40244 );
xor ( n48106 , n47977 , n40244 );
xor ( n48107 , n47965 , n40244 );
xor ( n48108 , n47953 , n40244 );
xor ( n48109 , n47941 , n40244 );
xor ( n48110 , n47929 , n40244 );
xor ( n48111 , n47918 , n40244 );
and ( n48112 , n48111 , n40244 );
and ( n48113 , n48110 , n48112 );
and ( n48114 , n48109 , n48113 );
and ( n48115 , n48108 , n48114 );
and ( n48116 , n48107 , n48115 );
and ( n48117 , n48106 , n48116 );
and ( n48118 , n48105 , n48117 );
xor ( n48119 , n48104 , n48118 );
and ( n48120 , n48119 , n48101 );
or ( n48121 , n48103 , n48120 );
and ( n48122 , n48121 , n47912 );
or ( n48123 , n47914 , n48122 );
and ( n48124 , n48123 , n32415 );
or ( n48125 , n35347 , n32419 );
or ( n48126 , n48125 , n32421 );
or ( n48127 , n48126 , n32423 );
or ( n48128 , n48127 , n32425 );
or ( n48129 , n48128 , n32427 );
or ( n48130 , n48129 , n32429 );
or ( n48131 , n48130 , n32431 );
or ( n48132 , n48131 , n32433 );
or ( n48133 , n48132 , n32435 );
and ( n48134 , n47900 , n48133 );
or ( n48135 , n47909 , n48124 , n48134 );
and ( n48136 , n48135 , n32456 );
and ( n48137 , n47900 , n47409 );
or ( n48138 , C0 , n48136 , n48137 );
buf ( n48139 , n48138 );
buf ( n48140 , n48139 );
buf ( n48141 , n31655 );
not ( n48142 , n34150 );
and ( n48143 , n48142 , n32838 );
not ( n48144 , n41392 );
and ( n48145 , n48144 , n32838 );
and ( n48146 , n32856 , n41392 );
or ( n48147 , n48145 , n48146 );
and ( n48148 , n48147 , n34150 );
or ( n48149 , n48143 , n48148 );
and ( n48150 , n48149 , n33381 );
not ( n48151 , n41402 );
not ( n48152 , n41392 );
and ( n48153 , n48152 , n32838 );
not ( n48154 , n34287 );
and ( n48155 , n48154 , n34270 );
xor ( n48156 , n34270 , n34193 );
and ( n48157 , n41460 , n41461 );
xor ( n48158 , n48156 , n48157 );
and ( n48159 , n48158 , n34287 );
or ( n48160 , n48155 , n48159 );
and ( n48161 , n48160 , n41392 );
or ( n48162 , n48153 , n48161 );
and ( n48163 , n48151 , n48162 );
and ( n48164 , n48160 , n41402 );
or ( n48165 , n48163 , n48164 );
and ( n48166 , n48165 , n33375 );
not ( n48167 , n32968 );
not ( n48168 , n41402 );
not ( n48169 , n41392 );
and ( n48170 , n48169 , n32838 );
and ( n48171 , n48160 , n41392 );
or ( n48172 , n48170 , n48171 );
and ( n48173 , n48168 , n48172 );
and ( n48174 , n48160 , n41402 );
or ( n48175 , n48173 , n48174 );
and ( n48176 , n48167 , n48175 );
not ( n48177 , n41424 );
not ( n48178 , n41428 );
and ( n48179 , n48178 , n48175 );
not ( n48180 , n34747 );
and ( n48181 , n48180 , n34726 );
xor ( n48182 , n34726 , n34625 );
and ( n48183 , n41486 , n41487 );
xor ( n48184 , n48182 , n48183 );
and ( n48185 , n48184 , n34747 );
or ( n48186 , n48181 , n48185 );
and ( n48187 , n48186 , n41428 );
or ( n48188 , n48179 , n48187 );
and ( n48189 , n48177 , n48188 );
not ( n48190 , n35036 );
and ( n48191 , n48190 , n35019 );
xor ( n48192 , n35019 , n34918 );
and ( n48193 , n41496 , n41497 );
xor ( n48194 , n48192 , n48193 );
and ( n48195 , n48194 , n35036 );
or ( n48196 , n48191 , n48195 );
and ( n48197 , n48196 , n41424 );
or ( n48198 , n48189 , n48197 );
and ( n48199 , n48198 , n32968 );
or ( n48200 , n48176 , n48199 );
and ( n48201 , n48200 , n33370 );
and ( n48202 , n32838 , n35062 );
or ( n48203 , C0 , n48150 , n48166 , n48201 , n48202 );
buf ( n48204 , n48203 );
buf ( n48205 , n48204 );
buf ( n48206 , n35539 );
buf ( n48207 , n31655 );
buf ( n48208 , n30987 );
buf ( n48209 , n30987 );
buf ( n48210 , n31655 );
not ( n48211 , n46356 );
and ( n48212 , n48211 , n31154 );
not ( n48213 , n31017 );
and ( n48214 , n46359 , n46360 , n48213 , n31013 , n46361 );
not ( n48215 , n48214 );
and ( n48216 , n48215 , n31154 );
and ( n48217 , n31172 , n48214 );
or ( n48218 , n48216 , n48217 );
and ( n48219 , n48218 , n46356 );
or ( n48220 , n48212 , n48219 );
and ( n48221 , n48220 , n31649 );
not ( n48222 , n46386 );
and ( n48223 , n46374 , n46380 , n48222 , n46392 , C1 );
not ( n48224 , n48223 );
not ( n48225 , n48214 );
and ( n48226 , n48225 , n31154 );
and ( n48227 , n46495 , n48214 );
or ( n48228 , n48226 , n48227 );
and ( n48229 , n48224 , n48228 );
and ( n48230 , n46495 , n48223 );
or ( n48231 , n48229 , n48230 );
and ( n48232 , n48231 , n31643 );
not ( n48233 , n31452 );
not ( n48234 , n48223 );
not ( n48235 , n48214 );
and ( n48236 , n48235 , n31154 );
and ( n48237 , n46495 , n48214 );
or ( n48238 , n48236 , n48237 );
and ( n48239 , n48234 , n48238 );
and ( n48240 , n46495 , n48223 );
or ( n48241 , n48239 , n48240 );
and ( n48242 , n48233 , n48241 );
not ( n48243 , n46539 );
and ( n48244 , n46520 , n46529 , n48243 , n46549 , C1 );
not ( n48245 , n48244 );
not ( n48246 , n46534 );
and ( n48247 , n46552 , n46553 , n48246 , n46544 , C1 );
not ( n48248 , n48247 );
and ( n48249 , n48248 , n48241 );
and ( n48250 , n46984 , n48247 );
or ( n48251 , n48249 , n48250 );
and ( n48252 , n48245 , n48251 );
and ( n48253 , n47267 , n48244 );
or ( n48254 , n48252 , n48253 );
and ( n48255 , n48254 , n31452 );
or ( n48256 , n48242 , n48255 );
and ( n48257 , n48256 , n31638 );
and ( n48258 , n31154 , n47277 );
or ( n48259 , C0 , n48221 , n48232 , n48257 , n48258 );
buf ( n48260 , n48259 );
buf ( n48261 , n48260 );
buf ( n48262 , n30987 );
buf ( n48263 , RI15b60738_1156);
and ( n48264 , n35291 , n48263 );
buf ( n48265 , RI15b3f9c0_35);
not ( n48266 , n48265 );
and ( n48267 , n48264 , n48266 );
not ( n48268 , n48267 );
and ( n48269 , n35292 , n48265 );
not ( n48270 , n48269 );
and ( n48271 , n35292 , n48266 );
and ( n48272 , n48271 , n48263 );
not ( n48273 , n48272 );
not ( n48274 , n48263 );
and ( n48275 , n48271 , n48274 );
not ( n48276 , n48275 );
and ( n48277 , n48273 , n48276 );
buf ( n48278 , n48277 );
and ( n48279 , n48270 , n48278 );
buf ( n48280 , n48269 );
or ( n48281 , n48279 , n48280 );
and ( n48282 , n48268 , n48281 );
buf ( n48283 , n48267 );
or ( n48284 , n48282 , n48283 );
and ( n48285 , n48284 , n39358 );
buf ( n48286 , n38450 );
and ( n48287 , n48263 , n48266 );
not ( n48288 , n48287 );
and ( n48289 , n48274 , n48266 );
not ( n48290 , n48289 );
and ( n48291 , n48288 , n48290 );
buf ( n48292 , n48291 );
and ( n48293 , n48292 , n39356 );
buf ( n48294 , RI15b3fa38_36);
not ( n48295 , n48294 );
and ( n48296 , n48295 , n48266 );
and ( n48297 , n48296 , n48263 );
not ( n48298 , n48297 );
or ( n48299 , n48265 , n48274 );
and ( n48300 , n48295 , n48299 );
not ( n48301 , n48300 );
not ( n48302 , n48294 );
and ( n48303 , n48301 , n48302 );
buf ( n48304 , n48300 );
or ( n48305 , n48303 , n48304 );
and ( n48306 , n48298 , n48305 );
buf ( n48307 , n48297 );
or ( n48308 , n48306 , n48307 );
and ( n48309 , n48308 , n39354 );
not ( n48310 , n48272 );
and ( n48311 , n35291 , n48294 );
not ( n48312 , n48311 );
or ( n48313 , n48263 , n48265 );
and ( n48314 , n35291 , n48295 );
and ( n48315 , n48313 , n48314 );
not ( n48316 , n48315 );
and ( n48317 , n48287 , n35291 );
and ( n48318 , n48317 , n48295 );
not ( n48319 , n48318 );
and ( n48320 , n48289 , n35292 );
not ( n48321 , n48320 );
and ( n48322 , n48265 , n35291 );
and ( n48323 , n48321 , n48322 );
buf ( n48324 , n48323 );
and ( n48325 , n48319 , n48324 );
buf ( n48326 , n48318 );
or ( n48327 , n48325 , n48326 );
and ( n48328 , n48316 , n48327 );
buf ( n48329 , n48315 );
or ( n48330 , n48328 , n48329 );
and ( n48331 , n48312 , n48330 );
and ( n48332 , n35284 , n48311 );
or ( n48333 , n48331 , n48332 );
and ( n48334 , n48310 , n48333 );
buf ( n48335 , n48334 );
and ( n48336 , n48335 , n39352 );
not ( n48337 , n48263 );
and ( n48338 , n48337 , n48265 );
buf ( n48339 , n48338 );
and ( n48340 , n48339 , n39349 );
or ( n48341 , n48285 , n48286 , n48293 , n48309 , n48336 , C0 , n48340 , C0 );
buf ( n48342 , n48341 );
buf ( n48343 , n48342 );
buf ( n48344 , n31655 );
buf ( n48345 , n30987 );
and ( n48346 , n31586 , n31007 );
not ( n48347 , n31077 );
and ( n48348 , n48347 , n34010 );
and ( n48349 , n31010 , n39816 );
and ( n48350 , n48349 , n31077 );
or ( n48351 , n48348 , n48350 );
and ( n48352 , n48351 , n31373 );
not ( n48353 , n31402 );
and ( n48354 , n48353 , n34010 );
and ( n48355 , n48349 , n31402 );
or ( n48356 , n48354 , n48355 );
and ( n48357 , n48356 , n31408 );
not ( n48358 , n31437 );
and ( n48359 , n48358 , n34010 );
not ( n48360 , n31455 );
and ( n48361 , n48360 , n34060 );
xor ( n48362 , n34010 , n34013 );
and ( n48363 , n48362 , n31455 );
or ( n48364 , n48361 , n48363 );
and ( n48365 , n48364 , n31437 );
or ( n48366 , n48359 , n48365 );
and ( n48367 , n48366 , n31468 );
not ( n48368 , n31497 );
and ( n48369 , n48368 , n34010 );
not ( n48370 , n31454 );
not ( n48371 , n31501 );
and ( n48372 , n48371 , n34060 );
xor ( n48373 , n34061 , n34065 );
and ( n48374 , n48373 , n31501 );
or ( n48375 , n48372 , n48374 );
and ( n48376 , n48370 , n48375 );
and ( n48377 , n48362 , n31454 );
or ( n48378 , n48376 , n48377 );
and ( n48379 , n48378 , n31497 );
or ( n48380 , n48369 , n48379 );
and ( n48381 , n48380 , n31521 );
and ( n48382 , n34010 , n31553 );
or ( n48383 , n48352 , n48357 , n48367 , n48381 , n48382 );
and ( n48384 , n48383 , n31557 );
not ( n48385 , n31452 );
not ( n48386 , n31619 );
and ( n48387 , n48386 , n34117 );
xor ( n48388 , n34118 , n34122 );
and ( n48389 , n48388 , n31619 );
or ( n48390 , n48387 , n48389 );
and ( n48391 , n48385 , n48390 );
and ( n48392 , n34010 , n31452 );
or ( n48393 , n48391 , n48392 );
and ( n48394 , n48393 , n31638 );
buf ( n48395 , n33973 );
and ( n48396 , n34010 , n31650 );
or ( n48397 , C0 , n48346 , n48384 , n48394 , n48395 , n48396 );
buf ( n48398 , n48397 );
buf ( n48399 , n48398 );
buf ( n48400 , n31655 );
buf ( n48401 , n31655 );
and ( n48402 , n31589 , n31007 );
not ( n48403 , n31077 );
and ( n48404 , n48403 , n31460 );
and ( n48405 , n33484 , n31077 );
or ( n48406 , n48404 , n48405 );
and ( n48407 , n48406 , n31373 );
not ( n48408 , n31402 );
and ( n48409 , n48408 , n31460 );
and ( n48410 , n33484 , n31402 );
or ( n48411 , n48409 , n48410 );
and ( n48412 , n48411 , n31408 );
not ( n48413 , n31437 );
and ( n48414 , n48413 , n31460 );
not ( n48415 , n31455 );
and ( n48416 , n48415 , n31507 );
not ( n48417 , n31460 );
and ( n48418 , n48417 , n31455 );
or ( n48419 , n48416 , n48418 );
and ( n48420 , n48419 , n31437 );
or ( n48421 , n48414 , n48420 );
and ( n48422 , n48421 , n31468 );
not ( n48423 , n31497 );
and ( n48424 , n48423 , n31460 );
not ( n48425 , n31454 );
not ( n48426 , n31501 );
and ( n48427 , n48426 , n31507 );
xor ( n48428 , n31508 , n31510 );
and ( n48429 , n48428 , n31501 );
or ( n48430 , n48427 , n48429 );
and ( n48431 , n48425 , n48430 );
and ( n48432 , n48417 , n31454 );
or ( n48433 , n48431 , n48432 );
and ( n48434 , n48433 , n31497 );
or ( n48435 , n48424 , n48434 );
and ( n48436 , n48435 , n31521 );
and ( n48437 , n31460 , n31553 );
or ( n48438 , n48407 , n48412 , n48422 , n48436 , n48437 );
and ( n48439 , n48438 , n31557 );
not ( n48440 , n31452 );
not ( n48441 , n31619 );
and ( n48442 , n48441 , n31626 );
xor ( n48443 , n31627 , n31629 );
and ( n48444 , n48443 , n31619 );
or ( n48445 , n48442 , n48444 );
and ( n48446 , n48440 , n48445 );
and ( n48447 , n31460 , n31452 );
or ( n48448 , n48446 , n48447 );
and ( n48449 , n48448 , n31638 );
and ( n48450 , n31460 , n31650 );
or ( n48451 , C0 , n48402 , n48439 , n48449 , C0 , n48450 );
buf ( n48452 , n48451 );
buf ( n48453 , n48452 );
buf ( n48454 , n30987 );
or ( n48455 , n31544 , n31546 );
and ( n48456 , n33763 , n48455 );
and ( n48457 , n31077 , n44703 );
not ( n48458 , n48457 );
and ( n48459 , n48458 , n33428 );
and ( n48460 , n33763 , n48457 );
or ( n48461 , n48459 , n48460 );
and ( n48462 , n48461 , n31373 );
not ( n48463 , n44807 );
and ( n48464 , n48463 , n33428 );
and ( n48465 , n33763 , n44807 );
or ( n48466 , n48464 , n48465 );
and ( n48467 , n48466 , n31408 );
and ( n48468 , n31437 , n44703 );
not ( n48469 , n48468 );
and ( n48470 , n48469 , n33428 );
and ( n48471 , n33763 , n48468 );
or ( n48472 , n48470 , n48471 );
and ( n48473 , n48472 , n31468 );
not ( n48474 , n44817 );
and ( n48475 , n48474 , n33428 );
and ( n48476 , n33763 , n44817 );
or ( n48477 , n48475 , n48476 );
and ( n48478 , n48477 , n31521 );
not ( n48479 , n39979 );
and ( n48480 , n48479 , n33428 );
and ( n48481 , n33470 , n39979 );
or ( n48482 , n48480 , n48481 );
and ( n48483 , n48482 , n31538 );
not ( n48484 , n45059 );
and ( n48485 , n48484 , n33428 );
and ( n48486 , n33470 , n45059 );
or ( n48487 , n48485 , n48486 );
and ( n48488 , n48487 , n31536 );
not ( n48489 , n33419 );
and ( n48490 , n48489 , n33428 );
xor ( n48491 , n33470 , n33695 );
and ( n48492 , n48491 , n33419 );
or ( n48493 , n48490 , n48492 );
and ( n48494 , n48493 , n31529 );
not ( n48495 , n33734 );
and ( n48496 , n48495 , n33428 );
not ( n48497 , n33533 );
xor ( n48498 , n33763 , n33813 );
and ( n48499 , n48497 , n48498 );
xnor ( n48500 , n33848 , n33915 );
and ( n48501 , n48500 , n33533 );
or ( n48502 , n48499 , n48501 );
and ( n48503 , n48502 , n33734 );
or ( n48504 , n48496 , n48503 );
and ( n48505 , n48504 , n31527 );
or ( n48506 , n31524 , n31523 );
or ( n48507 , n48506 , n31531 );
or ( n48508 , n48507 , n31534 );
or ( n48509 , n48508 , n31540 );
or ( n48510 , n48509 , n31542 );
or ( n48511 , n48510 , n31548 );
or ( n48512 , n48511 , n31550 );
or ( n48513 , n48512 , n31552 );
and ( n48514 , n33848 , n48513 );
or ( n48515 , n48456 , n48462 , n48467 , n48473 , n48478 , n48483 , n48488 , n48494 , n48505 , n48514 );
and ( n48516 , n48515 , n31557 );
and ( n48517 , n34000 , n33973 );
or ( n48518 , n31640 , n31638 );
or ( n48519 , n48518 , n31641 );
or ( n48520 , n48519 , n31643 );
or ( n48521 , n48520 , n31645 );
or ( n48522 , n48521 , n31647 );
or ( n48523 , n48522 , n31649 );
or ( n48524 , n48523 , n31007 );
and ( n48525 , n33428 , n48524 );
or ( n48526 , C0 , n48516 , n48517 , n48525 );
buf ( n48527 , n48526 );
buf ( n48528 , n48527 );
buf ( n48529 , n31655 );
buf ( n48530 , RI15b60828_1158);
or ( n48531 , n39346 , n38450 );
and ( n48532 , n48530 , n48531 );
buf ( n48533 , RI15b5e848_1090);
and ( n48534 , n48533 , n39359 );
or ( n48535 , n48532 , n48534 );
buf ( n48536 , n48535 );
buf ( n48537 , n48536 );
buf ( n48538 , n30987 );
buf ( n48539 , n31655 );
buf ( n48540 , n31655 );
buf ( n48541 , n30987 );
buf ( n48542 , n30987 );
buf ( n48543 , RI15b46950_273);
and ( n48544 , n48543 , n33377 );
and ( n48545 , n32598 , n32963 );
not ( n48546 , n48545 );
buf ( n48547 , RI15b470d0_289);
and ( n48548 , n48546 , n48547 );
not ( n48549 , n39572 );
and ( n48550 , n48549 , n39425 );
xor ( n48551 , n42624 , n42629 );
and ( n48552 , n48551 , n39572 );
or ( n48553 , n48550 , n48552 );
and ( n48554 , n48553 , n48545 );
or ( n48555 , n48548 , n48554 );
and ( n48556 , n48555 , n32890 );
and ( n48557 , n32953 , n32963 );
not ( n48558 , n48557 );
and ( n48559 , n48558 , n48547 );
and ( n48560 , n48553 , n48557 );
or ( n48561 , n48559 , n48560 );
and ( n48562 , n48561 , n33038 );
or ( n48563 , n33190 , n33172 );
or ( n48564 , n48563 , n32924 );
or ( n48565 , n48564 , n33191 );
or ( n48566 , n48565 , n33193 );
or ( n48567 , n48566 , n33195 );
or ( n48568 , n48567 , n33197 );
or ( n48569 , n48568 , n33199 );
or ( n48570 , n48569 , n33201 );
or ( n48571 , n48570 , n33203 );
and ( n48572 , n48547 , n48571 );
or ( n48573 , n48556 , n48562 , n48572 );
and ( n48574 , n48573 , n33208 );
or ( n48575 , n39801 , n33379 );
or ( n48576 , n48575 , n33381 );
or ( n48577 , n48576 , n32528 );
and ( n48578 , n48547 , n48577 );
or ( n48579 , C0 , n48544 , n48574 , n48578 );
buf ( n48580 , n48579 );
buf ( n48581 , n48580 );
buf ( n48582 , RI15b44880_203);
buf ( n48583 , RI15b44808_202);
buf ( n48584 , RI15b44790_201);
buf ( n48585 , RI15b44718_200);
buf ( n48586 , RI15b446a0_199);
buf ( n48587 , RI15b44628_198);
buf ( n48588 , RI15b445b0_197);
buf ( n48589 , RI15b44538_196);
buf ( n48590 , RI15b444c0_195);
buf ( n48591 , RI15b44448_194);
buf ( n48592 , RI15b443d0_193);
buf ( n48593 , RI15b44358_192);
buf ( n48594 , RI15b442e0_191);
buf ( n48595 , RI15b44268_190);
buf ( n48596 , RI15b441f0_189);
buf ( n48597 , RI15b44178_188);
buf ( n48598 , RI15b44100_187);
buf ( n48599 , RI15b44088_186);
buf ( n48600 , RI15b44010_185);
buf ( n48601 , RI15b43f98_184);
buf ( n48602 , RI15b43f20_183);
buf ( n48603 , RI15b43ea8_182);
buf ( n48604 , RI15b43e30_181);
buf ( n48605 , RI15b43db8_180);
buf ( n48606 , RI15b43d40_179);
buf ( n48607 , RI15b43cc8_178);
buf ( n48608 , RI15b43c50_177);
buf ( n48609 , RI15b43bd8_176);
buf ( n48610 , RI15b43b60_175);
and ( n48611 , n48609 , n48610 );
and ( n48612 , n48608 , n48611 );
and ( n48613 , n48607 , n48612 );
and ( n48614 , n48606 , n48613 );
and ( n48615 , n48605 , n48614 );
and ( n48616 , n48604 , n48615 );
and ( n48617 , n48603 , n48616 );
and ( n48618 , n48602 , n48617 );
and ( n48619 , n48601 , n48618 );
and ( n48620 , n48600 , n48619 );
and ( n48621 , n48599 , n48620 );
and ( n48622 , n48598 , n48621 );
and ( n48623 , n48597 , n48622 );
and ( n48624 , n48596 , n48623 );
and ( n48625 , n48595 , n48624 );
and ( n48626 , n48594 , n48625 );
and ( n48627 , n48593 , n48626 );
and ( n48628 , n48592 , n48627 );
and ( n48629 , n48591 , n48628 );
and ( n48630 , n48590 , n48629 );
and ( n48631 , n48589 , n48630 );
and ( n48632 , n48588 , n48631 );
and ( n48633 , n48587 , n48632 );
and ( n48634 , n48586 , n48633 );
and ( n48635 , n48585 , n48634 );
and ( n48636 , n48584 , n48635 );
and ( n48637 , n48583 , n48636 );
xor ( n48638 , n48582 , n48637 );
or ( n48639 , n33195 , n33197 );
and ( n48640 , n48638 , n48639 );
and ( n48641 , n32963 , n32967 );
and ( n48642 , n32598 , n48641 );
not ( n48643 , n48642 );
and ( n48644 , n48643 , n48582 );
and ( n48645 , n48638 , n48642 );
or ( n48646 , n48644 , n48645 );
and ( n48647 , n48646 , n32890 );
and ( n48648 , n32919 , n32967 );
not ( n48649 , n48648 );
and ( n48650 , n48649 , n48582 );
and ( n48651 , n48638 , n48648 );
or ( n48652 , n48650 , n48651 );
and ( n48653 , n48652 , n32924 );
and ( n48654 , n32953 , n48641 );
not ( n48655 , n48654 );
and ( n48656 , n48655 , n48582 );
and ( n48657 , n48638 , n48654 );
or ( n48658 , n48656 , n48657 );
and ( n48659 , n48658 , n33038 );
and ( n48660 , n33067 , n32967 );
not ( n48661 , n48660 );
and ( n48662 , n48661 , n48582 );
and ( n48663 , n48638 , n48660 );
or ( n48664 , n48662 , n48663 );
and ( n48665 , n48664 , n33172 );
not ( n48666 , n41576 );
and ( n48667 , n48666 , n48582 );
buf ( n48668 , RI15b43ae8_174);
and ( n48669 , n48610 , n48668 );
or ( n48670 , n48609 , n48669 );
and ( n48671 , n48608 , n48670 );
and ( n48672 , n48607 , n48671 );
and ( n48673 , n48606 , n48672 );
and ( n48674 , n48605 , n48673 );
and ( n48675 , n48604 , n48674 );
and ( n48676 , n48603 , n48675 );
and ( n48677 , n48602 , n48676 );
and ( n48678 , n48601 , n48677 );
and ( n48679 , n48600 , n48678 );
and ( n48680 , n48599 , n48679 );
and ( n48681 , n48598 , n48680 );
and ( n48682 , n48597 , n48681 );
and ( n48683 , n48596 , n48682 );
and ( n48684 , n48595 , n48683 );
and ( n48685 , n48594 , n48684 );
and ( n48686 , n48593 , n48685 );
and ( n48687 , n48592 , n48686 );
and ( n48688 , n48591 , n48687 );
and ( n48689 , n48590 , n48688 );
and ( n48690 , n48589 , n48689 );
and ( n48691 , n48588 , n48690 );
and ( n48692 , n48587 , n48691 );
and ( n48693 , n48586 , n48692 );
and ( n48694 , n48585 , n48693 );
and ( n48695 , n48584 , n48694 );
and ( n48696 , n48583 , n48695 );
xor ( n48697 , n48582 , n48696 );
and ( n48698 , n48697 , n41576 );
or ( n48699 , n48667 , n48698 );
and ( n48700 , n48699 , n33189 );
not ( n48701 , n32562 );
buf ( n48702 , n32562 );
buf ( n48703 , n32562 );
buf ( n48704 , n32562 );
buf ( n48705 , n32562 );
buf ( n48706 , n32562 );
buf ( n48707 , n32562 );
buf ( n48708 , n32562 );
buf ( n48709 , n32562 );
buf ( n48710 , n32562 );
buf ( n48711 , n32562 );
buf ( n48712 , n32562 );
buf ( n48713 , n32562 );
buf ( n48714 , n32562 );
buf ( n48715 , n32562 );
buf ( n48716 , n32562 );
buf ( n48717 , n32562 );
buf ( n48718 , n32562 );
buf ( n48719 , n32562 );
buf ( n48720 , n32562 );
buf ( n48721 , n32562 );
buf ( n48722 , n32562 );
buf ( n48723 , n32562 );
buf ( n48724 , n32562 );
buf ( n48725 , n32562 );
buf ( n48726 , n32562 );
or ( n48727 , n32596 , n41572 );
and ( n48728 , n32565 , n48727 );
or ( n48729 , n32567 , n32569 , n32562 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48728 );
and ( n48730 , n48701 , n48729 );
not ( n48731 , n48730 );
and ( n48732 , n48731 , n48582 );
and ( n48733 , n48697 , n48730 );
or ( n48734 , n48732 , n48733 );
and ( n48735 , n48734 , n33187 );
not ( n48736 , n32562 );
buf ( n48737 , n32562 );
buf ( n48738 , n32562 );
buf ( n48739 , n32562 );
buf ( n48740 , n32562 );
buf ( n48741 , n32562 );
buf ( n48742 , n32562 );
buf ( n48743 , n32562 );
buf ( n48744 , n32562 );
buf ( n48745 , n32562 );
buf ( n48746 , n32562 );
buf ( n48747 , n32562 );
buf ( n48748 , n32562 );
buf ( n48749 , n32562 );
buf ( n48750 , n32562 );
buf ( n48751 , n32562 );
buf ( n48752 , n32562 );
buf ( n48753 , n32562 );
buf ( n48754 , n32562 );
buf ( n48755 , n32562 );
buf ( n48756 , n32562 );
buf ( n48757 , n32562 );
buf ( n48758 , n32562 );
buf ( n48759 , n32562 );
buf ( n48760 , n32562 );
buf ( n48761 , n32562 );
or ( n48762 , n32596 , n41572 );
and ( n48763 , n32565 , n48762 );
or ( n48764 , n32567 , n32569 , n32562 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48763 );
and ( n48765 , n48736 , n48764 );
not ( n48766 , n48765 );
and ( n48767 , n48766 , n48582 );
xor ( n48768 , n48583 , n48695 );
xor ( n48769 , n48584 , n48694 );
xor ( n48770 , n48585 , n48693 );
xor ( n48771 , n48586 , n48692 );
xor ( n48772 , n48587 , n48691 );
xor ( n48773 , n48588 , n48690 );
xor ( n48774 , n48589 , n48689 );
xor ( n48775 , n48590 , n48688 );
xor ( n48776 , n48591 , n48687 );
xor ( n48777 , n48592 , n48686 );
xor ( n48778 , n48593 , n48685 );
xor ( n48779 , n48594 , n48684 );
xor ( n48780 , n48595 , n48683 );
xor ( n48781 , n48596 , n48682 );
xor ( n48782 , n48597 , n48681 );
xor ( n48783 , n48598 , n48680 );
xor ( n48784 , n48599 , n48679 );
xor ( n48785 , n48600 , n48678 );
xor ( n48786 , n48601 , n48677 );
xor ( n48787 , n48602 , n48676 );
xor ( n48788 , n48603 , n48675 );
xor ( n48789 , n48604 , n48674 );
not ( n48790 , n32547 );
not ( n48791 , n48790 );
buf ( n48792 , n48791 );
not ( n48793 , n48792 );
not ( n48794 , n48793 );
xor ( n48795 , n32543 , n32547 );
not ( n48796 , n48795 );
buf ( n48797 , n48796 );
buf ( n48798 , n48797 );
not ( n48799 , n48798 );
not ( n48800 , n48799 );
xor ( n48801 , n32539 , n45914 );
not ( n48802 , n48801 );
buf ( n48803 , n48802 );
buf ( n48804 , n48803 );
not ( n48805 , n48804 );
not ( n48806 , n48805 );
xor ( n48807 , n32535 , n45915 );
not ( n48808 , n48807 );
buf ( n48809 , n48808 );
buf ( n48810 , n48809 );
not ( n48811 , n48810 );
not ( n48812 , n48811 );
nor ( n48813 , n48794 , n48800 , n48806 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48814 , n32857 , n48813 );
nor ( n48815 , n48793 , n48800 , n48806 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48816 , n32859 , n48815 );
nor ( n48817 , n48794 , n48799 , n48806 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48818 , n32861 , n48817 );
nor ( n48819 , n48793 , n48799 , n48806 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48820 , n32863 , n48819 );
nor ( n48821 , n48794 , n48800 , n48805 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48822 , n32865 , n48821 );
nor ( n48823 , n48793 , n48800 , n48805 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48824 , n32867 , n48823 );
nor ( n48825 , n48794 , n48799 , n48805 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48826 , n32869 , n48825 );
nor ( n48827 , n48793 , n48799 , n48805 , n48812 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48828 , n32871 , n48827 );
nor ( n48829 , n48794 , n48800 , n48806 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48830 , n32873 , n48829 );
nor ( n48831 , n48793 , n48800 , n48806 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48832 , n32875 , n48831 );
nor ( n48833 , n48794 , n48799 , n48806 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48834 , n32877 , n48833 );
nor ( n48835 , n48793 , n48799 , n48806 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48836 , n32879 , n48835 );
nor ( n48837 , n48794 , n48800 , n48805 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48838 , n32881 , n48837 );
nor ( n48839 , n48793 , n48800 , n48805 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48840 , n32883 , n48839 );
nor ( n48841 , n48794 , n48799 , n48805 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48842 , n32885 , n48841 );
nor ( n48843 , n48793 , n48799 , n48805 , n48811 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n48844 , n32887 , n48843 );
or ( n48845 , n48814 , n48816 , n48818 , n48820 , n48822 , n48824 , n48826 , n48828 , n48830 , n48832 , n48834 , n48836 , n48838 , n48840 , n48842 , n48844 );
and ( n48846 , n48789 , n48845 );
xor ( n48847 , n48605 , n48673 );
and ( n48848 , n32824 , n48813 );
and ( n48849 , n32826 , n48815 );
and ( n48850 , n32828 , n48817 );
and ( n48851 , n32830 , n48819 );
and ( n48852 , n32832 , n48821 );
and ( n48853 , n32834 , n48823 );
and ( n48854 , n32836 , n48825 );
and ( n48855 , n32838 , n48827 );
and ( n48856 , n32840 , n48829 );
and ( n48857 , n32842 , n48831 );
and ( n48858 , n32844 , n48833 );
and ( n48859 , n32846 , n48835 );
and ( n48860 , n32848 , n48837 );
and ( n48861 , n32850 , n48839 );
and ( n48862 , n32852 , n48841 );
and ( n48863 , n32854 , n48843 );
or ( n48864 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 );
and ( n48865 , n48847 , n48864 );
xor ( n48866 , n48606 , n48672 );
and ( n48867 , n32791 , n48813 );
and ( n48868 , n32793 , n48815 );
and ( n48869 , n32795 , n48817 );
and ( n48870 , n32797 , n48819 );
and ( n48871 , n32799 , n48821 );
and ( n48872 , n32801 , n48823 );
and ( n48873 , n32803 , n48825 );
and ( n48874 , n32805 , n48827 );
and ( n48875 , n32807 , n48829 );
and ( n48876 , n32809 , n48831 );
and ( n48877 , n32811 , n48833 );
and ( n48878 , n32813 , n48835 );
and ( n48879 , n32815 , n48837 );
and ( n48880 , n32817 , n48839 );
and ( n48881 , n32819 , n48841 );
and ( n48882 , n32821 , n48843 );
or ( n48883 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 );
and ( n48884 , n48866 , n48883 );
xor ( n48885 , n48607 , n48671 );
and ( n48886 , n32757 , n48813 );
and ( n48887 , n32759 , n48815 );
and ( n48888 , n32761 , n48817 );
and ( n48889 , n32763 , n48819 );
and ( n48890 , n32765 , n48821 );
and ( n48891 , n32767 , n48823 );
and ( n48892 , n32769 , n48825 );
and ( n48893 , n32771 , n48827 );
and ( n48894 , n32773 , n48829 );
and ( n48895 , n32775 , n48831 );
and ( n48896 , n32777 , n48833 );
and ( n48897 , n32779 , n48835 );
and ( n48898 , n32781 , n48837 );
and ( n48899 , n32783 , n48839 );
and ( n48900 , n32785 , n48841 );
and ( n48901 , n32787 , n48843 );
or ( n48902 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 );
and ( n48903 , n48885 , n48902 );
xor ( n48904 , n48608 , n48670 );
and ( n48905 , n32723 , n48813 );
and ( n48906 , n32725 , n48815 );
and ( n48907 , n32727 , n48817 );
and ( n48908 , n32729 , n48819 );
and ( n48909 , n32731 , n48821 );
and ( n48910 , n32733 , n48823 );
and ( n48911 , n32735 , n48825 );
and ( n48912 , n32737 , n48827 );
and ( n48913 , n32739 , n48829 );
and ( n48914 , n32741 , n48831 );
and ( n48915 , n32743 , n48833 );
and ( n48916 , n32745 , n48835 );
and ( n48917 , n32747 , n48837 );
and ( n48918 , n32749 , n48839 );
and ( n48919 , n32751 , n48841 );
and ( n48920 , n32753 , n48843 );
or ( n48921 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 );
and ( n48922 , n48904 , n48921 );
xnor ( n48923 , n48609 , n48669 );
and ( n48924 , n32690 , n48813 );
and ( n48925 , n32692 , n48815 );
and ( n48926 , n32694 , n48817 );
and ( n48927 , n32696 , n48819 );
and ( n48928 , n32698 , n48821 );
and ( n48929 , n32700 , n48823 );
and ( n48930 , n32702 , n48825 );
and ( n48931 , n32704 , n48827 );
and ( n48932 , n32706 , n48829 );
and ( n48933 , n32708 , n48831 );
and ( n48934 , n32710 , n48833 );
and ( n48935 , n32712 , n48835 );
and ( n48936 , n32714 , n48837 );
and ( n48937 , n32716 , n48839 );
and ( n48938 , n32718 , n48841 );
and ( n48939 , n32720 , n48843 );
or ( n48940 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 );
and ( n48941 , n48923 , n48940 );
xor ( n48942 , n48610 , n48668 );
and ( n48943 , n32657 , n48813 );
and ( n48944 , n32659 , n48815 );
and ( n48945 , n32661 , n48817 );
and ( n48946 , n32663 , n48819 );
and ( n48947 , n32665 , n48821 );
and ( n48948 , n32667 , n48823 );
and ( n48949 , n32669 , n48825 );
and ( n48950 , n32671 , n48827 );
and ( n48951 , n32673 , n48829 );
and ( n48952 , n32675 , n48831 );
and ( n48953 , n32677 , n48833 );
and ( n48954 , n32679 , n48835 );
and ( n48955 , n32681 , n48837 );
and ( n48956 , n32683 , n48839 );
and ( n48957 , n32685 , n48841 );
and ( n48958 , n32687 , n48843 );
or ( n48959 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 );
and ( n48960 , n48942 , n48959 );
not ( n48961 , n48668 );
and ( n48962 , n32603 , n48813 );
and ( n48963 , n32607 , n48815 );
and ( n48964 , n32611 , n48817 );
and ( n48965 , n32615 , n48819 );
and ( n48966 , n32618 , n48821 );
and ( n48967 , n32622 , n48823 );
and ( n48968 , n32625 , n48825 );
and ( n48969 , n32628 , n48827 );
and ( n48970 , n32631 , n48829 );
and ( n48971 , n32634 , n48831 );
and ( n48972 , n32637 , n48833 );
and ( n48973 , n32640 , n48835 );
and ( n48974 , n32643 , n48837 );
and ( n48975 , n32646 , n48839 );
and ( n48976 , n32649 , n48841 );
and ( n48977 , n32652 , n48843 );
or ( n48978 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 );
and ( n48979 , n48961 , n48978 );
and ( n48980 , n48959 , n48979 );
and ( n48981 , n48942 , n48979 );
or ( n48982 , n48960 , n48980 , n48981 );
and ( n48983 , n48940 , n48982 );
and ( n48984 , n48923 , n48982 );
or ( n48985 , n48941 , n48983 , n48984 );
and ( n48986 , n48921 , n48985 );
and ( n48987 , n48904 , n48985 );
or ( n48988 , n48922 , n48986 , n48987 );
and ( n48989 , n48902 , n48988 );
and ( n48990 , n48885 , n48988 );
or ( n48991 , n48903 , n48989 , n48990 );
and ( n48992 , n48883 , n48991 );
and ( n48993 , n48866 , n48991 );
or ( n48994 , n48884 , n48992 , n48993 );
and ( n48995 , n48864 , n48994 );
and ( n48996 , n48847 , n48994 );
or ( n48997 , n48865 , n48995 , n48996 );
and ( n48998 , n48845 , n48997 );
and ( n48999 , n48789 , n48997 );
or ( n49000 , n48846 , n48998 , n48999 );
and ( n49001 , n48788 , n49000 );
and ( n49002 , n48787 , n49001 );
and ( n49003 , n48786 , n49002 );
and ( n49004 , n48785 , n49003 );
and ( n49005 , n48784 , n49004 );
and ( n49006 , n48783 , n49005 );
and ( n49007 , n48782 , n49006 );
and ( n49008 , n48781 , n49007 );
and ( n49009 , n48780 , n49008 );
and ( n49010 , n48779 , n49009 );
and ( n49011 , n48778 , n49010 );
and ( n49012 , n48777 , n49011 );
and ( n49013 , n48776 , n49012 );
and ( n49014 , n48775 , n49013 );
and ( n49015 , n48774 , n49014 );
and ( n49016 , n48773 , n49015 );
and ( n49017 , n48772 , n49016 );
and ( n49018 , n48771 , n49017 );
and ( n49019 , n48770 , n49018 );
and ( n49020 , n48769 , n49019 );
and ( n49021 , n48768 , n49020 );
xor ( n49022 , n48697 , n49021 );
and ( n49023 , n49022 , n48765 );
or ( n49024 , n48767 , n49023 );
and ( n49025 , n49024 , n33180 );
not ( n49026 , n32562 );
buf ( n49027 , n32562 );
buf ( n49028 , n32562 );
buf ( n49029 , n32562 );
buf ( n49030 , n32562 );
buf ( n49031 , n32562 );
buf ( n49032 , n32562 );
buf ( n49033 , n32562 );
buf ( n49034 , n32562 );
buf ( n49035 , n32562 );
buf ( n49036 , n32562 );
buf ( n49037 , n32562 );
buf ( n49038 , n32562 );
buf ( n49039 , n32562 );
buf ( n49040 , n32562 );
buf ( n49041 , n32562 );
buf ( n49042 , n32562 );
buf ( n49043 , n32562 );
buf ( n49044 , n32562 );
buf ( n49045 , n32562 );
buf ( n49046 , n32562 );
buf ( n49047 , n32562 );
buf ( n49048 , n32562 );
buf ( n49049 , n32562 );
buf ( n49050 , n32562 );
buf ( n49051 , n32562 );
and ( n49052 , n41572 , n32596 );
or ( n49053 , n32565 , n32567 , n32569 , n32562 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 );
and ( n49054 , n49026 , n49053 );
not ( n49055 , n49054 );
and ( n49056 , n49055 , n48582 );
not ( n49057 , n48845 );
xor ( n49058 , n48583 , n48636 );
xor ( n49059 , n48584 , n48635 );
xor ( n49060 , n48585 , n48634 );
xor ( n49061 , n48586 , n48633 );
xor ( n49062 , n48587 , n48632 );
xor ( n49063 , n48588 , n48631 );
xor ( n49064 , n48589 , n48630 );
xor ( n49065 , n48590 , n48629 );
xor ( n49066 , n48591 , n48628 );
xor ( n49067 , n48592 , n48627 );
xor ( n49068 , n48593 , n48626 );
xor ( n49069 , n48594 , n48625 );
xor ( n49070 , n48595 , n48624 );
xor ( n49071 , n48596 , n48623 );
xor ( n49072 , n48597 , n48622 );
xor ( n49073 , n48598 , n48621 );
xor ( n49074 , n48599 , n48620 );
xor ( n49075 , n48600 , n48619 );
xor ( n49076 , n48601 , n48618 );
xor ( n49077 , n48602 , n48617 );
xor ( n49078 , n48603 , n48616 );
xor ( n49079 , n48604 , n48615 );
and ( n49080 , n49079 , n48845 );
xor ( n49081 , n48605 , n48614 );
and ( n49082 , n49081 , n48864 );
xor ( n49083 , n48606 , n48613 );
and ( n49084 , n49083 , n48883 );
xor ( n49085 , n48607 , n48612 );
and ( n49086 , n49085 , n48902 );
xor ( n49087 , n48608 , n48611 );
and ( n49088 , n49087 , n48921 );
xor ( n49089 , n48609 , n48610 );
and ( n49090 , n49089 , n48940 );
not ( n49091 , n48610 );
and ( n49092 , n49091 , n48959 );
and ( n49093 , n48668 , n48978 );
and ( n49094 , n48959 , n49093 );
and ( n49095 , n49091 , n49093 );
or ( n49096 , n49092 , n49094 , n49095 );
and ( n49097 , n48940 , n49096 );
and ( n49098 , n49089 , n49096 );
or ( n49099 , n49090 , n49097 , n49098 );
and ( n49100 , n48921 , n49099 );
and ( n49101 , n49087 , n49099 );
or ( n49102 , n49088 , n49100 , n49101 );
and ( n49103 , n48902 , n49102 );
and ( n49104 , n49085 , n49102 );
or ( n49105 , n49086 , n49103 , n49104 );
and ( n49106 , n48883 , n49105 );
and ( n49107 , n49083 , n49105 );
or ( n49108 , n49084 , n49106 , n49107 );
and ( n49109 , n48864 , n49108 );
and ( n49110 , n49081 , n49108 );
or ( n49111 , n49082 , n49109 , n49110 );
and ( n49112 , n48845 , n49111 );
and ( n49113 , n49079 , n49111 );
or ( n49114 , n49080 , n49112 , n49113 );
and ( n49115 , n49078 , n49114 );
and ( n49116 , n49077 , n49115 );
and ( n49117 , n49076 , n49116 );
and ( n49118 , n49075 , n49117 );
and ( n49119 , n49074 , n49118 );
and ( n49120 , n49073 , n49119 );
and ( n49121 , n49072 , n49120 );
and ( n49122 , n49071 , n49121 );
and ( n49123 , n49070 , n49122 );
and ( n49124 , n49069 , n49123 );
and ( n49125 , n49068 , n49124 );
and ( n49126 , n49067 , n49125 );
and ( n49127 , n49066 , n49126 );
and ( n49128 , n49065 , n49127 );
and ( n49129 , n49064 , n49128 );
and ( n49130 , n49063 , n49129 );
and ( n49131 , n49062 , n49130 );
and ( n49132 , n49061 , n49131 );
and ( n49133 , n49060 , n49132 );
and ( n49134 , n49059 , n49133 );
and ( n49135 , n49058 , n49134 );
xor ( n49136 , n48638 , n49135 );
and ( n49137 , n49057 , n49136 );
and ( n49138 , n48610 , n48668 );
and ( n49139 , n48609 , n49138 );
and ( n49140 , n48608 , n49139 );
and ( n49141 , n48607 , n49140 );
and ( n49142 , n48606 , n49141 );
and ( n49143 , n48605 , n49142 );
and ( n49144 , n48604 , n49143 );
and ( n49145 , n48603 , n49144 );
and ( n49146 , n48602 , n49145 );
and ( n49147 , n48601 , n49146 );
and ( n49148 , n48600 , n49147 );
and ( n49149 , n48599 , n49148 );
and ( n49150 , n48598 , n49149 );
and ( n49151 , n48597 , n49150 );
and ( n49152 , n48596 , n49151 );
and ( n49153 , n48595 , n49152 );
and ( n49154 , n48594 , n49153 );
and ( n49155 , n48593 , n49154 );
and ( n49156 , n48592 , n49155 );
and ( n49157 , n48591 , n49156 );
and ( n49158 , n48590 , n49157 );
and ( n49159 , n48589 , n49158 );
and ( n49160 , n48588 , n49159 );
and ( n49161 , n48587 , n49160 );
and ( n49162 , n48586 , n49161 );
and ( n49163 , n48585 , n49162 );
and ( n49164 , n48584 , n49163 );
and ( n49165 , n48583 , n49164 );
xor ( n49166 , n48582 , n49165 );
xor ( n49167 , n48583 , n49164 );
xor ( n49168 , n48584 , n49163 );
xor ( n49169 , n48585 , n49162 );
xor ( n49170 , n48586 , n49161 );
xor ( n49171 , n48587 , n49160 );
xor ( n49172 , n48588 , n49159 );
xor ( n49173 , n48589 , n49158 );
xor ( n49174 , n48590 , n49157 );
xor ( n49175 , n48591 , n49156 );
xor ( n49176 , n48592 , n49155 );
xor ( n49177 , n48593 , n49154 );
xor ( n49178 , n48594 , n49153 );
xor ( n49179 , n48595 , n49152 );
xor ( n49180 , n48596 , n49151 );
xor ( n49181 , n48597 , n49150 );
xor ( n49182 , n48598 , n49149 );
xor ( n49183 , n48599 , n49148 );
xor ( n49184 , n48600 , n49147 );
xor ( n49185 , n48601 , n49146 );
xor ( n49186 , n48602 , n49145 );
xor ( n49187 , n48603 , n49144 );
xor ( n49188 , n48604 , n49143 );
not ( n49189 , n48845 );
not ( n49190 , n49189 );
and ( n49191 , n49188 , n49190 );
xor ( n49192 , n48605 , n49142 );
not ( n49193 , n48864 );
not ( n49194 , n49193 );
and ( n49195 , n49192 , n49194 );
xor ( n49196 , n48606 , n49141 );
not ( n49197 , n48883 );
not ( n49198 , n49197 );
and ( n49199 , n49196 , n49198 );
xor ( n49200 , n48607 , n49140 );
not ( n49201 , n48902 );
not ( n49202 , n49201 );
and ( n49203 , n49200 , n49202 );
xor ( n49204 , n48608 , n49139 );
not ( n49205 , n48921 );
not ( n49206 , n49205 );
and ( n49207 , n49204 , n49206 );
xor ( n49208 , n48609 , n49138 );
not ( n49209 , n48940 );
not ( n49210 , n49209 );
and ( n49211 , n49208 , n49210 );
xor ( n49212 , n48610 , n48668 );
not ( n49213 , n48959 );
not ( n49214 , n49213 );
and ( n49215 , n49212 , n49214 );
not ( n49216 , n48668 );
not ( n49217 , n48978 );
not ( n49218 , n49217 );
or ( n49219 , n49216 , n49218 );
and ( n49220 , n49214 , n49219 );
and ( n49221 , n49212 , n49219 );
or ( n49222 , n49215 , n49220 , n49221 );
and ( n49223 , n49210 , n49222 );
and ( n49224 , n49208 , n49222 );
or ( n49225 , n49211 , n49223 , n49224 );
and ( n49226 , n49206 , n49225 );
and ( n49227 , n49204 , n49225 );
or ( n49228 , n49207 , n49226 , n49227 );
and ( n49229 , n49202 , n49228 );
and ( n49230 , n49200 , n49228 );
or ( n49231 , n49203 , n49229 , n49230 );
and ( n49232 , n49198 , n49231 );
and ( n49233 , n49196 , n49231 );
or ( n49234 , n49199 , n49232 , n49233 );
and ( n49235 , n49194 , n49234 );
and ( n49236 , n49192 , n49234 );
or ( n49237 , n49195 , n49235 , n49236 );
and ( n49238 , n49190 , n49237 );
and ( n49239 , n49188 , n49237 );
or ( n49240 , n49191 , n49238 , n49239 );
or ( n49241 , n49187 , n49240 );
or ( n49242 , n49186 , n49241 );
or ( n49243 , n49185 , n49242 );
or ( n49244 , n49184 , n49243 );
or ( n49245 , n49183 , n49244 );
or ( n49246 , n49182 , n49245 );
or ( n49247 , n49181 , n49246 );
or ( n49248 , n49180 , n49247 );
or ( n49249 , n49179 , n49248 );
or ( n49250 , n49178 , n49249 );
or ( n49251 , n49177 , n49250 );
or ( n49252 , n49176 , n49251 );
or ( n49253 , n49175 , n49252 );
or ( n49254 , n49174 , n49253 );
or ( n49255 , n49173 , n49254 );
or ( n49256 , n49172 , n49255 );
or ( n49257 , n49171 , n49256 );
or ( n49258 , n49170 , n49257 );
or ( n49259 , n49169 , n49258 );
or ( n49260 , n49168 , n49259 );
or ( n49261 , n49167 , n49260 );
xnor ( n49262 , n49166 , n49261 );
and ( n49263 , n49262 , n48845 );
or ( n49264 , n49137 , n49263 );
and ( n49265 , n49264 , n49054 );
or ( n49266 , n49056 , n49265 );
and ( n49267 , n49266 , n33178 );
or ( n49268 , n33175 , n33174 );
or ( n49269 , n49268 , n33182 );
or ( n49270 , n49269 , n33185 );
or ( n49271 , n49270 , n33191 );
or ( n49272 , n49271 , n33193 );
or ( n49273 , n49272 , n33199 );
or ( n49274 , n49273 , n33201 );
or ( n49275 , n49274 , n33203 );
and ( n49276 , n49166 , n49275 );
or ( n49277 , n48640 , n48647 , n48653 , n48659 , n48665 , n48700 , n48735 , n49025 , n49267 , n49276 );
and ( n49278 , n49277 , n33208 );
and ( n49279 , n32975 , n35056 );
or ( n49280 , n33372 , n33370 );
or ( n49281 , n49280 , n33373 );
or ( n49282 , n49281 , n33375 );
or ( n49283 , n49282 , n33377 );
or ( n49284 , n49283 , n33379 );
or ( n49285 , n49284 , n33381 );
or ( n49286 , n49285 , n32528 );
and ( n49287 , n48582 , n49286 );
or ( n49288 , C0 , n49278 , n49279 , n49287 );
buf ( n49289 , n49288 );
buf ( n49290 , n49289 );
buf ( n49291 , n31655 );
buf ( n49292 , n30987 );
buf ( n49293 , n30987 );
buf ( n49294 , n31655 );
buf ( n49295 , n30987 );
not ( n49296 , n40163 );
and ( n49297 , n49296 , n32019 );
nor ( n49298 , n31673 , n42237 , n45160 , n31661 , n31657 );
not ( n49299 , n49298 );
and ( n49300 , n49299 , n32019 );
and ( n49301 , n32147 , n49298 );
or ( n49302 , n49300 , n49301 );
and ( n49303 , n49302 , n40163 );
or ( n49304 , n49297 , n49303 );
and ( n49305 , n49304 , n32498 );
nor ( n49306 , n40177 , n42246 , n45169 , n40194 , C0 );
not ( n49307 , n49306 );
not ( n49308 , n49298 );
and ( n49309 , n49308 , n32019 );
not ( n49310 , n40373 );
and ( n49311 , n49310 , n40261 );
xor ( n49312 , n40382 , n40384 );
and ( n49313 , n49312 , n40373 );
or ( n49314 , n49311 , n49313 );
and ( n49315 , n49314 , n49298 );
or ( n49316 , n49309 , n49315 );
and ( n49317 , n49307 , n49316 );
and ( n49318 , n49314 , n49306 );
or ( n49319 , n49317 , n49318 );
and ( n49320 , n49319 , n32473 );
not ( n49321 , n32475 );
not ( n49322 , n49306 );
not ( n49323 , n49298 );
and ( n49324 , n49323 , n32019 );
and ( n49325 , n49314 , n49298 );
or ( n49326 , n49324 , n49325 );
and ( n49327 , n49322 , n49326 );
and ( n49328 , n49314 , n49306 );
or ( n49329 , n49327 , n49328 );
and ( n49330 , n49321 , n49329 );
nor ( n49331 , n40417 , n42272 , n45195 , n40445 , C0 );
not ( n49332 , n49331 );
nor ( n49333 , n40413 , n42275 , n45198 , n40440 , C0 );
not ( n49334 , n49333 );
and ( n49335 , n49334 , n49329 );
not ( n49336 , n40952 );
and ( n49337 , n49336 , n40846 );
xor ( n49338 , n40961 , n40963 );
and ( n49339 , n49338 , n40952 );
or ( n49340 , n49337 , n49339 );
and ( n49341 , n49340 , n49333 );
or ( n49342 , n49335 , n49341 );
and ( n49343 , n49332 , n49342 );
not ( n49344 , n41247 );
and ( n49345 , n49344 , n41145 );
xor ( n49346 , n41256 , n41258 );
and ( n49347 , n49346 , n41247 );
or ( n49348 , n49345 , n49347 );
and ( n49349 , n49348 , n49331 );
or ( n49350 , n49343 , n49349 );
and ( n49351 , n49350 , n32475 );
or ( n49352 , n49330 , n49351 );
and ( n49353 , n49352 , n32486 );
and ( n49354 , n32019 , n41278 );
or ( n49355 , C0 , n49305 , n49320 , n49353 , n49354 );
buf ( n49356 , n49355 );
buf ( n49357 , n49356 );
buf ( n49358 , n30987 );
xor ( n49359 , n41795 , n44790 );
and ( n49360 , n49359 , n31548 );
not ( n49361 , n44807 );
and ( n49362 , n49361 , n41795 );
and ( n49363 , n42110 , n44807 );
or ( n49364 , n49362 , n49363 );
and ( n49365 , n49364 , n31408 );
not ( n49366 , n44817 );
and ( n49367 , n49366 , n41795 );
not ( n49368 , n41835 );
buf ( n49369 , RI15b532e0_703);
and ( n49370 , n49368 , n49369 );
not ( n49371 , n42124 );
and ( n49372 , n49371 , n42120 );
xor ( n49373 , n42120 , n41881 );
xor ( n49374 , n42104 , n41881 );
xor ( n49375 , n42088 , n41881 );
xor ( n49376 , n42072 , n41881 );
xor ( n49377 , n42056 , n41881 );
xor ( n49378 , n42040 , n41881 );
xor ( n49379 , n42024 , n41881 );
and ( n49380 , n42127 , n42143 );
and ( n49381 , n49379 , n49380 );
and ( n49382 , n49378 , n49381 );
and ( n49383 , n49377 , n49382 );
and ( n49384 , n49376 , n49383 );
and ( n49385 , n49375 , n49384 );
and ( n49386 , n49374 , n49385 );
xor ( n49387 , n49373 , n49386 );
and ( n49388 , n49387 , n42124 );
or ( n49389 , n49372 , n49388 );
and ( n49390 , n49389 , n41835 );
or ( n49391 , n49370 , n49390 );
and ( n49392 , n49391 , n44817 );
or ( n49393 , n49367 , n49392 );
and ( n49394 , n49393 , n31521 );
not ( n49395 , n45059 );
and ( n49396 , n49395 , n41795 );
and ( n49397 , n31340 , n42330 );
and ( n49398 , n31342 , n42332 );
and ( n49399 , n31344 , n42334 );
and ( n49400 , n31346 , n42336 );
and ( n49401 , n31348 , n42338 );
and ( n49402 , n31350 , n42340 );
and ( n49403 , n31352 , n42342 );
and ( n49404 , n31354 , n42344 );
and ( n49405 , n31356 , n42346 );
and ( n49406 , n31358 , n42348 );
and ( n49407 , n31360 , n42350 );
and ( n49408 , n31362 , n42352 );
and ( n49409 , n31364 , n42354 );
and ( n49410 , n31366 , n42356 );
and ( n49411 , n31368 , n42358 );
and ( n49412 , n31370 , n42360 );
or ( n49413 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 );
and ( n49414 , n49413 , n45059 );
or ( n49415 , n49396 , n49414 );
and ( n49416 , n49415 , n31536 );
and ( n49417 , n41795 , n45148 );
or ( n49418 , n49360 , n49365 , n49394 , n49416 , n49417 );
and ( n49419 , n49418 , n31557 );
and ( n49420 , n41795 , n40154 );
or ( n49421 , C0 , n49419 , n49420 );
buf ( n49422 , n49421 );
buf ( n49423 , n49422 );
buf ( n49424 , n31655 );
not ( n49425 , n46356 );
and ( n49426 , n49425 , n31264 );
nor ( n49427 , n46359 , n46360 , n31017 , n31013 , n31009 );
not ( n49428 , n49427 );
and ( n49429 , n49428 , n31264 );
and ( n49430 , n31272 , n49427 );
or ( n49431 , n49429 , n49430 );
and ( n49432 , n49431 , n46356 );
or ( n49433 , n49426 , n49432 );
and ( n49434 , n49433 , n31649 );
nor ( n49435 , n46374 , n46380 , n46386 , n46392 , C0 );
not ( n49436 , n49435 );
not ( n49437 , n49427 );
and ( n49438 , n49437 , n31264 );
not ( n49439 , n46487 );
and ( n49440 , n49439 , n46447 );
xor ( n49441 , n47439 , n47444 );
and ( n49442 , n49441 , n46487 );
or ( n49443 , n49440 , n49442 );
and ( n49444 , n49443 , n49427 );
or ( n49445 , n49438 , n49444 );
and ( n49446 , n49436 , n49445 );
and ( n49447 , n49443 , n49435 );
or ( n49448 , n49446 , n49447 );
and ( n49449 , n49448 , n31643 );
not ( n49450 , n31452 );
not ( n49451 , n49435 );
not ( n49452 , n49427 );
and ( n49453 , n49452 , n31264 );
and ( n49454 , n49443 , n49427 );
or ( n49455 , n49453 , n49454 );
and ( n49456 , n49451 , n49455 );
and ( n49457 , n49443 , n49435 );
or ( n49458 , n49456 , n49457 );
and ( n49459 , n49450 , n49458 );
nor ( n49460 , n46520 , n46529 , n46539 , n46549 , C0 );
not ( n49461 , n49460 );
nor ( n49462 , n46552 , n46553 , n46534 , n46544 , C0 );
not ( n49463 , n49462 );
and ( n49464 , n49463 , n49458 );
not ( n49465 , n46976 );
and ( n49466 , n49465 , n46921 );
xor ( n49467 , n47475 , n47480 );
and ( n49468 , n49467 , n46976 );
or ( n49469 , n49466 , n49468 );
and ( n49470 , n49469 , n49462 );
or ( n49471 , n49464 , n49470 );
and ( n49472 , n49461 , n49471 );
not ( n49473 , n47259 );
and ( n49474 , n49473 , n47208 );
xor ( n49475 , n47493 , n47498 );
and ( n49476 , n49475 , n47259 );
or ( n49477 , n49474 , n49476 );
and ( n49478 , n49477 , n49460 );
or ( n49479 , n49472 , n49478 );
and ( n49480 , n49479 , n31452 );
or ( n49481 , n49459 , n49480 );
and ( n49482 , n49481 , n31638 );
and ( n49483 , n31264 , n47277 );
or ( n49484 , C0 , n49434 , n49449 , n49482 , n49483 );
buf ( n49485 , n49484 );
buf ( n49486 , n49485 );
buf ( n49487 , n40201 );
xor ( n49488 , n47289 , n47293 );
and ( n49489 , n49488 , n32433 );
not ( n49490 , n47331 );
and ( n49491 , n49490 , n47289 );
buf ( n49492 , n31926 );
and ( n49493 , n49492 , n47331 );
or ( n49494 , n49491 , n49493 );
and ( n49495 , n49494 , n32413 );
and ( n49496 , n47289 , n47402 );
or ( n49497 , n49489 , n49495 , n49496 );
and ( n49498 , n49497 , n32456 );
and ( n49499 , n47289 , n47409 );
or ( n49500 , C0 , n49498 , n49499 );
buf ( n49501 , n49500 );
buf ( n49502 , n49501 );
buf ( n49503 , n31655 );
buf ( n49504 , n31655 );
buf ( n49505 , n30987 );
buf ( n49506 , n31655 );
buf ( n49507 , n30987 );
buf ( n49508 , n30987 );
and ( n49509 , n46017 , n32500 );
not ( n49510 , n35211 );
and ( n49511 , n49510 , n37531 );
buf ( n49512 , n49511 );
and ( n49513 , n49512 , n32421 );
not ( n49514 , n35245 );
and ( n49515 , n49514 , n37531 );
buf ( n49516 , n49515 );
and ( n49517 , n49516 , n32419 );
not ( n49518 , n35278 );
and ( n49519 , n49518 , n37531 );
not ( n49520 , n35295 );
buf ( n49521 , RI15b62a60_1231);
and ( n49522 , n49520 , n49521 );
and ( n49523 , n37585 , n37514 );
and ( n49524 , n37583 , n49523 );
and ( n49525 , n37581 , n49524 );
and ( n49526 , n37579 , n49525 );
and ( n49527 , n37577 , n49526 );
and ( n49528 , n35677 , n49527 );
and ( n49529 , n32488 , n49528 );
and ( n49530 , n37573 , n49529 );
and ( n49531 , n37571 , n49530 );
and ( n49532 , n37569 , n49531 );
and ( n49533 , n37567 , n49532 );
and ( n49534 , n37565 , n49533 );
and ( n49535 , n37563 , n49534 );
and ( n49536 , n37561 , n49535 );
and ( n49537 , n37559 , n49536 );
and ( n49538 , n37557 , n49537 );
and ( n49539 , n37555 , n49538 );
and ( n49540 , n37553 , n49539 );
and ( n49541 , n37551 , n49540 );
and ( n49542 , n37549 , n49541 );
and ( n49543 , n37547 , n49542 );
and ( n49544 , n37545 , n49543 );
and ( n49545 , n37543 , n49544 );
and ( n49546 , n37541 , n49545 );
and ( n49547 , n37539 , n49546 );
and ( n49548 , n37537 , n49547 );
and ( n49549 , n37535 , n49548 );
and ( n49550 , n37533 , n49549 );
xor ( n49551 , n37531 , n49550 );
and ( n49552 , n49551 , n35295 );
or ( n49553 , n49522 , n49552 );
and ( n49554 , n49553 , n35278 );
or ( n49555 , n49519 , n49554 );
and ( n49556 , n49555 , n32417 );
not ( n49557 , n35331 );
and ( n49558 , n49557 , n37531 );
not ( n49559 , n35294 );
not ( n49560 , n45995 );
and ( n49561 , n49560 , n49521 );
not ( n49562 , n49521 );
buf ( n49563 , RI15b629e8_1230);
not ( n49564 , n49563 );
buf ( n49565 , RI15b62970_1229);
not ( n49566 , n49565 );
buf ( n49567 , RI15b628f8_1228);
not ( n49568 , n49567 );
buf ( n49569 , RI15b62880_1227);
not ( n49570 , n49569 );
buf ( n49571 , RI15b62808_1226);
not ( n49572 , n49571 );
buf ( n49573 , RI15b62790_1225);
not ( n49574 , n49573 );
buf ( n49575 , RI15b62718_1224);
not ( n49576 , n49575 );
buf ( n49577 , RI15b626a0_1223);
not ( n49578 , n49577 );
buf ( n49579 , RI15b62628_1222);
not ( n49580 , n49579 );
buf ( n49581 , RI15b625b0_1221);
not ( n49582 , n49581 );
buf ( n49583 , RI15b62538_1220);
not ( n49584 , n49583 );
buf ( n49585 , RI15b624c0_1219);
not ( n49586 , n49585 );
buf ( n49587 , RI15b62448_1218);
not ( n49588 , n49587 );
buf ( n49589 , RI15b623d0_1217);
not ( n49590 , n49589 );
buf ( n49591 , RI15b62358_1216);
not ( n49592 , n49591 );
buf ( n49593 , RI15b622e0_1215);
not ( n49594 , n49593 );
buf ( n49595 , RI15b62268_1214);
not ( n49596 , n49595 );
buf ( n49597 , RI15b621f0_1213);
not ( n49598 , n49597 );
buf ( n49599 , RI15b62178_1212);
not ( n49600 , n49599 );
not ( n49601 , n47283 );
not ( n49602 , n47284 );
not ( n49603 , n47285 );
not ( n49604 , n47286 );
not ( n49605 , n47287 );
not ( n49606 , n47288 );
not ( n49607 , n47289 );
not ( n49608 , n47290 );
and ( n49609 , n45998 , n46002 );
and ( n49610 , n49608 , n49609 );
and ( n49611 , n49607 , n49610 );
and ( n49612 , n49606 , n49611 );
and ( n49613 , n49605 , n49612 );
and ( n49614 , n49604 , n49613 );
and ( n49615 , n49603 , n49614 );
and ( n49616 , n49602 , n49615 );
and ( n49617 , n49601 , n49616 );
and ( n49618 , n49600 , n49617 );
and ( n49619 , n49598 , n49618 );
and ( n49620 , n49596 , n49619 );
and ( n49621 , n49594 , n49620 );
and ( n49622 , n49592 , n49621 );
and ( n49623 , n49590 , n49622 );
and ( n49624 , n49588 , n49623 );
and ( n49625 , n49586 , n49624 );
and ( n49626 , n49584 , n49625 );
and ( n49627 , n49582 , n49626 );
and ( n49628 , n49580 , n49627 );
and ( n49629 , n49578 , n49628 );
and ( n49630 , n49576 , n49629 );
and ( n49631 , n49574 , n49630 );
and ( n49632 , n49572 , n49631 );
and ( n49633 , n49570 , n49632 );
and ( n49634 , n49568 , n49633 );
and ( n49635 , n49566 , n49634 );
and ( n49636 , n49564 , n49635 );
xor ( n49637 , n49562 , n49636 );
and ( n49638 , n49637 , n45995 );
or ( n49639 , n49561 , n49638 );
and ( n49640 , n49559 , n49639 );
and ( n49641 , n49551 , n35294 );
or ( n49642 , n49640 , n49641 );
and ( n49643 , n49642 , n35331 );
or ( n49644 , n49558 , n49643 );
and ( n49645 , n49644 , n32415 );
and ( n49646 , n37531 , n35354 );
or ( n49647 , n49513 , n49517 , n49556 , n49645 , n49646 );
and ( n49648 , n49647 , n32456 );
not ( n49649 , n32475 );
not ( n49650 , n46060 );
xor ( n49651 , n46017 , n46058 );
and ( n49652 , n49650 , n49651 );
not ( n49653 , n49651 );
xor ( n49654 , n46018 , n46057 );
not ( n49655 , n49654 );
xor ( n49656 , n46019 , n46056 );
not ( n49657 , n49656 );
xor ( n49658 , n46020 , n46055 );
not ( n49659 , n49658 );
xor ( n49660 , n46021 , n46054 );
not ( n49661 , n49660 );
not ( n49662 , n47745 );
xor ( n49663 , n46023 , n46052 );
not ( n49664 , n49663 );
xor ( n49665 , n46024 , n46051 );
not ( n49666 , n49665 );
xor ( n49667 , n46025 , n46050 );
not ( n49668 , n49667 );
xor ( n49669 , n46026 , n46049 );
not ( n49670 , n49669 );
xor ( n49671 , n46027 , n46048 );
not ( n49672 , n49671 );
xor ( n49673 , n46028 , n46047 );
not ( n49674 , n49673 );
xor ( n49675 , n46029 , n46046 );
not ( n49676 , n49675 );
xor ( n49677 , n46030 , n46045 );
not ( n49678 , n49677 );
xor ( n49679 , n46031 , n46044 );
not ( n49680 , n49679 );
xor ( n49681 , n46032 , n46043 );
not ( n49682 , n49681 );
xor ( n49683 , n46033 , n46042 );
not ( n49684 , n49683 );
xor ( n49685 , n46034 , n46041 );
not ( n49686 , n49685 );
xor ( n49687 , n46035 , n46040 );
not ( n49688 , n49687 );
xor ( n49689 , n46036 , n46039 );
not ( n49690 , n49689 );
xor ( n49691 , n46037 , n46038 );
not ( n49692 , n49691 );
not ( n49693 , n41315 );
not ( n49694 , n32471 );
not ( n49695 , n35669 );
not ( n49696 , n44750 );
xor ( n49697 , n32460 , n32467 );
not ( n49698 , n49697 );
xor ( n49699 , n32461 , n32466 );
not ( n49700 , n49699 );
xor ( n49701 , n32462 , n32465 );
not ( n49702 , n49701 );
and ( n49703 , n46064 , n46068 );
and ( n49704 , n49702 , n49703 );
and ( n49705 , n49700 , n49704 );
and ( n49706 , n49698 , n49705 );
and ( n49707 , n49696 , n49706 );
and ( n49708 , n49695 , n49707 );
and ( n49709 , n49694 , n49708 );
and ( n49710 , n49693 , n49709 );
and ( n49711 , n49692 , n49710 );
and ( n49712 , n49690 , n49711 );
and ( n49713 , n49688 , n49712 );
and ( n49714 , n49686 , n49713 );
and ( n49715 , n49684 , n49714 );
and ( n49716 , n49682 , n49715 );
and ( n49717 , n49680 , n49716 );
and ( n49718 , n49678 , n49717 );
and ( n49719 , n49676 , n49718 );
and ( n49720 , n49674 , n49719 );
and ( n49721 , n49672 , n49720 );
and ( n49722 , n49670 , n49721 );
and ( n49723 , n49668 , n49722 );
and ( n49724 , n49666 , n49723 );
and ( n49725 , n49664 , n49724 );
and ( n49726 , n49662 , n49725 );
and ( n49727 , n49661 , n49726 );
and ( n49728 , n49659 , n49727 );
and ( n49729 , n49657 , n49728 );
and ( n49730 , n49655 , n49729 );
xor ( n49731 , n49653 , n49730 );
and ( n49732 , n49731 , n46060 );
or ( n49733 , n49652 , n49732 );
and ( n49734 , n49649 , n49733 );
and ( n49735 , n37531 , n32475 );
or ( n49736 , n49734 , n49735 );
and ( n49737 , n49736 , n32486 );
and ( n49738 , n37531 , n35367 );
or ( n49739 , C0 , n49509 , n49648 , n49737 , C0 , n49738 );
buf ( n49740 , n49739 );
buf ( n49741 , n49740 );
buf ( n49742 , n31655 );
not ( n49743 , n48765 );
and ( n49744 , n49743 , n33233 );
xor ( n49745 , n48788 , n49000 );
and ( n49746 , n49745 , n48765 );
or ( n49747 , n49744 , n49746 );
and ( n49748 , n49747 , n33180 );
not ( n49749 , n49054 );
and ( n49750 , n49749 , n33233 );
not ( n49751 , n48845 );
xor ( n49752 , n49078 , n49114 );
and ( n49753 , n49751 , n49752 );
xnor ( n49754 , n49187 , n49240 );
and ( n49755 , n49754 , n48845 );
or ( n49756 , n49753 , n49755 );
and ( n49757 , n49756 , n49054 );
or ( n49758 , n49750 , n49757 );
and ( n49759 , n49758 , n33178 );
or ( n49760 , n33176 , n33182 );
or ( n49761 , n49760 , n33185 );
or ( n49762 , n49761 , n33187 );
or ( n49763 , n49762 , n33189 );
or ( n49764 , n49763 , n33172 );
or ( n49765 , n49764 , n33038 );
or ( n49766 , n49765 , n32924 );
or ( n49767 , n49766 , n32890 );
or ( n49768 , n49767 , n33191 );
or ( n49769 , n49768 , n33193 );
or ( n49770 , n49769 , n33195 );
or ( n49771 , n49770 , n33197 );
or ( n49772 , n49771 , n33199 );
or ( n49773 , n49772 , n33201 );
or ( n49774 , n49773 , n33203 );
and ( n49775 , n33233 , n49774 );
or ( n49776 , n49748 , n49759 , n49775 );
and ( n49777 , n49776 , n33208 );
and ( n49778 , n33317 , n33375 );
not ( n49779 , n32968 );
and ( n49780 , n49779 , n33317 );
and ( n49781 , n33238 , n33239 );
and ( n49782 , n33237 , n49781 );
and ( n49783 , n33236 , n49782 );
and ( n49784 , n33235 , n49783 );
and ( n49785 , n33234 , n49784 );
xor ( n49786 , n33233 , n49785 );
and ( n49787 , n49786 , n32968 );
or ( n49788 , n49780 , n49787 );
and ( n49789 , n49788 , n33370 );
and ( n49790 , n32996 , n35056 );
or ( n49791 , n33374 , n33377 );
or ( n49792 , n49791 , n33379 );
or ( n49793 , n49792 , n33381 );
or ( n49794 , n49793 , n32528 );
and ( n49795 , n33233 , n49794 );
or ( n49796 , C0 , n49777 , n49778 , n49789 , n49790 , n49795 );
buf ( n49797 , n49796 );
buf ( n49798 , n49797 );
not ( n49799 , n31728 );
and ( n49800 , n49799 , n46037 );
xor ( n49801 , n47614 , n47615 );
and ( n49802 , n49801 , n31728 );
or ( n49803 , n49800 , n49802 );
and ( n49804 , n49803 , n32253 );
not ( n49805 , n32283 );
and ( n49806 , n49805 , n46037 );
not ( n49807 , n31823 );
xor ( n49808 , n47669 , n47670 );
and ( n49809 , n49807 , n49808 );
xnor ( n49810 , n47719 , n47720 );
and ( n49811 , n49810 , n31823 );
or ( n49812 , n49809 , n49811 );
and ( n49813 , n49812 , n32283 );
or ( n49814 , n49806 , n49813 );
and ( n49815 , n49814 , n32398 );
and ( n49816 , n46037 , n32436 );
or ( n49817 , n49804 , n49815 , n49816 );
and ( n49818 , n49817 , n32456 );
and ( n49819 , n49691 , n32473 );
not ( n49820 , n32475 );
and ( n49821 , n49820 , n49691 );
xor ( n49822 , n46037 , n47749 );
and ( n49823 , n49822 , n32475 );
or ( n49824 , n49821 , n49823 );
and ( n49825 , n49824 , n32486 );
and ( n49826 , n37571 , n32489 );
and ( n49827 , n46037 , n32501 );
or ( n49828 , C0 , n49818 , n49819 , n49825 , n49826 , n49827 );
buf ( n49829 , n49828 );
buf ( n49830 , n49829 );
buf ( n49831 , n31655 );
buf ( n49832 , n30987 );
and ( n49833 , n33213 , n32528 );
not ( n49834 , n32598 );
and ( n49835 , n49834 , n32976 );
buf ( n49836 , n49835 );
and ( n49837 , n49836 , n32890 );
not ( n49838 , n32919 );
and ( n49839 , n49838 , n32976 );
buf ( n49840 , n49839 );
and ( n49841 , n49840 , n32924 );
not ( n49842 , n32953 );
and ( n49843 , n49842 , n32976 );
not ( n49844 , n32971 );
and ( n49845 , n49844 , n33077 );
xor ( n49846 , n32976 , n33029 );
and ( n49847 , n49846 , n32971 );
or ( n49848 , n49845 , n49847 );
and ( n49849 , n49848 , n32953 );
or ( n49850 , n49843 , n49849 );
and ( n49851 , n49850 , n33038 );
not ( n49852 , n33067 );
and ( n49853 , n49852 , n32976 );
not ( n49854 , n32970 );
not ( n49855 , n33071 );
and ( n49856 , n49855 , n33077 );
xor ( n49857 , n33078 , n33161 );
and ( n49858 , n49857 , n33071 );
or ( n49859 , n49856 , n49858 );
and ( n49860 , n49854 , n49859 );
and ( n49861 , n49846 , n32970 );
or ( n49862 , n49860 , n49861 );
and ( n49863 , n49862 , n33067 );
or ( n49864 , n49853 , n49863 );
and ( n49865 , n49864 , n33172 );
and ( n49866 , n32976 , n33204 );
or ( n49867 , n49837 , n49841 , n49851 , n49865 , n49866 );
and ( n49868 , n49867 , n33208 );
not ( n49869 , n32968 );
not ( n49870 , n33270 );
and ( n49871 , n49870 , n33277 );
xor ( n49872 , n33278 , n33361 );
and ( n49873 , n49872 , n33270 );
or ( n49874 , n49871 , n49873 );
and ( n49875 , n49869 , n49874 );
and ( n49876 , n32976 , n32968 );
or ( n49877 , n49875 , n49876 );
and ( n49878 , n49877 , n33370 );
and ( n49879 , n32976 , n33382 );
or ( n49880 , C0 , n49833 , n49868 , n49878 , C0 , n49879 );
buf ( n49881 , n49880 );
buf ( n49882 , n49881 );
buf ( n49883 , n30987 );
buf ( n49884 , n31655 );
not ( n49885 , n46356 );
and ( n49886 , n49885 , n31220 );
not ( n49887 , n48214 );
and ( n49888 , n49887 , n31220 );
and ( n49889 , n31238 , n48214 );
or ( n49890 , n49888 , n49889 );
and ( n49891 , n49890 , n46356 );
or ( n49892 , n49886 , n49891 );
and ( n49893 , n49892 , n31649 );
not ( n49894 , n48223 );
not ( n49895 , n48214 );
and ( n49896 , n49895 , n31220 );
not ( n49897 , n46487 );
and ( n49898 , n49897 , n46435 );
xor ( n49899 , n47440 , n47443 );
and ( n49900 , n49899 , n46487 );
or ( n49901 , n49898 , n49900 );
and ( n49902 , n49901 , n48214 );
or ( n49903 , n49896 , n49902 );
and ( n49904 , n49894 , n49903 );
and ( n49905 , n49901 , n48223 );
or ( n49906 , n49904 , n49905 );
and ( n49907 , n49906 , n31643 );
not ( n49908 , n31452 );
not ( n49909 , n48223 );
not ( n49910 , n48214 );
and ( n49911 , n49910 , n31220 );
and ( n49912 , n49901 , n48214 );
or ( n49913 , n49911 , n49912 );
and ( n49914 , n49909 , n49913 );
and ( n49915 , n49901 , n48223 );
or ( n49916 , n49914 , n49915 );
and ( n49917 , n49908 , n49916 );
not ( n49918 , n48244 );
not ( n49919 , n48247 );
and ( n49920 , n49919 , n49916 );
not ( n49921 , n46976 );
and ( n49922 , n49921 , n46904 );
xor ( n49923 , n47476 , n47479 );
and ( n49924 , n49923 , n46976 );
or ( n49925 , n49922 , n49924 );
and ( n49926 , n49925 , n48247 );
or ( n49927 , n49920 , n49926 );
and ( n49928 , n49918 , n49927 );
not ( n49929 , n47259 );
and ( n49930 , n49929 , n47191 );
xor ( n49931 , n47494 , n47497 );
and ( n49932 , n49931 , n47259 );
or ( n49933 , n49930 , n49932 );
and ( n49934 , n49933 , n48244 );
or ( n49935 , n49928 , n49934 );
and ( n49936 , n49935 , n31452 );
or ( n49937 , n49917 , n49936 );
and ( n49938 , n49937 , n31638 );
and ( n49939 , n31220 , n47277 );
or ( n49940 , C0 , n49893 , n49907 , n49938 , n49939 );
buf ( n49941 , n49940 );
buf ( n49942 , n49941 );
buf ( n49943 , n31655 );
buf ( n49944 , n30987 );
buf ( n49945 , n31655 );
not ( n49946 , n48267 );
not ( n49947 , n48269 );
not ( n49948 , n48272 );
and ( n49949 , n49947 , n49948 );
buf ( n49950 , n48269 );
or ( n49951 , n49949 , n49950 );
and ( n49952 , n49946 , n49951 );
buf ( n49953 , n49952 );
and ( n49954 , n49953 , n39358 );
not ( n49955 , n48287 );
and ( n49956 , n49955 , n39356 );
not ( n49957 , n48297 );
not ( n49958 , n48300 );
and ( n49959 , n49958 , n48294 );
buf ( n49960 , n48300 );
or ( n49961 , n49959 , n49960 );
and ( n49962 , n49957 , n49961 );
buf ( n49963 , n49962 );
and ( n49964 , n49963 , n39354 );
not ( n49965 , n48272 );
not ( n49966 , n48311 );
not ( n49967 , n48315 );
not ( n49968 , n48318 );
and ( n49969 , n49967 , n49968 );
buf ( n49970 , n48315 );
or ( n49971 , n49969 , n49970 );
and ( n49972 , n49966 , n49971 );
and ( n49973 , n35281 , n48311 );
or ( n49974 , n49972 , n49973 );
and ( n49975 , n49965 , n49974 );
buf ( n49976 , n49975 );
and ( n49977 , n49976 , n39352 );
buf ( n49978 , n39346 );
not ( n49979 , n48263 );
and ( n49980 , n49979 , n39349 );
buf ( n49981 , n39350 );
or ( n49982 , n49954 , C0 , n49956 , n49964 , n49977 , n49978 , n49980 , n49981 );
buf ( n49983 , n49982 );
buf ( n49984 , n49983 );
buf ( n49985 , n31655 );
buf ( n49986 , n30987 );
and ( n49987 , n46094 , n46087 );
and ( n49988 , n46107 , n49987 );
and ( n49989 , n46120 , n49988 );
and ( n49990 , n46133 , n49989 );
and ( n49991 , n46146 , n49990 );
and ( n49992 , n46159 , n49991 );
and ( n49993 , n46172 , n49992 );
and ( n49994 , n46185 , n49993 );
and ( n49995 , n46198 , n49994 );
and ( n49996 , n46211 , n49995 );
and ( n49997 , n46224 , n49996 );
and ( n49998 , n46237 , n49997 );
and ( n49999 , n46250 , n49998 );
xor ( n50000 , n46263 , n49999 );
and ( n50001 , n50000 , n32431 );
and ( n50002 , n35245 , n35292 );
not ( n50003 , n50002 );
and ( n50004 , n50003 , n46263 );
and ( n50005 , n40472 , n50002 );
or ( n50006 , n50004 , n50005 );
and ( n50007 , n50006 , n32419 );
and ( n50008 , n35331 , n35292 );
not ( n50009 , n50008 );
and ( n50010 , n50009 , n46263 );
not ( n50011 , n47910 );
buf ( n50012 , RI15b5f6d0_1121);
and ( n50013 , n50011 , n50012 );
not ( n50014 , n48101 );
and ( n50015 , n50014 , n48085 );
xor ( n50016 , n48085 , n40244 );
xor ( n50017 , n48073 , n40244 );
xor ( n50018 , n48061 , n40244 );
xor ( n50019 , n48049 , n40244 );
xor ( n50020 , n48037 , n40244 );
xor ( n50021 , n48025 , n40244 );
xor ( n50022 , n48013 , n40244 );
and ( n50023 , n48104 , n48118 );
and ( n50024 , n50022 , n50023 );
and ( n50025 , n50021 , n50024 );
and ( n50026 , n50020 , n50025 );
and ( n50027 , n50019 , n50026 );
and ( n50028 , n50018 , n50027 );
and ( n50029 , n50017 , n50028 );
xor ( n50030 , n50016 , n50029 );
and ( n50031 , n50030 , n48101 );
or ( n50032 , n50015 , n50031 );
and ( n50033 , n50032 , n47910 );
or ( n50034 , n50013 , n50033 );
and ( n50035 , n50034 , n50008 );
or ( n50036 , n50010 , n50035 );
and ( n50037 , n50036 , n32415 );
not ( n50038 , n31689 );
buf ( n50039 , n31689 );
buf ( n50040 , n31689 );
buf ( n50041 , n31689 );
buf ( n50042 , n31689 );
buf ( n50043 , n31689 );
buf ( n50044 , n31689 );
buf ( n50045 , n31689 );
buf ( n50046 , n31689 );
buf ( n50047 , n31689 );
buf ( n50048 , n31689 );
buf ( n50049 , n31689 );
buf ( n50050 , n31689 );
buf ( n50051 , n31689 );
buf ( n50052 , n31689 );
buf ( n50053 , n31689 );
buf ( n50054 , n31689 );
buf ( n50055 , n31689 );
buf ( n50056 , n31689 );
buf ( n50057 , n31689 );
buf ( n50058 , n31689 );
buf ( n50059 , n31689 );
buf ( n50060 , n31689 );
buf ( n50061 , n31689 );
buf ( n50062 , n31689 );
buf ( n50063 , n31689 );
or ( n50064 , n31723 , n31724 );
and ( n50065 , n31721 , n50064 );
or ( n50066 , n31692 , n31694 , n31689 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50065 );
and ( n50067 , n50038 , n50066 );
not ( n50068 , n50067 );
and ( n50069 , n50068 , n46263 );
and ( n50070 , n31826 , n47357 );
and ( n50071 , n31828 , n47359 );
and ( n50072 , n31830 , n47361 );
and ( n50073 , n31832 , n47363 );
and ( n50074 , n31834 , n47365 );
and ( n50075 , n31836 , n47367 );
and ( n50076 , n31838 , n47369 );
and ( n50077 , n31840 , n47371 );
and ( n50078 , n31842 , n47373 );
and ( n50079 , n31844 , n47375 );
and ( n50080 , n31846 , n47377 );
and ( n50081 , n31848 , n47379 );
and ( n50082 , n31850 , n47381 );
and ( n50083 , n31852 , n47383 );
and ( n50084 , n31854 , n47385 );
and ( n50085 , n31856 , n47387 );
or ( n50086 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 );
and ( n50087 , n50086 , n50067 );
or ( n50088 , n50069 , n50087 );
and ( n50089 , n50088 , n32411 );
or ( n50090 , n35345 , n32413 );
or ( n50091 , n50090 , n32417 );
or ( n50092 , n50091 , n32421 );
or ( n50093 , n50092 , n32423 );
or ( n50094 , n50093 , n32425 );
or ( n50095 , n50094 , n32427 );
or ( n50096 , n50095 , n32429 );
or ( n50097 , n50096 , n32433 );
or ( n50098 , n50097 , n32435 );
and ( n50099 , n46263 , n50098 );
or ( n50100 , n50001 , n50007 , n50037 , n50089 , n50099 );
and ( n50101 , n50100 , n32456 );
and ( n50102 , n46263 , n47409 );
or ( n50103 , C0 , n50101 , n50102 );
buf ( n50104 , n50103 );
buf ( n50105 , n50104 );
buf ( n50106 , n31655 );
not ( n50107 , n46356 );
and ( n50108 , n50107 , n31191 );
nor ( n50109 , n31025 , n46360 , n48213 , n31013 , n31009 );
not ( n50110 , n50109 );
and ( n50111 , n50110 , n31191 );
and ( n50112 , n31205 , n50109 );
or ( n50113 , n50111 , n50112 );
and ( n50114 , n50113 , n46356 );
or ( n50115 , n50108 , n50114 );
and ( n50116 , n50115 , n31649 );
nor ( n50117 , n46373 , n46380 , n48222 , n46392 , C0 );
not ( n50118 , n50117 );
not ( n50119 , n50109 );
and ( n50120 , n50119 , n31191 );
not ( n50121 , n46487 );
and ( n50122 , n50121 , n46423 );
xor ( n50123 , n47441 , n47442 );
and ( n50124 , n50123 , n46487 );
or ( n50125 , n50122 , n50124 );
and ( n50126 , n50125 , n50109 );
or ( n50127 , n50120 , n50126 );
and ( n50128 , n50118 , n50127 );
and ( n50129 , n50125 , n50117 );
or ( n50130 , n50128 , n50129 );
and ( n50131 , n50130 , n31643 );
not ( n50132 , n31452 );
not ( n50133 , n50117 );
not ( n50134 , n50109 );
and ( n50135 , n50134 , n31191 );
and ( n50136 , n50125 , n50109 );
or ( n50137 , n50135 , n50136 );
and ( n50138 , n50133 , n50137 );
and ( n50139 , n50125 , n50117 );
or ( n50140 , n50138 , n50139 );
and ( n50141 , n50132 , n50140 );
nor ( n50142 , n46519 , n46529 , n48243 , n46549 , C0 );
not ( n50143 , n50142 );
nor ( n50144 , n46515 , n46553 , n48246 , n46544 , C0 );
not ( n50145 , n50144 );
and ( n50146 , n50145 , n50140 );
not ( n50147 , n46976 );
and ( n50148 , n50147 , n46887 );
xor ( n50149 , n47477 , n47478 );
and ( n50150 , n50149 , n46976 );
or ( n50151 , n50148 , n50150 );
and ( n50152 , n50151 , n50144 );
or ( n50153 , n50146 , n50152 );
and ( n50154 , n50143 , n50153 );
not ( n50155 , n47259 );
and ( n50156 , n50155 , n47174 );
xor ( n50157 , n47495 , n47496 );
and ( n50158 , n50157 , n47259 );
or ( n50159 , n50156 , n50158 );
and ( n50160 , n50159 , n50142 );
or ( n50161 , n50154 , n50160 );
and ( n50162 , n50161 , n31452 );
or ( n50163 , n50141 , n50162 );
and ( n50164 , n50163 , n31638 );
and ( n50165 , n31191 , n47277 );
or ( n50166 , C0 , n50116 , n50131 , n50164 , n50165 );
buf ( n50167 , n50166 );
buf ( n50168 , n50167 );
buf ( n50169 , n30987 );
not ( n50170 , n36587 );
and ( n50171 , n50170 , n36481 );
xor ( n50172 , n36481 , n36091 );
xor ( n50173 , n36464 , n36091 );
xor ( n50174 , n36447 , n36091 );
xor ( n50175 , n36430 , n36091 );
xor ( n50176 , n36413 , n36091 );
xor ( n50177 , n36396 , n36091 );
xor ( n50178 , n36379 , n36091 );
xor ( n50179 , n36362 , n36091 );
xor ( n50180 , n36345 , n36091 );
xor ( n50181 , n36328 , n36091 );
xor ( n50182 , n36311 , n36091 );
xor ( n50183 , n36294 , n36091 );
xor ( n50184 , n36277 , n36091 );
xor ( n50185 , n36260 , n36091 );
xor ( n50186 , n36243 , n36091 );
xor ( n50187 , n36226 , n36091 );
xor ( n50188 , n36209 , n36091 );
xor ( n50189 , n36192 , n36091 );
xor ( n50190 , n36175 , n36091 );
xor ( n50191 , n36158 , n36091 );
xor ( n50192 , n36141 , n36091 );
xor ( n50193 , n36124 , n36091 );
and ( n50194 , n36590 , n36592 );
and ( n50195 , n50193 , n50194 );
and ( n50196 , n50192 , n50195 );
and ( n50197 , n50191 , n50196 );
and ( n50198 , n50190 , n50197 );
and ( n50199 , n50189 , n50198 );
and ( n50200 , n50188 , n50199 );
and ( n50201 , n50187 , n50200 );
and ( n50202 , n50186 , n50201 );
and ( n50203 , n50185 , n50202 );
and ( n50204 , n50184 , n50203 );
and ( n50205 , n50183 , n50204 );
and ( n50206 , n50182 , n50205 );
and ( n50207 , n50181 , n50206 );
and ( n50208 , n50180 , n50207 );
and ( n50209 , n50179 , n50208 );
and ( n50210 , n50178 , n50209 );
and ( n50211 , n50177 , n50210 );
and ( n50212 , n50176 , n50211 );
and ( n50213 , n50175 , n50212 );
and ( n50214 , n50174 , n50213 );
and ( n50215 , n50173 , n50214 );
xor ( n50216 , n50172 , n50215 );
and ( n50217 , n50216 , n36587 );
or ( n50218 , n50171 , n50217 );
and ( n50219 , n50218 , n36596 );
not ( n50220 , n37485 );
and ( n50221 , n50220 , n37383 );
xor ( n50222 , n37383 , n36993 );
xor ( n50223 , n37366 , n36993 );
xor ( n50224 , n37349 , n36993 );
xor ( n50225 , n37332 , n36993 );
xor ( n50226 , n37315 , n36993 );
xor ( n50227 , n37298 , n36993 );
xor ( n50228 , n37281 , n36993 );
xor ( n50229 , n37264 , n36993 );
xor ( n50230 , n37247 , n36993 );
xor ( n50231 , n37230 , n36993 );
xor ( n50232 , n37213 , n36993 );
xor ( n50233 , n37196 , n36993 );
xor ( n50234 , n37179 , n36993 );
xor ( n50235 , n37162 , n36993 );
xor ( n50236 , n37145 , n36993 );
xor ( n50237 , n37128 , n36993 );
xor ( n50238 , n37111 , n36993 );
xor ( n50239 , n37094 , n36993 );
xor ( n50240 , n37077 , n36993 );
xor ( n50241 , n37060 , n36993 );
xor ( n50242 , n37043 , n36993 );
xor ( n50243 , n37026 , n36993 );
and ( n50244 , n37488 , n37490 );
and ( n50245 , n50243 , n50244 );
and ( n50246 , n50242 , n50245 );
and ( n50247 , n50241 , n50246 );
and ( n50248 , n50240 , n50247 );
and ( n50249 , n50239 , n50248 );
and ( n50250 , n50238 , n50249 );
and ( n50251 , n50237 , n50250 );
and ( n50252 , n50236 , n50251 );
and ( n50253 , n50235 , n50252 );
and ( n50254 , n50234 , n50253 );
and ( n50255 , n50233 , n50254 );
and ( n50256 , n50232 , n50255 );
and ( n50257 , n50231 , n50256 );
and ( n50258 , n50230 , n50257 );
and ( n50259 , n50229 , n50258 );
and ( n50260 , n50228 , n50259 );
and ( n50261 , n50227 , n50260 );
and ( n50262 , n50226 , n50261 );
and ( n50263 , n50225 , n50262 );
and ( n50264 , n50224 , n50263 );
and ( n50265 , n50223 , n50264 );
xor ( n50266 , n50222 , n50265 );
and ( n50267 , n50266 , n37485 );
or ( n50268 , n50221 , n50267 );
and ( n50269 , n50268 , n37494 );
and ( n50270 , n41862 , n37506 );
or ( n50271 , n50219 , n50269 , n50270 );
buf ( n50272 , n50271 );
buf ( n50273 , n50272 );
buf ( n50274 , n31655 );
or ( n50275 , n32427 , n32429 );
and ( n50276 , n47655 , n50275 );
and ( n50277 , n35288 , n35292 );
and ( n50278 , n35211 , n50277 );
not ( n50279 , n50278 );
and ( n50280 , n50279 , n47568 );
and ( n50281 , n47655 , n50278 );
or ( n50282 , n50280 , n50281 );
and ( n50283 , n50282 , n32421 );
not ( n50284 , n50002 );
and ( n50285 , n50284 , n47568 );
and ( n50286 , n47655 , n50002 );
or ( n50287 , n50285 , n50286 );
and ( n50288 , n50287 , n32419 );
and ( n50289 , n35278 , n50277 );
not ( n50290 , n50289 );
and ( n50291 , n50290 , n47568 );
and ( n50292 , n47655 , n50289 );
or ( n50293 , n50291 , n50292 );
and ( n50294 , n50293 , n32417 );
not ( n50295 , n50008 );
and ( n50296 , n50295 , n47568 );
and ( n50297 , n47655 , n50008 );
or ( n50298 , n50296 , n50297 );
and ( n50299 , n50298 , n32415 );
not ( n50300 , n47331 );
and ( n50301 , n50300 , n47568 );
and ( n50302 , n47600 , n47331 );
or ( n50303 , n50301 , n50302 );
and ( n50304 , n50303 , n32413 );
not ( n50305 , n50067 );
and ( n50306 , n50305 , n47568 );
and ( n50307 , n47600 , n50067 );
or ( n50308 , n50306 , n50307 );
and ( n50309 , n50308 , n32411 );
not ( n50310 , n31728 );
and ( n50311 , n50310 , n47568 );
xor ( n50312 , n47600 , n47629 );
and ( n50313 , n50312 , n31728 );
or ( n50314 , n50311 , n50313 );
and ( n50315 , n50314 , n32253 );
not ( n50316 , n32283 );
and ( n50317 , n50316 , n47568 );
not ( n50318 , n31823 );
xor ( n50319 , n47655 , n47684 );
and ( n50320 , n50318 , n50319 );
xnor ( n50321 , n47705 , n47734 );
and ( n50322 , n50321 , n31823 );
or ( n50323 , n50320 , n50322 );
and ( n50324 , n50323 , n32283 );
or ( n50325 , n50317 , n50324 );
and ( n50326 , n50325 , n32398 );
or ( n50327 , n32404 , n32403 );
or ( n50328 , n50327 , n32406 );
or ( n50329 , n50328 , n32409 );
or ( n50330 , n50329 , n32423 );
or ( n50331 , n50330 , n32425 );
or ( n50332 , n50331 , n32431 );
or ( n50333 , n50332 , n32433 );
or ( n50334 , n50333 , n32435 );
and ( n50335 , n47705 , n50334 );
or ( n50336 , n50276 , n50283 , n50288 , n50294 , n50299 , n50304 , n50309 , n50315 , n50326 , n50335 );
and ( n50337 , n50336 , n32456 );
and ( n50338 , n37543 , n32489 );
or ( n50339 , n32491 , n32486 );
or ( n50340 , n50339 , n32492 );
or ( n50341 , n50340 , n32473 );
or ( n50342 , n50341 , n32494 );
or ( n50343 , n50342 , n32496 );
or ( n50344 , n50343 , n32498 );
or ( n50345 , n50344 , n32500 );
and ( n50346 , n47568 , n50345 );
or ( n50347 , C0 , n50337 , n50338 , n50346 );
buf ( n50348 , n50347 );
buf ( n50349 , n50348 );
and ( n50350 , n33233 , n32528 );
not ( n50351 , n32598 );
and ( n50352 , n50351 , n32996 );
buf ( n50353 , n50352 );
and ( n50354 , n50353 , n32890 );
not ( n50355 , n32919 );
and ( n50356 , n50355 , n32996 );
buf ( n50357 , n50356 );
and ( n50358 , n50357 , n32924 );
not ( n50359 , n32953 );
and ( n50360 , n50359 , n32996 );
not ( n50361 , n32971 );
and ( n50362 , n50361 , n33117 );
xor ( n50363 , n32996 , n33009 );
and ( n50364 , n50363 , n32971 );
or ( n50365 , n50362 , n50364 );
and ( n50366 , n50365 , n32953 );
or ( n50367 , n50360 , n50366 );
and ( n50368 , n50367 , n33038 );
not ( n50369 , n33067 );
and ( n50370 , n50369 , n32996 );
not ( n50371 , n32970 );
not ( n50372 , n33071 );
and ( n50373 , n50372 , n33117 );
xor ( n50374 , n33118 , n33141 );
and ( n50375 , n50374 , n33071 );
or ( n50376 , n50373 , n50375 );
and ( n50377 , n50371 , n50376 );
and ( n50378 , n50363 , n32970 );
or ( n50379 , n50377 , n50378 );
and ( n50380 , n50379 , n33067 );
or ( n50381 , n50370 , n50380 );
and ( n50382 , n50381 , n33172 );
and ( n50383 , n32996 , n33204 );
or ( n50384 , n50354 , n50358 , n50368 , n50382 , n50383 );
and ( n50385 , n50384 , n33208 );
not ( n50386 , n32968 );
not ( n50387 , n33270 );
and ( n50388 , n50387 , n33317 );
xor ( n50389 , n33318 , n33341 );
and ( n50390 , n50389 , n33270 );
or ( n50391 , n50388 , n50390 );
and ( n50392 , n50386 , n50391 );
and ( n50393 , n32996 , n32968 );
or ( n50394 , n50392 , n50393 );
and ( n50395 , n50394 , n33370 );
buf ( n50396 , n35056 );
and ( n50397 , n32996 , n33382 );
or ( n50398 , C0 , n50350 , n50385 , n50395 , n50396 , n50397 );
buf ( n50399 , n50398 );
buf ( n50400 , n50399 );
buf ( n50401 , n31655 );
buf ( n50402 , n30987 );
buf ( n50403 , n30987 );
buf ( n50404 , n31655 );
not ( n50405 , n31728 );
and ( n50406 , n50405 , n46017 );
buf ( n50407 , RI15b5d1c8_1042);
buf ( n50408 , RI15b5d150_1041);
buf ( n50409 , RI15b5d0d8_1040);
buf ( n50410 , RI15b5d060_1039);
buf ( n50411 , RI15b5cfe8_1038);
and ( n50412 , n47567 , n47598 );
and ( n50413 , n50411 , n50412 );
and ( n50414 , n50410 , n50413 );
and ( n50415 , n50409 , n50414 );
and ( n50416 , n50408 , n50415 );
xor ( n50417 , n50407 , n50416 );
xor ( n50418 , n50408 , n50415 );
xor ( n50419 , n50409 , n50414 );
xor ( n50420 , n50410 , n50413 );
xor ( n50421 , n50411 , n50412 );
and ( n50422 , n47599 , n47630 );
and ( n50423 , n50421 , n50422 );
and ( n50424 , n50420 , n50423 );
and ( n50425 , n50419 , n50424 );
and ( n50426 , n50418 , n50425 );
xor ( n50427 , n50417 , n50426 );
and ( n50428 , n50427 , n31728 );
or ( n50429 , n50406 , n50428 );
and ( n50430 , n50429 , n32253 );
not ( n50431 , n32283 );
and ( n50432 , n50431 , n46017 );
not ( n50433 , n31823 );
and ( n50434 , n47567 , n47653 );
and ( n50435 , n50411 , n50434 );
and ( n50436 , n50410 , n50435 );
and ( n50437 , n50409 , n50436 );
and ( n50438 , n50408 , n50437 );
xor ( n50439 , n50407 , n50438 );
xor ( n50440 , n50408 , n50437 );
xor ( n50441 , n50409 , n50436 );
xor ( n50442 , n50410 , n50435 );
xor ( n50443 , n50411 , n50434 );
and ( n50444 , n47654 , n47685 );
and ( n50445 , n50443 , n50444 );
and ( n50446 , n50442 , n50445 );
and ( n50447 , n50441 , n50446 );
and ( n50448 , n50440 , n50447 );
xor ( n50449 , n50439 , n50448 );
and ( n50450 , n50433 , n50449 );
and ( n50451 , n47567 , n47703 );
and ( n50452 , n50411 , n50451 );
and ( n50453 , n50410 , n50452 );
and ( n50454 , n50409 , n50453 );
and ( n50455 , n50408 , n50454 );
xor ( n50456 , n50407 , n50455 );
xor ( n50457 , n50408 , n50454 );
xor ( n50458 , n50409 , n50453 );
xor ( n50459 , n50410 , n50452 );
xor ( n50460 , n50411 , n50451 );
or ( n50461 , n47704 , n47735 );
or ( n50462 , n50460 , n50461 );
or ( n50463 , n50459 , n50462 );
or ( n50464 , n50458 , n50463 );
or ( n50465 , n50457 , n50464 );
xnor ( n50466 , n50456 , n50465 );
and ( n50467 , n50466 , n31823 );
or ( n50468 , n50450 , n50467 );
and ( n50469 , n50468 , n32283 );
or ( n50470 , n50432 , n50469 );
and ( n50471 , n50470 , n32398 );
and ( n50472 , n46017 , n32436 );
or ( n50473 , n50430 , n50471 , n50472 );
and ( n50474 , n50473 , n32456 );
and ( n50475 , n49651 , n32473 );
not ( n50476 , n32475 );
and ( n50477 , n50476 , n49651 );
and ( n50478 , n46022 , n47764 );
and ( n50479 , n46021 , n50478 );
and ( n50480 , n46020 , n50479 );
and ( n50481 , n46019 , n50480 );
and ( n50482 , n46018 , n50481 );
xor ( n50483 , n46017 , n50482 );
and ( n50484 , n50483 , n32475 );
or ( n50485 , n50477 , n50484 );
and ( n50486 , n50485 , n32486 );
and ( n50487 , n37531 , n32489 );
and ( n50488 , n46017 , n32501 );
or ( n50489 , C0 , n50474 , n50475 , n50486 , n50487 , n50488 );
buf ( n50490 , n50489 );
buf ( n50491 , n50490 );
buf ( n50492 , n30987 );
buf ( n50493 , n31655 );
buf ( n50494 , n31655 );
not ( n50495 , n43755 );
and ( n50496 , n50495 , n43462 );
xor ( n50497 , n43462 , n43259 );
xor ( n50498 , n43445 , n43259 );
xor ( n50499 , n43428 , n43259 );
xor ( n50500 , n43411 , n43259 );
xor ( n50501 , n43394 , n43259 );
xor ( n50502 , n43377 , n43259 );
and ( n50503 , n43758 , n43770 );
and ( n50504 , n50502 , n50503 );
and ( n50505 , n50501 , n50504 );
and ( n50506 , n50500 , n50505 );
and ( n50507 , n50499 , n50506 );
and ( n50508 , n50498 , n50507 );
xor ( n50509 , n50497 , n50508 );
and ( n50510 , n50509 , n43755 );
or ( n50511 , n50496 , n50510 );
and ( n50512 , n50511 , n43774 );
not ( n50513 , n44663 );
and ( n50514 , n50513 , n44374 );
xor ( n50515 , n44374 , n44171 );
xor ( n50516 , n44357 , n44171 );
xor ( n50517 , n44340 , n44171 );
xor ( n50518 , n44323 , n44171 );
xor ( n50519 , n44306 , n44171 );
xor ( n50520 , n44289 , n44171 );
and ( n50521 , n44666 , n44678 );
and ( n50522 , n50520 , n50521 );
and ( n50523 , n50519 , n50522 );
and ( n50524 , n50518 , n50523 );
and ( n50525 , n50517 , n50524 );
and ( n50526 , n50516 , n50525 );
xor ( n50527 , n50515 , n50526 );
and ( n50528 , n50527 , n44663 );
or ( n50529 , n50514 , n50528 );
and ( n50530 , n50529 , n44682 );
buf ( n50531 , RI15b45618_232);
and ( n50532 , n50531 , n44695 );
or ( n50533 , n50512 , n50530 , n50532 );
buf ( n50534 , n50533 );
buf ( n50535 , n50534 );
buf ( n50536 , n30987 );
buf ( n50537 , n30987 );
not ( n50538 , n40163 );
and ( n50539 , n50538 , n31799 );
nor ( n50540 , n42169 , n42237 , n45160 , n31661 , n31657 );
not ( n50541 , n50540 );
and ( n50542 , n50541 , n31799 );
and ( n50543 , n32252 , n50540 );
or ( n50544 , n50542 , n50543 );
and ( n50545 , n50544 , n40163 );
or ( n50546 , n50539 , n50545 );
and ( n50547 , n50546 , n32498 );
nor ( n50548 , n42179 , n42246 , n45169 , n40194 , C0 );
not ( n50549 , n50548 );
not ( n50550 , n50540 );
and ( n50551 , n50550 , n31799 );
and ( n50552 , n40393 , n50540 );
or ( n50553 , n50551 , n50552 );
and ( n50554 , n50549 , n50553 );
and ( n50555 , n40393 , n50548 );
or ( n50556 , n50554 , n50555 );
and ( n50557 , n50556 , n32473 );
not ( n50558 , n32475 );
not ( n50559 , n50548 );
not ( n50560 , n50540 );
and ( n50561 , n50560 , n31799 );
and ( n50562 , n40393 , n50540 );
or ( n50563 , n50561 , n50562 );
and ( n50564 , n50559 , n50563 );
and ( n50565 , n40393 , n50548 );
or ( n50566 , n50564 , n50565 );
and ( n50567 , n50558 , n50566 );
nor ( n50568 , n42205 , n42272 , n45195 , n40445 , C0 );
not ( n50569 , n50568 );
nor ( n50570 , n42208 , n42275 , n45198 , n40440 , C0 );
not ( n50571 , n50570 );
and ( n50572 , n50571 , n50566 );
and ( n50573 , n40972 , n50570 );
or ( n50574 , n50572 , n50573 );
and ( n50575 , n50569 , n50574 );
and ( n50576 , n41267 , n50568 );
or ( n50577 , n50575 , n50576 );
and ( n50578 , n50577 , n32475 );
or ( n50579 , n50567 , n50578 );
and ( n50580 , n50579 , n32486 );
and ( n50581 , n31799 , n41278 );
or ( n50582 , C0 , n50547 , n50557 , n50580 , n50581 );
buf ( n50583 , n50582 );
buf ( n50584 , n50583 );
buf ( n50585 , n30987 );
xor ( n50586 , n41613 , n41606 );
and ( n50587 , n50586 , n31548 );
not ( n50588 , n44807 );
and ( n50589 , n50588 , n41613 );
and ( n50590 , n41886 , n44807 );
or ( n50591 , n50589 , n50590 );
and ( n50592 , n50591 , n31408 );
not ( n50593 , n44817 );
and ( n50594 , n50593 , n41613 );
not ( n50595 , n41835 );
buf ( n50596 , RI15b52c50_689);
and ( n50597 , n50595 , n50596 );
not ( n50598 , n42124 );
and ( n50599 , n50598 , n41896 );
xor ( n50600 , n42134 , n42136 );
and ( n50601 , n50600 , n42124 );
or ( n50602 , n50599 , n50601 );
and ( n50603 , n50602 , n41835 );
or ( n50604 , n50597 , n50603 );
and ( n50605 , n50604 , n44817 );
or ( n50606 , n50594 , n50605 );
and ( n50607 , n50606 , n31521 );
not ( n50608 , n45059 );
and ( n50609 , n50608 , n41613 );
and ( n50610 , n33647 , n45059 );
or ( n50611 , n50609 , n50610 );
and ( n50612 , n50611 , n31536 );
and ( n50613 , n41613 , n45148 );
or ( n50614 , n50587 , n50592 , n50607 , n50612 , n50613 );
and ( n50615 , n50614 , n31557 );
and ( n50616 , n41613 , n40154 );
or ( n50617 , C0 , n50615 , n50616 );
buf ( n50618 , n50617 );
buf ( n50619 , n50618 );
buf ( n50620 , n31655 );
buf ( n50621 , n31655 );
buf ( n50622 , n30987 );
not ( n50623 , n34150 );
and ( n50624 , n50623 , n32850 );
not ( n50625 , n34154 );
and ( n50626 , n50625 , n32850 );
and ( n50627 , n32856 , n34154 );
or ( n50628 , n50626 , n50627 );
and ( n50629 , n50628 , n34150 );
or ( n50630 , n50624 , n50629 );
and ( n50631 , n50630 , n33381 );
not ( n50632 , n34184 );
not ( n50633 , n34154 );
and ( n50634 , n50633 , n32850 );
and ( n50635 , n48160 , n34154 );
or ( n50636 , n50634 , n50635 );
and ( n50637 , n50632 , n50636 );
and ( n50638 , n48160 , n34184 );
or ( n50639 , n50637 , n50638 );
and ( n50640 , n50639 , n33375 );
not ( n50641 , n32968 );
not ( n50642 , n34184 );
not ( n50643 , n34154 );
and ( n50644 , n50643 , n32850 );
and ( n50645 , n48160 , n34154 );
or ( n50646 , n50644 , n50645 );
and ( n50647 , n50642 , n50646 );
and ( n50648 , n48160 , n34184 );
or ( n50649 , n50647 , n50648 );
and ( n50650 , n50641 , n50649 );
not ( n50651 , n34355 );
not ( n50652 , n34358 );
and ( n50653 , n50652 , n50649 );
and ( n50654 , n48186 , n34358 );
or ( n50655 , n50653 , n50654 );
and ( n50656 , n50651 , n50655 );
and ( n50657 , n48196 , n34355 );
or ( n50658 , n50656 , n50657 );
and ( n50659 , n50658 , n32968 );
or ( n50660 , n50650 , n50659 );
and ( n50661 , n50660 , n33370 );
and ( n50662 , n32850 , n35062 );
or ( n50663 , C0 , n50631 , n50640 , n50661 , n50662 );
buf ( n50664 , n50663 );
buf ( n50665 , n50664 );
not ( n50666 , n34150 );
and ( n50667 , n50666 , n32683 );
not ( n50668 , n34154 );
and ( n50669 , n50668 , n32683 );
and ( n50670 , n32689 , n34154 );
or ( n50671 , n50669 , n50670 );
and ( n50672 , n50671 , n34150 );
or ( n50673 , n50667 , n50672 );
and ( n50674 , n50673 , n33381 );
not ( n50675 , n34184 );
not ( n50676 , n34154 );
and ( n50677 , n50676 , n32683 );
not ( n50678 , n34287 );
and ( n50679 , n50678 , n34205 );
xor ( n50680 , n34293 , n34295 );
and ( n50681 , n50680 , n34287 );
or ( n50682 , n50679 , n50681 );
and ( n50683 , n50682 , n34154 );
or ( n50684 , n50677 , n50683 );
and ( n50685 , n50675 , n50684 );
and ( n50686 , n50682 , n34184 );
or ( n50687 , n50685 , n50686 );
and ( n50688 , n50687 , n33375 );
not ( n50689 , n32968 );
not ( n50690 , n34184 );
not ( n50691 , n34154 );
and ( n50692 , n50691 , n32683 );
and ( n50693 , n50682 , n34154 );
or ( n50694 , n50692 , n50693 );
and ( n50695 , n50690 , n50694 );
and ( n50696 , n50682 , n34184 );
or ( n50697 , n50695 , n50696 );
and ( n50698 , n50689 , n50697 );
not ( n50699 , n34355 );
not ( n50700 , n34358 );
and ( n50701 , n50700 , n50697 );
not ( n50702 , n34747 );
and ( n50703 , n50702 , n34641 );
xor ( n50704 , n34753 , n34755 );
and ( n50705 , n50704 , n34747 );
or ( n50706 , n50703 , n50705 );
and ( n50707 , n50706 , n34358 );
or ( n50708 , n50701 , n50707 );
and ( n50709 , n50699 , n50708 );
not ( n50710 , n35036 );
and ( n50711 , n50710 , n34934 );
xor ( n50712 , n35042 , n35044 );
and ( n50713 , n50712 , n35036 );
or ( n50714 , n50711 , n50713 );
and ( n50715 , n50714 , n34355 );
or ( n50716 , n50709 , n50715 );
and ( n50717 , n50716 , n32968 );
or ( n50718 , n50698 , n50717 );
and ( n50719 , n50718 , n33370 );
and ( n50720 , n32683 , n35062 );
or ( n50721 , C0 , n50674 , n50688 , n50719 , n50720 );
buf ( n50722 , n50721 );
buf ( n50723 , n50722 );
buf ( n50724 , n30987 );
buf ( n50725 , n31655 );
buf ( n50726 , n31655 );
buf ( n50727 , n30987 );
buf ( n50728 , n31655 );
not ( n50729 , n34150 );
and ( n50730 , n50729 , n32793 );
and ( n50731 , n41389 , n32542 , n32538 , n32534 , n41391 );
not ( n50732 , n50731 );
and ( n50733 , n50732 , n32793 );
and ( n50734 , n32823 , n50731 );
or ( n50735 , n50733 , n50734 );
and ( n50736 , n50735 , n34150 );
or ( n50737 , n50730 , n50736 );
and ( n50738 , n50737 , n33381 );
and ( n50739 , n41400 , n34170 , n34177 , n34183 , C1 );
not ( n50740 , n50739 );
not ( n50741 , n50731 );
and ( n50742 , n50741 , n32793 );
and ( n50743 , n41464 , n50731 );
or ( n50744 , n50742 , n50743 );
and ( n50745 , n50740 , n50744 );
and ( n50746 , n41464 , n50739 );
or ( n50747 , n50745 , n50746 );
and ( n50748 , n50747 , n33375 );
not ( n50749 , n32968 );
not ( n50750 , n50739 );
not ( n50751 , n50731 );
and ( n50752 , n50751 , n32793 );
and ( n50753 , n41464 , n50731 );
or ( n50754 , n50752 , n50753 );
and ( n50755 , n50750 , n50754 );
and ( n50756 , n41464 , n50739 );
or ( n50757 , n50755 , n50756 );
and ( n50758 , n50749 , n50757 );
and ( n50759 , n41422 , n34333 , n34344 , n34354 , C1 );
not ( n50760 , n50759 );
and ( n50761 , n41426 , n34329 , n34339 , n34349 , C1 );
not ( n50762 , n50761 );
and ( n50763 , n50762 , n50757 );
and ( n50764 , n41490 , n50761 );
or ( n50765 , n50763 , n50764 );
and ( n50766 , n50760 , n50765 );
and ( n50767 , n41500 , n50759 );
or ( n50768 , n50766 , n50767 );
and ( n50769 , n50768 , n32968 );
or ( n50770 , n50758 , n50769 );
and ( n50771 , n50770 , n33370 );
and ( n50772 , n32793 , n35062 );
or ( n50773 , C0 , n50738 , n50748 , n50771 , n50772 );
buf ( n50774 , n50773 );
buf ( n50775 , n50774 );
buf ( n50776 , n30987 );
not ( n50777 , n48765 );
and ( n50778 , n50777 , n33239 );
xor ( n50779 , n48923 , n48940 );
xor ( n50780 , n50779 , n48982 );
and ( n50781 , n50780 , n48765 );
or ( n50782 , n50778 , n50781 );
and ( n50783 , n50782 , n33180 );
not ( n50784 , n49054 );
and ( n50785 , n50784 , n33239 );
not ( n50786 , n48845 );
xor ( n50787 , n49089 , n48940 );
xor ( n50788 , n50787 , n49096 );
and ( n50789 , n50786 , n50788 );
xor ( n50790 , n49208 , n49210 );
xor ( n50791 , n50790 , n49222 );
and ( n50792 , n50791 , n48845 );
or ( n50793 , n50789 , n50792 );
and ( n50794 , n50793 , n49054 );
or ( n50795 , n50785 , n50794 );
and ( n50796 , n50795 , n33178 );
and ( n50797 , n33239 , n49774 );
or ( n50798 , n50783 , n50796 , n50797 );
and ( n50799 , n50798 , n33208 );
and ( n50800 , n33329 , n33375 );
not ( n50801 , n32968 );
and ( n50802 , n50801 , n33329 );
not ( n50803 , n33239 );
and ( n50804 , n50803 , n32968 );
or ( n50805 , n50802 , n50804 );
and ( n50806 , n50805 , n33370 );
and ( n50807 , n33002 , n35056 );
and ( n50808 , n33239 , n49794 );
or ( n50809 , C0 , n50799 , n50800 , n50806 , n50807 , n50808 );
buf ( n50810 , n50809 );
buf ( n50811 , n50810 );
buf ( n50812 , n30987 );
buf ( n50813 , n31655 );
buf ( n50814 , RI15b5e8c0_1091);
not ( n50815 , n50814 );
and ( n50816 , n40228 , n50815 );
and ( n50817 , n50816 , n48533 );
buf ( n50818 , RI15b5e7d0_1089);
not ( n50819 , n50818 );
and ( n50820 , n50817 , n50819 );
buf ( n50821 , RI15b5e758_1088);
and ( n50822 , n50820 , n50821 );
buf ( n50823 , RI15b5d768_1054);
buf ( n50824 , RI15b5d7e0_1055);
buf ( n50825 , RI15b5d858_1056);
buf ( n50826 , RI15b5d8d0_1057);
nor ( n50827 , n50823 , n50824 , n50825 , n50826 );
and ( n50828 , n50822 , n50827 );
not ( n50829 , n50828 );
and ( n50830 , n41869 , n41518 );
and ( n50831 , n50830 , n41520 );
and ( n50832 , n50831 , n41523 );
and ( n50833 , n50832 , n41525 );
and ( n50834 , n50833 , n41531 );
not ( n50835 , n50834 );
and ( n50836 , n50835 , n40303 );
buf ( n50837 , RI15b53538_708);
and ( n50838 , n50837 , n50834 );
or ( n50839 , n50836 , n50838 );
and ( n50840 , n50829 , n50839 );
buf ( n50841 , RI15b5f9a0_1127);
and ( n50842 , n50841 , n50828 );
or ( n50843 , n50840 , n50842 );
buf ( n50844 , n50843 );
buf ( n50845 , n50844 );
buf ( n50846 , n31655 );
buf ( n50847 , n30987 );
buf ( n50848 , n31655 );
buf ( n50849 , n30987 );
not ( n50850 , n34150 );
and ( n50851 , n50850 , n32826 );
not ( n50852 , n50731 );
and ( n50853 , n50852 , n32826 );
and ( n50854 , n32856 , n50731 );
or ( n50855 , n50853 , n50854 );
and ( n50856 , n50855 , n34150 );
or ( n50857 , n50851 , n50856 );
and ( n50858 , n50857 , n33381 );
not ( n50859 , n50739 );
not ( n50860 , n50731 );
and ( n50861 , n50860 , n32826 );
and ( n50862 , n48160 , n50731 );
or ( n50863 , n50861 , n50862 );
and ( n50864 , n50859 , n50863 );
and ( n50865 , n48160 , n50739 );
or ( n50866 , n50864 , n50865 );
and ( n50867 , n50866 , n33375 );
not ( n50868 , n32968 );
not ( n50869 , n50739 );
not ( n50870 , n50731 );
and ( n50871 , n50870 , n32826 );
and ( n50872 , n48160 , n50731 );
or ( n50873 , n50871 , n50872 );
and ( n50874 , n50869 , n50873 );
and ( n50875 , n48160 , n50739 );
or ( n50876 , n50874 , n50875 );
and ( n50877 , n50868 , n50876 );
not ( n50878 , n50759 );
not ( n50879 , n50761 );
and ( n50880 , n50879 , n50876 );
and ( n50881 , n48186 , n50761 );
or ( n50882 , n50880 , n50881 );
and ( n50883 , n50878 , n50882 );
and ( n50884 , n48196 , n50759 );
or ( n50885 , n50883 , n50884 );
and ( n50886 , n50885 , n32968 );
or ( n50887 , n50877 , n50886 );
and ( n50888 , n50887 , n33370 );
and ( n50889 , n32826 , n35062 );
or ( n50890 , C0 , n50858 , n50867 , n50888 , n50889 );
buf ( n50891 , n50890 );
buf ( n50892 , n50891 );
buf ( n50893 , n30987 );
buf ( n50894 , n31655 );
buf ( n50895 , n30987 );
not ( n50896 , n35278 );
buf ( n50897 , RI15b5ec08_1098);
and ( n50898 , n50896 , n50897 );
not ( n50899 , n46092 );
buf ( n50900 , RI15b614d0_1185);
and ( n50901 , n50899 , n50900 );
not ( n50902 , n50900 );
not ( n50903 , n46276 );
not ( n50904 , n46263 );
not ( n50905 , n46250 );
not ( n50906 , n46237 );
not ( n50907 , n46224 );
not ( n50908 , n46211 );
not ( n50909 , n46198 );
not ( n50910 , n46185 );
not ( n50911 , n46172 );
not ( n50912 , n46159 );
not ( n50913 , n46146 );
not ( n50914 , n46133 );
not ( n50915 , n46120 );
not ( n50916 , n46107 );
not ( n50917 , n46094 );
not ( n50918 , n46087 );
and ( n50919 , n50917 , n50918 );
and ( n50920 , n50916 , n50919 );
and ( n50921 , n50915 , n50920 );
and ( n50922 , n50914 , n50921 );
and ( n50923 , n50913 , n50922 );
and ( n50924 , n50912 , n50923 );
and ( n50925 , n50911 , n50924 );
and ( n50926 , n50910 , n50925 );
and ( n50927 , n50909 , n50926 );
and ( n50928 , n50908 , n50927 );
and ( n50929 , n50907 , n50928 );
and ( n50930 , n50906 , n50929 );
and ( n50931 , n50905 , n50930 );
and ( n50932 , n50904 , n50931 );
and ( n50933 , n50903 , n50932 );
xor ( n50934 , n50902 , n50933 );
and ( n50935 , n50934 , n46092 );
or ( n50936 , n50901 , n50935 );
not ( n50937 , n50936 );
buf ( n50938 , n50937 );
buf ( n50939 , n50938 );
not ( n50940 , n50939 );
buf ( n50941 , n50940 );
buf ( n50942 , n50941 );
not ( n50943 , n50942 );
buf ( n50944 , n50943 );
not ( n50945 , n50944 );
not ( n50946 , n46092 );
buf ( n50947 , RI15b61b60_1199);
not ( n50948 , n50947 );
buf ( n50949 , RI15b61ae8_1198);
not ( n50950 , n50949 );
buf ( n50951 , RI15b61a70_1197);
not ( n50952 , n50951 );
buf ( n50953 , RI15b619f8_1196);
not ( n50954 , n50953 );
buf ( n50955 , RI15b61980_1195);
not ( n50956 , n50955 );
buf ( n50957 , RI15b61908_1194);
not ( n50958 , n50957 );
buf ( n50959 , RI15b61890_1193);
not ( n50960 , n50959 );
buf ( n50961 , RI15b61818_1192);
not ( n50962 , n50961 );
buf ( n50963 , RI15b617a0_1191);
not ( n50964 , n50963 );
buf ( n50965 , RI15b61728_1190);
not ( n50966 , n50965 );
buf ( n50967 , RI15b616b0_1189);
not ( n50968 , n50967 );
buf ( n50969 , RI15b61638_1188);
not ( n50970 , n50969 );
buf ( n50971 , RI15b615c0_1187);
not ( n50972 , n50971 );
buf ( n50973 , RI15b61548_1186);
not ( n50974 , n50973 );
and ( n50975 , n50902 , n50933 );
and ( n50976 , n50974 , n50975 );
and ( n50977 , n50972 , n50976 );
and ( n50978 , n50970 , n50977 );
and ( n50979 , n50968 , n50978 );
and ( n50980 , n50966 , n50979 );
and ( n50981 , n50964 , n50980 );
and ( n50982 , n50962 , n50981 );
and ( n50983 , n50960 , n50982 );
and ( n50984 , n50958 , n50983 );
and ( n50985 , n50956 , n50984 );
and ( n50986 , n50954 , n50985 );
and ( n50987 , n50952 , n50986 );
and ( n50988 , n50950 , n50987 );
and ( n50989 , n50948 , n50988 );
xor ( n50990 , n50946 , n50989 );
buf ( n50991 , n46092 );
and ( n50992 , n50990 , n50991 );
buf ( n50993 , n50992 );
not ( n50994 , n50993 );
not ( n50995 , n50994 );
not ( n50996 , n50995 );
not ( n50997 , n46092 );
and ( n50998 , n50997 , n50947 );
xor ( n50999 , n50948 , n50988 );
and ( n51000 , n50999 , n46092 );
or ( n51001 , n50998 , n51000 );
not ( n51002 , n51001 );
buf ( n51003 , n51002 );
buf ( n51004 , n51003 );
not ( n51005 , n51004 );
not ( n51006 , n51005 );
not ( n51007 , n46092 );
and ( n51008 , n51007 , n50949 );
xor ( n51009 , n50950 , n50987 );
and ( n51010 , n51009 , n46092 );
or ( n51011 , n51008 , n51010 );
not ( n51012 , n51011 );
buf ( n51013 , n51012 );
buf ( n51014 , n51013 );
not ( n51015 , n51014 );
not ( n51016 , n51015 );
not ( n51017 , n46092 );
and ( n51018 , n51017 , n50951 );
xor ( n51019 , n50952 , n50986 );
and ( n51020 , n51019 , n46092 );
or ( n51021 , n51018 , n51020 );
not ( n51022 , n51021 );
buf ( n51023 , n51022 );
buf ( n51024 , n51023 );
not ( n51025 , n51024 );
not ( n51026 , n51025 );
not ( n51027 , n46092 );
and ( n51028 , n51027 , n50953 );
xor ( n51029 , n50954 , n50985 );
and ( n51030 , n51029 , n46092 );
or ( n51031 , n51028 , n51030 );
not ( n51032 , n51031 );
buf ( n51033 , n51032 );
buf ( n51034 , n51033 );
not ( n51035 , n51034 );
not ( n51036 , n51035 );
not ( n51037 , n46092 );
and ( n51038 , n51037 , n50955 );
xor ( n51039 , n50956 , n50984 );
and ( n51040 , n51039 , n46092 );
or ( n51041 , n51038 , n51040 );
not ( n51042 , n51041 );
buf ( n51043 , n51042 );
buf ( n51044 , n51043 );
not ( n51045 , n51044 );
not ( n51046 , n51045 );
not ( n51047 , n46092 );
and ( n51048 , n51047 , n50957 );
xor ( n51049 , n50958 , n50983 );
and ( n51050 , n51049 , n46092 );
or ( n51051 , n51048 , n51050 );
not ( n51052 , n51051 );
buf ( n51053 , n51052 );
buf ( n51054 , n51053 );
not ( n51055 , n51054 );
not ( n51056 , n51055 );
not ( n51057 , n46092 );
and ( n51058 , n51057 , n50959 );
xor ( n51059 , n50960 , n50982 );
and ( n51060 , n51059 , n46092 );
or ( n51061 , n51058 , n51060 );
not ( n51062 , n51061 );
buf ( n51063 , n51062 );
buf ( n51064 , n51063 );
not ( n51065 , n51064 );
not ( n51066 , n51065 );
not ( n51067 , n46092 );
and ( n51068 , n51067 , n50961 );
xor ( n51069 , n50962 , n50981 );
and ( n51070 , n51069 , n46092 );
or ( n51071 , n51068 , n51070 );
not ( n51072 , n51071 );
buf ( n51073 , n51072 );
buf ( n51074 , n51073 );
not ( n51075 , n51074 );
not ( n51076 , n51075 );
not ( n51077 , n46092 );
and ( n51078 , n51077 , n50963 );
xor ( n51079 , n50964 , n50980 );
and ( n51080 , n51079 , n46092 );
or ( n51081 , n51078 , n51080 );
not ( n51082 , n51081 );
buf ( n51083 , n51082 );
buf ( n51084 , n51083 );
not ( n51085 , n51084 );
not ( n51086 , n51085 );
not ( n51087 , n46092 );
and ( n51088 , n51087 , n50965 );
xor ( n51089 , n50966 , n50979 );
and ( n51090 , n51089 , n46092 );
or ( n51091 , n51088 , n51090 );
not ( n51092 , n51091 );
buf ( n51093 , n51092 );
buf ( n51094 , n51093 );
not ( n51095 , n51094 );
not ( n51096 , n51095 );
not ( n51097 , n46092 );
and ( n51098 , n51097 , n50967 );
xor ( n51099 , n50968 , n50978 );
and ( n51100 , n51099 , n46092 );
or ( n51101 , n51098 , n51100 );
not ( n51102 , n51101 );
buf ( n51103 , n51102 );
buf ( n51104 , n51103 );
not ( n51105 , n51104 );
not ( n51106 , n51105 );
not ( n51107 , n46092 );
and ( n51108 , n51107 , n50969 );
xor ( n51109 , n50970 , n50977 );
and ( n51110 , n51109 , n46092 );
or ( n51111 , n51108 , n51110 );
not ( n51112 , n51111 );
buf ( n51113 , n51112 );
buf ( n51114 , n51113 );
not ( n51115 , n51114 );
not ( n51116 , n51115 );
not ( n51117 , n46092 );
and ( n51118 , n51117 , n50971 );
xor ( n51119 , n50972 , n50976 );
and ( n51120 , n51119 , n46092 );
or ( n51121 , n51118 , n51120 );
not ( n51122 , n51121 );
buf ( n51123 , n51122 );
buf ( n51124 , n51123 );
not ( n51125 , n51124 );
not ( n51126 , n51125 );
not ( n51127 , n46092 );
and ( n51128 , n51127 , n50973 );
xor ( n51129 , n50974 , n50975 );
and ( n51130 , n51129 , n46092 );
or ( n51131 , n51128 , n51130 );
not ( n51132 , n51131 );
buf ( n51133 , n51132 );
buf ( n51134 , n51133 );
not ( n51135 , n51134 );
not ( n51136 , n51135 );
not ( n51137 , n50940 );
and ( n51138 , n51136 , n51137 );
and ( n51139 , n51126 , n51138 );
and ( n51140 , n51116 , n51139 );
and ( n51141 , n51106 , n51140 );
and ( n51142 , n51096 , n51141 );
and ( n51143 , n51086 , n51142 );
and ( n51144 , n51076 , n51143 );
and ( n51145 , n51066 , n51144 );
and ( n51146 , n51056 , n51145 );
and ( n51147 , n51046 , n51146 );
and ( n51148 , n51036 , n51147 );
and ( n51149 , n51026 , n51148 );
and ( n51150 , n51016 , n51149 );
and ( n51151 , n51006 , n51150 );
and ( n51152 , n50996 , n51151 );
not ( n51153 , n51152 );
and ( n51154 , n51153 , n46092 );
buf ( n51155 , n51154 );
not ( n51156 , n51155 );
not ( n51157 , n46092 );
and ( n51158 , n51157 , n51135 );
xor ( n51159 , n51136 , n51137 );
and ( n51160 , n51159 , n46092 );
or ( n51161 , n51158 , n51160 );
and ( n51162 , n51156 , n51161 );
not ( n51163 , n51161 );
not ( n51164 , n50941 );
xor ( n51165 , n51163 , n51164 );
and ( n51166 , n51165 , n51155 );
or ( n51167 , n51162 , n51166 );
not ( n51168 , n51167 );
buf ( n51169 , n51168 );
buf ( n51170 , n51169 );
not ( n51171 , n51170 );
or ( n51172 , n50945 , n51171 );
not ( n51173 , n51155 );
not ( n51174 , n46092 );
and ( n51175 , n51174 , n51125 );
xor ( n51176 , n51126 , n51138 );
and ( n51177 , n51176 , n46092 );
or ( n51178 , n51175 , n51177 );
and ( n51179 , n51173 , n51178 );
not ( n51180 , n51178 );
and ( n51181 , n51163 , n51164 );
xor ( n51182 , n51180 , n51181 );
and ( n51183 , n51182 , n51155 );
or ( n51184 , n51179 , n51183 );
not ( n51185 , n51184 );
buf ( n51186 , n51185 );
buf ( n51187 , n51186 );
not ( n51188 , n51187 );
or ( n51189 , n51172 , n51188 );
not ( n51190 , n51155 );
not ( n51191 , n46092 );
and ( n51192 , n51191 , n51115 );
xor ( n51193 , n51116 , n51139 );
and ( n51194 , n51193 , n46092 );
or ( n51195 , n51192 , n51194 );
and ( n51196 , n51190 , n51195 );
not ( n51197 , n51195 );
and ( n51198 , n51180 , n51181 );
xor ( n51199 , n51197 , n51198 );
and ( n51200 , n51199 , n51155 );
or ( n51201 , n51196 , n51200 );
not ( n51202 , n51201 );
buf ( n51203 , n51202 );
buf ( n51204 , n51203 );
not ( n51205 , n51204 );
or ( n51206 , n51189 , n51205 );
not ( n51207 , n51155 );
not ( n51208 , n46092 );
and ( n51209 , n51208 , n51105 );
xor ( n51210 , n51106 , n51140 );
and ( n51211 , n51210 , n46092 );
or ( n51212 , n51209 , n51211 );
and ( n51213 , n51207 , n51212 );
not ( n51214 , n51212 );
and ( n51215 , n51197 , n51198 );
xor ( n51216 , n51214 , n51215 );
and ( n51217 , n51216 , n51155 );
or ( n51218 , n51213 , n51217 );
not ( n51219 , n51218 );
buf ( n51220 , n51219 );
buf ( n51221 , n51220 );
not ( n51222 , n51221 );
or ( n51223 , n51206 , n51222 );
not ( n51224 , n51155 );
not ( n51225 , n46092 );
and ( n51226 , n51225 , n51095 );
xor ( n51227 , n51096 , n51141 );
and ( n51228 , n51227 , n46092 );
or ( n51229 , n51226 , n51228 );
and ( n51230 , n51224 , n51229 );
not ( n51231 , n51229 );
and ( n51232 , n51214 , n51215 );
xor ( n51233 , n51231 , n51232 );
and ( n51234 , n51233 , n51155 );
or ( n51235 , n51230 , n51234 );
not ( n51236 , n51235 );
buf ( n51237 , n51236 );
buf ( n51238 , n51237 );
not ( n51239 , n51238 );
or ( n51240 , n51223 , n51239 );
not ( n51241 , n51155 );
not ( n51242 , n46092 );
and ( n51243 , n51242 , n51085 );
xor ( n51244 , n51086 , n51142 );
and ( n51245 , n51244 , n46092 );
or ( n51246 , n51243 , n51245 );
and ( n51247 , n51241 , n51246 );
not ( n51248 , n51246 );
and ( n51249 , n51231 , n51232 );
xor ( n51250 , n51248 , n51249 );
and ( n51251 , n51250 , n51155 );
or ( n51252 , n51247 , n51251 );
not ( n51253 , n51252 );
buf ( n51254 , n51253 );
buf ( n51255 , n51254 );
not ( n51256 , n51255 );
or ( n51257 , n51240 , n51256 );
not ( n51258 , n51155 );
not ( n51259 , n46092 );
and ( n51260 , n51259 , n51075 );
xor ( n51261 , n51076 , n51143 );
and ( n51262 , n51261 , n46092 );
or ( n51263 , n51260 , n51262 );
and ( n51264 , n51258 , n51263 );
not ( n51265 , n51263 );
and ( n51266 , n51248 , n51249 );
xor ( n51267 , n51265 , n51266 );
and ( n51268 , n51267 , n51155 );
or ( n51269 , n51264 , n51268 );
not ( n51270 , n51269 );
buf ( n51271 , n51270 );
buf ( n51272 , n51271 );
not ( n51273 , n51272 );
or ( n51274 , n51257 , n51273 );
not ( n51275 , n51155 );
not ( n51276 , n46092 );
and ( n51277 , n51276 , n51065 );
xor ( n51278 , n51066 , n51144 );
and ( n51279 , n51278 , n46092 );
or ( n51280 , n51277 , n51279 );
and ( n51281 , n51275 , n51280 );
not ( n51282 , n51280 );
and ( n51283 , n51265 , n51266 );
xor ( n51284 , n51282 , n51283 );
and ( n51285 , n51284 , n51155 );
or ( n51286 , n51281 , n51285 );
not ( n51287 , n51286 );
buf ( n51288 , n51287 );
buf ( n51289 , n51288 );
not ( n51290 , n51289 );
or ( n51291 , n51274 , n51290 );
not ( n51292 , n51155 );
not ( n51293 , n46092 );
and ( n51294 , n51293 , n51055 );
xor ( n51295 , n51056 , n51145 );
and ( n51296 , n51295 , n46092 );
or ( n51297 , n51294 , n51296 );
and ( n51298 , n51292 , n51297 );
not ( n51299 , n51297 );
and ( n51300 , n51282 , n51283 );
xor ( n51301 , n51299 , n51300 );
and ( n51302 , n51301 , n51155 );
or ( n51303 , n51298 , n51302 );
not ( n51304 , n51303 );
buf ( n51305 , n51304 );
buf ( n51306 , n51305 );
not ( n51307 , n51306 );
or ( n51308 , n51291 , n51307 );
not ( n51309 , n51155 );
not ( n51310 , n46092 );
and ( n51311 , n51310 , n51045 );
xor ( n51312 , n51046 , n51146 );
and ( n51313 , n51312 , n46092 );
or ( n51314 , n51311 , n51313 );
and ( n51315 , n51309 , n51314 );
not ( n51316 , n51314 );
and ( n51317 , n51299 , n51300 );
xor ( n51318 , n51316 , n51317 );
and ( n51319 , n51318 , n51155 );
or ( n51320 , n51315 , n51319 );
not ( n51321 , n51320 );
buf ( n51322 , n51321 );
buf ( n51323 , n51322 );
not ( n51324 , n51323 );
or ( n51325 , n51308 , n51324 );
not ( n51326 , n51155 );
not ( n51327 , n46092 );
and ( n51328 , n51327 , n51035 );
xor ( n51329 , n51036 , n51147 );
and ( n51330 , n51329 , n46092 );
or ( n51331 , n51328 , n51330 );
and ( n51332 , n51326 , n51331 );
not ( n51333 , n51331 );
and ( n51334 , n51316 , n51317 );
xor ( n51335 , n51333 , n51334 );
and ( n51336 , n51335 , n51155 );
or ( n51337 , n51332 , n51336 );
not ( n51338 , n51337 );
buf ( n51339 , n51338 );
buf ( n51340 , n51339 );
not ( n51341 , n51340 );
or ( n51342 , n51325 , n51341 );
not ( n51343 , n51155 );
not ( n51344 , n46092 );
and ( n51345 , n51344 , n51025 );
xor ( n51346 , n51026 , n51148 );
and ( n51347 , n51346 , n46092 );
or ( n51348 , n51345 , n51347 );
and ( n51349 , n51343 , n51348 );
not ( n51350 , n51348 );
and ( n51351 , n51333 , n51334 );
xor ( n51352 , n51350 , n51351 );
and ( n51353 , n51352 , n51155 );
or ( n51354 , n51349 , n51353 );
not ( n51355 , n51354 );
buf ( n51356 , n51355 );
buf ( n51357 , n51356 );
not ( n51358 , n51357 );
or ( n51359 , n51342 , n51358 );
not ( n51360 , n51155 );
not ( n51361 , n46092 );
and ( n51362 , n51361 , n51015 );
xor ( n51363 , n51016 , n51149 );
and ( n51364 , n51363 , n46092 );
or ( n51365 , n51362 , n51364 );
and ( n51366 , n51360 , n51365 );
not ( n51367 , n51365 );
and ( n51368 , n51350 , n51351 );
xor ( n51369 , n51367 , n51368 );
and ( n51370 , n51369 , n51155 );
or ( n51371 , n51366 , n51370 );
not ( n51372 , n51371 );
buf ( n51373 , n51372 );
buf ( n51374 , n51373 );
not ( n51375 , n51374 );
or ( n51376 , n51359 , n51375 );
not ( n51377 , n51155 );
not ( n51378 , n46092 );
and ( n51379 , n51378 , n51005 );
xor ( n51380 , n51006 , n51150 );
and ( n51381 , n51380 , n46092 );
or ( n51382 , n51379 , n51381 );
and ( n51383 , n51377 , n51382 );
not ( n51384 , n51382 );
and ( n51385 , n51367 , n51368 );
xor ( n51386 , n51384 , n51385 );
and ( n51387 , n51386 , n51155 );
or ( n51388 , n51383 , n51387 );
not ( n51389 , n51388 );
buf ( n51390 , n51389 );
buf ( n51391 , n51390 );
not ( n51392 , n51391 );
or ( n51393 , n51376 , n51392 );
buf ( n51394 , n51393 );
buf ( n51395 , n51394 );
and ( n51396 , n51395 , n51155 );
not ( n51397 , n51396 );
and ( n51398 , n51397 , n51256 );
xor ( n51399 , n51256 , n51155 );
xor ( n51400 , n51239 , n51155 );
xor ( n51401 , n51222 , n51155 );
xor ( n51402 , n51205 , n51155 );
xor ( n51403 , n51188 , n51155 );
xor ( n51404 , n51171 , n51155 );
xor ( n51405 , n50945 , n51155 );
and ( n51406 , n51405 , n51155 );
and ( n51407 , n51404 , n51406 );
and ( n51408 , n51403 , n51407 );
and ( n51409 , n51402 , n51408 );
and ( n51410 , n51401 , n51409 );
and ( n51411 , n51400 , n51410 );
xor ( n51412 , n51399 , n51411 );
and ( n51413 , n51412 , n51396 );
or ( n51414 , n51398 , n51413 );
and ( n51415 , n51414 , n35278 );
or ( n51416 , n50898 , n51415 );
and ( n51417 , n51416 , n32417 );
not ( n51418 , n50008 );
and ( n51419 , n51418 , n50897 );
buf ( n51420 , n40234 );
not ( n51421 , n51420 );
buf ( n51422 , n51421 );
not ( n51423 , n51422 );
not ( n51424 , n40244 );
and ( n51425 , n51424 , n40251 );
not ( n51426 , n40251 );
not ( n51427 , n40234 );
xor ( n51428 , n51426 , n51427 );
and ( n51429 , n51428 , n40244 );
or ( n51430 , n51425 , n51429 );
not ( n51431 , n51430 );
buf ( n51432 , n51431 );
buf ( n51433 , n51432 );
not ( n51434 , n51433 );
or ( n51435 , n51423 , n51434 );
not ( n51436 , n40244 );
and ( n51437 , n51436 , n40269 );
not ( n51438 , n40269 );
and ( n51439 , n51426 , n51427 );
xor ( n51440 , n51438 , n51439 );
and ( n51441 , n51440 , n40244 );
or ( n51442 , n51437 , n51441 );
not ( n51443 , n51442 );
buf ( n51444 , n51443 );
buf ( n51445 , n51444 );
not ( n51446 , n51445 );
or ( n51447 , n51435 , n51446 );
not ( n51448 , n40244 );
and ( n51449 , n51448 , n40287 );
not ( n51450 , n40287 );
and ( n51451 , n51438 , n51439 );
xor ( n51452 , n51450 , n51451 );
and ( n51453 , n51452 , n40244 );
or ( n51454 , n51449 , n51453 );
not ( n51455 , n51454 );
buf ( n51456 , n51455 );
buf ( n51457 , n51456 );
not ( n51458 , n51457 );
or ( n51459 , n51447 , n51458 );
not ( n51460 , n40244 );
and ( n51461 , n51460 , n40305 );
not ( n51462 , n40305 );
and ( n51463 , n51450 , n51451 );
xor ( n51464 , n51462 , n51463 );
and ( n51465 , n51464 , n40244 );
or ( n51466 , n51461 , n51465 );
not ( n51467 , n51466 );
buf ( n51468 , n51467 );
buf ( n51469 , n51468 );
not ( n51470 , n51469 );
or ( n51471 , n51459 , n51470 );
not ( n51472 , n40244 );
and ( n51473 , n51472 , n40323 );
not ( n51474 , n40323 );
and ( n51475 , n51462 , n51463 );
xor ( n51476 , n51474 , n51475 );
and ( n51477 , n51476 , n40244 );
or ( n51478 , n51473 , n51477 );
not ( n51479 , n51478 );
buf ( n51480 , n51479 );
buf ( n51481 , n51480 );
not ( n51482 , n51481 );
or ( n51483 , n51471 , n51482 );
not ( n51484 , n40244 );
and ( n51485 , n51484 , n40341 );
not ( n51486 , n40341 );
and ( n51487 , n51474 , n51475 );
xor ( n51488 , n51486 , n51487 );
and ( n51489 , n51488 , n40244 );
or ( n51490 , n51485 , n51489 );
not ( n51491 , n51490 );
buf ( n51492 , n51491 );
buf ( n51493 , n51492 );
not ( n51494 , n51493 );
or ( n51495 , n51483 , n51494 );
not ( n51496 , n40244 );
and ( n51497 , n51496 , n40359 );
not ( n51498 , n40359 );
and ( n51499 , n51486 , n51487 );
xor ( n51500 , n51498 , n51499 );
and ( n51501 , n51500 , n40244 );
or ( n51502 , n51497 , n51501 );
not ( n51503 , n51502 );
buf ( n51504 , n51503 );
buf ( n51505 , n51504 );
not ( n51506 , n51505 );
or ( n51507 , n51495 , n51506 );
not ( n51508 , n40244 );
and ( n51509 , n51508 , n40514 );
not ( n51510 , n40514 );
and ( n51511 , n51498 , n51499 );
xor ( n51512 , n51510 , n51511 );
and ( n51513 , n51512 , n40244 );
or ( n51514 , n51509 , n51513 );
not ( n51515 , n51514 );
buf ( n51516 , n51515 );
buf ( n51517 , n51516 );
not ( n51518 , n51517 );
or ( n51519 , n51507 , n51518 );
not ( n51520 , n40244 );
and ( n51521 , n51520 , n40507 );
not ( n51522 , n40507 );
and ( n51523 , n51510 , n51511 );
xor ( n51524 , n51522 , n51523 );
and ( n51525 , n51524 , n40244 );
or ( n51526 , n51521 , n51525 );
not ( n51527 , n51526 );
buf ( n51528 , n51527 );
buf ( n51529 , n51528 );
not ( n51530 , n51529 );
or ( n51531 , n51519 , n51530 );
not ( n51532 , n40244 );
and ( n51533 , n51532 , n40500 );
not ( n51534 , n40500 );
and ( n51535 , n51522 , n51523 );
xor ( n51536 , n51534 , n51535 );
and ( n51537 , n51536 , n40244 );
or ( n51538 , n51533 , n51537 );
not ( n51539 , n51538 );
buf ( n51540 , n51539 );
buf ( n51541 , n51540 );
not ( n51542 , n51541 );
or ( n51543 , n51531 , n51542 );
not ( n51544 , n40244 );
and ( n51545 , n51544 , n40493 );
not ( n51546 , n40493 );
and ( n51547 , n51534 , n51535 );
xor ( n51548 , n51546 , n51547 );
and ( n51549 , n51548 , n40244 );
or ( n51550 , n51545 , n51549 );
not ( n51551 , n51550 );
buf ( n51552 , n51551 );
buf ( n51553 , n51552 );
not ( n51554 , n51553 );
or ( n51555 , n51543 , n51554 );
not ( n51556 , n40244 );
and ( n51557 , n51556 , n40486 );
not ( n51558 , n40486 );
and ( n51559 , n51546 , n51547 );
xor ( n51560 , n51558 , n51559 );
and ( n51561 , n51560 , n40244 );
or ( n51562 , n51557 , n51561 );
not ( n51563 , n51562 );
buf ( n51564 , n51563 );
buf ( n51565 , n51564 );
not ( n51566 , n51565 );
or ( n51567 , n51555 , n51566 );
not ( n51568 , n40244 );
and ( n51569 , n51568 , n40479 );
not ( n51570 , n40479 );
and ( n51571 , n51558 , n51559 );
xor ( n51572 , n51570 , n51571 );
and ( n51573 , n51572 , n40244 );
or ( n51574 , n51569 , n51573 );
not ( n51575 , n51574 );
buf ( n51576 , n51575 );
buf ( n51577 , n51576 );
not ( n51578 , n51577 );
or ( n51579 , n51567 , n51578 );
not ( n51580 , n40244 );
and ( n51581 , n51580 , n40472 );
not ( n51582 , n40472 );
and ( n51583 , n51570 , n51571 );
xor ( n51584 , n51582 , n51583 );
and ( n51585 , n51584 , n40244 );
or ( n51586 , n51581 , n51585 );
not ( n51587 , n51586 );
buf ( n51588 , n51587 );
buf ( n51589 , n51588 );
not ( n51590 , n51589 );
or ( n51591 , n51579 , n51590 );
buf ( n51592 , n51591 );
buf ( n51593 , n51592 );
and ( n51594 , n51593 , n40244 );
not ( n51595 , n51594 );
and ( n51596 , n51595 , n51494 );
xor ( n51597 , n51494 , n40244 );
xor ( n51598 , n51482 , n40244 );
xor ( n51599 , n51470 , n40244 );
xor ( n51600 , n51458 , n40244 );
xor ( n51601 , n51446 , n40244 );
xor ( n51602 , n51434 , n40244 );
xor ( n51603 , n51423 , n40244 );
and ( n51604 , n51603 , n40244 );
and ( n51605 , n51602 , n51604 );
and ( n51606 , n51601 , n51605 );
and ( n51607 , n51600 , n51606 );
and ( n51608 , n51599 , n51607 );
and ( n51609 , n51598 , n51608 );
xor ( n51610 , n51597 , n51609 );
and ( n51611 , n51610 , n51594 );
or ( n51612 , n51596 , n51611 );
and ( n51613 , n51612 , n50008 );
or ( n51614 , n51419 , n51613 );
and ( n51615 , n51614 , n32415 );
and ( n51616 , n50897 , n48133 );
or ( n51617 , n51417 , n51615 , n51616 );
and ( n51618 , n51617 , n32456 );
and ( n51619 , n50897 , n47409 );
or ( n51620 , C0 , n51618 , n51619 );
buf ( n51621 , n51620 );
buf ( n51622 , n51621 );
buf ( n51623 , n31655 );
and ( n51624 , n33771 , n48455 );
not ( n51625 , n48457 );
and ( n51626 , n51625 , n33436 );
and ( n51627 , n33771 , n48457 );
or ( n51628 , n51626 , n51627 );
and ( n51629 , n51628 , n31373 );
not ( n51630 , n44807 );
and ( n51631 , n51630 , n33436 );
and ( n51632 , n33771 , n44807 );
or ( n51633 , n51631 , n51632 );
and ( n51634 , n51633 , n31408 );
not ( n51635 , n48468 );
and ( n51636 , n51635 , n33436 );
and ( n51637 , n33771 , n48468 );
or ( n51638 , n51636 , n51637 );
and ( n51639 , n51638 , n31468 );
not ( n51640 , n44817 );
and ( n51641 , n51640 , n33436 );
and ( n51642 , n33771 , n44817 );
or ( n51643 , n51641 , n51642 );
and ( n51644 , n51643 , n31521 );
not ( n51645 , n39979 );
and ( n51646 , n51645 , n33436 );
and ( n51647 , n33478 , n39979 );
or ( n51648 , n51646 , n51647 );
and ( n51649 , n51648 , n31538 );
not ( n51650 , n45059 );
and ( n51651 , n51650 , n33436 );
and ( n51652 , n33478 , n45059 );
or ( n51653 , n51651 , n51652 );
and ( n51654 , n51653 , n31536 );
not ( n51655 , n33419 );
and ( n51656 , n51655 , n33436 );
and ( n51657 , n35556 , n33419 );
or ( n51658 , n51656 , n51657 );
and ( n51659 , n51658 , n31529 );
not ( n51660 , n33734 );
and ( n51661 , n51660 , n33436 );
and ( n51662 , n35569 , n33734 );
or ( n51663 , n51661 , n51662 );
and ( n51664 , n51663 , n31527 );
and ( n51665 , n33856 , n48513 );
or ( n51666 , n51624 , n51629 , n51634 , n51639 , n51644 , n51649 , n51654 , n51659 , n51664 , n51665 );
and ( n51667 , n51666 , n31557 );
and ( n51668 , n34008 , n33973 );
and ( n51669 , n33436 , n48524 );
or ( n51670 , C0 , n51667 , n51668 , n51669 );
buf ( n51671 , n51670 );
buf ( n51672 , n51671 );
and ( n51673 , n41298 , n50275 );
not ( n51674 , n50278 );
and ( n51675 , n51674 , n41286 );
and ( n51676 , n41298 , n50278 );
or ( n51677 , n51675 , n51676 );
and ( n51678 , n51677 , n32421 );
not ( n51679 , n50002 );
and ( n51680 , n51679 , n41286 );
and ( n51681 , n41298 , n50002 );
or ( n51682 , n51680 , n51681 );
and ( n51683 , n51682 , n32419 );
not ( n51684 , n50289 );
and ( n51685 , n51684 , n41286 );
and ( n51686 , n41298 , n50289 );
or ( n51687 , n51685 , n51686 );
and ( n51688 , n51687 , n32417 );
not ( n51689 , n50008 );
and ( n51690 , n51689 , n41286 );
and ( n51691 , n41298 , n50008 );
or ( n51692 , n51690 , n51691 );
and ( n51693 , n51692 , n32415 );
not ( n51694 , n47331 );
and ( n51695 , n51694 , n41286 );
and ( n51696 , n41288 , n47331 );
or ( n51697 , n51695 , n51696 );
and ( n51698 , n51697 , n32413 );
not ( n51699 , n50067 );
and ( n51700 , n51699 , n41286 );
and ( n51701 , n41288 , n50067 );
or ( n51702 , n51700 , n51701 );
and ( n51703 , n51702 , n32411 );
not ( n51704 , n31728 );
and ( n51705 , n51704 , n41286 );
and ( n51706 , n41290 , n31728 );
or ( n51707 , n51705 , n51706 );
and ( n51708 , n51707 , n32253 );
not ( n51709 , n32283 );
and ( n51710 , n51709 , n41286 );
and ( n51711 , n41307 , n32283 );
or ( n51712 , n51710 , n51711 );
and ( n51713 , n51712 , n32398 );
and ( n51714 , n41303 , n50334 );
or ( n51715 , n51673 , n51678 , n51683 , n51688 , n51693 , n51698 , n51703 , n51708 , n51713 , n51714 );
and ( n51716 , n51715 , n32456 );
and ( n51717 , n37573 , n32489 );
and ( n51718 , n41286 , n50345 );
or ( n51719 , C0 , n51716 , n51717 , n51718 );
buf ( n51720 , n51719 );
buf ( n51721 , n51720 );
buf ( n51722 , n30987 );
buf ( n51723 , n31655 );
not ( n51724 , n31437 );
buf ( n51725 , RI15b526b0_677);
and ( n51726 , n51724 , n51725 );
not ( n51727 , n45766 );
and ( n51728 , n51727 , n45592 );
xor ( n51729 , n45774 , n45782 );
and ( n51730 , n51729 , n45766 );
or ( n51731 , n51728 , n51730 );
and ( n51732 , n51731 , n31437 );
or ( n51733 , n51726 , n51732 );
and ( n51734 , n51733 , n31468 );
not ( n51735 , n44817 );
and ( n51736 , n51735 , n51725 );
not ( n51737 , n44994 );
and ( n51738 , n51737 , n44870 );
xor ( n51739 , n45006 , n45014 );
and ( n51740 , n51739 , n44994 );
or ( n51741 , n51738 , n51740 );
and ( n51742 , n51741 , n44817 );
or ( n51743 , n51736 , n51742 );
and ( n51744 , n51743 , n31521 );
and ( n51745 , n51725 , n42158 );
or ( n51746 , n51734 , n51744 , n51745 );
and ( n51747 , n51746 , n31557 );
and ( n51748 , n51725 , n40154 );
or ( n51749 , C0 , n51747 , n51748 );
buf ( n51750 , n51749 );
buf ( n51751 , n51750 );
not ( n51752 , n40163 );
and ( n51753 , n51752 , n31879 );
not ( n51754 , n49298 );
and ( n51755 , n51754 , n31879 );
and ( n51756 , n32218 , n49298 );
or ( n51757 , n51755 , n51756 );
and ( n51758 , n51757 , n40163 );
or ( n51759 , n51753 , n51758 );
and ( n51760 , n51759 , n32498 );
not ( n51761 , n49306 );
not ( n51762 , n49298 );
and ( n51763 , n51762 , n31879 );
and ( n51764 , n42255 , n49298 );
or ( n51765 , n51763 , n51764 );
and ( n51766 , n51761 , n51765 );
and ( n51767 , n42255 , n49306 );
or ( n51768 , n51766 , n51767 );
and ( n51769 , n51768 , n32473 );
not ( n51770 , n32475 );
not ( n51771 , n49306 );
not ( n51772 , n49298 );
and ( n51773 , n51772 , n31879 );
and ( n51774 , n42255 , n49298 );
or ( n51775 , n51773 , n51774 );
and ( n51776 , n51771 , n51775 );
and ( n51777 , n42255 , n49306 );
or ( n51778 , n51776 , n51777 );
and ( n51779 , n51770 , n51778 );
not ( n51780 , n49331 );
not ( n51781 , n49333 );
and ( n51782 , n51781 , n51778 );
and ( n51783 , n42283 , n49333 );
or ( n51784 , n51782 , n51783 );
and ( n51785 , n51780 , n51784 );
and ( n51786 , n42291 , n49331 );
or ( n51787 , n51785 , n51786 );
and ( n51788 , n51787 , n32475 );
or ( n51789 , n51779 , n51788 );
and ( n51790 , n51789 , n32486 );
and ( n51791 , n31879 , n41278 );
or ( n51792 , C0 , n51760 , n51769 , n51790 , n51791 );
buf ( n51793 , n51792 );
buf ( n51794 , n51793 );
buf ( n51795 , n30987 );
buf ( n51796 , n30987 );
xor ( n51797 , n41743 , n44786 );
and ( n51798 , n51797 , n31548 );
not ( n51799 , n44807 );
and ( n51800 , n51799 , n41743 );
and ( n51801 , n42046 , n44807 );
or ( n51802 , n51800 , n51801 );
and ( n51803 , n51802 , n31408 );
not ( n51804 , n44817 );
and ( n51805 , n51804 , n41743 );
not ( n51806 , n41835 );
buf ( n51807 , RI15b53100_699);
and ( n51808 , n51806 , n51807 );
not ( n51809 , n42124 );
and ( n51810 , n51809 , n42056 );
xor ( n51811 , n49377 , n49382 );
and ( n51812 , n51811 , n42124 );
or ( n51813 , n51810 , n51812 );
and ( n51814 , n51813 , n41835 );
or ( n51815 , n51808 , n51814 );
and ( n51816 , n51815 , n44817 );
or ( n51817 , n51805 , n51816 );
and ( n51818 , n51817 , n31521 );
not ( n51819 , n45059 );
and ( n51820 , n51819 , n41743 );
and ( n51821 , n42362 , n45059 );
or ( n51822 , n51820 , n51821 );
and ( n51823 , n51822 , n31536 );
and ( n51824 , n41743 , n45148 );
or ( n51825 , n51798 , n51803 , n51818 , n51823 , n51824 );
and ( n51826 , n51825 , n31557 );
and ( n51827 , n41743 , n40154 );
or ( n51828 , C0 , n51826 , n51827 );
buf ( n51829 , n51828 );
buf ( n51830 , n51829 );
buf ( n51831 , n31655 );
buf ( n51832 , n30987 );
xor ( n51833 , n41626 , n44777 );
and ( n51834 , n51833 , n31548 );
not ( n51835 , n44807 );
and ( n51836 , n51835 , n41626 );
and ( n51837 , n41902 , n44807 );
or ( n51838 , n51836 , n51837 );
and ( n51839 , n51838 , n31408 );
not ( n51840 , n44817 );
and ( n51841 , n51840 , n41626 );
not ( n51842 , n41835 );
buf ( n51843 , RI15b52cc8_690);
and ( n51844 , n51842 , n51843 );
not ( n51845 , n42124 );
and ( n51846 , n51845 , n41912 );
xor ( n51847 , n42133 , n42137 );
and ( n51848 , n51847 , n42124 );
or ( n51849 , n51846 , n51848 );
and ( n51850 , n51849 , n41835 );
or ( n51851 , n51844 , n51850 );
and ( n51852 , n51851 , n44817 );
or ( n51853 , n51841 , n51852 );
and ( n51854 , n51853 , n31521 );
not ( n51855 , n45059 );
and ( n51856 , n51855 , n41626 );
and ( n51857 , n33628 , n45059 );
or ( n51858 , n51856 , n51857 );
and ( n51859 , n51858 , n31536 );
and ( n51860 , n41626 , n45148 );
or ( n51861 , n51834 , n51839 , n51854 , n51859 , n51860 );
and ( n51862 , n51861 , n31557 );
and ( n51863 , n41626 , n40154 );
or ( n51864 , C0 , n51862 , n51863 );
buf ( n51865 , n51864 );
buf ( n51866 , n51865 );
buf ( n51867 , n31655 );
not ( n51868 , n40163 );
and ( n51869 , n51868 , n31842 );
not ( n51870 , n50540 );
and ( n51871 , n51870 , n31842 );
and ( n51872 , n32235 , n50540 );
or ( n51873 , n51871 , n51872 );
and ( n51874 , n51873 , n40163 );
or ( n51875 , n51869 , n51874 );
and ( n51876 , n51875 , n32498 );
not ( n51877 , n50548 );
not ( n51878 , n50540 );
and ( n51879 , n51878 , n31842 );
and ( n51880 , n42188 , n50540 );
or ( n51881 , n51879 , n51880 );
and ( n51882 , n51877 , n51881 );
and ( n51883 , n42188 , n50548 );
or ( n51884 , n51882 , n51883 );
and ( n51885 , n51884 , n32473 );
not ( n51886 , n32475 );
not ( n51887 , n50548 );
not ( n51888 , n50540 );
and ( n51889 , n51888 , n31842 );
and ( n51890 , n42188 , n50540 );
or ( n51891 , n51889 , n51890 );
and ( n51892 , n51887 , n51891 );
and ( n51893 , n42188 , n50548 );
or ( n51894 , n51892 , n51893 );
and ( n51895 , n51886 , n51894 );
not ( n51896 , n50568 );
not ( n51897 , n50570 );
and ( n51898 , n51897 , n51894 );
and ( n51899 , n42216 , n50570 );
or ( n51900 , n51898 , n51899 );
and ( n51901 , n51896 , n51900 );
and ( n51902 , n42224 , n50568 );
or ( n51903 , n51901 , n51902 );
and ( n51904 , n51903 , n32475 );
or ( n51905 , n51895 , n51904 );
and ( n51906 , n51905 , n32486 );
and ( n51907 , n31842 , n41278 );
or ( n51908 , C0 , n51876 , n51885 , n51906 , n51907 );
buf ( n51909 , n51908 );
buf ( n51910 , n51909 );
buf ( n51911 , n30987 );
not ( n51912 , n32953 );
buf ( n51913 , RI15b46ba8_278);
and ( n51914 , n51912 , n51913 );
not ( n51915 , n39572 );
and ( n51916 , n51915 , n39490 );
xor ( n51917 , n42619 , n42634 );
and ( n51918 , n51917 , n39572 );
or ( n51919 , n51916 , n51918 );
and ( n51920 , n51919 , n32953 );
or ( n51921 , n51914 , n51920 );
and ( n51922 , n51921 , n33038 );
not ( n51923 , n39586 );
and ( n51924 , n51923 , n51913 );
not ( n51925 , n39775 );
and ( n51926 , n51925 , n39699 );
xor ( n51927 , n42655 , n42670 );
and ( n51928 , n51927 , n39775 );
or ( n51929 , n51926 , n51928 );
and ( n51930 , n51929 , n39586 );
or ( n51931 , n51924 , n51930 );
and ( n51932 , n51931 , n33172 );
and ( n51933 , n51913 , n39795 );
or ( n51934 , n51922 , n51932 , n51933 );
and ( n51935 , n51934 , n33208 );
and ( n51936 , n51913 , n39805 );
or ( n51937 , C0 , n51935 , n51936 );
buf ( n51938 , n51937 );
buf ( n51939 , n51938 );
buf ( n51940 , n30987 );
buf ( n51941 , n31655 );
buf ( n51942 , n31655 );
buf ( n51943 , n30987 );
and ( n51944 , n33221 , n32528 );
not ( n51945 , n32598 );
and ( n51946 , n51945 , n32984 );
buf ( n51947 , n51946 );
and ( n51948 , n51947 , n32890 );
not ( n51949 , n32919 );
and ( n51950 , n51949 , n32984 );
buf ( n51951 , n51950 );
and ( n51952 , n51951 , n32924 );
not ( n51953 , n32953 );
and ( n51954 , n51953 , n32984 );
not ( n51955 , n32971 );
and ( n51956 , n51955 , n33093 );
xor ( n51957 , n32984 , n33021 );
and ( n51958 , n51957 , n32971 );
or ( n51959 , n51956 , n51958 );
and ( n51960 , n51959 , n32953 );
or ( n51961 , n51954 , n51960 );
and ( n51962 , n51961 , n33038 );
not ( n51963 , n33067 );
and ( n51964 , n51963 , n32984 );
not ( n51965 , n32970 );
not ( n51966 , n33071 );
and ( n51967 , n51966 , n33093 );
xor ( n51968 , n33094 , n33153 );
and ( n51969 , n51968 , n33071 );
or ( n51970 , n51967 , n51969 );
and ( n51971 , n51965 , n51970 );
and ( n51972 , n51957 , n32970 );
or ( n51973 , n51971 , n51972 );
and ( n51974 , n51973 , n33067 );
or ( n51975 , n51964 , n51974 );
and ( n51976 , n51975 , n33172 );
and ( n51977 , n32984 , n33204 );
or ( n51978 , n51948 , n51952 , n51962 , n51976 , n51977 );
and ( n51979 , n51978 , n33208 );
not ( n51980 , n32968 );
not ( n51981 , n33270 );
and ( n51982 , n51981 , n33293 );
xor ( n51983 , n33294 , n33353 );
and ( n51984 , n51983 , n33270 );
or ( n51985 , n51982 , n51984 );
and ( n51986 , n51980 , n51985 );
and ( n51987 , n32984 , n32968 );
or ( n51988 , n51986 , n51987 );
and ( n51989 , n51988 , n33370 );
and ( n51990 , n32984 , n33382 );
or ( n51991 , C0 , n51944 , n51979 , n51989 , C0 , n51990 );
buf ( n51992 , n51991 );
buf ( n51993 , n51992 );
buf ( n51994 , n30987 );
buf ( n51995 , n31655 );
not ( n51996 , n31728 );
and ( n51997 , n51996 , n46029 );
xor ( n51998 , n47606 , n47623 );
and ( n51999 , n51998 , n31728 );
or ( n52000 , n51997 , n51999 );
and ( n52001 , n52000 , n32253 );
not ( n52002 , n32283 );
and ( n52003 , n52002 , n46029 );
not ( n52004 , n31823 );
xor ( n52005 , n47661 , n47678 );
and ( n52006 , n52004 , n52005 );
xnor ( n52007 , n47711 , n47728 );
and ( n52008 , n52007 , n31823 );
or ( n52009 , n52006 , n52008 );
and ( n52010 , n52009 , n32283 );
or ( n52011 , n52003 , n52010 );
and ( n52012 , n52011 , n32398 );
and ( n52013 , n46029 , n32436 );
or ( n52014 , n52001 , n52012 , n52013 );
and ( n52015 , n52014 , n32456 );
and ( n52016 , n49675 , n32473 );
not ( n52017 , n32475 );
and ( n52018 , n52017 , n49675 );
xor ( n52019 , n46029 , n47757 );
and ( n52020 , n52019 , n32475 );
or ( n52021 , n52018 , n52020 );
and ( n52022 , n52021 , n32486 );
and ( n52023 , n37555 , n32489 );
and ( n52024 , n46029 , n32501 );
or ( n52025 , C0 , n52015 , n52016 , n52022 , n52023 , n52024 );
buf ( n52026 , n52025 );
buf ( n52027 , n52026 );
buf ( n52028 , n31655 );
buf ( n52029 , n30987 );
and ( n52030 , n33225 , n32528 );
not ( n52031 , n32598 );
and ( n52032 , n52031 , n32988 );
buf ( n52033 , n52032 );
and ( n52034 , n52033 , n32890 );
not ( n52035 , n32919 );
and ( n52036 , n52035 , n32988 );
buf ( n52037 , n52036 );
and ( n52038 , n52037 , n32924 );
not ( n52039 , n32953 );
and ( n52040 , n52039 , n32988 );
not ( n52041 , n32971 );
and ( n52042 , n52041 , n33101 );
xor ( n52043 , n32988 , n33017 );
and ( n52044 , n52043 , n32971 );
or ( n52045 , n52042 , n52044 );
and ( n52046 , n52045 , n32953 );
or ( n52047 , n52040 , n52046 );
and ( n52048 , n52047 , n33038 );
not ( n52049 , n33067 );
and ( n52050 , n52049 , n32988 );
not ( n52051 , n32970 );
not ( n52052 , n33071 );
and ( n52053 , n52052 , n33101 );
xor ( n52054 , n33102 , n33149 );
and ( n52055 , n52054 , n33071 );
or ( n52056 , n52053 , n52055 );
and ( n52057 , n52051 , n52056 );
and ( n52058 , n52043 , n32970 );
or ( n52059 , n52057 , n52058 );
and ( n52060 , n52059 , n33067 );
or ( n52061 , n52050 , n52060 );
and ( n52062 , n52061 , n33172 );
and ( n52063 , n32988 , n33204 );
or ( n52064 , n52034 , n52038 , n52048 , n52062 , n52063 );
and ( n52065 , n52064 , n33208 );
not ( n52066 , n32968 );
not ( n52067 , n33270 );
and ( n52068 , n52067 , n33301 );
xor ( n52069 , n33302 , n33349 );
and ( n52070 , n52069 , n33270 );
or ( n52071 , n52068 , n52070 );
and ( n52072 , n52066 , n52071 );
and ( n52073 , n32988 , n32968 );
or ( n52074 , n52072 , n52073 );
and ( n52075 , n52074 , n33370 );
buf ( n52076 , n35056 );
and ( n52077 , n32988 , n33382 );
or ( n52078 , C0 , n52030 , n52065 , n52075 , n52076 , n52077 );
buf ( n52079 , n52078 );
buf ( n52080 , n52079 );
not ( n52081 , n31728 );
and ( n52082 , n52081 , n46025 );
xor ( n52083 , n47602 , n47627 );
and ( n52084 , n52083 , n31728 );
or ( n52085 , n52082 , n52084 );
and ( n52086 , n52085 , n32253 );
not ( n52087 , n32283 );
and ( n52088 , n52087 , n46025 );
not ( n52089 , n31823 );
xor ( n52090 , n47657 , n47682 );
and ( n52091 , n52089 , n52090 );
xnor ( n52092 , n47707 , n47732 );
and ( n52093 , n52092 , n31823 );
or ( n52094 , n52091 , n52093 );
and ( n52095 , n52094 , n32283 );
or ( n52096 , n52088 , n52095 );
and ( n52097 , n52096 , n32398 );
and ( n52098 , n46025 , n32436 );
or ( n52099 , n52086 , n52097 , n52098 );
and ( n52100 , n52099 , n32456 );
and ( n52101 , n49667 , n32473 );
not ( n52102 , n32475 );
and ( n52103 , n52102 , n49667 );
xor ( n52104 , n46025 , n47761 );
and ( n52105 , n52104 , n32475 );
or ( n52106 , n52103 , n52105 );
and ( n52107 , n52106 , n32486 );
and ( n52108 , n37547 , n32489 );
and ( n52109 , n46025 , n32501 );
or ( n52110 , C0 , n52100 , n52101 , n52107 , n52108 , n52109 );
buf ( n52111 , n52110 );
buf ( n52112 , n52111 );
buf ( n52113 , n30987 );
buf ( n52114 , n31655 );
buf ( n52115 , n31655 );
buf ( n52116 , n30987 );
buf ( n52117 , n30987 );
not ( n52118 , n40163 );
and ( n52119 , n52118 , n32050 );
and ( n52120 , n42169 , n42237 , n45160 , n31661 , n42170 );
not ( n52121 , n52120 );
and ( n52122 , n52121 , n32050 );
and ( n52123 , n32130 , n52120 );
or ( n52124 , n52122 , n52123 );
and ( n52125 , n52124 , n40163 );
or ( n52126 , n52119 , n52125 );
and ( n52127 , n52126 , n32498 );
and ( n52128 , n42179 , n42246 , n45169 , n40194 , C1 );
not ( n52129 , n52128 );
not ( n52130 , n52120 );
and ( n52131 , n52130 , n32050 );
and ( n52132 , n45833 , n52120 );
or ( n52133 , n52131 , n52132 );
and ( n52134 , n52129 , n52133 );
and ( n52135 , n45833 , n52128 );
or ( n52136 , n52134 , n52135 );
and ( n52137 , n52136 , n32473 );
not ( n52138 , n32475 );
not ( n52139 , n52128 );
not ( n52140 , n52120 );
and ( n52141 , n52140 , n32050 );
and ( n52142 , n45833 , n52120 );
or ( n52143 , n52141 , n52142 );
and ( n52144 , n52139 , n52143 );
and ( n52145 , n45833 , n52128 );
or ( n52146 , n52144 , n52145 );
and ( n52147 , n52138 , n52146 );
and ( n52148 , n42205 , n42272 , n45195 , n40445 , C1 );
not ( n52149 , n52148 );
and ( n52150 , n42208 , n42275 , n45198 , n40440 , C1 );
not ( n52151 , n52150 );
and ( n52152 , n52151 , n52146 );
and ( n52153 , n45857 , n52150 );
or ( n52154 , n52152 , n52153 );
and ( n52155 , n52149 , n52154 );
and ( n52156 , n45865 , n52148 );
or ( n52157 , n52155 , n52156 );
and ( n52158 , n52157 , n32475 );
or ( n52159 , n52147 , n52158 );
and ( n52160 , n52159 , n32486 );
and ( n52161 , n32050 , n41278 );
or ( n52162 , C0 , n52127 , n52137 , n52160 , n52161 );
buf ( n52163 , n52162 );
buf ( n52164 , n52163 );
buf ( n52165 , n31655 );
not ( n52166 , n41606 );
and ( n52167 , n52166 , n31548 );
not ( n52168 , n44807 );
and ( n52169 , n52168 , n41606 );
and ( n52170 , n41873 , n44807 );
or ( n52171 , n52169 , n52170 );
and ( n52172 , n52171 , n31408 );
not ( n52173 , n44817 );
and ( n52174 , n52173 , n41606 );
not ( n52175 , n41835 );
buf ( n52176 , RI15b52bd8_688);
and ( n52177 , n52175 , n52176 );
not ( n52178 , n42124 );
and ( n52179 , n52178 , n41877 );
xor ( n52180 , n42135 , n41881 );
and ( n52181 , n52180 , n42124 );
or ( n52182 , n52179 , n52181 );
and ( n52183 , n52182 , n41835 );
or ( n52184 , n52177 , n52183 );
and ( n52185 , n52184 , n44817 );
or ( n52186 , n52174 , n52185 );
and ( n52187 , n52186 , n31521 );
not ( n52188 , n45059 );
and ( n52189 , n52188 , n41606 );
and ( n52190 , n33666 , n45059 );
or ( n52191 , n52189 , n52190 );
and ( n52192 , n52191 , n31536 );
and ( n52193 , n41606 , n45148 );
or ( n52194 , n52167 , n52172 , n52187 , n52192 , n52193 );
and ( n52195 , n52194 , n31557 );
and ( n52196 , n41606 , n40154 );
or ( n52197 , C0 , n52195 , n52196 );
buf ( n52198 , n52197 );
buf ( n52199 , n52198 );
buf ( n52200 , n30987 );
buf ( n52201 , n31655 );
buf ( n52202 , n31655 );
buf ( n52203 , n30987 );
not ( n52204 , n50828 );
not ( n52205 , n50834 );
and ( n52206 , n52205 , n40583 );
buf ( n52207 , RI15b53f88_730);
and ( n52208 , n52207 , n50834 );
or ( n52209 , n52206 , n52208 );
and ( n52210 , n52204 , n52209 );
buf ( n52211 , RI15b603f0_1149);
and ( n52212 , n52211 , n50828 );
or ( n52213 , n52210 , n52212 );
buf ( n52214 , n52213 );
buf ( n52215 , n52214 );
and ( n52216 , n33127 , n41543 );
and ( n52217 , n33125 , n52216 );
and ( n52218 , n33123 , n52217 );
and ( n52219 , n33121 , n52218 );
and ( n52220 , n33119 , n52219 );
and ( n52221 , n33117 , n52220 );
and ( n52222 , n33115 , n52221 );
and ( n52223 , n33113 , n52222 );
and ( n52224 , n33111 , n52223 );
xor ( n52225 , n33109 , n52224 );
and ( n52226 , n52225 , n33201 );
not ( n52227 , n41576 );
and ( n52228 , n52227 , n33109 );
not ( n52229 , n32547 );
buf ( n52230 , n52229 );
not ( n52231 , n52230 );
not ( n52232 , n52231 );
not ( n52233 , n32543 );
not ( n52234 , n52233 );
buf ( n52235 , n52234 );
buf ( n52236 , n52235 );
not ( n52237 , n52236 );
not ( n52238 , n52237 );
xor ( n52239 , n32539 , n32543 );
not ( n52240 , n52239 );
buf ( n52241 , n52240 );
buf ( n52242 , n52241 );
not ( n52243 , n52242 );
not ( n52244 , n52243 );
and ( n52245 , n32539 , n32543 );
xor ( n52246 , n32535 , n52245 );
not ( n52247 , n52246 );
buf ( n52248 , n52247 );
buf ( n52249 , n52248 );
not ( n52250 , n52249 );
not ( n52251 , n52250 );
nor ( n52252 , n52232 , n52238 , n52244 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52253 , n32757 , n52252 );
nor ( n52254 , n52231 , n52238 , n52244 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52255 , n32759 , n52254 );
nor ( n52256 , n52232 , n52237 , n52244 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52257 , n32761 , n52256 );
nor ( n52258 , n52231 , n52237 , n52244 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52259 , n32763 , n52258 );
nor ( n52260 , n52232 , n52238 , n52243 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52261 , n32765 , n52260 );
nor ( n52262 , n52231 , n52238 , n52243 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52263 , n32767 , n52262 );
nor ( n52264 , n52232 , n52237 , n52243 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52265 , n32769 , n52264 );
nor ( n52266 , n52231 , n52237 , n52243 , n52251 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52267 , n32771 , n52266 );
nor ( n52268 , n52232 , n52238 , n52244 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52269 , n32773 , n52268 );
nor ( n52270 , n52231 , n52238 , n52244 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52271 , n32775 , n52270 );
nor ( n52272 , n52232 , n52237 , n52244 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52273 , n32777 , n52272 );
nor ( n52274 , n52231 , n52237 , n52244 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52275 , n32779 , n52274 );
nor ( n52276 , n52232 , n52238 , n52243 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52277 , n32781 , n52276 );
nor ( n52278 , n52231 , n52238 , n52243 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52279 , n32783 , n52278 );
nor ( n52280 , n52232 , n52237 , n52243 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52281 , n32785 , n52280 );
nor ( n52282 , n52231 , n52237 , n52243 , n52250 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n52283 , n32787 , n52282 );
or ( n52284 , n52253 , n52255 , n52257 , n52259 , n52261 , n52263 , n52265 , n52267 , n52269 , n52271 , n52273 , n52275 , n52277 , n52279 , n52281 , n52283 );
and ( n52285 , n52284 , n41576 );
or ( n52286 , n52228 , n52285 );
and ( n52287 , n52286 , n33189 );
and ( n52288 , n33109 , n41592 );
or ( n52289 , n52226 , n52287 , n52288 );
and ( n52290 , n52289 , n33208 );
and ( n52291 , n33109 , n39805 );
or ( n52292 , C0 , n52290 , n52291 );
buf ( n52293 , n52292 );
buf ( n52294 , n52293 );
buf ( n52295 , n30987 );
buf ( n52296 , n30987 );
not ( n52297 , n43755 );
and ( n52298 , n52297 , n43734 );
xor ( n52299 , n43734 , n43259 );
xor ( n52300 , n43717 , n43259 );
xor ( n52301 , n43700 , n43259 );
xor ( n52302 , n43683 , n43259 );
xor ( n52303 , n43666 , n43259 );
xor ( n52304 , n43649 , n43259 );
xor ( n52305 , n43632 , n43259 );
xor ( n52306 , n43615 , n43259 );
xor ( n52307 , n43598 , n43259 );
xor ( n52308 , n43581 , n43259 );
xor ( n52309 , n43564 , n43259 );
xor ( n52310 , n43547 , n43259 );
xor ( n52311 , n43530 , n43259 );
xor ( n52312 , n43513 , n43259 );
xor ( n52313 , n43496 , n43259 );
xor ( n52314 , n43479 , n43259 );
and ( n52315 , n50497 , n50508 );
and ( n52316 , n52314 , n52315 );
and ( n52317 , n52313 , n52316 );
and ( n52318 , n52312 , n52317 );
and ( n52319 , n52311 , n52318 );
and ( n52320 , n52310 , n52319 );
and ( n52321 , n52309 , n52320 );
and ( n52322 , n52308 , n52321 );
and ( n52323 , n52307 , n52322 );
and ( n52324 , n52306 , n52323 );
and ( n52325 , n52305 , n52324 );
and ( n52326 , n52304 , n52325 );
and ( n52327 , n52303 , n52326 );
and ( n52328 , n52302 , n52327 );
and ( n52329 , n52301 , n52328 );
and ( n52330 , n52300 , n52329 );
xor ( n52331 , n52299 , n52330 );
and ( n52332 , n52331 , n43755 );
or ( n52333 , n52298 , n52332 );
and ( n52334 , n52333 , n43774 );
not ( n52335 , n44663 );
and ( n52336 , n52335 , n44646 );
xor ( n52337 , n44646 , n44171 );
xor ( n52338 , n44629 , n44171 );
xor ( n52339 , n44612 , n44171 );
xor ( n52340 , n44595 , n44171 );
xor ( n52341 , n44578 , n44171 );
xor ( n52342 , n44561 , n44171 );
xor ( n52343 , n44544 , n44171 );
xor ( n52344 , n44527 , n44171 );
xor ( n52345 , n44510 , n44171 );
xor ( n52346 , n44493 , n44171 );
xor ( n52347 , n44476 , n44171 );
xor ( n52348 , n44459 , n44171 );
xor ( n52349 , n44442 , n44171 );
xor ( n52350 , n44425 , n44171 );
xor ( n52351 , n44408 , n44171 );
xor ( n52352 , n44391 , n44171 );
and ( n52353 , n50515 , n50526 );
and ( n52354 , n52352 , n52353 );
and ( n52355 , n52351 , n52354 );
and ( n52356 , n52350 , n52355 );
and ( n52357 , n52349 , n52356 );
and ( n52358 , n52348 , n52357 );
and ( n52359 , n52347 , n52358 );
and ( n52360 , n52346 , n52359 );
and ( n52361 , n52345 , n52360 );
and ( n52362 , n52344 , n52361 );
and ( n52363 , n52343 , n52362 );
and ( n52364 , n52342 , n52363 );
and ( n52365 , n52341 , n52364 );
and ( n52366 , n52340 , n52365 );
and ( n52367 , n52339 , n52366 );
and ( n52368 , n52338 , n52367 );
xor ( n52369 , n52337 , n52368 );
and ( n52370 , n52369 , n44663 );
or ( n52371 , n52336 , n52370 );
and ( n52372 , n52371 , n44682 );
buf ( n52373 , RI15b45d98_248);
and ( n52374 , n52373 , n44695 );
or ( n52375 , n52334 , n52372 , n52374 );
buf ( n52376 , n52375 );
buf ( n52377 , n52376 );
buf ( n52378 , n30987 );
buf ( n52379 , n31655 );
buf ( n52380 , n31655 );
buf ( n52381 , n31655 );
buf ( n52382 , n30987 );
not ( n52383 , n46356 );
and ( n52384 , n52383 , n31025 );
and ( n52385 , n46373 , n46356 );
or ( n52386 , n52384 , n52385 );
and ( n52387 , n52386 , n31649 );
not ( n52388 , n44702 );
and ( n52389 , n52388 , n31010 );
buf ( n52390 , n52389 );
not ( n52391 , n52390 );
not ( n52392 , n44702 );
and ( n52393 , n52392 , n31018 );
buf ( n52394 , RI15b50dd8_624);
not ( n52395 , n52394 );
buf ( n52396 , RI15b50d60_623);
not ( n52397 , n52396 );
buf ( n52398 , RI15b50ce8_622);
not ( n52399 , n52398 );
buf ( n52400 , RI15b50c70_621);
not ( n52401 , n52400 );
buf ( n52402 , RI15b50bf8_620);
not ( n52403 , n52402 );
buf ( n52404 , RI15b50b80_619);
not ( n52405 , n52404 );
not ( n52406 , n42376 );
not ( n52407 , n42377 );
not ( n52408 , n42378 );
not ( n52409 , n42379 );
not ( n52410 , n33422 );
not ( n52411 , n33423 );
not ( n52412 , n33424 );
not ( n52413 , n33425 );
not ( n52414 , n33426 );
not ( n52415 , n33427 );
not ( n52416 , n33428 );
not ( n52417 , n33429 );
not ( n52418 , n33430 );
not ( n52419 , n33431 );
not ( n52420 , n33432 );
not ( n52421 , n33433 );
not ( n52422 , n33434 );
not ( n52423 , n33435 );
not ( n52424 , n33436 );
not ( n52425 , n33437 );
not ( n52426 , n33438 );
not ( n52427 , n33439 );
not ( n52428 , n33440 );
not ( n52429 , n33441 );
not ( n52430 , n33442 );
not ( n52431 , n33443 );
and ( n52432 , n52430 , n52431 );
and ( n52433 , n52429 , n52432 );
and ( n52434 , n52428 , n52433 );
and ( n52435 , n52427 , n52434 );
and ( n52436 , n52426 , n52435 );
and ( n52437 , n52425 , n52436 );
and ( n52438 , n52424 , n52437 );
and ( n52439 , n52423 , n52438 );
and ( n52440 , n52422 , n52439 );
and ( n52441 , n52421 , n52440 );
and ( n52442 , n52420 , n52441 );
and ( n52443 , n52419 , n52442 );
and ( n52444 , n52418 , n52443 );
and ( n52445 , n52417 , n52444 );
and ( n52446 , n52416 , n52445 );
and ( n52447 , n52415 , n52446 );
and ( n52448 , n52414 , n52447 );
and ( n52449 , n52413 , n52448 );
and ( n52450 , n52412 , n52449 );
and ( n52451 , n52411 , n52450 );
and ( n52452 , n52410 , n52451 );
and ( n52453 , n52409 , n52452 );
and ( n52454 , n52408 , n52453 );
and ( n52455 , n52407 , n52454 );
and ( n52456 , n52406 , n52455 );
and ( n52457 , n52405 , n52456 );
and ( n52458 , n52403 , n52457 );
and ( n52459 , n52401 , n52458 );
and ( n52460 , n52399 , n52459 );
and ( n52461 , n52397 , n52460 );
xor ( n52462 , n52395 , n52461 );
buf ( n52463 , n52394 );
and ( n52464 , n52462 , n52463 );
buf ( n52465 , n52464 );
not ( n52466 , n52465 );
not ( n52467 , n52394 );
and ( n52468 , n52467 , n33442 );
xor ( n52469 , n52430 , n52431 );
and ( n52470 , n52469 , n52394 );
or ( n52471 , n52468 , n52470 );
and ( n52472 , n52466 , n52471 );
not ( n52473 , n52471 );
buf ( n52474 , n33443 );
not ( n52475 , n52474 );
xor ( n52476 , n52473 , n52475 );
and ( n52477 , n52476 , n52465 );
or ( n52478 , n52472 , n52477 );
not ( n52479 , n52478 );
buf ( n52480 , n52479 );
buf ( n52481 , n52480 );
not ( n52482 , n52481 );
xor ( n52483 , n52482 , n52465 );
buf ( n52484 , n52474 );
not ( n52485 , n52484 );
buf ( n52486 , n52485 );
not ( n52487 , n52486 );
xor ( n52488 , n52487 , n52465 );
and ( n52489 , n52488 , n52465 );
and ( n52490 , n52483 , n52489 );
buf ( n52491 , n52490 );
or ( n52492 , n52487 , n52482 );
buf ( n52493 , n52492 );
buf ( n52494 , n52493 );
and ( n52495 , n52494 , n52465 );
and ( n52496 , n52491 , n52495 );
buf ( n52497 , n52496 );
not ( n52498 , n52495 );
and ( n52499 , n52498 , n52482 );
xor ( n52500 , n52483 , n52489 );
and ( n52501 , n52500 , n52495 );
or ( n52502 , n52499 , n52501 );
not ( n52503 , n52495 );
and ( n52504 , n52503 , n52487 );
xor ( n52505 , n52488 , n52465 );
and ( n52506 , n52505 , n52495 );
or ( n52507 , n52504 , n52506 );
and ( n52508 , n52502 , n52507 );
xor ( n52509 , n52497 , n52508 );
buf ( n52510 , n52509 );
buf ( n52511 , n52510 );
not ( n52512 , n52511 );
buf ( n52513 , n52512 );
buf ( n52514 , n52513 );
not ( n52515 , n52514 );
buf ( n52516 , n52515 );
buf ( n52517 , n52516 );
buf ( n52518 , n52474 );
not ( n52519 , n52518 );
buf ( n52520 , n52519 );
not ( n52521 , n52520 );
buf ( n52522 , n52521 );
buf ( n52523 , n52522 );
and ( n52524 , n52523 , n52465 );
not ( n52525 , n52524 );
and ( n52526 , n52525 , n52521 );
xor ( n52527 , n52521 , n52465 );
xor ( n52528 , n52527 , n52465 );
and ( n52529 , n52528 , n52524 );
or ( n52530 , n52526 , n52529 );
not ( n52531 , n52530 );
not ( n52532 , n52531 );
and ( n52533 , n52517 , n52532 );
buf ( n52534 , n52533 );
and ( n52535 , n52534 , n44702 );
or ( n52536 , n52393 , n52535 );
not ( n52537 , n52536 );
not ( n52538 , n44702 );
and ( n52539 , n52538 , n31014 );
and ( n52540 , n52497 , n52508 );
buf ( n52541 , n52540 );
buf ( n52542 , n52541 );
not ( n52543 , n52542 );
buf ( n52544 , n52543 );
buf ( n52545 , n52544 );
not ( n52546 , n52545 );
buf ( n52547 , n52546 );
buf ( n52548 , n52547 );
and ( n52549 , n52548 , n52532 );
buf ( n52550 , n52549 );
and ( n52551 , n52550 , n44702 );
or ( n52552 , n52539 , n52551 );
not ( n52553 , n52552 );
buf ( n52554 , n52390 );
buf ( n52555 , n52390 );
buf ( n52556 , n52390 );
buf ( n52557 , n52390 );
buf ( n52558 , n52390 );
buf ( n52559 , n52390 );
buf ( n52560 , n52390 );
buf ( n52561 , n52390 );
buf ( n52562 , n52390 );
buf ( n52563 , n52390 );
buf ( n52564 , n52390 );
buf ( n52565 , n52390 );
buf ( n52566 , n52390 );
buf ( n52567 , n52390 );
buf ( n52568 , n52390 );
buf ( n52569 , n52390 );
buf ( n52570 , n52390 );
buf ( n52571 , n52390 );
buf ( n52572 , n52390 );
buf ( n52573 , n52390 );
buf ( n52574 , n52390 );
buf ( n52575 , n52390 );
buf ( n52576 , n52390 );
buf ( n52577 , n52390 );
buf ( n52578 , n52390 );
buf ( n52579 , n52390 );
not ( n52580 , n44702 );
and ( n52581 , n52580 , n31026 );
not ( n52582 , n52532 );
buf ( n52583 , n52582 );
not ( n52584 , n52507 );
buf ( n52585 , n52584 );
not ( n52586 , n52585 );
buf ( n52587 , n52586 );
not ( n52588 , n52587 );
buf ( n52589 , n52588 );
buf ( n52590 , n52589 );
and ( n52591 , n52590 , n52532 );
or ( n52592 , n52583 , n52591 );
and ( n52593 , n52592 , n44702 );
or ( n52594 , n52581 , n52593 );
not ( n52595 , n52594 );
not ( n52596 , n44702 );
and ( n52597 , n52596 , n31022 );
xor ( n52598 , n52502 , n52507 );
buf ( n52599 , n52598 );
buf ( n52600 , n52599 );
not ( n52601 , n52600 );
buf ( n52602 , n52601 );
buf ( n52603 , n52602 );
not ( n52604 , n52603 );
buf ( n52605 , n52604 );
buf ( n52606 , n52605 );
and ( n52607 , n52606 , n52532 );
buf ( n52608 , n52607 );
and ( n52609 , n52608 , n44702 );
or ( n52610 , n52597 , n52609 );
not ( n52611 , n52610 );
and ( n52612 , n52595 , n52611 );
or ( n52613 , n52537 , n52553 , n52390 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52612 );
nand ( n52614 , n52391 , n52613 );
not ( n52615 , n52614 );
not ( n52616 , n44702 );
and ( n52617 , n52616 , n31025 );
buf ( n52618 , n44702 );
or ( n52619 , n52617 , n52618 );
and ( n52620 , n52615 , n52619 );
buf ( n52621 , n52620 );
and ( n52622 , n52621 , n31647 );
and ( n52623 , n46515 , n31643 );
buf ( n52624 , n46515 );
and ( n52625 , n52624 , n31638 );
or ( n52626 , n47275 , n31007 );
and ( n52627 , n31025 , n52626 );
or ( n52628 , C0 , n52387 , n52622 , n52623 , n52625 , n52627 );
buf ( n52629 , n52628 );
buf ( n52630 , n52629 );
buf ( n52631 , n30987 );
buf ( n52632 , n31655 );
not ( n52633 , n31728 );
and ( n52634 , n52633 , n32460 );
xor ( n52635 , n31860 , n31893 );
xor ( n52636 , n52635 , n32081 );
and ( n52637 , n52636 , n31728 );
or ( n52638 , n52634 , n52637 );
and ( n52639 , n52638 , n32253 );
not ( n52640 , n32283 );
and ( n52641 , n52640 , n32460 );
not ( n52642 , n31823 );
xor ( n52643 , n32298 , n31893 );
xor ( n52644 , n52643 , n32320 );
and ( n52645 , n52642 , n52644 );
xor ( n52646 , n32348 , n32350 );
xor ( n52647 , n52646 , n32383 );
and ( n52648 , n52647 , n31823 );
or ( n52649 , n52645 , n52648 );
and ( n52650 , n52649 , n32283 );
or ( n52651 , n52641 , n52650 );
and ( n52652 , n52651 , n32398 );
and ( n52653 , n32460 , n32436 );
or ( n52654 , n52639 , n52652 , n52653 );
and ( n52655 , n52654 , n32456 );
and ( n52656 , n49697 , n32473 );
not ( n52657 , n32475 );
and ( n52658 , n52657 , n49697 );
xor ( n52659 , n32460 , n32479 );
and ( n52660 , n52659 , n32475 );
or ( n52661 , n52658 , n52660 );
and ( n52662 , n52661 , n32486 );
and ( n52663 , n37579 , n32489 );
and ( n52664 , n32460 , n32501 );
or ( n52665 , C0 , n52655 , n52656 , n52662 , n52663 , n52664 );
buf ( n52666 , n52665 );
buf ( n52667 , n52666 );
buf ( n52668 , n31655 );
buf ( n52669 , RI15b475f8_300);
buf ( n52670 , n52669 );
not ( n52671 , n34150 );
and ( n52672 , n52671 , n32704 );
not ( n52673 , n41392 );
and ( n52674 , n52673 , n32704 );
and ( n52675 , n32722 , n41392 );
or ( n52676 , n52674 , n52675 );
and ( n52677 , n52676 , n34150 );
or ( n52678 , n52672 , n52677 );
and ( n52679 , n52678 , n33381 );
not ( n52680 , n41402 );
not ( n52681 , n41392 );
and ( n52682 , n52681 , n32704 );
and ( n52683 , n42565 , n41392 );
or ( n52684 , n52682 , n52683 );
and ( n52685 , n52680 , n52684 );
and ( n52686 , n42565 , n41402 );
or ( n52687 , n52685 , n52686 );
and ( n52688 , n52687 , n33375 );
not ( n52689 , n32968 );
not ( n52690 , n41402 );
not ( n52691 , n41392 );
and ( n52692 , n52691 , n32704 );
and ( n52693 , n42565 , n41392 );
or ( n52694 , n52692 , n52693 );
and ( n52695 , n52690 , n52694 );
and ( n52696 , n42565 , n41402 );
or ( n52697 , n52695 , n52696 );
and ( n52698 , n52689 , n52697 );
not ( n52699 , n41424 );
not ( n52700 , n41428 );
and ( n52701 , n52700 , n52697 );
and ( n52702 , n42589 , n41428 );
or ( n52703 , n52701 , n52702 );
and ( n52704 , n52699 , n52703 );
and ( n52705 , n42597 , n41424 );
or ( n52706 , n52704 , n52705 );
and ( n52707 , n52706 , n32968 );
or ( n52708 , n52698 , n52707 );
and ( n52709 , n52708 , n33370 );
and ( n52710 , n32704 , n35062 );
or ( n52711 , C0 , n52679 , n52688 , n52709 , n52710 );
buf ( n52712 , n52711 );
buf ( n52713 , n52712 );
buf ( n52714 , n31655 );
buf ( n52715 , n30987 );
buf ( n52716 , n30987 );
buf ( n52717 , n30987 );
buf ( n52718 , n31655 );
buf ( n52719 , RI15b3fab0_37);
or ( n52720 , n39352 , n39354 );
and ( n52721 , n52719 , n52720 );
buf ( n52722 , n39350 );
or ( n52723 , n39349 , n39346 );
or ( n52724 , n52723 , n39356 );
or ( n52725 , n52724 , n38450 );
or ( n52726 , n52725 , n39358 );
and ( n52727 , n32475 , n52726 );
or ( n52728 , n52721 , n52722 , n52727 );
buf ( n52729 , n52728 );
buf ( n52730 , n52729 );
buf ( n52731 , n31655 );
not ( n52732 , n46356 );
and ( n52733 , n52732 , n31319 );
and ( n52734 , n31025 , n46360 , n48213 , n31013 , n46361 );
not ( n52735 , n52734 );
and ( n52736 , n52735 , n31319 );
and ( n52737 , n31339 , n52734 );
or ( n52738 , n52736 , n52737 );
and ( n52739 , n52738 , n46356 );
or ( n52740 , n52733 , n52739 );
and ( n52741 , n52740 , n31649 );
and ( n52742 , n46373 , n46380 , n48222 , n46392 , C1 );
not ( n52743 , n52742 );
not ( n52744 , n52734 );
and ( n52745 , n52744 , n31319 );
and ( n52746 , n47449 , n52734 );
or ( n52747 , n52745 , n52746 );
and ( n52748 , n52743 , n52747 );
and ( n52749 , n47449 , n52742 );
or ( n52750 , n52748 , n52749 );
and ( n52751 , n52750 , n31643 );
not ( n52752 , n31452 );
not ( n52753 , n52742 );
not ( n52754 , n52734 );
and ( n52755 , n52754 , n31319 );
and ( n52756 , n47449 , n52734 );
or ( n52757 , n52755 , n52756 );
and ( n52758 , n52753 , n52757 );
and ( n52759 , n47449 , n52742 );
or ( n52760 , n52758 , n52759 );
and ( n52761 , n52752 , n52760 );
and ( n52762 , n46519 , n46529 , n48243 , n46549 , C1 );
not ( n52763 , n52762 );
and ( n52764 , n46515 , n46553 , n48246 , n46544 , C1 );
not ( n52765 , n52764 );
and ( n52766 , n52765 , n52760 );
and ( n52767 , n47485 , n52764 );
or ( n52768 , n52766 , n52767 );
and ( n52769 , n52763 , n52768 );
and ( n52770 , n47503 , n52762 );
or ( n52771 , n52769 , n52770 );
and ( n52772 , n52771 , n31452 );
or ( n52773 , n52761 , n52772 );
and ( n52774 , n52773 , n31638 );
and ( n52775 , n31319 , n47277 );
or ( n52776 , C0 , n52741 , n52751 , n52774 , n52775 );
buf ( n52777 , n52776 );
buf ( n52778 , n52777 );
buf ( n52779 , n31655 );
buf ( n52780 , n30987 );
buf ( n52781 , n31655 );
buf ( n52782 , n30987 );
not ( n52783 , n43755 );
and ( n52784 , n52783 , n43292 );
xor ( n52785 , n43762 , n43766 );
and ( n52786 , n52785 , n43755 );
or ( n52787 , n52784 , n52786 );
and ( n52788 , n52787 , n43774 );
not ( n52789 , n44663 );
and ( n52790 , n52789 , n44204 );
xor ( n52791 , n44670 , n44674 );
and ( n52792 , n52791 , n44663 );
or ( n52793 , n52790 , n52792 );
and ( n52794 , n52793 , n44682 );
buf ( n52795 , RI15b45168_222);
and ( n52796 , n52795 , n44695 );
or ( n52797 , n52788 , n52794 , n52796 );
buf ( n52798 , n52797 );
buf ( n52799 , n52798 );
buf ( n52800 , n31655 );
not ( n52801 , n34150 );
and ( n52802 , n52801 , n32871 );
not ( n52803 , n41392 );
and ( n52804 , n52803 , n32871 );
and ( n52805 , n32889 , n41392 );
or ( n52806 , n52804 , n52805 );
and ( n52807 , n52806 , n34150 );
or ( n52808 , n52802 , n52807 );
and ( n52809 , n52808 , n33381 );
not ( n52810 , n41402 );
not ( n52811 , n41392 );
and ( n52812 , n52811 , n32871 );
not ( n52813 , n34287 );
and ( n52814 , n52813 , n34283 );
xor ( n52815 , n34283 , n34193 );
and ( n52816 , n48156 , n48157 );
xor ( n52817 , n52815 , n52816 );
and ( n52818 , n52817 , n34287 );
or ( n52819 , n52814 , n52818 );
and ( n52820 , n52819 , n41392 );
or ( n52821 , n52812 , n52820 );
and ( n52822 , n52810 , n52821 );
and ( n52823 , n52819 , n41402 );
or ( n52824 , n52822 , n52823 );
and ( n52825 , n52824 , n33375 );
not ( n52826 , n32968 );
not ( n52827 , n41402 );
not ( n52828 , n41392 );
and ( n52829 , n52828 , n32871 );
and ( n52830 , n52819 , n41392 );
or ( n52831 , n52829 , n52830 );
and ( n52832 , n52827 , n52831 );
and ( n52833 , n52819 , n41402 );
or ( n52834 , n52832 , n52833 );
and ( n52835 , n52826 , n52834 );
not ( n52836 , n41424 );
not ( n52837 , n41428 );
and ( n52838 , n52837 , n52834 );
not ( n52839 , n34747 );
and ( n52840 , n52839 , n34743 );
xor ( n52841 , n34743 , n34625 );
and ( n52842 , n48182 , n48183 );
xor ( n52843 , n52841 , n52842 );
and ( n52844 , n52843 , n34747 );
or ( n52845 , n52840 , n52844 );
and ( n52846 , n52845 , n41428 );
or ( n52847 , n52838 , n52846 );
and ( n52848 , n52836 , n52847 );
not ( n52849 , n35036 );
and ( n52850 , n52849 , n35032 );
xor ( n52851 , n35032 , n34918 );
and ( n52852 , n48192 , n48193 );
xor ( n52853 , n52851 , n52852 );
and ( n52854 , n52853 , n35036 );
or ( n52855 , n52850 , n52854 );
and ( n52856 , n52855 , n41424 );
or ( n52857 , n52848 , n52856 );
and ( n52858 , n52857 , n32968 );
or ( n52859 , n52835 , n52858 );
and ( n52860 , n52859 , n33370 );
and ( n52861 , n32871 , n35062 );
or ( n52862 , C0 , n52809 , n52825 , n52860 , n52861 );
buf ( n52863 , n52862 );
buf ( n52864 , n52863 );
buf ( n52865 , n31655 );
buf ( n52866 , n30987 );
buf ( n52867 , n30987 );
buf ( n52868 , n30987 );
buf ( n52869 , RI15b542d0_737);
not ( n52870 , n31077 );
and ( n52871 , n52869 , n52870 );
and ( n52872 , n52871 , n31373 );
not ( n52873 , n31402 );
and ( n52874 , n52873 , n52869 );
buf ( n52875 , n31402 );
or ( n52876 , n52874 , n52875 );
and ( n52877 , n52876 , n31408 );
not ( n52878 , n31437 );
and ( n52879 , n52869 , n52878 );
and ( n52880 , n52879 , n31468 );
not ( n52881 , n31497 );
and ( n52882 , n52881 , n52869 );
buf ( n52883 , n31497 );
or ( n52884 , n52882 , n52883 );
and ( n52885 , n52884 , n31521 );
and ( n52886 , n52869 , n31553 );
or ( n52887 , n52872 , n52877 , n52880 , n52885 , n52886 );
and ( n52888 , n52887 , n31557 );
or ( n52889 , n31638 , n31641 );
or ( n52890 , n52889 , n31643 );
or ( n52891 , n52890 , n31645 );
or ( n52892 , n52891 , n31647 );
or ( n52893 , n52892 , n31649 );
or ( n52894 , n52893 , n31007 );
and ( n52895 , n52869 , n52894 );
or ( n52896 , n33973 , n31640 );
buf ( n52897 , n52896 );
or ( n52898 , C0 , n52888 , n52895 , n52897 );
buf ( n52899 , n52898 );
buf ( n52900 , n52899 );
not ( n52901 , n40163 );
and ( n52902 , n52901 , n31873 );
and ( n52903 , n31673 , n42237 , n45160 , n31661 , n42170 );
not ( n52904 , n52903 );
and ( n52905 , n52904 , n31873 );
and ( n52906 , n32218 , n52903 );
or ( n52907 , n52905 , n52906 );
and ( n52908 , n52907 , n40163 );
or ( n52909 , n52902 , n52908 );
and ( n52910 , n52909 , n32498 );
and ( n52911 , n40177 , n42246 , n45169 , n40194 , C1 );
not ( n52912 , n52911 );
not ( n52913 , n52903 );
and ( n52914 , n52913 , n31873 );
and ( n52915 , n42255 , n52903 );
or ( n52916 , n52914 , n52915 );
and ( n52917 , n52912 , n52916 );
and ( n52918 , n42255 , n52911 );
or ( n52919 , n52917 , n52918 );
and ( n52920 , n52919 , n32473 );
not ( n52921 , n32475 );
not ( n52922 , n52911 );
not ( n52923 , n52903 );
and ( n52924 , n52923 , n31873 );
and ( n52925 , n42255 , n52903 );
or ( n52926 , n52924 , n52925 );
and ( n52927 , n52922 , n52926 );
and ( n52928 , n42255 , n52911 );
or ( n52929 , n52927 , n52928 );
and ( n52930 , n52921 , n52929 );
and ( n52931 , n40417 , n42272 , n45195 , n40445 , C1 );
not ( n52932 , n52931 );
and ( n52933 , n40413 , n42275 , n45198 , n40440 , C1 );
not ( n52934 , n52933 );
and ( n52935 , n52934 , n52929 );
and ( n52936 , n42283 , n52933 );
or ( n52937 , n52935 , n52936 );
and ( n52938 , n52932 , n52937 );
and ( n52939 , n42291 , n52931 );
or ( n52940 , n52938 , n52939 );
and ( n52941 , n52940 , n32475 );
or ( n52942 , n52930 , n52941 );
and ( n52943 , n52942 , n32486 );
and ( n52944 , n31873 , n41278 );
or ( n52945 , C0 , n52910 , n52920 , n52943 , n52944 );
buf ( n52946 , n52945 );
buf ( n52947 , n52946 );
buf ( n52948 , n30987 );
buf ( n52949 , n31655 );
buf ( n52950 , n31655 );
buf ( n52951 , n30987 );
not ( n52952 , n43755 );
and ( n52953 , n52952 , n43632 );
xor ( n52954 , n52305 , n52324 );
and ( n52955 , n52954 , n43755 );
or ( n52956 , n52953 , n52955 );
and ( n52957 , n52956 , n43774 );
not ( n52958 , n44663 );
and ( n52959 , n52958 , n44544 );
xor ( n52960 , n52343 , n52362 );
and ( n52961 , n52960 , n44663 );
or ( n52962 , n52959 , n52961 );
and ( n52963 , n52962 , n44682 );
buf ( n52964 , RI15b45ac8_242);
and ( n52965 , n52964 , n44695 );
or ( n52966 , n52957 , n52963 , n52965 );
buf ( n52967 , n52966 );
buf ( n52968 , n52967 );
buf ( n52969 , n30987 );
buf ( n52970 , n31655 );
buf ( n52971 , n31655 );
buf ( n52972 , n30987 );
not ( n52973 , n34150 );
and ( n52974 , n52973 , n32759 );
not ( n52975 , n50731 );
and ( n52976 , n52975 , n32759 );
and ( n52977 , n32789 , n50731 );
or ( n52978 , n52976 , n52977 );
and ( n52979 , n52978 , n34150 );
or ( n52980 , n52974 , n52979 );
and ( n52981 , n52980 , n33381 );
not ( n52982 , n50739 );
not ( n52983 , n50731 );
and ( n52984 , n52983 , n32759 );
and ( n52985 , n34301 , n50731 );
or ( n52986 , n52984 , n52985 );
and ( n52987 , n52982 , n52986 );
and ( n52988 , n34301 , n50739 );
or ( n52989 , n52987 , n52988 );
and ( n52990 , n52989 , n33375 );
not ( n52991 , n32968 );
not ( n52992 , n50739 );
not ( n52993 , n50731 );
and ( n52994 , n52993 , n32759 );
and ( n52995 , n34301 , n50731 );
or ( n52996 , n52994 , n52995 );
and ( n52997 , n52992 , n52996 );
and ( n52998 , n34301 , n50739 );
or ( n52999 , n52997 , n52998 );
and ( n53000 , n52991 , n52999 );
not ( n53001 , n50759 );
not ( n53002 , n50761 );
and ( n53003 , n53002 , n52999 );
and ( n53004 , n34761 , n50761 );
or ( n53005 , n53003 , n53004 );
and ( n53006 , n53001 , n53005 );
and ( n53007 , n35050 , n50759 );
or ( n53008 , n53006 , n53007 );
and ( n53009 , n53008 , n32968 );
or ( n53010 , n53000 , n53009 );
and ( n53011 , n53010 , n33370 );
and ( n53012 , n32759 , n35062 );
or ( n53013 , C0 , n52981 , n52990 , n53011 , n53012 );
buf ( n53014 , n53013 );
buf ( n53015 , n53014 );
buf ( n53016 , n30987 );
buf ( n53017 , n31655 );
buf ( n53018 , n31655 );
and ( n53019 , n31568 , n31007 );
not ( n53020 , n31077 );
and ( n53021 , n53020 , n35394 );
buf ( n53022 , n53021 );
and ( n53023 , n53022 , n31373 );
not ( n53024 , n31402 );
and ( n53025 , n53024 , n35394 );
buf ( n53026 , n53025 );
and ( n53027 , n53026 , n31408 );
not ( n53028 , n31437 );
and ( n53029 , n53028 , n35394 );
not ( n53030 , n31455 );
and ( n53031 , n53030 , n35437 );
xor ( n53032 , n35394 , n35404 );
and ( n53033 , n53032 , n31455 );
or ( n53034 , n53031 , n53033 );
and ( n53035 , n53034 , n31437 );
or ( n53036 , n53029 , n53035 );
and ( n53037 , n53036 , n31468 );
not ( n53038 , n31497 );
and ( n53039 , n53038 , n35394 );
not ( n53040 , n31454 );
not ( n53041 , n31501 );
and ( n53042 , n53041 , n35437 );
xor ( n53043 , n35438 , n35454 );
and ( n53044 , n53043 , n31501 );
or ( n53045 , n53042 , n53044 );
and ( n53046 , n53040 , n53045 );
and ( n53047 , n53032 , n31454 );
or ( n53048 , n53046 , n53047 );
and ( n53049 , n53048 , n31497 );
or ( n53050 , n53039 , n53049 );
and ( n53051 , n53050 , n31521 );
and ( n53052 , n35394 , n31553 );
or ( n53053 , n53023 , n53027 , n53037 , n53051 , n53052 );
and ( n53054 , n53053 , n31557 );
not ( n53055 , n31452 );
not ( n53056 , n31619 );
and ( n53057 , n53056 , n35492 );
xor ( n53058 , n35493 , n35508 );
and ( n53059 , n53058 , n31619 );
or ( n53060 , n53057 , n53059 );
and ( n53061 , n53055 , n53060 );
and ( n53062 , n35394 , n31452 );
or ( n53063 , n53061 , n53062 );
and ( n53064 , n53063 , n31638 );
and ( n53065 , n35394 , n31650 );
or ( n53066 , C0 , n53019 , n53054 , n53064 , C0 , n53065 );
buf ( n53067 , n53066 );
buf ( n53068 , n53067 );
not ( n53069 , n33419 );
and ( n53070 , n53069 , n31576 );
and ( n53071 , n48491 , n33419 );
or ( n53072 , n53070 , n53071 );
and ( n53073 , n53072 , n31529 );
not ( n53074 , n33734 );
and ( n53075 , n53074 , n31576 );
and ( n53076 , n48502 , n33734 );
or ( n53077 , n53075 , n53076 );
and ( n53078 , n53077 , n31527 );
and ( n53079 , n31576 , n33942 );
or ( n53080 , n53073 , n53078 , n53079 );
and ( n53081 , n53080 , n31557 );
and ( n53082 , n34097 , n31643 );
not ( n53083 , n31452 );
and ( n53084 , n53083 , n34097 );
xor ( n53085 , n31576 , n33961 );
and ( n53086 , n53085 , n31452 );
or ( n53087 , n53084 , n53086 );
and ( n53088 , n53087 , n31638 );
and ( n53089 , n34000 , n33973 );
and ( n53090 , n31576 , n33978 );
or ( n53091 , C0 , n53081 , n53082 , n53088 , n53089 , n53090 );
buf ( n53092 , n53091 );
buf ( n53093 , n53092 );
buf ( n53094 , n31655 );
buf ( n53095 , n30987 );
buf ( n53096 , n30987 );
and ( n53097 , n32294 , n50275 );
not ( n53098 , n50278 );
and ( n53099 , n53098 , n31733 );
and ( n53100 , n32294 , n50278 );
or ( n53101 , n53099 , n53100 );
and ( n53102 , n53101 , n32421 );
not ( n53103 , n50002 );
and ( n53104 , n53103 , n31733 );
and ( n53105 , n32294 , n50002 );
or ( n53106 , n53104 , n53105 );
and ( n53107 , n53106 , n32419 );
not ( n53108 , n50289 );
and ( n53109 , n53108 , n31733 );
and ( n53110 , n32294 , n50289 );
or ( n53111 , n53109 , n53110 );
and ( n53112 , n53111 , n32417 );
not ( n53113 , n50008 );
and ( n53114 , n53113 , n31733 );
and ( n53115 , n32294 , n50008 );
or ( n53116 , n53114 , n53115 );
and ( n53117 , n53116 , n32415 );
not ( n53118 , n47331 );
and ( n53119 , n53118 , n31733 );
and ( n53120 , n31749 , n47331 );
or ( n53121 , n53119 , n53120 );
and ( n53122 , n53121 , n32413 );
not ( n53123 , n50067 );
and ( n53124 , n53123 , n31733 );
and ( n53125 , n31749 , n50067 );
or ( n53126 , n53124 , n53125 );
and ( n53127 , n53126 , n32411 );
not ( n53128 , n31728 );
and ( n53129 , n53128 , n31733 );
and ( n53130 , n35649 , n31728 );
or ( n53131 , n53129 , n53130 );
and ( n53132 , n53131 , n32253 );
not ( n53133 , n32283 );
and ( n53134 , n53133 , n31733 );
and ( n53135 , n35662 , n32283 );
or ( n53136 , n53134 , n53135 );
and ( n53137 , n53136 , n32398 );
and ( n53138 , n32340 , n50334 );
or ( n53139 , n53097 , n53102 , n53107 , n53112 , n53117 , n53122 , n53127 , n53132 , n53137 , n53138 );
and ( n53140 , n53139 , n32456 );
and ( n53141 , n35677 , n32489 );
and ( n53142 , n31733 , n50345 );
or ( n53143 , C0 , n53140 , n53141 , n53142 );
buf ( n53144 , n53143 );
buf ( n53145 , n53144 );
buf ( n53146 , n30987 );
not ( n53147 , n31437 );
buf ( n53148 , RI15b527a0_679);
and ( n53149 , n53147 , n53148 );
not ( n53150 , n45766 );
and ( n53151 , n53150 , n45626 );
xor ( n53152 , n45772 , n45784 );
and ( n53153 , n53152 , n45766 );
or ( n53154 , n53151 , n53153 );
and ( n53155 , n53154 , n31437 );
or ( n53156 , n53149 , n53155 );
and ( n53157 , n53156 , n31468 );
not ( n53158 , n44817 );
and ( n53159 , n53158 , n53148 );
not ( n53160 , n44994 );
and ( n53161 , n53160 , n44894 );
xor ( n53162 , n45004 , n45016 );
and ( n53163 , n53162 , n44994 );
or ( n53164 , n53161 , n53163 );
and ( n53165 , n53164 , n44817 );
or ( n53166 , n53159 , n53165 );
and ( n53167 , n53166 , n31521 );
and ( n53168 , n53148 , n42158 );
or ( n53169 , n53157 , n53167 , n53168 );
and ( n53170 , n53169 , n31557 );
and ( n53171 , n53148 , n40154 );
or ( n53172 , C0 , n53170 , n53171 );
buf ( n53173 , n53172 );
buf ( n53174 , n53173 );
buf ( n53175 , n31655 );
buf ( n53176 , n31655 );
buf ( n53177 , n30987 );
not ( n53178 , n34150 );
and ( n53179 , n53178 , n32859 );
not ( n53180 , n50731 );
and ( n53181 , n53180 , n32859 );
and ( n53182 , n32889 , n50731 );
or ( n53183 , n53181 , n53182 );
and ( n53184 , n53183 , n34150 );
or ( n53185 , n53179 , n53184 );
and ( n53186 , n53185 , n33381 );
not ( n53187 , n50739 );
not ( n53188 , n50731 );
and ( n53189 , n53188 , n32859 );
and ( n53190 , n52819 , n50731 );
or ( n53191 , n53189 , n53190 );
and ( n53192 , n53187 , n53191 );
and ( n53193 , n52819 , n50739 );
or ( n53194 , n53192 , n53193 );
and ( n53195 , n53194 , n33375 );
not ( n53196 , n32968 );
not ( n53197 , n50739 );
not ( n53198 , n50731 );
and ( n53199 , n53198 , n32859 );
and ( n53200 , n52819 , n50731 );
or ( n53201 , n53199 , n53200 );
and ( n53202 , n53197 , n53201 );
and ( n53203 , n52819 , n50739 );
or ( n53204 , n53202 , n53203 );
and ( n53205 , n53196 , n53204 );
not ( n53206 , n50759 );
not ( n53207 , n50761 );
and ( n53208 , n53207 , n53204 );
and ( n53209 , n52845 , n50761 );
or ( n53210 , n53208 , n53209 );
and ( n53211 , n53206 , n53210 );
and ( n53212 , n52855 , n50759 );
or ( n53213 , n53211 , n53212 );
and ( n53214 , n53213 , n32968 );
or ( n53215 , n53205 , n53214 );
and ( n53216 , n53215 , n33370 );
and ( n53217 , n32859 , n35062 );
or ( n53218 , C0 , n53186 , n53195 , n53216 , n53217 );
buf ( n53219 , n53218 );
buf ( n53220 , n53219 );
buf ( n53221 , n30987 );
buf ( n53222 , n31655 );
buf ( n53223 , n30987 );
buf ( n53224 , n31655 );
not ( n53225 , n40163 );
and ( n53226 , n53225 , n31902 );
and ( n53227 , n42169 , n42237 , n31665 , n31661 , n42170 );
not ( n53228 , n53227 );
and ( n53229 , n53228 , n31902 );
and ( n53230 , n32200 , n53227 );
or ( n53231 , n53229 , n53230 );
and ( n53232 , n53231 , n40163 );
or ( n53233 , n53226 , n53232 );
and ( n53234 , n53233 , n32498 );
and ( n53235 , n42179 , n42246 , n40188 , n40194 , C1 );
not ( n53236 , n53235 );
not ( n53237 , n53227 );
and ( n53238 , n53237 , n31902 );
not ( n53239 , n40373 );
and ( n53240 , n53239 , n40315 );
xor ( n53241 , n40379 , n40387 );
and ( n53242 , n53241 , n40373 );
or ( n53243 , n53240 , n53242 );
and ( n53244 , n53243 , n53227 );
or ( n53245 , n53238 , n53244 );
and ( n53246 , n53236 , n53245 );
and ( n53247 , n53243 , n53235 );
or ( n53248 , n53246 , n53247 );
and ( n53249 , n53248 , n32473 );
not ( n53250 , n32475 );
not ( n53251 , n53235 );
not ( n53252 , n53227 );
and ( n53253 , n53252 , n31902 );
and ( n53254 , n53243 , n53227 );
or ( n53255 , n53253 , n53254 );
and ( n53256 , n53251 , n53255 );
and ( n53257 , n53243 , n53235 );
or ( n53258 , n53256 , n53257 );
and ( n53259 , n53250 , n53258 );
and ( n53260 , n42205 , n42272 , n40435 , n40445 , C1 );
not ( n53261 , n53260 );
and ( n53262 , n42208 , n42275 , n40430 , n40440 , C1 );
not ( n53263 , n53262 );
and ( n53264 , n53263 , n53258 );
not ( n53265 , n40952 );
and ( n53266 , n53265 , n40897 );
xor ( n53267 , n40958 , n40966 );
and ( n53268 , n53267 , n40952 );
or ( n53269 , n53266 , n53268 );
and ( n53270 , n53269 , n53262 );
or ( n53271 , n53264 , n53270 );
and ( n53272 , n53261 , n53271 );
not ( n53273 , n41247 );
and ( n53274 , n53273 , n41196 );
xor ( n53275 , n41253 , n41261 );
and ( n53276 , n53275 , n41247 );
or ( n53277 , n53274 , n53276 );
and ( n53278 , n53277 , n53260 );
or ( n53279 , n53272 , n53278 );
and ( n53280 , n53279 , n32475 );
or ( n53281 , n53259 , n53280 );
and ( n53282 , n53281 , n32486 );
and ( n53283 , n31902 , n41278 );
or ( n53284 , C0 , n53234 , n53249 , n53282 , n53283 );
buf ( n53285 , n53284 );
buf ( n53286 , n53285 );
buf ( n53287 , RI15b53088_698);
and ( n53288 , n53287 , n31645 );
not ( n53289 , n45274 );
buf ( n53290 , RI15b53808_714);
and ( n53291 , n53289 , n53290 );
not ( n53292 , n41809 );
and ( n53293 , n53292 , n41740 );
xor ( n53294 , n41740 , n41611 );
xor ( n53295 , n41727 , n41611 );
and ( n53296 , n41812 , n41828 );
and ( n53297 , n53295 , n53296 );
xor ( n53298 , n53294 , n53297 );
and ( n53299 , n53298 , n41809 );
or ( n53300 , n53293 , n53299 );
and ( n53301 , n53300 , n45274 );
or ( n53302 , n53291 , n53301 );
and ( n53303 , n53302 , n31373 );
not ( n53304 , n45280 );
and ( n53305 , n53304 , n53290 );
and ( n53306 , n53300 , n45280 );
or ( n53307 , n53305 , n53306 );
and ( n53308 , n53307 , n31468 );
and ( n53309 , n53290 , n45802 );
or ( n53310 , n53303 , n53308 , n53309 );
and ( n53311 , n53310 , n31557 );
and ( n53312 , n53290 , n45808 );
or ( n53313 , C0 , n53288 , n53311 , n53312 );
buf ( n53314 , n53313 );
buf ( n53315 , n53314 );
buf ( n53316 , RI15b5ee60_1103);
and ( n53317 , n53316 , n32494 );
not ( n53318 , n46083 );
buf ( n53319 , RI15b60468_1150);
and ( n53320 , n53318 , n53319 );
buf ( n53321 , n53320 );
and ( n53322 , n53321 , n32421 );
not ( n53323 , n46326 );
and ( n53324 , n53323 , n53319 );
not ( n53325 , n51396 );
and ( n53326 , n53325 , n51341 );
xor ( n53327 , n51341 , n51155 );
xor ( n53328 , n51324 , n51155 );
xor ( n53329 , n51307 , n51155 );
xor ( n53330 , n51290 , n51155 );
xor ( n53331 , n51273 , n51155 );
and ( n53332 , n51399 , n51411 );
and ( n53333 , n53331 , n53332 );
and ( n53334 , n53330 , n53333 );
and ( n53335 , n53329 , n53334 );
and ( n53336 , n53328 , n53335 );
xor ( n53337 , n53327 , n53336 );
and ( n53338 , n53337 , n51396 );
or ( n53339 , n53326 , n53338 );
and ( n53340 , n53339 , n46326 );
or ( n53341 , n53324 , n53340 );
and ( n53342 , n53341 , n32417 );
and ( n53343 , n53319 , n46340 );
or ( n53344 , n53322 , n53342 , n53343 );
and ( n53345 , n53344 , n32456 );
and ( n53346 , n53319 , n46349 );
or ( n53347 , C0 , n53317 , n53345 , n53346 );
buf ( n53348 , n53347 );
buf ( n53349 , n53348 );
buf ( n53350 , n31655 );
not ( n53351 , n46356 );
and ( n53352 , n53351 , n31216 );
and ( n53353 , n46359 , n31021 , n48213 , n31013 , n46361 );
not ( n53354 , n53353 );
and ( n53355 , n53354 , n31216 );
and ( n53356 , n31238 , n53353 );
or ( n53357 , n53355 , n53356 );
and ( n53358 , n53357 , n46356 );
or ( n53359 , n53352 , n53358 );
and ( n53360 , n53359 , n31649 );
and ( n53361 , n46374 , n46379 , n48222 , n46392 , C1 );
not ( n53362 , n53361 );
not ( n53363 , n53353 );
and ( n53364 , n53363 , n31216 );
and ( n53365 , n49901 , n53353 );
or ( n53366 , n53364 , n53365 );
and ( n53367 , n53362 , n53366 );
and ( n53368 , n49901 , n53361 );
or ( n53369 , n53367 , n53368 );
and ( n53370 , n53369 , n31643 );
not ( n53371 , n31452 );
not ( n53372 , n53361 );
not ( n53373 , n53353 );
and ( n53374 , n53373 , n31216 );
and ( n53375 , n49901 , n53353 );
or ( n53376 , n53374 , n53375 );
and ( n53377 , n53372 , n53376 );
and ( n53378 , n49901 , n53361 );
or ( n53379 , n53377 , n53378 );
and ( n53380 , n53371 , n53379 );
and ( n53381 , n46520 , n46528 , n48243 , n46549 , C1 );
not ( n53382 , n53381 );
and ( n53383 , n46552 , n46524 , n48246 , n46544 , C1 );
not ( n53384 , n53383 );
and ( n53385 , n53384 , n53379 );
and ( n53386 , n49925 , n53383 );
or ( n53387 , n53385 , n53386 );
and ( n53388 , n53382 , n53387 );
and ( n53389 , n49933 , n53381 );
or ( n53390 , n53388 , n53389 );
and ( n53391 , n53390 , n31452 );
or ( n53392 , n53380 , n53391 );
and ( n53393 , n53392 , n31638 );
and ( n53394 , n31216 , n47277 );
or ( n53395 , C0 , n53360 , n53370 , n53393 , n53394 );
buf ( n53396 , n53395 );
buf ( n53397 , n53396 );
buf ( n53398 , n30987 );
buf ( n53399 , n31655 );
and ( n53400 , n42406 , n48455 );
not ( n53401 , n48457 );
and ( n53402 , n53401 , n42379 );
and ( n53403 , n42406 , n48457 );
or ( n53404 , n53402 , n53403 );
and ( n53405 , n53404 , n31373 );
not ( n53406 , n44807 );
and ( n53407 , n53406 , n42379 );
and ( n53408 , n42406 , n44807 );
or ( n53409 , n53407 , n53408 );
and ( n53410 , n53409 , n31408 );
not ( n53411 , n48468 );
and ( n53412 , n53411 , n42379 );
and ( n53413 , n42406 , n48468 );
or ( n53414 , n53412 , n53413 );
and ( n53415 , n53414 , n31468 );
not ( n53416 , n44817 );
and ( n53417 , n53416 , n42379 );
and ( n53418 , n42406 , n44817 );
or ( n53419 , n53417 , n53418 );
and ( n53420 , n53419 , n31521 );
not ( n53421 , n39979 );
and ( n53422 , n53421 , n42379 );
and ( n53423 , n42387 , n39979 );
or ( n53424 , n53422 , n53423 );
and ( n53425 , n53424 , n31538 );
not ( n53426 , n45059 );
and ( n53427 , n53426 , n42379 );
and ( n53428 , n42387 , n45059 );
or ( n53429 , n53427 , n53428 );
and ( n53430 , n53429 , n31536 );
not ( n53431 , n33419 );
and ( n53432 , n53431 , n42379 );
xor ( n53433 , n42387 , n42388 );
and ( n53434 , n53433 , n33419 );
or ( n53435 , n53432 , n53434 );
and ( n53436 , n53435 , n31529 );
not ( n53437 , n33734 );
and ( n53438 , n53437 , n42379 );
not ( n53439 , n33533 );
xor ( n53440 , n42406 , n42407 );
and ( n53441 , n53439 , n53440 );
xnor ( n53442 , n42420 , n42421 );
and ( n53443 , n53442 , n33533 );
or ( n53444 , n53441 , n53443 );
and ( n53445 , n53444 , n33734 );
or ( n53446 , n53438 , n53445 );
and ( n53447 , n53446 , n31527 );
and ( n53448 , n42420 , n48513 );
or ( n53449 , n53400 , n53405 , n53410 , n53415 , n53420 , n53425 , n53430 , n53436 , n53447 , n53448 );
and ( n53450 , n53449 , n31557 );
and ( n53451 , n35395 , n33973 );
and ( n53452 , n42379 , n48524 );
or ( n53453 , C0 , n53450 , n53451 , n53452 );
buf ( n53454 , n53453 );
buf ( n53455 , n53454 );
buf ( n53456 , n30987 );
buf ( n53457 , n31655 );
not ( n53458 , n38443 );
and ( n53459 , n53458 , n38371 );
xor ( n53460 , n38371 , n37947 );
xor ( n53461 , n38354 , n37947 );
xor ( n53462 , n38337 , n37947 );
xor ( n53463 , n38320 , n37947 );
xor ( n53464 , n38303 , n37947 );
xor ( n53465 , n38286 , n37947 );
xor ( n53466 , n38269 , n37947 );
xor ( n53467 , n38252 , n37947 );
xor ( n53468 , n38235 , n37947 );
xor ( n53469 , n38218 , n37947 );
xor ( n53470 , n38201 , n37947 );
xor ( n53471 , n38184 , n37947 );
xor ( n53472 , n38167 , n37947 );
xor ( n53473 , n38150 , n37947 );
xor ( n53474 , n38133 , n37947 );
xor ( n53475 , n38116 , n37947 );
xor ( n53476 , n38099 , n37947 );
xor ( n53477 , n38082 , n37947 );
xor ( n53478 , n38065 , n37947 );
xor ( n53479 , n38048 , n37947 );
xor ( n53480 , n38031 , n37947 );
xor ( n53481 , n38014 , n37947 );
xor ( n53482 , n37997 , n37947 );
xor ( n53483 , n37980 , n37947 );
xor ( n53484 , n37963 , n37947 );
and ( n53485 , n38446 , n37947 );
and ( n53486 , n53484 , n53485 );
and ( n53487 , n53483 , n53486 );
and ( n53488 , n53482 , n53487 );
and ( n53489 , n53481 , n53488 );
and ( n53490 , n53480 , n53489 );
and ( n53491 , n53479 , n53490 );
and ( n53492 , n53478 , n53491 );
and ( n53493 , n53477 , n53492 );
and ( n53494 , n53476 , n53493 );
and ( n53495 , n53475 , n53494 );
and ( n53496 , n53474 , n53495 );
and ( n53497 , n53473 , n53496 );
and ( n53498 , n53472 , n53497 );
and ( n53499 , n53471 , n53498 );
and ( n53500 , n53470 , n53499 );
and ( n53501 , n53469 , n53500 );
and ( n53502 , n53468 , n53501 );
and ( n53503 , n53467 , n53502 );
and ( n53504 , n53466 , n53503 );
and ( n53505 , n53465 , n53504 );
and ( n53506 , n53464 , n53505 );
and ( n53507 , n53463 , n53506 );
and ( n53508 , n53462 , n53507 );
and ( n53509 , n53461 , n53508 );
xor ( n53510 , n53460 , n53509 );
and ( n53511 , n53510 , n38443 );
or ( n53512 , n53459 , n53511 );
and ( n53513 , n53512 , n38450 );
not ( n53514 , n39339 );
and ( n53515 , n53514 , n39271 );
xor ( n53516 , n39271 , n38847 );
xor ( n53517 , n39254 , n38847 );
xor ( n53518 , n39237 , n38847 );
xor ( n53519 , n39220 , n38847 );
xor ( n53520 , n39203 , n38847 );
xor ( n53521 , n39186 , n38847 );
xor ( n53522 , n39169 , n38847 );
xor ( n53523 , n39152 , n38847 );
xor ( n53524 , n39135 , n38847 );
xor ( n53525 , n39118 , n38847 );
xor ( n53526 , n39101 , n38847 );
xor ( n53527 , n39084 , n38847 );
xor ( n53528 , n39067 , n38847 );
xor ( n53529 , n39050 , n38847 );
xor ( n53530 , n39033 , n38847 );
xor ( n53531 , n39016 , n38847 );
xor ( n53532 , n38999 , n38847 );
xor ( n53533 , n38982 , n38847 );
xor ( n53534 , n38965 , n38847 );
xor ( n53535 , n38948 , n38847 );
xor ( n53536 , n38931 , n38847 );
xor ( n53537 , n38914 , n38847 );
xor ( n53538 , n38897 , n38847 );
xor ( n53539 , n38880 , n38847 );
xor ( n53540 , n38863 , n38847 );
and ( n53541 , n39342 , n38847 );
and ( n53542 , n53540 , n53541 );
and ( n53543 , n53539 , n53542 );
and ( n53544 , n53538 , n53543 );
and ( n53545 , n53537 , n53544 );
and ( n53546 , n53536 , n53545 );
and ( n53547 , n53535 , n53546 );
and ( n53548 , n53534 , n53547 );
and ( n53549 , n53533 , n53548 );
and ( n53550 , n53532 , n53549 );
and ( n53551 , n53531 , n53550 );
and ( n53552 , n53530 , n53551 );
and ( n53553 , n53529 , n53552 );
and ( n53554 , n53528 , n53553 );
and ( n53555 , n53527 , n53554 );
and ( n53556 , n53526 , n53555 );
and ( n53557 , n53525 , n53556 );
and ( n53558 , n53524 , n53557 );
and ( n53559 , n53523 , n53558 );
and ( n53560 , n53522 , n53559 );
and ( n53561 , n53521 , n53560 );
and ( n53562 , n53520 , n53561 );
and ( n53563 , n53519 , n53562 );
and ( n53564 , n53518 , n53563 );
and ( n53565 , n53517 , n53564 );
xor ( n53566 , n53516 , n53565 );
and ( n53567 , n53566 , n39339 );
or ( n53568 , n53515 , n53567 );
and ( n53569 , n53568 , n39346 );
and ( n53570 , n40224 , n39359 );
or ( n53571 , n53513 , n53569 , n53570 );
buf ( n53572 , n53571 );
buf ( n53573 , n53572 );
buf ( n53574 , n30987 );
and ( n53575 , n31585 , n31007 );
not ( n53576 , n31077 );
and ( n53577 , n53576 , n34009 );
buf ( n53578 , n53577 );
and ( n53579 , n53578 , n31373 );
not ( n53580 , n31402 );
and ( n53581 , n53580 , n34009 );
buf ( n53582 , n53581 );
and ( n53583 , n53582 , n31408 );
not ( n53584 , n31437 );
and ( n53585 , n53584 , n34009 );
not ( n53586 , n31455 );
and ( n53587 , n53586 , n34058 );
xor ( n53588 , n34009 , n34014 );
and ( n53589 , n53588 , n31455 );
or ( n53590 , n53587 , n53589 );
and ( n53591 , n53590 , n31437 );
or ( n53592 , n53585 , n53591 );
and ( n53593 , n53592 , n31468 );
not ( n53594 , n31497 );
and ( n53595 , n53594 , n34009 );
not ( n53596 , n31454 );
not ( n53597 , n31501 );
and ( n53598 , n53597 , n34058 );
xor ( n53599 , n34059 , n34066 );
and ( n53600 , n53599 , n31501 );
or ( n53601 , n53598 , n53600 );
and ( n53602 , n53596 , n53601 );
and ( n53603 , n53588 , n31454 );
or ( n53604 , n53602 , n53603 );
and ( n53605 , n53604 , n31497 );
or ( n53606 , n53595 , n53605 );
and ( n53607 , n53606 , n31521 );
and ( n53608 , n34009 , n31553 );
or ( n53609 , n53579 , n53583 , n53593 , n53607 , n53608 );
and ( n53610 , n53609 , n31557 );
not ( n53611 , n31452 );
not ( n53612 , n31619 );
and ( n53613 , n53612 , n34115 );
xor ( n53614 , n34116 , n34123 );
and ( n53615 , n53614 , n31619 );
or ( n53616 , n53613 , n53615 );
and ( n53617 , n53611 , n53616 );
and ( n53618 , n34009 , n31452 );
or ( n53619 , n53617 , n53618 );
and ( n53620 , n53619 , n31638 );
buf ( n53621 , n33973 );
and ( n53622 , n34009 , n31650 );
or ( n53623 , C0 , n53575 , n53610 , n53620 , n53621 , n53622 );
buf ( n53624 , n53623 );
buf ( n53625 , n53624 );
buf ( n53626 , n31655 );
buf ( n53627 , n31655 );
and ( n53628 , n31628 , n31007 );
not ( n53629 , n31077 );
and ( n53630 , n53629 , n35687 );
and ( n53631 , n33479 , n31077 );
or ( n53632 , n53630 , n53631 );
and ( n53633 , n53632 , n31373 );
not ( n53634 , n31402 );
and ( n53635 , n53634 , n35687 );
and ( n53636 , n33479 , n31402 );
or ( n53637 , n53635 , n53636 );
and ( n53638 , n53637 , n31408 );
not ( n53639 , n31437 );
and ( n53640 , n53639 , n35687 );
not ( n53641 , n31455 );
and ( n53642 , n53641 , n31509 );
and ( n53643 , n35687 , n31455 );
or ( n53644 , n53642 , n53643 );
and ( n53645 , n53644 , n31437 );
or ( n53646 , n53640 , n53645 );
and ( n53647 , n53646 , n31468 );
not ( n53648 , n31497 );
and ( n53649 , n53648 , n35687 );
not ( n53650 , n31454 );
buf ( n53651 , n31509 );
and ( n53652 , n53650 , n53651 );
and ( n53653 , n35687 , n31454 );
or ( n53654 , n53652 , n53653 );
and ( n53655 , n53654 , n31497 );
or ( n53656 , n53649 , n53655 );
and ( n53657 , n53656 , n31521 );
and ( n53658 , n35687 , n31553 );
or ( n53659 , n53633 , n53638 , n53647 , n53657 , n53658 );
and ( n53660 , n53659 , n31557 );
not ( n53661 , n31452 );
buf ( n53662 , n31628 );
and ( n53663 , n53661 , n53662 );
and ( n53664 , n35687 , n31452 );
or ( n53665 , n53663 , n53664 );
and ( n53666 , n53665 , n31638 );
and ( n53667 , n35687 , n31650 );
or ( n53668 , C0 , n53628 , n53660 , n53666 , C0 , n53667 );
buf ( n53669 , n53668 );
buf ( n53670 , n53669 );
buf ( n53671 , n30987 );
buf ( n53672 , n30987 );
buf ( n53673 , n30987 );
not ( n53674 , n40163 );
and ( n53675 , n53674 , n32013 );
not ( n53676 , n52903 );
and ( n53677 , n53676 , n32013 );
and ( n53678 , n32147 , n52903 );
or ( n53679 , n53677 , n53678 );
and ( n53680 , n53679 , n40163 );
or ( n53681 , n53675 , n53680 );
and ( n53682 , n53681 , n32498 );
not ( n53683 , n52911 );
not ( n53684 , n52903 );
and ( n53685 , n53684 , n32013 );
and ( n53686 , n49314 , n52903 );
or ( n53687 , n53685 , n53686 );
and ( n53688 , n53683 , n53687 );
and ( n53689 , n49314 , n52911 );
or ( n53690 , n53688 , n53689 );
and ( n53691 , n53690 , n32473 );
not ( n53692 , n32475 );
not ( n53693 , n52911 );
not ( n53694 , n52903 );
and ( n53695 , n53694 , n32013 );
and ( n53696 , n49314 , n52903 );
or ( n53697 , n53695 , n53696 );
and ( n53698 , n53693 , n53697 );
and ( n53699 , n49314 , n52911 );
or ( n53700 , n53698 , n53699 );
and ( n53701 , n53692 , n53700 );
not ( n53702 , n52931 );
not ( n53703 , n52933 );
and ( n53704 , n53703 , n53700 );
and ( n53705 , n49340 , n52933 );
or ( n53706 , n53704 , n53705 );
and ( n53707 , n53702 , n53706 );
and ( n53708 , n49348 , n52931 );
or ( n53709 , n53707 , n53708 );
and ( n53710 , n53709 , n32475 );
or ( n53711 , n53701 , n53710 );
and ( n53712 , n53711 , n32486 );
and ( n53713 , n32013 , n41278 );
or ( n53714 , C0 , n53682 , n53691 , n53712 , n53713 );
buf ( n53715 , n53714 );
buf ( n53716 , n53715 );
buf ( n53717 , n31655 );
buf ( n53718 , n35687 );
not ( n53719 , n53718 );
buf ( n53720 , n53719 );
not ( n53721 , n53720 );
not ( n53722 , n35375 );
and ( n53723 , n53722 , n31460 );
not ( n53724 , n31460 );
not ( n53725 , n35687 );
xor ( n53726 , n53724 , n53725 );
and ( n53727 , n53726 , n35375 );
or ( n53728 , n53723 , n53727 );
not ( n53729 , n53728 );
buf ( n53730 , n53729 );
buf ( n53731 , n53730 );
not ( n53732 , n53731 );
or ( n53733 , n53721 , n53732 );
buf ( n53734 , n53733 );
buf ( n53735 , n53734 );
and ( n53736 , n53735 , n35375 );
not ( n53737 , n53736 );
and ( n53738 , n53737 , n53721 );
xor ( n53739 , n53721 , n35375 );
xor ( n53740 , n53739 , n35375 );
and ( n53741 , n53740 , n53736 );
or ( n53742 , n53738 , n53741 );
not ( n53743 , n53742 );
not ( n53744 , n53736 );
and ( n53745 , n53744 , n53732 );
xor ( n53746 , n53732 , n35375 );
and ( n53747 , n53739 , n35375 );
xor ( n53748 , n53746 , n53747 );
and ( n53749 , n53748 , n53736 );
or ( n53750 , n53745 , n53749 );
not ( n53751 , n53750 );
and ( n53752 , n53746 , n53747 );
buf ( n53753 , n53752 );
and ( n53754 , n53753 , n53736 );
buf ( n53755 , n53754 );
nor ( n53756 , n53743 , n53751 , n53755 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n53757 , n53756 );
nor ( n53758 , n53742 , n53751 , n53755 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n53759 , n53758 );
or ( n53760 , n53757 , n53759 , C0 , C0 );
buf ( n53761 , RI15b54618_744);
not ( n53762 , n31452 );
buf ( n53763 , RI15b54708_746);
buf ( n53764 , n53763 );
buf ( n53765 , n53763 );
buf ( n53766 , n53763 );
buf ( n53767 , n53763 );
buf ( n53768 , n53763 );
buf ( n53769 , n53763 );
buf ( n53770 , n53763 );
buf ( n53771 , n53763 );
buf ( n53772 , n53763 );
buf ( n53773 , n53763 );
buf ( n53774 , n53763 );
buf ( n53775 , n53763 );
buf ( n53776 , n53763 );
buf ( n53777 , n53763 );
buf ( n53778 , n53763 );
buf ( n53779 , n53763 );
buf ( n53780 , n53763 );
buf ( n53781 , n53763 );
buf ( n53782 , n53763 );
buf ( n53783 , n53763 );
buf ( n53784 , n53763 );
buf ( n53785 , n53763 );
buf ( n53786 , n53763 );
buf ( n53787 , n53763 );
buf ( n53788 , n53763 );
buf ( n53789 , n53763 );
buf ( n53790 , n53763 );
buf ( n53791 , n53763 );
buf ( n53792 , n53763 );
nor ( n53793 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 );
and ( n53794 , n53760 , n53793 );
buf ( n53795 , n53756 );
buf ( n53796 , n53758 );
or ( n53797 , C0 , n53795 , n53796 , C0 , C0 );
not ( n53798 , n53761 );
buf ( n53799 , n53763 );
buf ( n53800 , n53763 );
buf ( n53801 , n53763 );
buf ( n53802 , n53763 );
buf ( n53803 , n53763 );
buf ( n53804 , n53763 );
buf ( n53805 , n53763 );
buf ( n53806 , n53763 );
buf ( n53807 , n53763 );
buf ( n53808 , n53763 );
buf ( n53809 , n53763 );
buf ( n53810 , n53763 );
buf ( n53811 , n53763 );
buf ( n53812 , n53763 );
buf ( n53813 , n53763 );
buf ( n53814 , n53763 );
buf ( n53815 , n53763 );
buf ( n53816 , n53763 );
buf ( n53817 , n53763 );
buf ( n53818 , n53763 );
buf ( n53819 , n53763 );
buf ( n53820 , n53763 );
buf ( n53821 , n53763 );
buf ( n53822 , n53763 );
buf ( n53823 , n53763 );
buf ( n53824 , n53763 );
buf ( n53825 , n53763 );
buf ( n53826 , n53763 );
buf ( n53827 , n53763 );
nor ( n53828 , n53798 , n31452 , n53763 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 );
and ( n53829 , n53797 , n53828 );
buf ( n53830 , n53756 );
buf ( n53831 , n53758 );
nor ( n53832 , n53742 , n53750 , n53755 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n53833 , n53832 );
or ( n53834 , C0 , n53830 , n53831 , C0 , n53833 );
buf ( n53835 , n53763 );
buf ( n53836 , n53763 );
buf ( n53837 , n53763 );
buf ( n53838 , n53763 );
buf ( n53839 , n53763 );
buf ( n53840 , n53763 );
buf ( n53841 , n53763 );
buf ( n53842 , n53763 );
buf ( n53843 , n53763 );
buf ( n53844 , n53763 );
buf ( n53845 , n53763 );
buf ( n53846 , n53763 );
buf ( n53847 , n53763 );
buf ( n53848 , n53763 );
buf ( n53849 , n53763 );
buf ( n53850 , n53763 );
buf ( n53851 , n53763 );
buf ( n53852 , n53763 );
buf ( n53853 , n53763 );
buf ( n53854 , n53763 );
buf ( n53855 , n53763 );
buf ( n53856 , n53763 );
buf ( n53857 , n53763 );
buf ( n53858 , n53763 );
buf ( n53859 , n53763 );
buf ( n53860 , n53763 );
buf ( n53861 , n53763 );
buf ( n53862 , n53763 );
buf ( n53863 , n53763 );
nor ( n53864 , n53761 , n31452 , n53763 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 );
and ( n53865 , n53834 , n53864 );
or ( n53866 , C0 , n53794 , n53829 , n53865 );
buf ( n53867 , n53866 );
buf ( n53868 , n53867 );
buf ( n53869 , n30987 );
buf ( n53870 , RI15b46fe0_287);
buf ( n53871 , n53870 );
buf ( n53872 , n30987 );
buf ( n53873 , n31655 );
not ( n53874 , n48765 );
and ( n53875 , n53874 , n33222 );
xor ( n53876 , n48777 , n49011 );
and ( n53877 , n53876 , n48765 );
or ( n53878 , n53875 , n53877 );
and ( n53879 , n53878 , n33180 );
not ( n53880 , n49054 );
and ( n53881 , n53880 , n33222 );
not ( n53882 , n48845 );
xor ( n53883 , n49067 , n49125 );
and ( n53884 , n53882 , n53883 );
xnor ( n53885 , n49176 , n49251 );
and ( n53886 , n53885 , n48845 );
or ( n53887 , n53884 , n53886 );
and ( n53888 , n53887 , n49054 );
or ( n53889 , n53881 , n53888 );
and ( n53890 , n53889 , n33178 );
and ( n53891 , n33222 , n49774 );
or ( n53892 , n53879 , n53890 , n53891 );
and ( n53893 , n53892 , n33208 );
and ( n53894 , n33295 , n33375 );
not ( n53895 , n32968 );
and ( n53896 , n53895 , n33295 );
and ( n53897 , n33233 , n49785 );
and ( n53898 , n33232 , n53897 );
and ( n53899 , n33231 , n53898 );
and ( n53900 , n33230 , n53899 );
and ( n53901 , n33229 , n53900 );
and ( n53902 , n33228 , n53901 );
and ( n53903 , n33227 , n53902 );
and ( n53904 , n33226 , n53903 );
and ( n53905 , n33225 , n53904 );
and ( n53906 , n33224 , n53905 );
and ( n53907 , n33223 , n53906 );
xor ( n53908 , n33222 , n53907 );
and ( n53909 , n53908 , n32968 );
or ( n53910 , n53896 , n53909 );
and ( n53911 , n53910 , n33370 );
and ( n53912 , n32985 , n35056 );
and ( n53913 , n33222 , n49794 );
or ( n53914 , C0 , n53893 , n53894 , n53911 , n53912 , n53913 );
buf ( n53915 , n53914 );
buf ( n53916 , n53915 );
buf ( n53917 , n31655 );
and ( n53918 , n46028 , n32500 );
not ( n53919 , n35211 );
and ( n53920 , n53919 , n37553 );
buf ( n53921 , n53920 );
and ( n53922 , n53921 , n32421 );
not ( n53923 , n35245 );
and ( n53924 , n53923 , n37553 );
buf ( n53925 , n53924 );
and ( n53926 , n53925 , n32419 );
not ( n53927 , n35278 );
and ( n53928 , n53927 , n37553 );
not ( n53929 , n35295 );
and ( n53930 , n53929 , n49583 );
xor ( n53931 , n37553 , n49539 );
and ( n53932 , n53931 , n35295 );
or ( n53933 , n53930 , n53932 );
and ( n53934 , n53933 , n35278 );
or ( n53935 , n53928 , n53934 );
and ( n53936 , n53935 , n32417 );
not ( n53937 , n35331 );
and ( n53938 , n53937 , n37553 );
not ( n53939 , n35294 );
not ( n53940 , n45995 );
and ( n53941 , n53940 , n49583 );
xor ( n53942 , n49584 , n49625 );
and ( n53943 , n53942 , n45995 );
or ( n53944 , n53941 , n53943 );
and ( n53945 , n53939 , n53944 );
and ( n53946 , n53931 , n35294 );
or ( n53947 , n53945 , n53946 );
and ( n53948 , n53947 , n35331 );
or ( n53949 , n53938 , n53948 );
and ( n53950 , n53949 , n32415 );
and ( n53951 , n37553 , n35354 );
or ( n53952 , n53922 , n53926 , n53936 , n53950 , n53951 );
and ( n53953 , n53952 , n32456 );
not ( n53954 , n32475 );
not ( n53955 , n46060 );
and ( n53956 , n53955 , n49673 );
xor ( n53957 , n49674 , n49719 );
and ( n53958 , n53957 , n46060 );
or ( n53959 , n53956 , n53958 );
and ( n53960 , n53954 , n53959 );
and ( n53961 , n37553 , n32475 );
or ( n53962 , n53960 , n53961 );
and ( n53963 , n53962 , n32486 );
buf ( n53964 , n32489 );
and ( n53965 , n37553 , n35367 );
or ( n53966 , C0 , n53918 , n53953 , n53963 , n53964 , n53965 );
buf ( n53967 , n53966 );
buf ( n53968 , n53967 );
buf ( n53969 , n31655 );
not ( n53970 , n36587 );
and ( n53971 , n53970 , n36175 );
xor ( n53972 , n50190 , n50197 );
and ( n53973 , n53972 , n36587 );
or ( n53974 , n53971 , n53973 );
and ( n53975 , n53974 , n36596 );
not ( n53976 , n37485 );
and ( n53977 , n53976 , n37077 );
xor ( n53978 , n50240 , n50247 );
and ( n53979 , n53978 , n37485 );
or ( n53980 , n53977 , n53979 );
and ( n53981 , n53980 , n37494 );
and ( n53982 , n41844 , n37506 );
or ( n53983 , n53975 , n53981 , n53982 );
buf ( n53984 , n53983 );
buf ( n53985 , n53984 );
buf ( n53986 , n30987 );
buf ( n53987 , RI15b60918_1160);
and ( n53988 , n53987 , n48531 );
and ( n53989 , n50823 , n39359 );
or ( n53990 , n53988 , n53989 );
buf ( n53991 , n53990 );
buf ( n53992 , n53991 );
buf ( n53993 , n30987 );
xor ( n53994 , n41639 , n44778 );
and ( n53995 , n53994 , n31548 );
not ( n53996 , n44807 );
and ( n53997 , n53996 , n41639 );
and ( n53998 , n41918 , n44807 );
or ( n53999 , n53997 , n53998 );
and ( n54000 , n53999 , n31408 );
not ( n54001 , n44817 );
and ( n54002 , n54001 , n41639 );
not ( n54003 , n41835 );
buf ( n54004 , RI15b52d40_691);
and ( n54005 , n54003 , n54004 );
not ( n54006 , n42124 );
and ( n54007 , n54006 , n41928 );
xor ( n54008 , n42132 , n42138 );
and ( n54009 , n54008 , n42124 );
or ( n54010 , n54007 , n54009 );
and ( n54011 , n54010 , n41835 );
or ( n54012 , n54005 , n54011 );
and ( n54013 , n54012 , n44817 );
or ( n54014 , n54002 , n54013 );
and ( n54015 , n54014 , n31521 );
not ( n54016 , n45059 );
and ( n54017 , n54016 , n41639 );
and ( n54018 , n33609 , n45059 );
or ( n54019 , n54017 , n54018 );
and ( n54020 , n54019 , n31536 );
and ( n54021 , n41639 , n45148 );
or ( n54022 , n53995 , n54000 , n54015 , n54020 , n54021 );
and ( n54023 , n54022 , n31557 );
and ( n54024 , n41639 , n40154 );
or ( n54025 , C0 , n54023 , n54024 );
buf ( n54026 , n54025 );
buf ( n54027 , n54026 );
buf ( n54028 , n31655 );
not ( n54029 , n40163 );
and ( n54030 , n54029 , n31877 );
not ( n54031 , n50540 );
and ( n54032 , n54031 , n31877 );
and ( n54033 , n32218 , n50540 );
or ( n54034 , n54032 , n54033 );
and ( n54035 , n54034 , n40163 );
or ( n54036 , n54030 , n54035 );
and ( n54037 , n54036 , n32498 );
not ( n54038 , n50548 );
not ( n54039 , n50540 );
and ( n54040 , n54039 , n31877 );
and ( n54041 , n42255 , n50540 );
or ( n54042 , n54040 , n54041 );
and ( n54043 , n54038 , n54042 );
and ( n54044 , n42255 , n50548 );
or ( n54045 , n54043 , n54044 );
and ( n54046 , n54045 , n32473 );
not ( n54047 , n32475 );
not ( n54048 , n50548 );
not ( n54049 , n50540 );
and ( n54050 , n54049 , n31877 );
and ( n54051 , n42255 , n50540 );
or ( n54052 , n54050 , n54051 );
and ( n54053 , n54048 , n54052 );
and ( n54054 , n42255 , n50548 );
or ( n54055 , n54053 , n54054 );
and ( n54056 , n54047 , n54055 );
not ( n54057 , n50568 );
not ( n54058 , n50570 );
and ( n54059 , n54058 , n54055 );
and ( n54060 , n42283 , n50570 );
or ( n54061 , n54059 , n54060 );
and ( n54062 , n54057 , n54061 );
and ( n54063 , n42291 , n50568 );
or ( n54064 , n54062 , n54063 );
and ( n54065 , n54064 , n32475 );
or ( n54066 , n54056 , n54065 );
and ( n54067 , n54066 , n32486 );
and ( n54068 , n31877 , n41278 );
or ( n54069 , C0 , n54037 , n54046 , n54067 , n54068 );
buf ( n54070 , n54069 );
buf ( n54071 , n54070 );
buf ( n54072 , n30987 );
buf ( n54073 , n30987 );
buf ( n54074 , n31655 );
buf ( n54075 , RI15b460e0_255);
and ( n54076 , n54075 , n33377 );
not ( n54077 , n48545 );
buf ( n54078 , RI15b476e8_302);
and ( n54079 , n54077 , n54078 );
buf ( n54080 , n54079 );
and ( n54081 , n54080 , n32890 );
not ( n54082 , n48557 );
and ( n54083 , n54082 , n54078 );
not ( n54084 , n39374 );
buf ( n54085 , RI15b48c00_347);
and ( n54086 , n54084 , n54085 );
not ( n54087 , n54085 );
not ( n54088 , n39558 );
not ( n54089 , n39545 );
not ( n54090 , n39532 );
not ( n54091 , n39519 );
not ( n54092 , n39506 );
not ( n54093 , n39493 );
not ( n54094 , n39480 );
not ( n54095 , n39467 );
not ( n54096 , n39454 );
not ( n54097 , n39441 );
not ( n54098 , n39428 );
not ( n54099 , n39415 );
not ( n54100 , n39402 );
not ( n54101 , n39389 );
not ( n54102 , n39376 );
not ( n54103 , n39369 );
and ( n54104 , n54102 , n54103 );
and ( n54105 , n54101 , n54104 );
and ( n54106 , n54100 , n54105 );
and ( n54107 , n54099 , n54106 );
and ( n54108 , n54098 , n54107 );
and ( n54109 , n54097 , n54108 );
and ( n54110 , n54096 , n54109 );
and ( n54111 , n54095 , n54110 );
and ( n54112 , n54094 , n54111 );
and ( n54113 , n54093 , n54112 );
and ( n54114 , n54092 , n54113 );
and ( n54115 , n54091 , n54114 );
and ( n54116 , n54090 , n54115 );
and ( n54117 , n54089 , n54116 );
and ( n54118 , n54088 , n54117 );
xor ( n54119 , n54087 , n54118 );
and ( n54120 , n54119 , n39374 );
or ( n54121 , n54086 , n54120 );
not ( n54122 , n54121 );
buf ( n54123 , n54122 );
buf ( n54124 , n54123 );
not ( n54125 , n54124 );
buf ( n54126 , n54125 );
buf ( n54127 , n54126 );
not ( n54128 , n54127 );
buf ( n54129 , n54128 );
not ( n54130 , n54129 );
not ( n54131 , n39374 );
buf ( n54132 , RI15b49290_361);
not ( n54133 , n54132 );
buf ( n54134 , RI15b49218_360);
not ( n54135 , n54134 );
buf ( n54136 , RI15b491a0_359);
not ( n54137 , n54136 );
buf ( n54138 , RI15b49128_358);
not ( n54139 , n54138 );
buf ( n54140 , RI15b490b0_357);
not ( n54141 , n54140 );
buf ( n54142 , RI15b49038_356);
not ( n54143 , n54142 );
buf ( n54144 , RI15b48fc0_355);
not ( n54145 , n54144 );
buf ( n54146 , RI15b48f48_354);
not ( n54147 , n54146 );
buf ( n54148 , RI15b48ed0_353);
not ( n54149 , n54148 );
buf ( n54150 , RI15b48e58_352);
not ( n54151 , n54150 );
buf ( n54152 , RI15b48de0_351);
not ( n54153 , n54152 );
buf ( n54154 , RI15b48d68_350);
not ( n54155 , n54154 );
buf ( n54156 , RI15b48cf0_349);
not ( n54157 , n54156 );
buf ( n54158 , RI15b48c78_348);
not ( n54159 , n54158 );
and ( n54160 , n54087 , n54118 );
and ( n54161 , n54159 , n54160 );
and ( n54162 , n54157 , n54161 );
and ( n54163 , n54155 , n54162 );
and ( n54164 , n54153 , n54163 );
and ( n54165 , n54151 , n54164 );
and ( n54166 , n54149 , n54165 );
and ( n54167 , n54147 , n54166 );
and ( n54168 , n54145 , n54167 );
and ( n54169 , n54143 , n54168 );
and ( n54170 , n54141 , n54169 );
and ( n54171 , n54139 , n54170 );
and ( n54172 , n54137 , n54171 );
and ( n54173 , n54135 , n54172 );
and ( n54174 , n54133 , n54173 );
xor ( n54175 , n54131 , n54174 );
buf ( n54176 , n39374 );
and ( n54177 , n54175 , n54176 );
buf ( n54178 , n54177 );
not ( n54179 , n54178 );
not ( n54180 , n54179 );
not ( n54181 , n54180 );
not ( n54182 , n39374 );
and ( n54183 , n54182 , n54132 );
xor ( n54184 , n54133 , n54173 );
and ( n54185 , n54184 , n39374 );
or ( n54186 , n54183 , n54185 );
not ( n54187 , n54186 );
buf ( n54188 , n54187 );
buf ( n54189 , n54188 );
not ( n54190 , n54189 );
not ( n54191 , n54190 );
not ( n54192 , n39374 );
and ( n54193 , n54192 , n54134 );
xor ( n54194 , n54135 , n54172 );
and ( n54195 , n54194 , n39374 );
or ( n54196 , n54193 , n54195 );
not ( n54197 , n54196 );
buf ( n54198 , n54197 );
buf ( n54199 , n54198 );
not ( n54200 , n54199 );
not ( n54201 , n54200 );
not ( n54202 , n39374 );
and ( n54203 , n54202 , n54136 );
xor ( n54204 , n54137 , n54171 );
and ( n54205 , n54204 , n39374 );
or ( n54206 , n54203 , n54205 );
not ( n54207 , n54206 );
buf ( n54208 , n54207 );
buf ( n54209 , n54208 );
not ( n54210 , n54209 );
not ( n54211 , n54210 );
not ( n54212 , n39374 );
and ( n54213 , n54212 , n54138 );
xor ( n54214 , n54139 , n54170 );
and ( n54215 , n54214 , n39374 );
or ( n54216 , n54213 , n54215 );
not ( n54217 , n54216 );
buf ( n54218 , n54217 );
buf ( n54219 , n54218 );
not ( n54220 , n54219 );
not ( n54221 , n54220 );
not ( n54222 , n39374 );
and ( n54223 , n54222 , n54140 );
xor ( n54224 , n54141 , n54169 );
and ( n54225 , n54224 , n39374 );
or ( n54226 , n54223 , n54225 );
not ( n54227 , n54226 );
buf ( n54228 , n54227 );
buf ( n54229 , n54228 );
not ( n54230 , n54229 );
not ( n54231 , n54230 );
not ( n54232 , n39374 );
and ( n54233 , n54232 , n54142 );
xor ( n54234 , n54143 , n54168 );
and ( n54235 , n54234 , n39374 );
or ( n54236 , n54233 , n54235 );
not ( n54237 , n54236 );
buf ( n54238 , n54237 );
buf ( n54239 , n54238 );
not ( n54240 , n54239 );
not ( n54241 , n54240 );
not ( n54242 , n39374 );
and ( n54243 , n54242 , n54144 );
xor ( n54244 , n54145 , n54167 );
and ( n54245 , n54244 , n39374 );
or ( n54246 , n54243 , n54245 );
not ( n54247 , n54246 );
buf ( n54248 , n54247 );
buf ( n54249 , n54248 );
not ( n54250 , n54249 );
not ( n54251 , n54250 );
not ( n54252 , n39374 );
and ( n54253 , n54252 , n54146 );
xor ( n54254 , n54147 , n54166 );
and ( n54255 , n54254 , n39374 );
or ( n54256 , n54253 , n54255 );
not ( n54257 , n54256 );
buf ( n54258 , n54257 );
buf ( n54259 , n54258 );
not ( n54260 , n54259 );
not ( n54261 , n54260 );
not ( n54262 , n39374 );
and ( n54263 , n54262 , n54148 );
xor ( n54264 , n54149 , n54165 );
and ( n54265 , n54264 , n39374 );
or ( n54266 , n54263 , n54265 );
not ( n54267 , n54266 );
buf ( n54268 , n54267 );
buf ( n54269 , n54268 );
not ( n54270 , n54269 );
not ( n54271 , n54270 );
not ( n54272 , n39374 );
and ( n54273 , n54272 , n54150 );
xor ( n54274 , n54151 , n54164 );
and ( n54275 , n54274 , n39374 );
or ( n54276 , n54273 , n54275 );
not ( n54277 , n54276 );
buf ( n54278 , n54277 );
buf ( n54279 , n54278 );
not ( n54280 , n54279 );
not ( n54281 , n54280 );
not ( n54282 , n39374 );
and ( n54283 , n54282 , n54152 );
xor ( n54284 , n54153 , n54163 );
and ( n54285 , n54284 , n39374 );
or ( n54286 , n54283 , n54285 );
not ( n54287 , n54286 );
buf ( n54288 , n54287 );
buf ( n54289 , n54288 );
not ( n54290 , n54289 );
not ( n54291 , n54290 );
not ( n54292 , n39374 );
and ( n54293 , n54292 , n54154 );
xor ( n54294 , n54155 , n54162 );
and ( n54295 , n54294 , n39374 );
or ( n54296 , n54293 , n54295 );
not ( n54297 , n54296 );
buf ( n54298 , n54297 );
buf ( n54299 , n54298 );
not ( n54300 , n54299 );
not ( n54301 , n54300 );
not ( n54302 , n39374 );
and ( n54303 , n54302 , n54156 );
xor ( n54304 , n54157 , n54161 );
and ( n54305 , n54304 , n39374 );
or ( n54306 , n54303 , n54305 );
not ( n54307 , n54306 );
buf ( n54308 , n54307 );
buf ( n54309 , n54308 );
not ( n54310 , n54309 );
not ( n54311 , n54310 );
not ( n54312 , n39374 );
and ( n54313 , n54312 , n54158 );
xor ( n54314 , n54159 , n54160 );
and ( n54315 , n54314 , n39374 );
or ( n54316 , n54313 , n54315 );
not ( n54317 , n54316 );
buf ( n54318 , n54317 );
buf ( n54319 , n54318 );
not ( n54320 , n54319 );
not ( n54321 , n54320 );
not ( n54322 , n54125 );
and ( n54323 , n54321 , n54322 );
and ( n54324 , n54311 , n54323 );
and ( n54325 , n54301 , n54324 );
and ( n54326 , n54291 , n54325 );
and ( n54327 , n54281 , n54326 );
and ( n54328 , n54271 , n54327 );
and ( n54329 , n54261 , n54328 );
and ( n54330 , n54251 , n54329 );
and ( n54331 , n54241 , n54330 );
and ( n54332 , n54231 , n54331 );
and ( n54333 , n54221 , n54332 );
and ( n54334 , n54211 , n54333 );
and ( n54335 , n54201 , n54334 );
and ( n54336 , n54191 , n54335 );
and ( n54337 , n54181 , n54336 );
not ( n54338 , n54337 );
and ( n54339 , n54338 , n39374 );
buf ( n54340 , n54339 );
not ( n54341 , n54340 );
not ( n54342 , n39374 );
and ( n54343 , n54342 , n54320 );
xor ( n54344 , n54321 , n54322 );
and ( n54345 , n54344 , n39374 );
or ( n54346 , n54343 , n54345 );
and ( n54347 , n54341 , n54346 );
not ( n54348 , n54346 );
not ( n54349 , n54126 );
xor ( n54350 , n54348 , n54349 );
and ( n54351 , n54350 , n54340 );
or ( n54352 , n54347 , n54351 );
not ( n54353 , n54352 );
buf ( n54354 , n54353 );
buf ( n54355 , n54354 );
not ( n54356 , n54355 );
or ( n54357 , n54130 , n54356 );
not ( n54358 , n54340 );
not ( n54359 , n39374 );
and ( n54360 , n54359 , n54310 );
xor ( n54361 , n54311 , n54323 );
and ( n54362 , n54361 , n39374 );
or ( n54363 , n54360 , n54362 );
and ( n54364 , n54358 , n54363 );
not ( n54365 , n54363 );
and ( n54366 , n54348 , n54349 );
xor ( n54367 , n54365 , n54366 );
and ( n54368 , n54367 , n54340 );
or ( n54369 , n54364 , n54368 );
not ( n54370 , n54369 );
buf ( n54371 , n54370 );
buf ( n54372 , n54371 );
not ( n54373 , n54372 );
or ( n54374 , n54357 , n54373 );
not ( n54375 , n54340 );
not ( n54376 , n39374 );
and ( n54377 , n54376 , n54300 );
xor ( n54378 , n54301 , n54324 );
and ( n54379 , n54378 , n39374 );
or ( n54380 , n54377 , n54379 );
and ( n54381 , n54375 , n54380 );
not ( n54382 , n54380 );
and ( n54383 , n54365 , n54366 );
xor ( n54384 , n54382 , n54383 );
and ( n54385 , n54384 , n54340 );
or ( n54386 , n54381 , n54385 );
not ( n54387 , n54386 );
buf ( n54388 , n54387 );
buf ( n54389 , n54388 );
not ( n54390 , n54389 );
or ( n54391 , n54374 , n54390 );
not ( n54392 , n54340 );
not ( n54393 , n39374 );
and ( n54394 , n54393 , n54290 );
xor ( n54395 , n54291 , n54325 );
and ( n54396 , n54395 , n39374 );
or ( n54397 , n54394 , n54396 );
and ( n54398 , n54392 , n54397 );
not ( n54399 , n54397 );
and ( n54400 , n54382 , n54383 );
xor ( n54401 , n54399 , n54400 );
and ( n54402 , n54401 , n54340 );
or ( n54403 , n54398 , n54402 );
not ( n54404 , n54403 );
buf ( n54405 , n54404 );
buf ( n54406 , n54405 );
not ( n54407 , n54406 );
or ( n54408 , n54391 , n54407 );
not ( n54409 , n54340 );
not ( n54410 , n39374 );
and ( n54411 , n54410 , n54280 );
xor ( n54412 , n54281 , n54326 );
and ( n54413 , n54412 , n39374 );
or ( n54414 , n54411 , n54413 );
and ( n54415 , n54409 , n54414 );
not ( n54416 , n54414 );
and ( n54417 , n54399 , n54400 );
xor ( n54418 , n54416 , n54417 );
and ( n54419 , n54418 , n54340 );
or ( n54420 , n54415 , n54419 );
not ( n54421 , n54420 );
buf ( n54422 , n54421 );
buf ( n54423 , n54422 );
not ( n54424 , n54423 );
or ( n54425 , n54408 , n54424 );
not ( n54426 , n54340 );
not ( n54427 , n39374 );
and ( n54428 , n54427 , n54270 );
xor ( n54429 , n54271 , n54327 );
and ( n54430 , n54429 , n39374 );
or ( n54431 , n54428 , n54430 );
and ( n54432 , n54426 , n54431 );
not ( n54433 , n54431 );
and ( n54434 , n54416 , n54417 );
xor ( n54435 , n54433 , n54434 );
and ( n54436 , n54435 , n54340 );
or ( n54437 , n54432 , n54436 );
not ( n54438 , n54437 );
buf ( n54439 , n54438 );
buf ( n54440 , n54439 );
not ( n54441 , n54440 );
or ( n54442 , n54425 , n54441 );
not ( n54443 , n54340 );
not ( n54444 , n39374 );
and ( n54445 , n54444 , n54260 );
xor ( n54446 , n54261 , n54328 );
and ( n54447 , n54446 , n39374 );
or ( n54448 , n54445 , n54447 );
and ( n54449 , n54443 , n54448 );
not ( n54450 , n54448 );
and ( n54451 , n54433 , n54434 );
xor ( n54452 , n54450 , n54451 );
and ( n54453 , n54452 , n54340 );
or ( n54454 , n54449 , n54453 );
not ( n54455 , n54454 );
buf ( n54456 , n54455 );
buf ( n54457 , n54456 );
not ( n54458 , n54457 );
or ( n54459 , n54442 , n54458 );
not ( n54460 , n54340 );
not ( n54461 , n39374 );
and ( n54462 , n54461 , n54250 );
xor ( n54463 , n54251 , n54329 );
and ( n54464 , n54463 , n39374 );
or ( n54465 , n54462 , n54464 );
and ( n54466 , n54460 , n54465 );
not ( n54467 , n54465 );
and ( n54468 , n54450 , n54451 );
xor ( n54469 , n54467 , n54468 );
and ( n54470 , n54469 , n54340 );
or ( n54471 , n54466 , n54470 );
not ( n54472 , n54471 );
buf ( n54473 , n54472 );
buf ( n54474 , n54473 );
not ( n54475 , n54474 );
or ( n54476 , n54459 , n54475 );
not ( n54477 , n54340 );
not ( n54478 , n39374 );
and ( n54479 , n54478 , n54240 );
xor ( n54480 , n54241 , n54330 );
and ( n54481 , n54480 , n39374 );
or ( n54482 , n54479 , n54481 );
and ( n54483 , n54477 , n54482 );
not ( n54484 , n54482 );
and ( n54485 , n54467 , n54468 );
xor ( n54486 , n54484 , n54485 );
and ( n54487 , n54486 , n54340 );
or ( n54488 , n54483 , n54487 );
not ( n54489 , n54488 );
buf ( n54490 , n54489 );
buf ( n54491 , n54490 );
not ( n54492 , n54491 );
or ( n54493 , n54476 , n54492 );
not ( n54494 , n54340 );
not ( n54495 , n39374 );
and ( n54496 , n54495 , n54230 );
xor ( n54497 , n54231 , n54331 );
and ( n54498 , n54497 , n39374 );
or ( n54499 , n54496 , n54498 );
and ( n54500 , n54494 , n54499 );
not ( n54501 , n54499 );
and ( n54502 , n54484 , n54485 );
xor ( n54503 , n54501 , n54502 );
and ( n54504 , n54503 , n54340 );
or ( n54505 , n54500 , n54504 );
not ( n54506 , n54505 );
buf ( n54507 , n54506 );
buf ( n54508 , n54507 );
not ( n54509 , n54508 );
or ( n54510 , n54493 , n54509 );
not ( n54511 , n54340 );
not ( n54512 , n39374 );
and ( n54513 , n54512 , n54220 );
xor ( n54514 , n54221 , n54332 );
and ( n54515 , n54514 , n39374 );
or ( n54516 , n54513 , n54515 );
and ( n54517 , n54511 , n54516 );
not ( n54518 , n54516 );
and ( n54519 , n54501 , n54502 );
xor ( n54520 , n54518 , n54519 );
and ( n54521 , n54520 , n54340 );
or ( n54522 , n54517 , n54521 );
not ( n54523 , n54522 );
buf ( n54524 , n54523 );
buf ( n54525 , n54524 );
not ( n54526 , n54525 );
or ( n54527 , n54510 , n54526 );
not ( n54528 , n54340 );
not ( n54529 , n39374 );
and ( n54530 , n54529 , n54210 );
xor ( n54531 , n54211 , n54333 );
and ( n54532 , n54531 , n39374 );
or ( n54533 , n54530 , n54532 );
and ( n54534 , n54528 , n54533 );
not ( n54535 , n54533 );
and ( n54536 , n54518 , n54519 );
xor ( n54537 , n54535 , n54536 );
and ( n54538 , n54537 , n54340 );
or ( n54539 , n54534 , n54538 );
not ( n54540 , n54539 );
buf ( n54541 , n54540 );
buf ( n54542 , n54541 );
not ( n54543 , n54542 );
or ( n54544 , n54527 , n54543 );
not ( n54545 , n54340 );
not ( n54546 , n39374 );
and ( n54547 , n54546 , n54200 );
xor ( n54548 , n54201 , n54334 );
and ( n54549 , n54548 , n39374 );
or ( n54550 , n54547 , n54549 );
and ( n54551 , n54545 , n54550 );
not ( n54552 , n54550 );
and ( n54553 , n54535 , n54536 );
xor ( n54554 , n54552 , n54553 );
and ( n54555 , n54554 , n54340 );
or ( n54556 , n54551 , n54555 );
not ( n54557 , n54556 );
buf ( n54558 , n54557 );
buf ( n54559 , n54558 );
not ( n54560 , n54559 );
or ( n54561 , n54544 , n54560 );
not ( n54562 , n54340 );
not ( n54563 , n39374 );
and ( n54564 , n54563 , n54190 );
xor ( n54565 , n54191 , n54335 );
and ( n54566 , n54565 , n39374 );
or ( n54567 , n54564 , n54566 );
and ( n54568 , n54562 , n54567 );
not ( n54569 , n54567 );
and ( n54570 , n54552 , n54553 );
xor ( n54571 , n54569 , n54570 );
and ( n54572 , n54571 , n54340 );
or ( n54573 , n54568 , n54572 );
not ( n54574 , n54573 );
buf ( n54575 , n54574 );
buf ( n54576 , n54575 );
not ( n54577 , n54576 );
or ( n54578 , n54561 , n54577 );
buf ( n54579 , n54578 );
buf ( n54580 , n54579 );
and ( n54581 , n54580 , n54340 );
not ( n54582 , n54581 );
and ( n54583 , n54582 , n54356 );
xor ( n54584 , n54356 , n54340 );
xor ( n54585 , n54130 , n54340 );
and ( n54586 , n54585 , n54340 );
xor ( n54587 , n54584 , n54586 );
and ( n54588 , n54587 , n54581 );
or ( n54589 , n54583 , n54588 );
and ( n54590 , n54589 , n48557 );
or ( n54591 , n54083 , n54590 );
and ( n54592 , n54591 , n33038 );
and ( n54593 , n54078 , n48571 );
or ( n54594 , n54081 , n54592 , n54593 );
and ( n54595 , n54594 , n33208 );
and ( n54596 , n54078 , n48577 );
or ( n54597 , C0 , n54076 , n54595 , n54596 );
buf ( n54598 , n54597 );
buf ( n54599 , n54598 );
buf ( n54600 , n31655 );
buf ( n54601 , n30987 );
buf ( n54602 , n31655 );
buf ( n54603 , RI15b52638_676);
and ( n54604 , n54603 , n31645 );
not ( n54605 , n45274 );
buf ( n54606 , RI15b53c40_723);
and ( n54607 , n54605 , n54606 );
buf ( n54608 , n54607 );
and ( n54609 , n54608 , n31373 );
not ( n54610 , n45280 );
and ( n54611 , n54610 , n54606 );
not ( n54612 , n45766 );
and ( n54613 , n54612 , n45575 );
xor ( n54614 , n45775 , n45781 );
and ( n54615 , n54614 , n45766 );
or ( n54616 , n54613 , n54615 );
and ( n54617 , n54616 , n45280 );
or ( n54618 , n54611 , n54617 );
and ( n54619 , n54618 , n31468 );
and ( n54620 , n54606 , n45802 );
or ( n54621 , n54609 , n54619 , n54620 );
and ( n54622 , n54621 , n31557 );
and ( n54623 , n54606 , n45808 );
or ( n54624 , C0 , n54604 , n54622 , n54623 );
buf ( n54625 , n54624 );
buf ( n54626 , n54625 );
not ( n54627 , n40163 );
and ( n54628 , n54627 , n31939 );
and ( n54629 , n31673 , n31669 , n45160 , n31661 , n42170 );
not ( n54630 , n54629 );
and ( n54631 , n54630 , n31939 );
and ( n54632 , n32183 , n54629 );
or ( n54633 , n54631 , n54632 );
and ( n54634 , n54633 , n40163 );
or ( n54635 , n54628 , n54634 );
and ( n54636 , n54635 , n32498 );
and ( n54637 , n40177 , n40182 , n45169 , n40194 , C1 );
not ( n54638 , n54637 );
not ( n54639 , n54629 );
and ( n54640 , n54639 , n31939 );
and ( n54641 , n45178 , n54629 );
or ( n54642 , n54640 , n54641 );
and ( n54643 , n54638 , n54642 );
and ( n54644 , n45178 , n54637 );
or ( n54645 , n54643 , n54644 );
and ( n54646 , n54645 , n32473 );
not ( n54647 , n32475 );
not ( n54648 , n54637 );
not ( n54649 , n54629 );
and ( n54650 , n54649 , n31939 );
and ( n54651 , n45178 , n54629 );
or ( n54652 , n54650 , n54651 );
and ( n54653 , n54648 , n54652 );
and ( n54654 , n45178 , n54637 );
or ( n54655 , n54653 , n54654 );
and ( n54656 , n54647 , n54655 );
and ( n54657 , n40417 , n40425 , n45195 , n40445 , C1 );
not ( n54658 , n54657 );
and ( n54659 , n40413 , n40421 , n45198 , n40440 , C1 );
not ( n54660 , n54659 );
and ( n54661 , n54660 , n54655 );
and ( n54662 , n45206 , n54659 );
or ( n54663 , n54661 , n54662 );
and ( n54664 , n54658 , n54663 );
and ( n54665 , n45214 , n54657 );
or ( n54666 , n54664 , n54665 );
and ( n54667 , n54666 , n32475 );
or ( n54668 , n54656 , n54667 );
and ( n54669 , n54668 , n32486 );
and ( n54670 , n31939 , n41278 );
or ( n54671 , C0 , n54636 , n54646 , n54669 , n54670 );
buf ( n54672 , n54671 );
buf ( n54673 , n54672 );
buf ( n54674 , n30987 );
buf ( n54675 , n31655 );
and ( n54676 , n39376 , n39369 );
and ( n54677 , n39389 , n54676 );
xor ( n54678 , n39402 , n54677 );
and ( n54679 , n54678 , n33199 );
not ( n54680 , n48648 );
and ( n54681 , n54680 , n39402 );
and ( n54682 , n34221 , n48648 );
or ( n54683 , n54681 , n54682 );
and ( n54684 , n54683 , n32924 );
not ( n54685 , n48660 );
and ( n54686 , n54685 , n39402 );
not ( n54687 , n39584 );
buf ( n54688 , RI15b468d8_272);
and ( n54689 , n54687 , n54688 );
not ( n54690 , n39775 );
and ( n54691 , n54690 , n39627 );
xor ( n54692 , n42661 , n42664 );
and ( n54693 , n54692 , n39775 );
or ( n54694 , n54691 , n54693 );
and ( n54695 , n54694 , n39584 );
or ( n54696 , n54689 , n54695 );
and ( n54697 , n54696 , n48660 );
or ( n54698 , n54686 , n54697 );
and ( n54699 , n54698 , n33172 );
not ( n54700 , n48730 );
and ( n54701 , n54700 , n39402 );
and ( n54702 , n48921 , n48730 );
or ( n54703 , n54701 , n54702 );
and ( n54704 , n54703 , n33187 );
or ( n54705 , n33186 , n33189 );
or ( n54706 , n54705 , n33038 );
or ( n54707 , n54706 , n32890 );
or ( n54708 , n54707 , n33191 );
or ( n54709 , n54708 , n33193 );
or ( n54710 , n54709 , n33195 );
or ( n54711 , n54710 , n33197 );
or ( n54712 , n54711 , n33201 );
or ( n54713 , n54712 , n33203 );
and ( n54714 , n39402 , n54713 );
or ( n54715 , n54679 , n54684 , n54699 , n54704 , n54714 );
and ( n54716 , n54715 , n33208 );
and ( n54717 , n39402 , n39805 );
or ( n54718 , C0 , n54716 , n54717 );
buf ( n54719 , n54718 );
buf ( n54720 , n54719 );
buf ( n54721 , n30987 );
buf ( n54722 , n30987 );
not ( n54723 , n41532 );
buf ( n54724 , RI15b45ff0_253);
not ( n54725 , n54724 );
buf ( n54726 , RI15b45f78_252);
and ( n54727 , n54725 , n54726 );
buf ( n54728 , RI15b45f00_251);
not ( n54729 , n54728 );
and ( n54730 , n54727 , n54729 );
buf ( n54731 , RI15b45e88_250);
not ( n54732 , n54731 );
and ( n54733 , n54730 , n54732 );
buf ( n54734 , RI15b44e98_216);
buf ( n54735 , RI15b44f10_217);
buf ( n54736 , RI15b44f88_218);
buf ( n54737 , RI15b45000_219);
nor ( n54738 , n54734 , n54735 , n54736 , n54737 );
and ( n54739 , n54733 , n54738 );
not ( n54740 , n54739 );
and ( n54741 , n54723 , n54740 );
buf ( n54742 , n41532 );
or ( n54743 , n54741 , n54742 );
buf ( n54744 , n54743 );
buf ( n54745 , n54744 );
buf ( n54746 , n31655 );
buf ( n54747 , n30987 );
not ( n54748 , n40163 );
and ( n54749 , n54748 , n32015 );
not ( n54750 , n52120 );
and ( n54751 , n54750 , n32015 );
and ( n54752 , n32147 , n52120 );
or ( n54753 , n54751 , n54752 );
and ( n54754 , n54753 , n40163 );
or ( n54755 , n54749 , n54754 );
and ( n54756 , n54755 , n32498 );
not ( n54757 , n52128 );
not ( n54758 , n52120 );
and ( n54759 , n54758 , n32015 );
and ( n54760 , n49314 , n52120 );
or ( n54761 , n54759 , n54760 );
and ( n54762 , n54757 , n54761 );
and ( n54763 , n49314 , n52128 );
or ( n54764 , n54762 , n54763 );
and ( n54765 , n54764 , n32473 );
not ( n54766 , n32475 );
not ( n54767 , n52128 );
not ( n54768 , n52120 );
and ( n54769 , n54768 , n32015 );
and ( n54770 , n49314 , n52120 );
or ( n54771 , n54769 , n54770 );
and ( n54772 , n54767 , n54771 );
and ( n54773 , n49314 , n52128 );
or ( n54774 , n54772 , n54773 );
and ( n54775 , n54766 , n54774 );
not ( n54776 , n52148 );
not ( n54777 , n52150 );
and ( n54778 , n54777 , n54774 );
and ( n54779 , n49340 , n52150 );
or ( n54780 , n54778 , n54779 );
and ( n54781 , n54776 , n54780 );
and ( n54782 , n49348 , n52148 );
or ( n54783 , n54781 , n54782 );
and ( n54784 , n54783 , n32475 );
or ( n54785 , n54775 , n54784 );
and ( n54786 , n54785 , n32486 );
and ( n54787 , n32015 , n41278 );
or ( n54788 , C0 , n54756 , n54765 , n54786 , n54787 );
buf ( n54789 , n54788 );
buf ( n54790 , n54789 );
buf ( n54791 , n31655 );
buf ( n54792 , RI15b54258_736);
and ( n54793 , n31450 , n54792 );
not ( n54794 , n48265 );
and ( n54795 , n54793 , n54794 );
not ( n54796 , n54795 );
and ( n54797 , n31451 , n48265 );
not ( n54798 , n54797 );
and ( n54799 , n31451 , n54794 );
and ( n54800 , n54799 , n54792 );
not ( n54801 , n54800 );
not ( n54802 , n54792 );
and ( n54803 , n54799 , n54802 );
not ( n54804 , n54803 );
and ( n54805 , n54801 , n54804 );
buf ( n54806 , n54805 );
and ( n54807 , n54798 , n54806 );
buf ( n54808 , n54797 );
or ( n54809 , n54807 , n54808 );
and ( n54810 , n54796 , n54809 );
buf ( n54811 , n54795 );
or ( n54812 , n54810 , n54811 );
and ( n54813 , n54812 , n37505 );
buf ( n54814 , n36596 );
and ( n54815 , n54792 , n54794 );
not ( n54816 , n54815 );
and ( n54817 , n54802 , n54794 );
not ( n54818 , n54817 );
and ( n54819 , n54816 , n54818 );
buf ( n54820 , n54819 );
and ( n54821 , n54820 , n37503 );
not ( n54822 , n48294 );
and ( n54823 , n54822 , n54794 );
and ( n54824 , n54823 , n54792 );
not ( n54825 , n54824 );
or ( n54826 , n48265 , n54802 );
and ( n54827 , n54822 , n54826 );
not ( n54828 , n54827 );
not ( n54829 , n48294 );
and ( n54830 , n54828 , n54829 );
buf ( n54831 , n54827 );
or ( n54832 , n54830 , n54831 );
and ( n54833 , n54825 , n54832 );
buf ( n54834 , n54824 );
or ( n54835 , n54833 , n54834 );
and ( n54836 , n54835 , n37501 );
not ( n54837 , n54800 );
and ( n54838 , n31450 , n48294 );
not ( n54839 , n54838 );
or ( n54840 , n54792 , n48265 );
and ( n54841 , n31450 , n54822 );
and ( n54842 , n54840 , n54841 );
not ( n54843 , n54842 );
and ( n54844 , n54815 , n31450 );
and ( n54845 , n54844 , n54822 );
not ( n54846 , n54845 );
and ( n54847 , n54817 , n31451 );
not ( n54848 , n54847 );
and ( n54849 , n48265 , n31450 );
and ( n54850 , n54848 , n54849 );
buf ( n54851 , n54850 );
and ( n54852 , n54846 , n54851 );
buf ( n54853 , n54845 );
or ( n54854 , n54852 , n54853 );
and ( n54855 , n54843 , n54854 );
buf ( n54856 , n54842 );
or ( n54857 , n54855 , n54856 );
and ( n54858 , n54839 , n54857 );
and ( n54859 , n31443 , n54838 );
or ( n54860 , n54858 , n54859 );
and ( n54861 , n54837 , n54860 );
buf ( n54862 , n54861 );
and ( n54863 , n54862 , n37499 );
not ( n54864 , n54792 );
and ( n54865 , n54864 , n48265 );
buf ( n54866 , n54865 );
and ( n54867 , n54866 , n37496 );
or ( n54868 , n54813 , n54814 , n54821 , n54836 , n54863 , C0 , n54867 , C0 );
buf ( n54869 , n54868 );
buf ( n54870 , n54869 );
buf ( n54871 , n30987 );
not ( n54872 , n31728 );
and ( n54873 , n54872 , n46036 );
xor ( n54874 , n47613 , n47616 );
and ( n54875 , n54874 , n31728 );
or ( n54876 , n54873 , n54875 );
and ( n54877 , n54876 , n32253 );
not ( n54878 , n32283 );
and ( n54879 , n54878 , n46036 );
not ( n54880 , n31823 );
xor ( n54881 , n47668 , n47671 );
and ( n54882 , n54880 , n54881 );
xnor ( n54883 , n47718 , n47721 );
and ( n54884 , n54883 , n31823 );
or ( n54885 , n54882 , n54884 );
and ( n54886 , n54885 , n32283 );
or ( n54887 , n54879 , n54886 );
and ( n54888 , n54887 , n32398 );
and ( n54889 , n46036 , n32436 );
or ( n54890 , n54877 , n54888 , n54889 );
and ( n54891 , n54890 , n32456 );
and ( n54892 , n49689 , n32473 );
not ( n54893 , n32475 );
and ( n54894 , n54893 , n49689 );
xor ( n54895 , n46036 , n47750 );
and ( n54896 , n54895 , n32475 );
or ( n54897 , n54894 , n54896 );
and ( n54898 , n54897 , n32486 );
and ( n54899 , n37569 , n32489 );
and ( n54900 , n46036 , n32501 );
or ( n54901 , C0 , n54891 , n54892 , n54898 , n54899 , n54900 );
buf ( n54902 , n54901 );
buf ( n54903 , n54902 );
buf ( n54904 , n31655 );
buf ( n54905 , n30987 );
and ( n54906 , n33214 , n32528 );
not ( n54907 , n32598 );
and ( n54908 , n54907 , n32977 );
buf ( n54909 , n54908 );
and ( n54910 , n54909 , n32890 );
not ( n54911 , n32919 );
and ( n54912 , n54911 , n32977 );
buf ( n54913 , n54912 );
and ( n54914 , n54913 , n32924 );
not ( n54915 , n32953 );
and ( n54916 , n54915 , n32977 );
not ( n54917 , n32971 );
and ( n54918 , n54917 , n33079 );
xor ( n54919 , n32977 , n33028 );
and ( n54920 , n54919 , n32971 );
or ( n54921 , n54918 , n54920 );
and ( n54922 , n54921 , n32953 );
or ( n54923 , n54916 , n54922 );
and ( n54924 , n54923 , n33038 );
not ( n54925 , n33067 );
and ( n54926 , n54925 , n32977 );
not ( n54927 , n32970 );
not ( n54928 , n33071 );
and ( n54929 , n54928 , n33079 );
xor ( n54930 , n33080 , n33160 );
and ( n54931 , n54930 , n33071 );
or ( n54932 , n54929 , n54931 );
and ( n54933 , n54927 , n54932 );
and ( n54934 , n54919 , n32970 );
or ( n54935 , n54933 , n54934 );
and ( n54936 , n54935 , n33067 );
or ( n54937 , n54926 , n54936 );
and ( n54938 , n54937 , n33172 );
and ( n54939 , n32977 , n33204 );
or ( n54940 , n54910 , n54914 , n54924 , n54938 , n54939 );
and ( n54941 , n54940 , n33208 );
not ( n54942 , n32968 );
not ( n54943 , n33270 );
and ( n54944 , n54943 , n33279 );
xor ( n54945 , n33280 , n33360 );
and ( n54946 , n54945 , n33270 );
or ( n54947 , n54944 , n54946 );
and ( n54948 , n54942 , n54947 );
and ( n54949 , n32977 , n32968 );
or ( n54950 , n54948 , n54949 );
and ( n54951 , n54950 , n33370 );
and ( n54952 , n32977 , n33382 );
or ( n54953 , C0 , n54906 , n54941 , n54951 , C0 , n54952 );
buf ( n54954 , n54953 );
buf ( n54955 , n54954 );
buf ( n54956 , n30987 );
buf ( n54957 , n31655 );
not ( n54958 , n41532 );
and ( n54959 , n54958 , n34443 );
buf ( n54960 , RI15b53b50_721);
and ( n54961 , n54960 , n41532 );
or ( n54962 , n54959 , n54961 );
buf ( n54963 , n54962 );
buf ( n54964 , n54963 );
buf ( n54965 , n31655 );
buf ( n54966 , n30987 );
and ( n54967 , n39402 , n54677 );
and ( n54968 , n39415 , n54967 );
and ( n54969 , n39428 , n54968 );
and ( n54970 , n39441 , n54969 );
and ( n54971 , n39454 , n54970 );
and ( n54972 , n39467 , n54971 );
and ( n54973 , n39480 , n54972 );
and ( n54974 , n39493 , n54973 );
and ( n54975 , n39506 , n54974 );
and ( n54976 , n39519 , n54975 );
and ( n54977 , n39532 , n54976 );
and ( n54978 , n39545 , n54977 );
and ( n54979 , n39558 , n54978 );
and ( n54980 , n54085 , n54979 );
and ( n54981 , n54158 , n54980 );
and ( n54982 , n54156 , n54981 );
and ( n54983 , n54154 , n54982 );
and ( n54984 , n54152 , n54983 );
xor ( n54985 , n54150 , n54984 );
and ( n54986 , n54985 , n33199 );
not ( n54987 , n48648 );
and ( n54988 , n54987 , n54150 );
and ( n54989 , n34435 , n48648 );
or ( n54990 , n54988 , n54989 );
and ( n54991 , n54990 , n32924 );
not ( n54992 , n48660 );
and ( n54993 , n54992 , n54150 );
buf ( n54994 , n34188 );
not ( n54995 , n54994 );
buf ( n54996 , n54995 );
not ( n54997 , n54996 );
not ( n54998 , n34193 );
and ( n54999 , n54998 , n34195 );
not ( n55000 , n34195 );
not ( n55001 , n34188 );
xor ( n55002 , n55000 , n55001 );
and ( n55003 , n55002 , n34193 );
or ( n55004 , n54999 , n55003 );
not ( n55005 , n55004 );
buf ( n55006 , n55005 );
buf ( n55007 , n55006 );
not ( n55008 , n55007 );
or ( n55009 , n54997 , n55008 );
not ( n55010 , n34193 );
and ( n55011 , n55010 , n34208 );
not ( n55012 , n34208 );
and ( n55013 , n55000 , n55001 );
xor ( n55014 , n55012 , n55013 );
and ( n55015 , n55014 , n34193 );
or ( n55016 , n55011 , n55015 );
not ( n55017 , n55016 );
buf ( n55018 , n55017 );
buf ( n55019 , n55018 );
not ( n55020 , n55019 );
or ( n55021 , n55009 , n55020 );
not ( n55022 , n34193 );
and ( n55023 , n55022 , n34221 );
not ( n55024 , n34221 );
and ( n55025 , n55012 , n55013 );
xor ( n55026 , n55024 , n55025 );
and ( n55027 , n55026 , n34193 );
or ( n55028 , n55023 , n55027 );
not ( n55029 , n55028 );
buf ( n55030 , n55029 );
buf ( n55031 , n55030 );
not ( n55032 , n55031 );
or ( n55033 , n55021 , n55032 );
not ( n55034 , n34193 );
and ( n55035 , n55034 , n34234 );
not ( n55036 , n34234 );
and ( n55037 , n55024 , n55025 );
xor ( n55038 , n55036 , n55037 );
and ( n55039 , n55038 , n34193 );
or ( n55040 , n55035 , n55039 );
not ( n55041 , n55040 );
buf ( n55042 , n55041 );
buf ( n55043 , n55042 );
not ( n55044 , n55043 );
or ( n55045 , n55033 , n55044 );
not ( n55046 , n34193 );
and ( n55047 , n55046 , n34247 );
not ( n55048 , n34247 );
and ( n55049 , n55036 , n55037 );
xor ( n55050 , n55048 , n55049 );
and ( n55051 , n55050 , n34193 );
or ( n55052 , n55047 , n55051 );
not ( n55053 , n55052 );
buf ( n55054 , n55053 );
buf ( n55055 , n55054 );
not ( n55056 , n55055 );
or ( n55057 , n55045 , n55056 );
not ( n55058 , n34193 );
and ( n55059 , n55058 , n34260 );
not ( n55060 , n34260 );
and ( n55061 , n55048 , n55049 );
xor ( n55062 , n55060 , n55061 );
and ( n55063 , n55062 , n34193 );
or ( n55064 , n55059 , n55063 );
not ( n55065 , n55064 );
buf ( n55066 , n55065 );
buf ( n55067 , n55066 );
not ( n55068 , n55067 );
or ( n55069 , n55057 , n55068 );
not ( n55070 , n34193 );
and ( n55071 , n55070 , n34273 );
not ( n55072 , n34273 );
and ( n55073 , n55060 , n55061 );
xor ( n55074 , n55072 , n55073 );
and ( n55075 , n55074 , n34193 );
or ( n55076 , n55071 , n55075 );
not ( n55077 , n55076 );
buf ( n55078 , n55077 );
buf ( n55079 , n55078 );
not ( n55080 , n55079 );
or ( n55081 , n55069 , n55080 );
not ( n55082 , n34193 );
and ( n55083 , n55082 , n34379 );
not ( n55084 , n34379 );
and ( n55085 , n55072 , n55073 );
xor ( n55086 , n55084 , n55085 );
and ( n55087 , n55086 , n34193 );
or ( n55088 , n55083 , n55087 );
not ( n55089 , n55088 );
buf ( n55090 , n55089 );
buf ( n55091 , n55090 );
not ( n55092 , n55091 );
or ( n55093 , n55081 , n55092 );
not ( n55094 , n34193 );
and ( n55095 , n55094 , n34377 );
not ( n55096 , n34377 );
and ( n55097 , n55084 , n55085 );
xor ( n55098 , n55096 , n55097 );
and ( n55099 , n55098 , n34193 );
or ( n55100 , n55095 , n55099 );
not ( n55101 , n55100 );
buf ( n55102 , n55101 );
buf ( n55103 , n55102 );
not ( n55104 , n55103 );
or ( n55105 , n55093 , n55104 );
not ( n55106 , n34193 );
and ( n55107 , n55106 , n34375 );
not ( n55108 , n34375 );
and ( n55109 , n55096 , n55097 );
xor ( n55110 , n55108 , n55109 );
and ( n55111 , n55110 , n34193 );
or ( n55112 , n55107 , n55111 );
not ( n55113 , n55112 );
buf ( n55114 , n55113 );
buf ( n55115 , n55114 );
not ( n55116 , n55115 );
or ( n55117 , n55105 , n55116 );
not ( n55118 , n34193 );
and ( n55119 , n55118 , n34373 );
not ( n55120 , n34373 );
and ( n55121 , n55108 , n55109 );
xor ( n55122 , n55120 , n55121 );
and ( n55123 , n55122 , n34193 );
or ( n55124 , n55119 , n55123 );
not ( n55125 , n55124 );
buf ( n55126 , n55125 );
buf ( n55127 , n55126 );
not ( n55128 , n55127 );
or ( n55129 , n55117 , n55128 );
not ( n55130 , n34193 );
and ( n55131 , n55130 , n34371 );
not ( n55132 , n34371 );
and ( n55133 , n55120 , n55121 );
xor ( n55134 , n55132 , n55133 );
and ( n55135 , n55134 , n34193 );
or ( n55136 , n55131 , n55135 );
not ( n55137 , n55136 );
buf ( n55138 , n55137 );
buf ( n55139 , n55138 );
not ( n55140 , n55139 );
or ( n55141 , n55129 , n55140 );
not ( n55142 , n34193 );
and ( n55143 , n55142 , n34369 );
not ( n55144 , n34369 );
and ( n55145 , n55132 , n55133 );
xor ( n55146 , n55144 , n55145 );
and ( n55147 , n55146 , n34193 );
or ( n55148 , n55143 , n55147 );
not ( n55149 , n55148 );
buf ( n55150 , n55149 );
buf ( n55151 , n55150 );
not ( n55152 , n55151 );
or ( n55153 , n55141 , n55152 );
not ( n55154 , n34193 );
and ( n55155 , n55154 , n34367 );
not ( n55156 , n34367 );
and ( n55157 , n55144 , n55145 );
xor ( n55158 , n55156 , n55157 );
and ( n55159 , n55158 , n34193 );
or ( n55160 , n55155 , n55159 );
not ( n55161 , n55160 );
buf ( n55162 , n55161 );
buf ( n55163 , n55162 );
not ( n55164 , n55163 );
or ( n55165 , n55153 , n55164 );
buf ( n55166 , n55165 );
buf ( n55167 , n55166 );
and ( n55168 , n55167 , n34193 );
not ( n55169 , n55168 );
and ( n55170 , n55169 , n55056 );
xor ( n55171 , n55056 , n34193 );
xor ( n55172 , n55044 , n34193 );
xor ( n55173 , n55032 , n34193 );
xor ( n55174 , n55020 , n34193 );
xor ( n55175 , n55008 , n34193 );
xor ( n55176 , n54997 , n34193 );
and ( n55177 , n55176 , n34193 );
and ( n55178 , n55175 , n55177 );
and ( n55179 , n55174 , n55178 );
and ( n55180 , n55173 , n55179 );
and ( n55181 , n55172 , n55180 );
xor ( n55182 , n55171 , n55181 );
and ( n55183 , n55182 , n55168 );
or ( n55184 , n55170 , n55183 );
and ( n55185 , n55184 , n48660 );
or ( n55186 , n54993 , n55185 );
and ( n55187 , n55186 , n33172 );
not ( n55188 , n48730 );
and ( n55189 , n55188 , n54150 );
not ( n55190 , n32547 );
not ( n55191 , n55190 );
buf ( n55192 , n55191 );
not ( n55193 , n55192 );
not ( n55194 , n55193 );
xnor ( n55195 , n32543 , n32547 );
not ( n55196 , n55195 );
buf ( n55197 , n55196 );
buf ( n55198 , n55197 );
not ( n55199 , n55198 );
not ( n55200 , n55199 );
or ( n55201 , n32543 , n32547 );
xor ( n55202 , n32539 , n55201 );
not ( n55203 , n55202 );
buf ( n55204 , n55203 );
buf ( n55205 , n55204 );
not ( n55206 , n55205 );
not ( n55207 , n55206 );
and ( n55208 , n32539 , n55201 );
xor ( n55209 , n32535 , n55208 );
not ( n55210 , n55209 );
buf ( n55211 , n55210 );
buf ( n55212 , n55211 );
not ( n55213 , n55212 );
not ( n55214 , n55213 );
nor ( n55215 , n55194 , n55200 , n55207 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55216 , n32791 , n55215 );
nor ( n55217 , n55193 , n55200 , n55207 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55218 , n32793 , n55217 );
nor ( n55219 , n55194 , n55199 , n55207 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55220 , n32795 , n55219 );
nor ( n55221 , n55193 , n55199 , n55207 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55222 , n32797 , n55221 );
nor ( n55223 , n55194 , n55200 , n55206 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55224 , n32799 , n55223 );
nor ( n55225 , n55193 , n55200 , n55206 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55226 , n32801 , n55225 );
nor ( n55227 , n55194 , n55199 , n55206 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55228 , n32803 , n55227 );
nor ( n55229 , n55193 , n55199 , n55206 , n55214 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55230 , n32805 , n55229 );
nor ( n55231 , n55194 , n55200 , n55207 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55232 , n32807 , n55231 );
nor ( n55233 , n55193 , n55200 , n55207 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55234 , n32809 , n55233 );
nor ( n55235 , n55194 , n55199 , n55207 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55236 , n32811 , n55235 );
nor ( n55237 , n55193 , n55199 , n55207 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55238 , n32813 , n55237 );
nor ( n55239 , n55194 , n55200 , n55206 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55240 , n32815 , n55239 );
nor ( n55241 , n55193 , n55200 , n55206 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55242 , n32817 , n55241 );
nor ( n55243 , n55194 , n55199 , n55206 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55244 , n32819 , n55243 );
nor ( n55245 , n55193 , n55199 , n55206 , n55213 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n55246 , n32821 , n55245 );
or ( n55247 , n55216 , n55218 , n55220 , n55222 , n55224 , n55226 , n55228 , n55230 , n55232 , n55234 , n55236 , n55238 , n55240 , n55242 , n55244 , n55246 );
and ( n55248 , n55247 , n48730 );
or ( n55249 , n55189 , n55248 );
and ( n55250 , n55249 , n33187 );
and ( n55251 , n54150 , n54713 );
or ( n55252 , n54986 , n54991 , n55187 , n55250 , n55251 );
and ( n55253 , n55252 , n33208 );
and ( n55254 , n54150 , n39805 );
or ( n55255 , C0 , n55253 , n55254 );
buf ( n55256 , n55255 );
buf ( n55257 , n55256 );
buf ( n55258 , n30987 );
buf ( n55259 , n31655 );
buf ( n55260 , n31655 );
not ( n55261 , n46356 );
and ( n55262 , n55261 , n31356 );
nor ( n55263 , n46359 , n46360 , n48213 , n31013 , n31009 );
not ( n55264 , n55263 );
and ( n55265 , n55264 , n31356 );
and ( n55266 , n31372 , n55263 );
or ( n55267 , n55265 , n55266 );
and ( n55268 , n55267 , n46356 );
or ( n55269 , n55262 , n55268 );
and ( n55270 , n55269 , n31649 );
nor ( n55271 , n46374 , n46380 , n48222 , n46392 , C0 );
not ( n55272 , n55271 );
not ( n55273 , n55263 );
and ( n55274 , n55273 , n31356 );
and ( n55275 , n47849 , n55263 );
or ( n55276 , n55274 , n55275 );
and ( n55277 , n55272 , n55276 );
and ( n55278 , n47849 , n55271 );
or ( n55279 , n55277 , n55278 );
and ( n55280 , n55279 , n31643 );
not ( n55281 , n31452 );
not ( n55282 , n55271 );
not ( n55283 , n55263 );
and ( n55284 , n55283 , n31356 );
and ( n55285 , n47849 , n55263 );
or ( n55286 , n55284 , n55285 );
and ( n55287 , n55282 , n55286 );
and ( n55288 , n47849 , n55271 );
or ( n55289 , n55287 , n55288 );
and ( n55290 , n55281 , n55289 );
nor ( n55291 , n46520 , n46529 , n48243 , n46549 , C0 );
not ( n55292 , n55291 );
nor ( n55293 , n46552 , n46553 , n48246 , n46544 , C0 );
not ( n55294 , n55293 );
and ( n55295 , n55294 , n55289 );
and ( n55296 , n47877 , n55293 );
or ( n55297 , n55295 , n55296 );
and ( n55298 , n55292 , n55297 );
and ( n55299 , n47887 , n55291 );
or ( n55300 , n55298 , n55299 );
and ( n55301 , n55300 , n31452 );
or ( n55302 , n55290 , n55301 );
and ( n55303 , n55302 , n31638 );
and ( n55304 , n31356 , n47277 );
or ( n55305 , C0 , n55270 , n55280 , n55303 , n55304 );
buf ( n55306 , n55305 );
buf ( n55307 , n55306 );
buf ( n55308 , n30987 );
xor ( n55309 , n46094 , n46087 );
and ( n55310 , n55309 , n32431 );
not ( n55311 , n50002 );
and ( n55312 , n55311 , n46094 );
and ( n55313 , n40251 , n50002 );
or ( n55314 , n55312 , n55313 );
and ( n55315 , n55314 , n32419 );
not ( n55316 , n50008 );
and ( n55317 , n55316 , n46094 );
not ( n55318 , n47910 );
buf ( n55319 , RI15b5f0b8_1108);
and ( n55320 , n55318 , n55319 );
not ( n55321 , n48101 );
and ( n55322 , n55321 , n47929 );
xor ( n55323 , n48110 , n48112 );
and ( n55324 , n55323 , n48101 );
or ( n55325 , n55322 , n55324 );
and ( n55326 , n55325 , n47910 );
or ( n55327 , n55320 , n55326 );
and ( n55328 , n55327 , n50008 );
or ( n55329 , n55317 , n55328 );
and ( n55330 , n55329 , n32415 );
not ( n55331 , n50067 );
and ( n55332 , n55331 , n46094 );
and ( n55333 , n32033 , n50067 );
or ( n55334 , n55332 , n55333 );
and ( n55335 , n55334 , n32411 );
and ( n55336 , n46094 , n50098 );
or ( n55337 , n55310 , n55315 , n55330 , n55335 , n55336 );
and ( n55338 , n55337 , n32456 );
and ( n55339 , n46094 , n47409 );
or ( n55340 , C0 , n55338 , n55339 );
buf ( n55341 , n55340 );
buf ( n55342 , n55341 );
buf ( n55343 , n31655 );
not ( n55344 , n41532 );
and ( n55345 , n55344 , n34433 );
buf ( n55346 , RI15b53da8_726);
and ( n55347 , n55346 , n41532 );
or ( n55348 , n55345 , n55347 );
buf ( n55349 , n55348 );
buf ( n55350 , n55349 );
buf ( n55351 , n31655 );
buf ( n55352 , n31655 );
buf ( n55353 , n30987 );
xor ( n55354 , n54085 , n54979 );
and ( n55355 , n55354 , n33199 );
not ( n55356 , n48648 );
and ( n55357 , n55356 , n54085 );
and ( n55358 , n34362 , n48648 );
or ( n55359 , n55357 , n55358 );
and ( n55360 , n55359 , n32924 );
not ( n55361 , n48660 );
and ( n55362 , n55361 , n54085 );
not ( n55363 , n55168 );
and ( n55364 , n55363 , n54997 );
xor ( n55365 , n55176 , n34193 );
and ( n55366 , n55365 , n55168 );
or ( n55367 , n55364 , n55366 );
and ( n55368 , n55367 , n48660 );
or ( n55369 , n55362 , n55368 );
and ( n55370 , n55369 , n33172 );
not ( n55371 , n48730 );
and ( n55372 , n55371 , n54085 );
and ( n55373 , n32603 , n55215 );
and ( n55374 , n32607 , n55217 );
and ( n55375 , n32611 , n55219 );
and ( n55376 , n32615 , n55221 );
and ( n55377 , n32618 , n55223 );
and ( n55378 , n32622 , n55225 );
and ( n55379 , n32625 , n55227 );
and ( n55380 , n32628 , n55229 );
and ( n55381 , n32631 , n55231 );
and ( n55382 , n32634 , n55233 );
and ( n55383 , n32637 , n55235 );
and ( n55384 , n32640 , n55237 );
and ( n55385 , n32643 , n55239 );
and ( n55386 , n32646 , n55241 );
and ( n55387 , n32649 , n55243 );
and ( n55388 , n32652 , n55245 );
or ( n55389 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 );
and ( n55390 , n55389 , n48730 );
or ( n55391 , n55372 , n55390 );
and ( n55392 , n55391 , n33187 );
and ( n55393 , n54085 , n54713 );
or ( n55394 , n55355 , n55360 , n55370 , n55392 , n55393 );
and ( n55395 , n55394 , n33208 );
and ( n55396 , n54085 , n39805 );
or ( n55397 , C0 , n55395 , n55396 );
buf ( n55398 , n55397 );
buf ( n55399 , n55398 );
buf ( n55400 , n30987 );
xor ( n55401 , n39428 , n54968 );
and ( n55402 , n55401 , n33199 );
not ( n55403 , n48648 );
and ( n55404 , n55403 , n39428 );
and ( n55405 , n34247 , n48648 );
or ( n55406 , n55404 , n55405 );
and ( n55407 , n55406 , n32924 );
not ( n55408 , n48660 );
and ( n55409 , n55408 , n39428 );
not ( n55410 , n39584 );
buf ( n55411 , RI15b469c8_274);
and ( n55412 , n55410 , n55411 );
not ( n55413 , n39775 );
and ( n55414 , n55413 , n39651 );
xor ( n55415 , n42659 , n42666 );
and ( n55416 , n55415 , n39775 );
or ( n55417 , n55414 , n55416 );
and ( n55418 , n55417 , n39584 );
or ( n55419 , n55412 , n55418 );
and ( n55420 , n55419 , n48660 );
or ( n55421 , n55409 , n55420 );
and ( n55422 , n55421 , n33172 );
not ( n55423 , n48730 );
and ( n55424 , n55423 , n39428 );
and ( n55425 , n48883 , n48730 );
or ( n55426 , n55424 , n55425 );
and ( n55427 , n55426 , n33187 );
and ( n55428 , n39428 , n54713 );
or ( n55429 , n55402 , n55407 , n55422 , n55427 , n55428 );
and ( n55430 , n55429 , n33208 );
and ( n55431 , n39428 , n39805 );
or ( n55432 , C0 , n55430 , n55431 );
buf ( n55433 , n55432 );
buf ( n55434 , n55433 );
buf ( n55435 , n31655 );
buf ( n55436 , n30987 );
buf ( n55437 , n30987 );
buf ( n55438 , n31655 );
not ( n55439 , n50828 );
not ( n55440 , n50834 );
and ( n55441 , n55439 , n55440 );
buf ( n55442 , n50828 );
or ( n55443 , n55441 , n55442 );
buf ( n55444 , n55443 );
buf ( n55445 , n55444 );
buf ( n55446 , n30987 );
buf ( n55447 , RI15b5f220_1111);
and ( n55448 , n55447 , n32494 );
not ( n55449 , n46083 );
and ( n55450 , n55449 , n50841 );
not ( n55451 , n46290 );
and ( n55452 , n55451 , n46143 );
xor ( n55453 , n46302 , n46310 );
and ( n55454 , n55453 , n46290 );
or ( n55455 , n55452 , n55454 );
and ( n55456 , n55455 , n46083 );
or ( n55457 , n55450 , n55456 );
and ( n55458 , n55457 , n32421 );
not ( n55459 , n46326 );
and ( n55460 , n55459 , n50841 );
and ( n55461 , n55455 , n46326 );
or ( n55462 , n55460 , n55461 );
and ( n55463 , n55462 , n32417 );
and ( n55464 , n50841 , n46340 );
or ( n55465 , n55458 , n55463 , n55464 );
and ( n55466 , n55465 , n32456 );
and ( n55467 , n50841 , n46349 );
or ( n55468 , C0 , n55448 , n55466 , n55467 );
buf ( n55469 , n55468 );
buf ( n55470 , n55469 );
not ( n55471 , n46356 );
and ( n55472 , n55471 , n31177 );
and ( n55473 , n31025 , n46360 , n31017 , n31013 , n46361 );
not ( n55474 , n55473 );
and ( n55475 , n55474 , n31177 );
and ( n55476 , n31205 , n55473 );
or ( n55477 , n55475 , n55476 );
and ( n55478 , n55477 , n46356 );
or ( n55479 , n55472 , n55478 );
and ( n55480 , n55479 , n31649 );
and ( n55481 , n46373 , n46380 , n46386 , n46392 , C1 );
not ( n55482 , n55481 );
not ( n55483 , n55473 );
and ( n55484 , n55483 , n31177 );
and ( n55485 , n50125 , n55473 );
or ( n55486 , n55484 , n55485 );
and ( n55487 , n55482 , n55486 );
and ( n55488 , n50125 , n55481 );
or ( n55489 , n55487 , n55488 );
and ( n55490 , n55489 , n31643 );
not ( n55491 , n31452 );
not ( n55492 , n55481 );
not ( n55493 , n55473 );
and ( n55494 , n55493 , n31177 );
and ( n55495 , n50125 , n55473 );
or ( n55496 , n55494 , n55495 );
and ( n55497 , n55492 , n55496 );
and ( n55498 , n50125 , n55481 );
or ( n55499 , n55497 , n55498 );
and ( n55500 , n55491 , n55499 );
and ( n55501 , n46519 , n46529 , n46539 , n46549 , C1 );
not ( n55502 , n55501 );
and ( n55503 , n46515 , n46553 , n46534 , n46544 , C1 );
not ( n55504 , n55503 );
and ( n55505 , n55504 , n55499 );
and ( n55506 , n50151 , n55503 );
or ( n55507 , n55505 , n55506 );
and ( n55508 , n55502 , n55507 );
and ( n55509 , n50159 , n55501 );
or ( n55510 , n55508 , n55509 );
and ( n55511 , n55510 , n31452 );
or ( n55512 , n55500 , n55511 );
and ( n55513 , n55512 , n31638 );
and ( n55514 , n31177 , n47277 );
or ( n55515 , C0 , n55480 , n55490 , n55513 , n55514 );
buf ( n55516 , n55515 );
buf ( n55517 , n55516 );
buf ( n55518 , n31655 );
buf ( n55519 , n31655 );
buf ( n55520 , n31655 );
buf ( n55521 , n31655 );
buf ( n55522 , n30987 );
buf ( n55523 , n30987 );
and ( n55524 , n51913 , n33377 );
not ( n55525 , n48545 );
buf ( n55526 , RI15b47328_294);
and ( n55527 , n55525 , n55526 );
and ( n55528 , n51919 , n48545 );
or ( n55529 , n55527 , n55528 );
and ( n55530 , n55529 , n32890 );
not ( n55531 , n48557 );
and ( n55532 , n55531 , n55526 );
and ( n55533 , n51919 , n48557 );
or ( n55534 , n55532 , n55533 );
and ( n55535 , n55534 , n33038 );
and ( n55536 , n55526 , n48571 );
or ( n55537 , n55530 , n55535 , n55536 );
and ( n55538 , n55537 , n33208 );
and ( n55539 , n55526 , n48577 );
or ( n55540 , C0 , n55524 , n55538 , n55539 );
buf ( n55541 , n55540 );
buf ( n55542 , n55541 );
buf ( n55543 , n30987 );
not ( n55544 , n35542 );
and ( n55545 , n55544 , n41860 );
buf ( n55546 , RI15b45a50_241);
and ( n55547 , n55546 , n35542 );
or ( n55548 , n55545 , n55547 );
buf ( n55549 , n55548 );
buf ( n55550 , n55549 );
buf ( n55551 , n30987 );
buf ( n55552 , n31655 );
not ( n55553 , n40163 );
and ( n55554 , n55553 , n31661 );
and ( n55555 , n40194 , n40163 );
or ( n55556 , n55554 , n55555 );
and ( n55557 , n55556 , n32498 );
buf ( n55558 , RI15b584e8_878);
not ( n55559 , n55558 );
and ( n55560 , n55559 , n31658 );
buf ( n55561 , n55560 );
not ( n55562 , n55561 );
not ( n55563 , n55558 );
and ( n55564 , n55563 , n31666 );
buf ( n55565 , RI15b5d240_1043);
not ( n55566 , n55565 );
not ( n55567 , n50407 );
not ( n55568 , n50408 );
not ( n55569 , n50409 );
not ( n55570 , n50410 );
not ( n55571 , n50411 );
not ( n55572 , n47567 );
not ( n55573 , n47568 );
not ( n55574 , n47569 );
not ( n55575 , n47570 );
not ( n55576 , n47571 );
not ( n55577 , n47572 );
not ( n55578 , n47573 );
not ( n55579 , n47574 );
not ( n55580 , n47575 );
not ( n55581 , n47576 );
not ( n55582 , n47577 );
not ( n55583 , n47578 );
not ( n55584 , n47579 );
not ( n55585 , n47580 );
not ( n55586 , n47581 );
not ( n55587 , n47582 );
not ( n55588 , n41286 );
not ( n55589 , n31732 );
not ( n55590 , n31733 );
not ( n55591 , n31734 );
not ( n55592 , n31735 );
not ( n55593 , n31736 );
not ( n55594 , n31737 );
not ( n55595 , n31738 );
not ( n55596 , n31739 );
not ( n55597 , n31740 );
and ( n55598 , n55596 , n55597 );
and ( n55599 , n55595 , n55598 );
and ( n55600 , n55594 , n55599 );
and ( n55601 , n55593 , n55600 );
and ( n55602 , n55592 , n55601 );
and ( n55603 , n55591 , n55602 );
and ( n55604 , n55590 , n55603 );
and ( n55605 , n55589 , n55604 );
and ( n55606 , n55588 , n55605 );
and ( n55607 , n55587 , n55606 );
and ( n55608 , n55586 , n55607 );
and ( n55609 , n55585 , n55608 );
and ( n55610 , n55584 , n55609 );
and ( n55611 , n55583 , n55610 );
and ( n55612 , n55582 , n55611 );
and ( n55613 , n55581 , n55612 );
and ( n55614 , n55580 , n55613 );
and ( n55615 , n55579 , n55614 );
and ( n55616 , n55578 , n55615 );
and ( n55617 , n55577 , n55616 );
and ( n55618 , n55576 , n55617 );
and ( n55619 , n55575 , n55618 );
and ( n55620 , n55574 , n55619 );
and ( n55621 , n55573 , n55620 );
and ( n55622 , n55572 , n55621 );
and ( n55623 , n55571 , n55622 );
and ( n55624 , n55570 , n55623 );
and ( n55625 , n55569 , n55624 );
and ( n55626 , n55568 , n55625 );
and ( n55627 , n55567 , n55626 );
xor ( n55628 , n55566 , n55627 );
buf ( n55629 , n55565 );
and ( n55630 , n55628 , n55629 );
buf ( n55631 , n55630 );
not ( n55632 , n55631 );
not ( n55633 , n55565 );
and ( n55634 , n55633 , n31739 );
xor ( n55635 , n55596 , n55597 );
and ( n55636 , n55635 , n55565 );
or ( n55637 , n55634 , n55636 );
and ( n55638 , n55632 , n55637 );
not ( n55639 , n55637 );
buf ( n55640 , n31740 );
not ( n55641 , n55640 );
xor ( n55642 , n55639 , n55641 );
and ( n55643 , n55642 , n55631 );
or ( n55644 , n55638 , n55643 );
not ( n55645 , n55644 );
buf ( n55646 , n55645 );
buf ( n55647 , n55646 );
not ( n55648 , n55647 );
xor ( n55649 , n55648 , n55631 );
buf ( n55650 , n55640 );
not ( n55651 , n55650 );
buf ( n55652 , n55651 );
not ( n55653 , n55652 );
xor ( n55654 , n55653 , n55631 );
and ( n55655 , n55654 , n55631 );
and ( n55656 , n55649 , n55655 );
buf ( n55657 , n55656 );
or ( n55658 , n55653 , n55648 );
buf ( n55659 , n55658 );
buf ( n55660 , n55659 );
and ( n55661 , n55660 , n55631 );
and ( n55662 , n55657 , n55661 );
buf ( n55663 , n55662 );
not ( n55664 , n55661 );
and ( n55665 , n55664 , n55648 );
xor ( n55666 , n55649 , n55655 );
and ( n55667 , n55666 , n55661 );
or ( n55668 , n55665 , n55667 );
not ( n55669 , n55661 );
and ( n55670 , n55669 , n55653 );
xor ( n55671 , n55654 , n55631 );
and ( n55672 , n55671 , n55661 );
or ( n55673 , n55670 , n55672 );
and ( n55674 , n55668 , n55673 );
xor ( n55675 , n55663 , n55674 );
buf ( n55676 , n55675 );
buf ( n55677 , n55676 );
not ( n55678 , n55677 );
buf ( n55679 , n55678 );
buf ( n55680 , n55679 );
not ( n55681 , n55680 );
buf ( n55682 , n55681 );
buf ( n55683 , n55682 );
buf ( n55684 , n55640 );
not ( n55685 , n55684 );
buf ( n55686 , n55685 );
not ( n55687 , n55686 );
buf ( n55688 , n55687 );
buf ( n55689 , n55688 );
and ( n55690 , n55689 , n55631 );
not ( n55691 , n55690 );
and ( n55692 , n55691 , n55687 );
xor ( n55693 , n55687 , n55631 );
xor ( n55694 , n55693 , n55631 );
and ( n55695 , n55694 , n55690 );
or ( n55696 , n55692 , n55695 );
not ( n55697 , n55696 );
not ( n55698 , n55697 );
and ( n55699 , n55683 , n55698 );
buf ( n55700 , n55699 );
and ( n55701 , n55700 , n55558 );
or ( n55702 , n55564 , n55701 );
not ( n55703 , n55702 );
not ( n55704 , n55558 );
and ( n55705 , n55704 , n31662 );
and ( n55706 , n55663 , n55674 );
buf ( n55707 , n55706 );
buf ( n55708 , n55707 );
not ( n55709 , n55708 );
buf ( n55710 , n55709 );
buf ( n55711 , n55710 );
not ( n55712 , n55711 );
buf ( n55713 , n55712 );
buf ( n55714 , n55713 );
and ( n55715 , n55714 , n55698 );
buf ( n55716 , n55715 );
and ( n55717 , n55716 , n55558 );
or ( n55718 , n55705 , n55717 );
not ( n55719 , n55718 );
buf ( n55720 , n55561 );
buf ( n55721 , n55561 );
buf ( n55722 , n55561 );
buf ( n55723 , n55561 );
buf ( n55724 , n55561 );
buf ( n55725 , n55561 );
buf ( n55726 , n55561 );
buf ( n55727 , n55561 );
buf ( n55728 , n55561 );
buf ( n55729 , n55561 );
buf ( n55730 , n55561 );
buf ( n55731 , n55561 );
buf ( n55732 , n55561 );
buf ( n55733 , n55561 );
buf ( n55734 , n55561 );
buf ( n55735 , n55561 );
buf ( n55736 , n55561 );
buf ( n55737 , n55561 );
buf ( n55738 , n55561 );
buf ( n55739 , n55561 );
buf ( n55740 , n55561 );
buf ( n55741 , n55561 );
buf ( n55742 , n55561 );
buf ( n55743 , n55561 );
buf ( n55744 , n55561 );
buf ( n55745 , n55561 );
not ( n55746 , n55558 );
and ( n55747 , n55746 , n31674 );
not ( n55748 , n55698 );
buf ( n55749 , n55748 );
not ( n55750 , n55673 );
buf ( n55751 , n55750 );
not ( n55752 , n55751 );
buf ( n55753 , n55752 );
not ( n55754 , n55753 );
buf ( n55755 , n55754 );
buf ( n55756 , n55755 );
and ( n55757 , n55756 , n55698 );
or ( n55758 , n55749 , n55757 );
and ( n55759 , n55758 , n55558 );
or ( n55760 , n55747 , n55759 );
not ( n55761 , n55760 );
not ( n55762 , n55558 );
and ( n55763 , n55762 , n31670 );
xor ( n55764 , n55668 , n55673 );
buf ( n55765 , n55764 );
buf ( n55766 , n55765 );
not ( n55767 , n55766 );
buf ( n55768 , n55767 );
buf ( n55769 , n55768 );
not ( n55770 , n55769 );
buf ( n55771 , n55770 );
buf ( n55772 , n55771 );
and ( n55773 , n55772 , n55698 );
buf ( n55774 , n55773 );
and ( n55775 , n55774 , n55558 );
or ( n55776 , n55763 , n55775 );
not ( n55777 , n55776 );
and ( n55778 , n55761 , n55777 );
or ( n55779 , n55703 , n55719 , n55561 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55778 );
nand ( n55780 , n55562 , n55779 );
not ( n55781 , n55780 );
not ( n55782 , n55558 );
and ( n55783 , n55782 , n31661 );
buf ( n55784 , n55783 );
and ( n55785 , n55781 , n55784 );
buf ( n55786 , n55785 );
and ( n55787 , n55786 , n32496 );
and ( n55788 , n40440 , n32473 );
not ( n55789 , n32475 );
and ( n55790 , n55789 , n40440 );
and ( n55791 , n40425 , n40417 );
and ( n55792 , n40435 , n55791 );
xor ( n55793 , n40445 , n55792 );
not ( n55794 , n55793 );
buf ( n55795 , n55794 );
not ( n55796 , n55795 );
and ( n55797 , n55796 , n32475 );
or ( n55798 , n55790 , n55797 );
and ( n55799 , n55798 , n32486 );
or ( n55800 , n41276 , n32500 );
and ( n55801 , n31661 , n55800 );
or ( n55802 , C0 , n55557 , n55787 , n55788 , n55799 , n55801 );
buf ( n55803 , n55802 );
buf ( n55804 , n55803 );
not ( n55805 , n33419 );
and ( n55806 , n55805 , n31588 );
xor ( n55807 , n33611 , n33628 );
xor ( n55808 , n55807 , n33670 );
and ( n55809 , n55808 , n33419 );
or ( n55810 , n55806 , n55809 );
and ( n55811 , n55810 , n31529 );
not ( n55812 , n33734 );
and ( n55813 , n55812 , n31588 );
not ( n55814 , n33533 );
xor ( n55815 , n33781 , n33628 );
xor ( n55816 , n55815 , n33788 );
and ( n55817 , n55814 , n55816 );
xor ( n55818 , n33876 , n33878 );
xor ( n55819 , n55818 , n33890 );
and ( n55820 , n55819 , n33533 );
or ( n55821 , n55817 , n55820 );
and ( n55822 , n55821 , n33734 );
or ( n55823 , n55813 , n55822 );
and ( n55824 , n55823 , n31527 );
and ( n55825 , n31588 , n33942 );
or ( n55826 , n55811 , n55824 , n55825 );
and ( n55827 , n55826 , n31557 );
and ( n55828 , n31624 , n31643 );
not ( n55829 , n31452 );
and ( n55830 , n55829 , n31624 );
not ( n55831 , n31588 );
and ( n55832 , n55831 , n31452 );
or ( n55833 , n55830 , n55832 );
and ( n55834 , n55833 , n31638 );
and ( n55835 , n31459 , n33973 );
and ( n55836 , n31588 , n33978 );
or ( n55837 , C0 , n55827 , n55828 , n55834 , n55835 , n55836 );
buf ( n55838 , n55837 );
buf ( n55839 , n55838 );
xor ( n55840 , n44771 , n44796 );
and ( n55841 , n55840 , n31548 );
not ( n55842 , n44807 );
and ( n55843 , n55842 , n44771 );
and ( n55844 , n46652 , n44807 );
or ( n55845 , n55843 , n55844 );
and ( n55846 , n55845 , n31408 );
not ( n55847 , n44817 );
and ( n55848 , n55847 , n44771 );
not ( n55849 , n44994 );
and ( n55850 , n55849 , n44882 );
xor ( n55851 , n45005 , n45015 );
and ( n55852 , n55851 , n44994 );
or ( n55853 , n55850 , n55852 );
and ( n55854 , n55853 , n44817 );
or ( n55855 , n55848 , n55854 );
and ( n55856 , n55855 , n31521 );
not ( n55857 , n45059 );
and ( n55858 , n55857 , n44771 );
and ( n55859 , n31274 , n40095 );
and ( n55860 , n31276 , n40097 );
and ( n55861 , n31278 , n40099 );
and ( n55862 , n31280 , n40101 );
and ( n55863 , n31282 , n40103 );
and ( n55864 , n31284 , n40105 );
and ( n55865 , n31286 , n40107 );
and ( n55866 , n31288 , n40109 );
and ( n55867 , n31290 , n40111 );
and ( n55868 , n31292 , n40113 );
and ( n55869 , n31294 , n40115 );
and ( n55870 , n31296 , n40117 );
and ( n55871 , n31298 , n40119 );
and ( n55872 , n31300 , n40121 );
and ( n55873 , n31302 , n40123 );
and ( n55874 , n31304 , n40125 );
or ( n55875 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 );
and ( n55876 , n55875 , n45059 );
or ( n55877 , n55858 , n55876 );
and ( n55878 , n55877 , n31536 );
and ( n55879 , n44771 , n45148 );
or ( n55880 , n55841 , n55846 , n55856 , n55878 , n55879 );
and ( n55881 , n55880 , n31557 );
and ( n55882 , n44771 , n40154 );
or ( n55883 , C0 , n55881 , n55882 );
buf ( n55884 , n55883 );
buf ( n55885 , n55884 );
not ( n55886 , n40163 );
and ( n55887 , n55886 , n31951 );
nor ( n55888 , n42169 , n31669 , n45160 , n31661 , n31657 );
not ( n55889 , n55888 );
and ( n55890 , n55889 , n31951 );
and ( n55891 , n32183 , n55888 );
or ( n55892 , n55890 , n55891 );
and ( n55893 , n55892 , n40163 );
or ( n55894 , n55887 , n55893 );
and ( n55895 , n55894 , n32498 );
nor ( n55896 , n42179 , n40182 , n45169 , n40194 , C0 );
not ( n55897 , n55896 );
not ( n55898 , n55888 );
and ( n55899 , n55898 , n31951 );
and ( n55900 , n45178 , n55888 );
or ( n55901 , n55899 , n55900 );
and ( n55902 , n55897 , n55901 );
and ( n55903 , n45178 , n55896 );
or ( n55904 , n55902 , n55903 );
and ( n55905 , n55904 , n32473 );
not ( n55906 , n32475 );
not ( n55907 , n55896 );
not ( n55908 , n55888 );
and ( n55909 , n55908 , n31951 );
and ( n55910 , n45178 , n55888 );
or ( n55911 , n55909 , n55910 );
and ( n55912 , n55907 , n55911 );
and ( n55913 , n45178 , n55896 );
or ( n55914 , n55912 , n55913 );
and ( n55915 , n55906 , n55914 );
nor ( n55916 , n42205 , n40425 , n45195 , n40445 , C0 );
not ( n55917 , n55916 );
nor ( n55918 , n42208 , n40421 , n45198 , n40440 , C0 );
not ( n55919 , n55918 );
and ( n55920 , n55919 , n55914 );
and ( n55921 , n45206 , n55918 );
or ( n55922 , n55920 , n55921 );
and ( n55923 , n55917 , n55922 );
and ( n55924 , n45214 , n55916 );
or ( n55925 , n55923 , n55924 );
and ( n55926 , n55925 , n32475 );
or ( n55927 , n55915 , n55926 );
and ( n55928 , n55927 , n32486 );
and ( n55929 , n31951 , n41278 );
or ( n55930 , C0 , n55895 , n55905 , n55928 , n55929 );
buf ( n55931 , n55930 );
buf ( n55932 , n55931 );
buf ( n55933 , n30987 );
buf ( n55934 , n30987 );
buf ( n55935 , n31655 );
buf ( n55936 , n31655 );
buf ( n55937 , n30987 );
not ( n55938 , n34150 );
and ( n55939 , n55938 , n32725 );
not ( n55940 , n50731 );
and ( n55941 , n55940 , n32725 );
and ( n55942 , n32755 , n50731 );
or ( n55943 , n55941 , n55942 );
and ( n55944 , n55943 , n34150 );
or ( n55945 , n55939 , n55944 );
and ( n55946 , n55945 , n33381 );
not ( n55947 , n50739 );
not ( n55948 , n50731 );
and ( n55949 , n55948 , n32725 );
and ( n55950 , n35083 , n50731 );
or ( n55951 , n55949 , n55950 );
and ( n55952 , n55947 , n55951 );
and ( n55953 , n35083 , n50739 );
or ( n55954 , n55952 , n55953 );
and ( n55955 , n55954 , n33375 );
not ( n55956 , n32968 );
not ( n55957 , n50739 );
not ( n55958 , n50731 );
and ( n55959 , n55958 , n32725 );
and ( n55960 , n35083 , n50731 );
or ( n55961 , n55959 , n55960 );
and ( n55962 , n55957 , n55961 );
and ( n55963 , n35083 , n50739 );
or ( n55964 , n55962 , n55963 );
and ( n55965 , n55956 , n55964 );
not ( n55966 , n50759 );
not ( n55967 , n50761 );
and ( n55968 , n55967 , n55964 );
and ( n55969 , n35107 , n50761 );
or ( n55970 , n55968 , n55969 );
and ( n55971 , n55966 , n55970 );
and ( n55972 , n35115 , n50759 );
or ( n55973 , n55971 , n55972 );
and ( n55974 , n55973 , n32968 );
or ( n55975 , n55965 , n55974 );
and ( n55976 , n55975 , n33370 );
and ( n55977 , n32725 , n35062 );
or ( n55978 , C0 , n55946 , n55955 , n55976 , n55977 );
buf ( n55979 , n55978 );
buf ( n55980 , n55979 );
buf ( n55981 , n30987 );
buf ( n55982 , n31655 );
buf ( n55983 , n31655 );
buf ( n55984 , n30987 );
not ( n55985 , n34150 );
and ( n55986 , n55985 , n32883 );
not ( n55987 , n34154 );
and ( n55988 , n55987 , n32883 );
and ( n55989 , n32889 , n34154 );
or ( n55990 , n55988 , n55989 );
and ( n55991 , n55990 , n34150 );
or ( n55992 , n55986 , n55991 );
and ( n55993 , n55992 , n33381 );
not ( n55994 , n34184 );
not ( n55995 , n34154 );
and ( n55996 , n55995 , n32883 );
and ( n55997 , n52819 , n34154 );
or ( n55998 , n55996 , n55997 );
and ( n55999 , n55994 , n55998 );
and ( n56000 , n52819 , n34184 );
or ( n56001 , n55999 , n56000 );
and ( n56002 , n56001 , n33375 );
not ( n56003 , n32968 );
not ( n56004 , n34184 );
not ( n56005 , n34154 );
and ( n56006 , n56005 , n32883 );
and ( n56007 , n52819 , n34154 );
or ( n56008 , n56006 , n56007 );
and ( n56009 , n56004 , n56008 );
and ( n56010 , n52819 , n34184 );
or ( n56011 , n56009 , n56010 );
and ( n56012 , n56003 , n56011 );
not ( n56013 , n34355 );
not ( n56014 , n34358 );
and ( n56015 , n56014 , n56011 );
and ( n56016 , n52845 , n34358 );
or ( n56017 , n56015 , n56016 );
and ( n56018 , n56013 , n56017 );
and ( n56019 , n52855 , n34355 );
or ( n56020 , n56018 , n56019 );
and ( n56021 , n56020 , n32968 );
or ( n56022 , n56012 , n56021 );
and ( n56023 , n56022 , n33370 );
and ( n56024 , n32883 , n35062 );
or ( n56025 , C0 , n55993 , n56002 , n56023 , n56024 );
buf ( n56026 , n56025 );
buf ( n56027 , n56026 );
not ( n56028 , n34150 );
and ( n56029 , n56028 , n32646 );
not ( n56030 , n34154 );
and ( n56031 , n56030 , n32646 );
and ( n56032 , n32655 , n34154 );
or ( n56033 , n56031 , n56032 );
and ( n56034 , n56033 , n34150 );
or ( n56035 , n56029 , n56034 );
and ( n56036 , n56035 , n33381 );
not ( n56037 , n34184 );
not ( n56038 , n34154 );
and ( n56039 , n56038 , n32646 );
not ( n56040 , n34287 );
and ( n56041 , n56040 , n34192 );
xor ( n56042 , n34294 , n34193 );
and ( n56043 , n56042 , n34287 );
or ( n56044 , n56041 , n56043 );
and ( n56045 , n56044 , n34154 );
or ( n56046 , n56039 , n56045 );
and ( n56047 , n56037 , n56046 );
and ( n56048 , n56044 , n34184 );
or ( n56049 , n56047 , n56048 );
and ( n56050 , n56049 , n33375 );
not ( n56051 , n32968 );
not ( n56052 , n34184 );
not ( n56053 , n34154 );
and ( n56054 , n56053 , n32646 );
and ( n56055 , n56044 , n34154 );
or ( n56056 , n56054 , n56055 );
and ( n56057 , n56052 , n56056 );
and ( n56058 , n56044 , n34184 );
or ( n56059 , n56057 , n56058 );
and ( n56060 , n56051 , n56059 );
not ( n56061 , n34355 );
not ( n56062 , n34358 );
and ( n56063 , n56062 , n56059 );
not ( n56064 , n34747 );
and ( n56065 , n56064 , n34415 );
xor ( n56066 , n34754 , n34625 );
and ( n56067 , n56066 , n34747 );
or ( n56068 , n56065 , n56067 );
and ( n56069 , n56068 , n34358 );
or ( n56070 , n56063 , n56069 );
and ( n56071 , n56061 , n56070 );
not ( n56072 , n35036 );
and ( n56073 , n56072 , n34826 );
xor ( n56074 , n35043 , n34918 );
and ( n56075 , n56074 , n35036 );
or ( n56076 , n56073 , n56075 );
and ( n56077 , n56076 , n34355 );
or ( n56078 , n56071 , n56077 );
and ( n56079 , n56078 , n32968 );
or ( n56080 , n56060 , n56079 );
and ( n56081 , n56080 , n33370 );
and ( n56082 , n32646 , n35062 );
or ( n56083 , C0 , n56036 , n56050 , n56081 , n56082 );
buf ( n56084 , n56083 );
buf ( n56085 , n56084 );
buf ( n56086 , n30987 );
buf ( n56087 , n31655 );
buf ( n56088 , n31655 );
buf ( n56089 , n31655 );
buf ( n56090 , n30987 );
not ( n56091 , n34150 );
and ( n56092 , n56091 , n32848 );
nor ( n56093 , n41389 , n34153 , n32538 , n32534 , n32530 );
not ( n56094 , n56093 );
and ( n56095 , n56094 , n32848 );
and ( n56096 , n32856 , n56093 );
or ( n56097 , n56095 , n56096 );
and ( n56098 , n56097 , n34150 );
or ( n56099 , n56092 , n56098 );
and ( n56100 , n56099 , n33381 );
nor ( n56101 , n41400 , n34171 , n34177 , n34183 , C0 );
not ( n56102 , n56101 );
not ( n56103 , n56093 );
and ( n56104 , n56103 , n32848 );
and ( n56105 , n48160 , n56093 );
or ( n56106 , n56104 , n56105 );
and ( n56107 , n56102 , n56106 );
and ( n56108 , n48160 , n56101 );
or ( n56109 , n56107 , n56108 );
and ( n56110 , n56109 , n33375 );
not ( n56111 , n32968 );
not ( n56112 , n56101 );
not ( n56113 , n56093 );
and ( n56114 , n56113 , n32848 );
and ( n56115 , n48160 , n56093 );
or ( n56116 , n56114 , n56115 );
and ( n56117 , n56112 , n56116 );
and ( n56118 , n48160 , n56101 );
or ( n56119 , n56117 , n56118 );
and ( n56120 , n56111 , n56119 );
nor ( n56121 , n41422 , n34334 , n34344 , n34354 , C0 );
not ( n56122 , n56121 );
nor ( n56123 , n41426 , n34357 , n34339 , n34349 , C0 );
not ( n56124 , n56123 );
and ( n56125 , n56124 , n56119 );
and ( n56126 , n48186 , n56123 );
or ( n56127 , n56125 , n56126 );
and ( n56128 , n56122 , n56127 );
and ( n56129 , n48196 , n56121 );
or ( n56130 , n56128 , n56129 );
and ( n56131 , n56130 , n32968 );
or ( n56132 , n56120 , n56131 );
and ( n56133 , n56132 , n33370 );
and ( n56134 , n32848 , n35062 );
or ( n56135 , C0 , n56100 , n56110 , n56133 , n56134 );
buf ( n56136 , n56135 );
buf ( n56137 , n56136 );
not ( n56138 , n34150 );
and ( n56139 , n56138 , n32685 );
nor ( n56140 , n41389 , n32542 , n32538 , n32534 , n32530 );
not ( n56141 , n56140 );
and ( n56142 , n56141 , n32685 );
and ( n56143 , n32689 , n56140 );
or ( n56144 , n56142 , n56143 );
and ( n56145 , n56144 , n34150 );
or ( n56146 , n56139 , n56145 );
and ( n56147 , n56146 , n33381 );
nor ( n56148 , n41400 , n34170 , n34177 , n34183 , C0 );
not ( n56149 , n56148 );
not ( n56150 , n56140 );
and ( n56151 , n56150 , n32685 );
and ( n56152 , n50682 , n56140 );
or ( n56153 , n56151 , n56152 );
and ( n56154 , n56149 , n56153 );
and ( n56155 , n50682 , n56148 );
or ( n56156 , n56154 , n56155 );
and ( n56157 , n56156 , n33375 );
not ( n56158 , n32968 );
not ( n56159 , n56148 );
not ( n56160 , n56140 );
and ( n56161 , n56160 , n32685 );
and ( n56162 , n50682 , n56140 );
or ( n56163 , n56161 , n56162 );
and ( n56164 , n56159 , n56163 );
and ( n56165 , n50682 , n56148 );
or ( n56166 , n56164 , n56165 );
and ( n56167 , n56158 , n56166 );
nor ( n56168 , n41422 , n34333 , n34344 , n34354 , C0 );
not ( n56169 , n56168 );
nor ( n56170 , n41426 , n34329 , n34339 , n34349 , C0 );
not ( n56171 , n56170 );
and ( n56172 , n56171 , n56166 );
and ( n56173 , n50706 , n56170 );
or ( n56174 , n56172 , n56173 );
and ( n56175 , n56169 , n56174 );
and ( n56176 , n50714 , n56168 );
or ( n56177 , n56175 , n56176 );
and ( n56178 , n56177 , n32968 );
or ( n56179 , n56167 , n56178 );
and ( n56180 , n56179 , n33370 );
and ( n56181 , n32685 , n35062 );
or ( n56182 , C0 , n56147 , n56157 , n56180 , n56181 );
buf ( n56183 , n56182 );
buf ( n56184 , n56183 );
buf ( n56185 , n30987 );
buf ( n56186 , n30987 );
buf ( n56187 , n31655 );
buf ( n56188 , n31655 );
buf ( n56189 , n30987 );
not ( n56190 , n34150 );
and ( n56191 , n56190 , n32813 );
nor ( n56192 , n32546 , n32542 , n41390 , n32534 , n32530 );
not ( n56193 , n56192 );
and ( n56194 , n56193 , n32813 );
and ( n56195 , n32823 , n56192 );
or ( n56196 , n56194 , n56195 );
and ( n56197 , n56196 , n34150 );
or ( n56198 , n56191 , n56197 );
and ( n56199 , n56198 , n33381 );
nor ( n56200 , n34165 , n34170 , n41401 , n34183 , C0 );
not ( n56201 , n56200 );
not ( n56202 , n56192 );
and ( n56203 , n56202 , n32813 );
and ( n56204 , n41464 , n56192 );
or ( n56205 , n56203 , n56204 );
and ( n56206 , n56201 , n56205 );
and ( n56207 , n41464 , n56200 );
or ( n56208 , n56206 , n56207 );
and ( n56209 , n56208 , n33375 );
not ( n56210 , n32968 );
not ( n56211 , n56200 );
not ( n56212 , n56192 );
and ( n56213 , n56212 , n32813 );
and ( n56214 , n41464 , n56192 );
or ( n56215 , n56213 , n56214 );
and ( n56216 , n56211 , n56215 );
and ( n56217 , n41464 , n56200 );
or ( n56218 , n56216 , n56217 );
and ( n56219 , n56210 , n56218 );
nor ( n56220 , n34325 , n34333 , n41423 , n34354 , C0 );
not ( n56221 , n56220 );
nor ( n56222 , n34321 , n34329 , n41427 , n34349 , C0 );
not ( n56223 , n56222 );
and ( n56224 , n56223 , n56218 );
and ( n56225 , n41490 , n56222 );
or ( n56226 , n56224 , n56225 );
and ( n56227 , n56221 , n56226 );
and ( n56228 , n41500 , n56220 );
or ( n56229 , n56227 , n56228 );
and ( n56230 , n56229 , n32968 );
or ( n56231 , n56219 , n56230 );
and ( n56232 , n56231 , n33370 );
and ( n56233 , n32813 , n35062 );
or ( n56234 , C0 , n56199 , n56209 , n56232 , n56233 );
buf ( n56235 , n56234 );
buf ( n56236 , n56235 );
not ( n56237 , n34150 );
and ( n56238 , n56237 , n32720 );
nor ( n56239 , n32546 , n32542 , n32538 , n32534 , n32530 );
not ( n56240 , n56239 );
and ( n56241 , n56240 , n32720 );
and ( n56242 , n32722 , n56239 );
or ( n56243 , n56241 , n56242 );
and ( n56244 , n56243 , n34150 );
or ( n56245 , n56238 , n56244 );
and ( n56246 , n56245 , n33381 );
nor ( n56247 , n34165 , n34170 , n34177 , n34183 , C0 );
not ( n56248 , n56247 );
not ( n56249 , n56239 );
and ( n56250 , n56249 , n32720 );
and ( n56251 , n42565 , n56239 );
or ( n56252 , n56250 , n56251 );
and ( n56253 , n56248 , n56252 );
and ( n56254 , n42565 , n56247 );
or ( n56255 , n56253 , n56254 );
and ( n56256 , n56255 , n33375 );
not ( n56257 , n32968 );
not ( n56258 , n56247 );
not ( n56259 , n56239 );
and ( n56260 , n56259 , n32720 );
and ( n56261 , n42565 , n56239 );
or ( n56262 , n56260 , n56261 );
and ( n56263 , n56258 , n56262 );
and ( n56264 , n42565 , n56247 );
or ( n56265 , n56263 , n56264 );
and ( n56266 , n56257 , n56265 );
nor ( n56267 , n34325 , n34333 , n34344 , n34354 , C0 );
not ( n56268 , n56267 );
nor ( n56269 , n34321 , n34329 , n34339 , n34349 , C0 );
not ( n56270 , n56269 );
and ( n56271 , n56270 , n56265 );
and ( n56272 , n42589 , n56269 );
or ( n56273 , n56271 , n56272 );
and ( n56274 , n56268 , n56273 );
and ( n56275 , n42597 , n56267 );
or ( n56276 , n56274 , n56275 );
and ( n56277 , n56276 , n32968 );
or ( n56278 , n56266 , n56277 );
and ( n56279 , n56278 , n33370 );
and ( n56280 , n32720 , n35062 );
or ( n56281 , C0 , n56246 , n56256 , n56279 , n56280 );
buf ( n56282 , n56281 );
buf ( n56283 , n56282 );
buf ( n56284 , n31655 );
not ( n56285 , n40163 );
and ( n56286 , n56285 , n32005 );
and ( n56287 , n31673 , n42237 , n31665 , n31661 , n42170 );
not ( n56288 , n56287 );
and ( n56289 , n56288 , n32005 );
and ( n56290 , n32147 , n56287 );
or ( n56291 , n56289 , n56290 );
and ( n56292 , n56291 , n40163 );
or ( n56293 , n56286 , n56292 );
and ( n56294 , n56293 , n32498 );
and ( n56295 , n40177 , n42246 , n40188 , n40194 , C1 );
not ( n56296 , n56295 );
not ( n56297 , n56287 );
and ( n56298 , n56297 , n32005 );
and ( n56299 , n49314 , n56287 );
or ( n56300 , n56298 , n56299 );
and ( n56301 , n56296 , n56300 );
and ( n56302 , n49314 , n56295 );
or ( n56303 , n56301 , n56302 );
and ( n56304 , n56303 , n32473 );
not ( n56305 , n32475 );
not ( n56306 , n56295 );
not ( n56307 , n56287 );
and ( n56308 , n56307 , n32005 );
and ( n56309 , n49314 , n56287 );
or ( n56310 , n56308 , n56309 );
and ( n56311 , n56306 , n56310 );
and ( n56312 , n49314 , n56295 );
or ( n56313 , n56311 , n56312 );
and ( n56314 , n56305 , n56313 );
and ( n56315 , n40417 , n42272 , n40435 , n40445 , C1 );
not ( n56316 , n56315 );
and ( n56317 , n40413 , n42275 , n40430 , n40440 , C1 );
not ( n56318 , n56317 );
and ( n56319 , n56318 , n56313 );
and ( n56320 , n49340 , n56317 );
or ( n56321 , n56319 , n56320 );
and ( n56322 , n56316 , n56321 );
and ( n56323 , n49348 , n56315 );
or ( n56324 , n56322 , n56323 );
and ( n56325 , n56324 , n32475 );
or ( n56326 , n56314 , n56325 );
and ( n56327 , n56326 , n32486 );
and ( n56328 , n32005 , n41278 );
or ( n56329 , C0 , n56294 , n56304 , n56327 , n56328 );
buf ( n56330 , n56329 );
buf ( n56331 , n56330 );
buf ( n56332 , n30987 );
buf ( n56333 , RI15b52e30_693);
and ( n56334 , n56333 , n31645 );
not ( n56335 , n45274 );
buf ( n56336 , RI15b535b0_709);
and ( n56337 , n56335 , n56336 );
not ( n56338 , n41809 );
and ( n56339 , n56338 , n41675 );
xor ( n56340 , n41815 , n41825 );
and ( n56341 , n56340 , n41809 );
or ( n56342 , n56339 , n56341 );
and ( n56343 , n56342 , n45274 );
or ( n56344 , n56337 , n56343 );
and ( n56345 , n56344 , n31373 );
not ( n56346 , n45280 );
and ( n56347 , n56346 , n56336 );
and ( n56348 , n56342 , n45280 );
or ( n56349 , n56347 , n56348 );
and ( n56350 , n56349 , n31468 );
and ( n56351 , n56336 , n45802 );
or ( n56352 , n56345 , n56350 , n56351 );
and ( n56353 , n56352 , n31557 );
and ( n56354 , n56336 , n45808 );
or ( n56355 , C0 , n56334 , n56353 , n56354 );
buf ( n56356 , n56355 );
buf ( n56357 , n56356 );
buf ( n56358 , n31655 );
buf ( n56359 , n30987 );
and ( n56360 , n33109 , n52224 );
and ( n56361 , n33107 , n56360 );
and ( n56362 , n33105 , n56361 );
xor ( n56363 , n33103 , n56362 );
and ( n56364 , n56363 , n33201 );
not ( n56365 , n41576 );
and ( n56366 , n56365 , n33103 );
and ( n56367 , n32857 , n52252 );
and ( n56368 , n32859 , n52254 );
and ( n56369 , n32861 , n52256 );
and ( n56370 , n32863 , n52258 );
and ( n56371 , n32865 , n52260 );
and ( n56372 , n32867 , n52262 );
and ( n56373 , n32869 , n52264 );
and ( n56374 , n32871 , n52266 );
and ( n56375 , n32873 , n52268 );
and ( n56376 , n32875 , n52270 );
and ( n56377 , n32877 , n52272 );
and ( n56378 , n32879 , n52274 );
and ( n56379 , n32881 , n52276 );
and ( n56380 , n32883 , n52278 );
and ( n56381 , n32885 , n52280 );
and ( n56382 , n32887 , n52282 );
or ( n56383 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 );
and ( n56384 , n56383 , n41576 );
or ( n56385 , n56366 , n56384 );
and ( n56386 , n56385 , n33189 );
and ( n56387 , n33103 , n41592 );
or ( n56388 , n56364 , n56386 , n56387 );
and ( n56389 , n56388 , n33208 );
and ( n56390 , n33103 , n39805 );
or ( n56391 , C0 , n56389 , n56390 );
buf ( n56392 , n56391 );
buf ( n56393 , n56392 );
not ( n56394 , n50828 );
not ( n56395 , n50834 );
and ( n56396 , n56395 , n40604 );
buf ( n56397 , RI15b53e20_727);
and ( n56398 , n56397 , n50834 );
or ( n56399 , n56396 , n56398 );
and ( n56400 , n56394 , n56399 );
buf ( n56401 , RI15b60288_1146);
and ( n56402 , n56401 , n50828 );
or ( n56403 , n56400 , n56402 );
buf ( n56404 , n56403 );
buf ( n56405 , n56404 );
buf ( n56406 , n30987 );
buf ( n56407 , n31655 );
buf ( n56408 , n30987 );
buf ( n56409 , n30987 );
buf ( n56410 , n31655 );
not ( n56411 , n34150 );
and ( n56412 , n56411 , n32777 );
nor ( n56413 , n41389 , n32542 , n41390 , n32534 , n32530 );
not ( n56414 , n56413 );
and ( n56415 , n56414 , n32777 );
and ( n56416 , n32789 , n56413 );
or ( n56417 , n56415 , n56416 );
and ( n56418 , n56417 , n34150 );
or ( n56419 , n56412 , n56418 );
and ( n56420 , n56419 , n33381 );
nor ( n56421 , n41400 , n34170 , n41401 , n34183 , C0 );
not ( n56422 , n56421 );
not ( n56423 , n56413 );
and ( n56424 , n56423 , n32777 );
and ( n56425 , n34301 , n56413 );
or ( n56426 , n56424 , n56425 );
and ( n56427 , n56422 , n56426 );
and ( n56428 , n34301 , n56421 );
or ( n56429 , n56427 , n56428 );
and ( n56430 , n56429 , n33375 );
not ( n56431 , n32968 );
not ( n56432 , n56421 );
not ( n56433 , n56413 );
and ( n56434 , n56433 , n32777 );
and ( n56435 , n34301 , n56413 );
or ( n56436 , n56434 , n56435 );
and ( n56437 , n56432 , n56436 );
and ( n56438 , n34301 , n56421 );
or ( n56439 , n56437 , n56438 );
and ( n56440 , n56431 , n56439 );
nor ( n56441 , n41422 , n34333 , n41423 , n34354 , C0 );
not ( n56442 , n56441 );
nor ( n56443 , n41426 , n34329 , n41427 , n34349 , C0 );
not ( n56444 , n56443 );
and ( n56445 , n56444 , n56439 );
and ( n56446 , n34761 , n56443 );
or ( n56447 , n56445 , n56446 );
and ( n56448 , n56442 , n56447 );
and ( n56449 , n35050 , n56441 );
or ( n56450 , n56448 , n56449 );
and ( n56451 , n56450 , n32968 );
or ( n56452 , n56440 , n56451 );
and ( n56453 , n56452 , n33370 );
and ( n56454 , n32777 , n35062 );
or ( n56455 , C0 , n56420 , n56430 , n56453 , n56454 );
buf ( n56456 , n56455 );
buf ( n56457 , n56456 );
buf ( n56458 , n31655 );
not ( n56459 , n34150 );
and ( n56460 , n56459 , n32546 );
and ( n56461 , n34165 , n34150 );
or ( n56462 , n56460 , n56461 );
and ( n56463 , n56462 , n33381 );
buf ( n56464 , RI15b3fc18_40);
not ( n56465 , n56464 );
and ( n56466 , n56465 , n32531 );
buf ( n56467 , n56466 );
not ( n56468 , n56467 );
not ( n56469 , n56464 );
and ( n56470 , n56469 , n32539 );
buf ( n56471 , RI15b44970_205);
not ( n56472 , n56471 );
buf ( n56473 , RI15b448f8_204);
not ( n56474 , n56473 );
not ( n56475 , n48582 );
not ( n56476 , n48583 );
not ( n56477 , n48584 );
not ( n56478 , n48585 );
not ( n56479 , n48586 );
not ( n56480 , n48587 );
not ( n56481 , n48588 );
not ( n56482 , n48589 );
not ( n56483 , n48590 );
not ( n56484 , n48591 );
not ( n56485 , n48592 );
not ( n56486 , n48593 );
not ( n56487 , n48594 );
not ( n56488 , n48595 );
not ( n56489 , n48596 );
not ( n56490 , n48597 );
not ( n56491 , n48598 );
not ( n56492 , n48599 );
not ( n56493 , n48600 );
not ( n56494 , n48601 );
not ( n56495 , n48602 );
not ( n56496 , n48603 );
not ( n56497 , n48604 );
not ( n56498 , n48605 );
not ( n56499 , n48606 );
not ( n56500 , n48607 );
not ( n56501 , n48608 );
not ( n56502 , n48609 );
not ( n56503 , n48610 );
not ( n56504 , n48668 );
and ( n56505 , n56503 , n56504 );
and ( n56506 , n56502 , n56505 );
and ( n56507 , n56501 , n56506 );
and ( n56508 , n56500 , n56507 );
and ( n56509 , n56499 , n56508 );
and ( n56510 , n56498 , n56509 );
and ( n56511 , n56497 , n56510 );
and ( n56512 , n56496 , n56511 );
and ( n56513 , n56495 , n56512 );
and ( n56514 , n56494 , n56513 );
and ( n56515 , n56493 , n56514 );
and ( n56516 , n56492 , n56515 );
and ( n56517 , n56491 , n56516 );
and ( n56518 , n56490 , n56517 );
and ( n56519 , n56489 , n56518 );
and ( n56520 , n56488 , n56519 );
and ( n56521 , n56487 , n56520 );
and ( n56522 , n56486 , n56521 );
and ( n56523 , n56485 , n56522 );
and ( n56524 , n56484 , n56523 );
and ( n56525 , n56483 , n56524 );
and ( n56526 , n56482 , n56525 );
and ( n56527 , n56481 , n56526 );
and ( n56528 , n56480 , n56527 );
and ( n56529 , n56479 , n56528 );
and ( n56530 , n56478 , n56529 );
and ( n56531 , n56477 , n56530 );
and ( n56532 , n56476 , n56531 );
and ( n56533 , n56475 , n56532 );
and ( n56534 , n56474 , n56533 );
xor ( n56535 , n56472 , n56534 );
buf ( n56536 , n56471 );
and ( n56537 , n56535 , n56536 );
buf ( n56538 , n56537 );
not ( n56539 , n56538 );
not ( n56540 , n56471 );
and ( n56541 , n56540 , n48610 );
xor ( n56542 , n56503 , n56504 );
and ( n56543 , n56542 , n56471 );
or ( n56544 , n56541 , n56543 );
and ( n56545 , n56539 , n56544 );
not ( n56546 , n56544 );
buf ( n56547 , n48668 );
not ( n56548 , n56547 );
xor ( n56549 , n56546 , n56548 );
and ( n56550 , n56549 , n56538 );
or ( n56551 , n56545 , n56550 );
not ( n56552 , n56551 );
buf ( n56553 , n56552 );
buf ( n56554 , n56553 );
not ( n56555 , n56554 );
xor ( n56556 , n56555 , n56538 );
buf ( n56557 , n56547 );
not ( n56558 , n56557 );
buf ( n56559 , n56558 );
not ( n56560 , n56559 );
xor ( n56561 , n56560 , n56538 );
and ( n56562 , n56561 , n56538 );
and ( n56563 , n56556 , n56562 );
buf ( n56564 , n56563 );
or ( n56565 , n56560 , n56555 );
buf ( n56566 , n56565 );
buf ( n56567 , n56566 );
and ( n56568 , n56567 , n56538 );
and ( n56569 , n56564 , n56568 );
buf ( n56570 , n56569 );
not ( n56571 , n56568 );
and ( n56572 , n56571 , n56555 );
xor ( n56573 , n56556 , n56562 );
and ( n56574 , n56573 , n56568 );
or ( n56575 , n56572 , n56574 );
not ( n56576 , n56568 );
and ( n56577 , n56576 , n56560 );
xor ( n56578 , n56561 , n56538 );
and ( n56579 , n56578 , n56568 );
or ( n56580 , n56577 , n56579 );
and ( n56581 , n56575 , n56580 );
xor ( n56582 , n56570 , n56581 );
buf ( n56583 , n56582 );
buf ( n56584 , n56583 );
not ( n56585 , n56584 );
buf ( n56586 , n56585 );
buf ( n56587 , n56586 );
not ( n56588 , n56587 );
buf ( n56589 , n56588 );
buf ( n56590 , n56589 );
buf ( n56591 , n56547 );
not ( n56592 , n56591 );
buf ( n56593 , n56592 );
not ( n56594 , n56593 );
buf ( n56595 , n56594 );
buf ( n56596 , n56595 );
and ( n56597 , n56596 , n56538 );
not ( n56598 , n56597 );
and ( n56599 , n56598 , n56594 );
xor ( n56600 , n56594 , n56538 );
xor ( n56601 , n56600 , n56538 );
and ( n56602 , n56601 , n56597 );
or ( n56603 , n56599 , n56602 );
not ( n56604 , n56603 );
not ( n56605 , n56604 );
and ( n56606 , n56590 , n56605 );
buf ( n56607 , n56606 );
and ( n56608 , n56607 , n56464 );
or ( n56609 , n56470 , n56608 );
not ( n56610 , n56609 );
not ( n56611 , n56464 );
and ( n56612 , n56611 , n32535 );
and ( n56613 , n56570 , n56581 );
buf ( n56614 , n56613 );
buf ( n56615 , n56614 );
not ( n56616 , n56615 );
buf ( n56617 , n56616 );
buf ( n56618 , n56617 );
not ( n56619 , n56618 );
buf ( n56620 , n56619 );
buf ( n56621 , n56620 );
and ( n56622 , n56621 , n56605 );
buf ( n56623 , n56622 );
and ( n56624 , n56623 , n56464 );
or ( n56625 , n56612 , n56624 );
not ( n56626 , n56625 );
buf ( n56627 , n56467 );
buf ( n56628 , n56467 );
buf ( n56629 , n56467 );
buf ( n56630 , n56467 );
buf ( n56631 , n56467 );
buf ( n56632 , n56467 );
buf ( n56633 , n56467 );
buf ( n56634 , n56467 );
buf ( n56635 , n56467 );
buf ( n56636 , n56467 );
buf ( n56637 , n56467 );
buf ( n56638 , n56467 );
buf ( n56639 , n56467 );
buf ( n56640 , n56467 );
buf ( n56641 , n56467 );
buf ( n56642 , n56467 );
buf ( n56643 , n56467 );
buf ( n56644 , n56467 );
buf ( n56645 , n56467 );
buf ( n56646 , n56467 );
buf ( n56647 , n56467 );
buf ( n56648 , n56467 );
buf ( n56649 , n56467 );
buf ( n56650 , n56467 );
buf ( n56651 , n56467 );
buf ( n56652 , n56467 );
not ( n56653 , n56464 );
and ( n56654 , n56653 , n32547 );
not ( n56655 , n56605 );
buf ( n56656 , n56655 );
not ( n56657 , n56580 );
buf ( n56658 , n56657 );
not ( n56659 , n56658 );
buf ( n56660 , n56659 );
not ( n56661 , n56660 );
buf ( n56662 , n56661 );
buf ( n56663 , n56662 );
and ( n56664 , n56663 , n56605 );
or ( n56665 , n56656 , n56664 );
and ( n56666 , n56665 , n56464 );
or ( n56667 , n56654 , n56666 );
not ( n56668 , n56667 );
not ( n56669 , n56464 );
and ( n56670 , n56669 , n32543 );
xor ( n56671 , n56575 , n56580 );
buf ( n56672 , n56671 );
buf ( n56673 , n56672 );
not ( n56674 , n56673 );
buf ( n56675 , n56674 );
buf ( n56676 , n56675 );
not ( n56677 , n56676 );
buf ( n56678 , n56677 );
buf ( n56679 , n56678 );
and ( n56680 , n56679 , n56605 );
buf ( n56681 , n56680 );
and ( n56682 , n56681 , n56464 );
or ( n56683 , n56670 , n56682 );
not ( n56684 , n56683 );
and ( n56685 , n56668 , n56684 );
or ( n56686 , n56610 , n56626 , n56467 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56685 );
nand ( n56687 , n56468 , n56686 );
not ( n56688 , n56687 );
not ( n56689 , n56464 );
and ( n56690 , n56689 , n32546 );
buf ( n56691 , n56464 );
or ( n56692 , n56690 , n56691 );
and ( n56693 , n56688 , n56692 );
buf ( n56694 , n56693 );
and ( n56695 , n56694 , n33379 );
and ( n56696 , n34321 , n33375 );
buf ( n56697 , n34321 );
and ( n56698 , n56697 , n33370 );
or ( n56699 , n35060 , n32528 );
and ( n56700 , n32546 , n56699 );
or ( n56701 , C0 , n56463 , n56695 , n56696 , n56698 , n56700 );
buf ( n56702 , n56701 );
buf ( n56703 , n56702 );
buf ( n56704 , n31655 );
buf ( n56705 , n30987 );
not ( n56706 , n34150 );
and ( n56707 , n56706 , n32603 );
and ( n56708 , n32546 , n32542 , n32538 , n32534 , n41391 );
not ( n56709 , n56708 );
and ( n56710 , n56709 , n32603 );
and ( n56711 , n32655 , n56708 );
or ( n56712 , n56710 , n56711 );
and ( n56713 , n56712 , n34150 );
or ( n56714 , n56707 , n56713 );
and ( n56715 , n56714 , n33381 );
and ( n56716 , n34165 , n34170 , n34177 , n34183 , C1 );
not ( n56717 , n56716 );
not ( n56718 , n56708 );
and ( n56719 , n56718 , n32603 );
and ( n56720 , n56044 , n56708 );
or ( n56721 , n56719 , n56720 );
and ( n56722 , n56717 , n56721 );
and ( n56723 , n56044 , n56716 );
or ( n56724 , n56722 , n56723 );
and ( n56725 , n56724 , n33375 );
not ( n56726 , n32968 );
not ( n56727 , n56716 );
not ( n56728 , n56708 );
and ( n56729 , n56728 , n32603 );
and ( n56730 , n56044 , n56708 );
or ( n56731 , n56729 , n56730 );
and ( n56732 , n56727 , n56731 );
and ( n56733 , n56044 , n56716 );
or ( n56734 , n56732 , n56733 );
and ( n56735 , n56726 , n56734 );
and ( n56736 , n34325 , n34333 , n34344 , n34354 , C1 );
not ( n56737 , n56736 );
and ( n56738 , n34321 , n34329 , n34339 , n34349 , C1 );
not ( n56739 , n56738 );
and ( n56740 , n56739 , n56734 );
and ( n56741 , n56068 , n56738 );
or ( n56742 , n56740 , n56741 );
and ( n56743 , n56737 , n56742 );
and ( n56744 , n56076 , n56736 );
or ( n56745 , n56743 , n56744 );
and ( n56746 , n56745 , n32968 );
or ( n56747 , n56735 , n56746 );
and ( n56748 , n56747 , n33370 );
and ( n56749 , n32603 , n35062 );
or ( n56750 , C0 , n56715 , n56725 , n56748 , n56749 );
buf ( n56751 , n56750 );
buf ( n56752 , n56751 );
buf ( n56753 , n30987 );
buf ( n56754 , n31655 );
and ( n56755 , n33762 , n48455 );
not ( n56756 , n48457 );
and ( n56757 , n56756 , n33427 );
and ( n56758 , n33762 , n48457 );
or ( n56759 , n56757 , n56758 );
and ( n56760 , n56759 , n31373 );
not ( n56761 , n44807 );
and ( n56762 , n56761 , n33427 );
and ( n56763 , n33762 , n44807 );
or ( n56764 , n56762 , n56763 );
and ( n56765 , n56764 , n31408 );
not ( n56766 , n48468 );
and ( n56767 , n56766 , n33427 );
and ( n56768 , n33762 , n48468 );
or ( n56769 , n56767 , n56768 );
and ( n56770 , n56769 , n31468 );
not ( n56771 , n44817 );
and ( n56772 , n56771 , n33427 );
and ( n56773 , n33762 , n44817 );
or ( n56774 , n56772 , n56773 );
and ( n56775 , n56774 , n31521 );
not ( n56776 , n39979 );
and ( n56777 , n56776 , n33427 );
and ( n56778 , n33469 , n39979 );
or ( n56779 , n56777 , n56778 );
and ( n56780 , n56779 , n31538 );
not ( n56781 , n45059 );
and ( n56782 , n56781 , n33427 );
and ( n56783 , n33469 , n45059 );
or ( n56784 , n56782 , n56783 );
and ( n56785 , n56784 , n31536 );
not ( n56786 , n33419 );
and ( n56787 , n56786 , n33427 );
xor ( n56788 , n33469 , n33696 );
and ( n56789 , n56788 , n33419 );
or ( n56790 , n56787 , n56789 );
and ( n56791 , n56790 , n31529 );
not ( n56792 , n33734 );
and ( n56793 , n56792 , n33427 );
not ( n56794 , n33533 );
xor ( n56795 , n33762 , n33814 );
and ( n56796 , n56794 , n56795 );
xnor ( n56797 , n33847 , n33916 );
and ( n56798 , n56797 , n33533 );
or ( n56799 , n56796 , n56798 );
and ( n56800 , n56799 , n33734 );
or ( n56801 , n56793 , n56800 );
and ( n56802 , n56801 , n31527 );
and ( n56803 , n33847 , n48513 );
or ( n56804 , n56755 , n56760 , n56765 , n56770 , n56775 , n56780 , n56785 , n56791 , n56802 , n56803 );
and ( n56805 , n56804 , n31557 );
and ( n56806 , n33999 , n33973 );
and ( n56807 , n33427 , n48524 );
or ( n56808 , C0 , n56805 , n56806 , n56807 );
buf ( n56809 , n56808 );
buf ( n56810 , n56809 );
buf ( n56811 , n31655 );
buf ( n56812 , RI15b608a0_1159);
not ( n56813 , n56812 );
and ( n56814 , n56813 , n48531 );
buf ( n56815 , n39350 );
or ( n56816 , n39349 , n39352 );
or ( n56817 , n56816 , n39354 );
or ( n56818 , n56817 , n39356 );
or ( n56819 , n56818 , n39358 );
and ( n56820 , n50818 , n56819 );
or ( n56821 , n56814 , n56815 , n56820 );
buf ( n56822 , n56821 );
buf ( n56823 , n56822 );
buf ( n56824 , n30987 );
not ( n56825 , n35542 );
and ( n56826 , n56825 , n41854 );
buf ( n56827 , RI15b45780_235);
and ( n56828 , n56827 , n35542 );
or ( n56829 , n56826 , n56828 );
buf ( n56830 , n56829 );
buf ( n56831 , n56830 );
buf ( n56832 , n30987 );
buf ( n56833 , n30987 );
not ( n56834 , n34150 );
and ( n56835 , n56834 , n32741 );
nor ( n56836 , n32546 , n34153 , n41390 , n32534 , n32530 );
not ( n56837 , n56836 );
and ( n56838 , n56837 , n32741 );
and ( n56839 , n32755 , n56836 );
or ( n56840 , n56838 , n56839 );
and ( n56841 , n56840 , n34150 );
or ( n56842 , n56835 , n56841 );
and ( n56843 , n56842 , n33381 );
nor ( n56844 , n34165 , n34171 , n41401 , n34183 , C0 );
not ( n56845 , n56844 );
not ( n56846 , n56836 );
and ( n56847 , n56846 , n32741 );
and ( n56848 , n35083 , n56836 );
or ( n56849 , n56847 , n56848 );
and ( n56850 , n56845 , n56849 );
and ( n56851 , n35083 , n56844 );
or ( n56852 , n56850 , n56851 );
and ( n56853 , n56852 , n33375 );
not ( n56854 , n32968 );
not ( n56855 , n56844 );
not ( n56856 , n56836 );
and ( n56857 , n56856 , n32741 );
and ( n56858 , n35083 , n56836 );
or ( n56859 , n56857 , n56858 );
and ( n56860 , n56855 , n56859 );
and ( n56861 , n35083 , n56844 );
or ( n56862 , n56860 , n56861 );
and ( n56863 , n56854 , n56862 );
nor ( n56864 , n34325 , n34334 , n41423 , n34354 , C0 );
not ( n56865 , n56864 );
nor ( n56866 , n34321 , n34357 , n41427 , n34349 , C0 );
not ( n56867 , n56866 );
and ( n56868 , n56867 , n56862 );
and ( n56869 , n35107 , n56866 );
or ( n56870 , n56868 , n56869 );
and ( n56871 , n56865 , n56870 );
and ( n56872 , n35115 , n56864 );
or ( n56873 , n56871 , n56872 );
and ( n56874 , n56873 , n32968 );
or ( n56875 , n56863 , n56874 );
and ( n56876 , n56875 , n33370 );
and ( n56877 , n32741 , n35062 );
or ( n56878 , C0 , n56843 , n56853 , n56876 , n56877 );
buf ( n56879 , n56878 );
buf ( n56880 , n56879 );
buf ( n56881 , n31655 );
buf ( n56882 , n31655 );
buf ( n56883 , n31655 );
buf ( n56884 , n40217 );
not ( n56885 , n35297 );
and ( n56886 , n56885 , n32433 );
not ( n56887 , n47331 );
and ( n56888 , n56887 , n35297 );
buf ( n56889 , n32066 );
and ( n56890 , n56889 , n47331 );
or ( n56891 , n56888 , n56890 );
and ( n56892 , n56891 , n32413 );
and ( n56893 , n35297 , n47402 );
or ( n56894 , n56886 , n56892 , n56893 );
and ( n56895 , n56894 , n32456 );
and ( n56896 , n35297 , n47409 );
or ( n56897 , C0 , n56895 , n56896 );
buf ( n56898 , n56897 );
buf ( n56899 , n56898 );
buf ( n56900 , n30987 );
buf ( n56901 , n31655 );
not ( n56902 , n46356 );
and ( n56903 , n56902 , n31123 );
nor ( n56904 , n31025 , n31021 , n48213 , n31013 , n31009 );
not ( n56905 , n56904 );
and ( n56906 , n56905 , n31123 );
and ( n56907 , n31138 , n56904 );
or ( n56908 , n56906 , n56907 );
and ( n56909 , n56908 , n46356 );
or ( n56910 , n56903 , n56909 );
and ( n56911 , n56910 , n31649 );
nor ( n56912 , n46373 , n46379 , n48222 , n46392 , C0 );
not ( n56913 , n56912 );
not ( n56914 , n56904 );
and ( n56915 , n56914 , n31123 );
not ( n56916 , n46487 );
and ( n56917 , n56916 , n46400 );
xor ( n56918 , n46491 , n41881 );
and ( n56919 , n56918 , n46487 );
or ( n56920 , n56917 , n56919 );
and ( n56921 , n56920 , n56904 );
or ( n56922 , n56915 , n56921 );
and ( n56923 , n56913 , n56922 );
and ( n56924 , n56920 , n56912 );
or ( n56925 , n56923 , n56924 );
and ( n56926 , n56925 , n31643 );
not ( n56927 , n31452 );
not ( n56928 , n56912 );
not ( n56929 , n56904 );
and ( n56930 , n56929 , n31123 );
and ( n56931 , n56920 , n56904 );
or ( n56932 , n56930 , n56931 );
and ( n56933 , n56928 , n56932 );
and ( n56934 , n56920 , n56912 );
or ( n56935 , n56933 , n56934 );
and ( n56936 , n56927 , n56935 );
nor ( n56937 , n46519 , n46528 , n48243 , n46549 , C0 );
not ( n56938 , n56937 );
nor ( n56939 , n46515 , n46524 , n48246 , n46544 , C0 );
not ( n56940 , n56939 );
and ( n56941 , n56940 , n56935 );
not ( n56942 , n46976 );
and ( n56943 , n56942 , n46606 );
xor ( n56944 , n46980 , n46854 );
and ( n56945 , n56944 , n46976 );
or ( n56946 , n56943 , n56945 );
and ( n56947 , n56946 , n56939 );
or ( n56948 , n56941 , n56947 );
and ( n56949 , n56938 , n56948 );
not ( n56950 , n47259 );
and ( n56951 , n56950 , n47049 );
xor ( n56952 , n47263 , n47141 );
and ( n56953 , n56952 , n47259 );
or ( n56954 , n56951 , n56953 );
and ( n56955 , n56954 , n56937 );
or ( n56956 , n56949 , n56955 );
and ( n56957 , n56956 , n31452 );
or ( n56958 , n56936 , n56957 );
and ( n56959 , n56958 , n31638 );
and ( n56960 , n31123 , n47277 );
or ( n56961 , C0 , n56911 , n56926 , n56959 , n56960 );
buf ( n56962 , n56961 );
buf ( n56963 , n56962 );
not ( n56964 , n31437 );
and ( n56965 , n56964 , n51843 );
not ( n56966 , n41809 );
and ( n56967 , n56966 , n41636 );
xor ( n56968 , n41818 , n41822 );
and ( n56969 , n56968 , n41809 );
or ( n56970 , n56967 , n56969 );
and ( n56971 , n56970 , n31437 );
or ( n56972 , n56965 , n56971 );
and ( n56973 , n56972 , n31468 );
not ( n56974 , n41837 );
and ( n56975 , n56974 , n51843 );
and ( n56976 , n51849 , n41837 );
or ( n56977 , n56975 , n56976 );
and ( n56978 , n56977 , n31521 );
and ( n56979 , n51843 , n42158 );
or ( n56980 , n56973 , n56978 , n56979 );
and ( n56981 , n56980 , n31557 );
and ( n56982 , n51843 , n40154 );
or ( n56983 , C0 , n56981 , n56982 );
buf ( n56984 , n56983 );
buf ( n56985 , n56984 );
not ( n56986 , n40163 );
and ( n56987 , n56986 , n31896 );
and ( n56988 , n31673 , n31669 , n31665 , n31661 , n42170 );
not ( n56989 , n56988 );
and ( n56990 , n56989 , n31896 );
and ( n56991 , n32200 , n56988 );
or ( n56992 , n56990 , n56991 );
and ( n56993 , n56992 , n40163 );
or ( n56994 , n56987 , n56993 );
and ( n56995 , n56994 , n32498 );
and ( n56996 , n40177 , n40182 , n40188 , n40194 , C1 );
not ( n56997 , n56996 );
not ( n56998 , n56988 );
and ( n56999 , n56998 , n31896 );
and ( n57000 , n53243 , n56988 );
or ( n57001 , n56999 , n57000 );
and ( n57002 , n56997 , n57001 );
and ( n57003 , n53243 , n56996 );
or ( n57004 , n57002 , n57003 );
and ( n57005 , n57004 , n32473 );
not ( n57006 , n32475 );
not ( n57007 , n56996 );
not ( n57008 , n56988 );
and ( n57009 , n57008 , n31896 );
and ( n57010 , n53243 , n56988 );
or ( n57011 , n57009 , n57010 );
and ( n57012 , n57007 , n57011 );
and ( n57013 , n53243 , n56996 );
or ( n57014 , n57012 , n57013 );
and ( n57015 , n57006 , n57014 );
and ( n57016 , n40417 , n40425 , n40435 , n40445 , C1 );
not ( n57017 , n57016 );
and ( n57018 , n40413 , n40421 , n40430 , n40440 , C1 );
not ( n57019 , n57018 );
and ( n57020 , n57019 , n57014 );
and ( n57021 , n53269 , n57018 );
or ( n57022 , n57020 , n57021 );
and ( n57023 , n57017 , n57022 );
and ( n57024 , n53277 , n57016 );
or ( n57025 , n57023 , n57024 );
and ( n57026 , n57025 , n32475 );
or ( n57027 , n57015 , n57026 );
and ( n57028 , n57027 , n32486 );
and ( n57029 , n31896 , n41278 );
or ( n57030 , C0 , n56995 , n57005 , n57028 , n57029 );
buf ( n57031 , n57030 );
buf ( n57032 , n57031 );
buf ( n57033 , n31655 );
buf ( n57034 , n30987 );
buf ( n57035 , n40212 );
not ( n57036 , n34150 );
and ( n57037 , n57036 , n32706 );
nor ( n57038 , n41389 , n34153 , n41390 , n32534 , n32530 );
not ( n57039 , n57038 );
and ( n57040 , n57039 , n32706 );
and ( n57041 , n32722 , n57038 );
or ( n57042 , n57040 , n57041 );
and ( n57043 , n57042 , n34150 );
or ( n57044 , n57037 , n57043 );
and ( n57045 , n57044 , n33381 );
nor ( n57046 , n41400 , n34171 , n41401 , n34183 , C0 );
not ( n57047 , n57046 );
not ( n57048 , n57038 );
and ( n57049 , n57048 , n32706 );
and ( n57050 , n42565 , n57038 );
or ( n57051 , n57049 , n57050 );
and ( n57052 , n57047 , n57051 );
and ( n57053 , n42565 , n57046 );
or ( n57054 , n57052 , n57053 );
and ( n57055 , n57054 , n33375 );
not ( n57056 , n32968 );
not ( n57057 , n57046 );
not ( n57058 , n57038 );
and ( n57059 , n57058 , n32706 );
and ( n57060 , n42565 , n57038 );
or ( n57061 , n57059 , n57060 );
and ( n57062 , n57057 , n57061 );
and ( n57063 , n42565 , n57046 );
or ( n57064 , n57062 , n57063 );
and ( n57065 , n57056 , n57064 );
nor ( n57066 , n41422 , n34334 , n41423 , n34354 , C0 );
not ( n57067 , n57066 );
nor ( n57068 , n41426 , n34357 , n41427 , n34349 , C0 );
not ( n57069 , n57068 );
and ( n57070 , n57069 , n57064 );
and ( n57071 , n42589 , n57068 );
or ( n57072 , n57070 , n57071 );
and ( n57073 , n57067 , n57072 );
and ( n57074 , n42597 , n57066 );
or ( n57075 , n57073 , n57074 );
and ( n57076 , n57075 , n32968 );
or ( n57077 , n57065 , n57076 );
and ( n57078 , n57077 , n33370 );
and ( n57079 , n32706 , n35062 );
or ( n57080 , C0 , n57045 , n57055 , n57078 , n57079 );
buf ( n57081 , n57080 );
buf ( n57082 , n57081 );
buf ( n57083 , n30987 );
buf ( n57084 , n31655 );
buf ( n57085 , n31655 );
buf ( n57086 , n30987 );
buf ( n57087 , n30987 );
buf ( n57088 , n31655 );
not ( n57089 , n31437 );
buf ( n57090 , RI15b525c0_675);
and ( n57091 , n57089 , n57090 );
not ( n57092 , n45766 );
and ( n57093 , n57092 , n45558 );
xor ( n57094 , n45776 , n45780 );
and ( n57095 , n57094 , n45766 );
or ( n57096 , n57093 , n57095 );
and ( n57097 , n57096 , n31437 );
or ( n57098 , n57091 , n57097 );
and ( n57099 , n57098 , n31468 );
not ( n57100 , n44817 );
and ( n57101 , n57100 , n57090 );
not ( n57102 , n44994 );
and ( n57103 , n57102 , n44846 );
xor ( n57104 , n45008 , n45012 );
and ( n57105 , n57104 , n44994 );
or ( n57106 , n57103 , n57105 );
and ( n57107 , n57106 , n44817 );
or ( n57108 , n57101 , n57107 );
and ( n57109 , n57108 , n31521 );
and ( n57110 , n57090 , n42158 );
or ( n57111 , n57099 , n57109 , n57110 );
and ( n57112 , n57111 , n31557 );
and ( n57113 , n57090 , n40154 );
or ( n57114 , C0 , n57112 , n57113 );
buf ( n57115 , n57114 );
buf ( n57116 , n57115 );
and ( n57117 , n47668 , n50275 );
not ( n57118 , n50278 );
and ( n57119 , n57118 , n47581 );
and ( n57120 , n47668 , n50278 );
or ( n57121 , n57119 , n57120 );
and ( n57122 , n57121 , n32421 );
not ( n57123 , n50002 );
and ( n57124 , n57123 , n47581 );
and ( n57125 , n47668 , n50002 );
or ( n57126 , n57124 , n57125 );
and ( n57127 , n57126 , n32419 );
not ( n57128 , n50289 );
and ( n57129 , n57128 , n47581 );
and ( n57130 , n47668 , n50289 );
or ( n57131 , n57129 , n57130 );
and ( n57132 , n57131 , n32417 );
not ( n57133 , n50008 );
and ( n57134 , n57133 , n47581 );
and ( n57135 , n47668 , n50008 );
or ( n57136 , n57134 , n57135 );
and ( n57137 , n57136 , n32415 );
not ( n57138 , n47331 );
and ( n57139 , n57138 , n47581 );
and ( n57140 , n47613 , n47331 );
or ( n57141 , n57139 , n57140 );
and ( n57142 , n57141 , n32413 );
not ( n57143 , n50067 );
and ( n57144 , n57143 , n47581 );
and ( n57145 , n47613 , n50067 );
or ( n57146 , n57144 , n57145 );
and ( n57147 , n57146 , n32411 );
not ( n57148 , n31728 );
and ( n57149 , n57148 , n47581 );
and ( n57150 , n54874 , n31728 );
or ( n57151 , n57149 , n57150 );
and ( n57152 , n57151 , n32253 );
not ( n57153 , n32283 );
and ( n57154 , n57153 , n47581 );
and ( n57155 , n54885 , n32283 );
or ( n57156 , n57154 , n57155 );
and ( n57157 , n57156 , n32398 );
and ( n57158 , n47718 , n50334 );
or ( n57159 , n57117 , n57122 , n57127 , n57132 , n57137 , n57142 , n57147 , n57152 , n57157 , n57158 );
and ( n57160 , n57159 , n32456 );
and ( n57161 , n37569 , n32489 );
and ( n57162 , n47581 , n50345 );
or ( n57163 , C0 , n57160 , n57161 , n57162 );
buf ( n57164 , n57163 );
buf ( n57165 , n57164 );
buf ( n57166 , n31655 );
buf ( n57167 , RI15b47418_296);
buf ( n57168 , n57167 );
not ( n57169 , n34150 );
and ( n57170 , n57169 , n32671 );
not ( n57171 , n41392 );
and ( n57172 , n57171 , n32671 );
and ( n57173 , n32689 , n41392 );
or ( n57174 , n57172 , n57173 );
and ( n57175 , n57174 , n34150 );
or ( n57176 , n57170 , n57175 );
and ( n57177 , n57176 , n33381 );
not ( n57178 , n41402 );
not ( n57179 , n41392 );
and ( n57180 , n57179 , n32671 );
and ( n57181 , n50682 , n41392 );
or ( n57182 , n57180 , n57181 );
and ( n57183 , n57178 , n57182 );
and ( n57184 , n50682 , n41402 );
or ( n57185 , n57183 , n57184 );
and ( n57186 , n57185 , n33375 );
not ( n57187 , n32968 );
not ( n57188 , n41402 );
not ( n57189 , n41392 );
and ( n57190 , n57189 , n32671 );
and ( n57191 , n50682 , n41392 );
or ( n57192 , n57190 , n57191 );
and ( n57193 , n57188 , n57192 );
and ( n57194 , n50682 , n41402 );
or ( n57195 , n57193 , n57194 );
and ( n57196 , n57187 , n57195 );
not ( n57197 , n41424 );
not ( n57198 , n41428 );
and ( n57199 , n57198 , n57195 );
and ( n57200 , n50706 , n41428 );
or ( n57201 , n57199 , n57200 );
and ( n57202 , n57197 , n57201 );
and ( n57203 , n50714 , n41424 );
or ( n57204 , n57202 , n57203 );
and ( n57205 , n57204 , n32968 );
or ( n57206 , n57196 , n57205 );
and ( n57207 , n57206 , n33370 );
and ( n57208 , n32671 , n35062 );
or ( n57209 , C0 , n57177 , n57186 , n57207 , n57208 );
buf ( n57210 , n57209 );
buf ( n57211 , n57210 );
buf ( n57212 , n31655 );
buf ( n57213 , n30987 );
buf ( n57214 , n30987 );
buf ( n57215 , n30987 );
xor ( n57216 , n31505 , n39924 );
and ( n57217 , n57216 , n31550 );
not ( n57218 , n39979 );
and ( n57219 , n57218 , n31505 );
buf ( n57220 , n31203 );
and ( n57221 , n57220 , n39979 );
or ( n57222 , n57219 , n57221 );
and ( n57223 , n57222 , n31538 );
and ( n57224 , n31505 , n40143 );
or ( n57225 , n57217 , n57223 , n57224 );
and ( n57226 , n57225 , n31557 );
and ( n57227 , n31505 , n40154 );
or ( n57228 , C0 , n57226 , n57227 );
buf ( n57229 , n57228 );
buf ( n57230 , n57229 );
not ( n57231 , n40163 );
and ( n57232 , n57231 , n31850 );
nor ( n57233 , n42169 , n42237 , n31665 , n31661 , n31657 );
not ( n57234 , n57233 );
and ( n57235 , n57234 , n31850 );
and ( n57236 , n32235 , n57233 );
or ( n57237 , n57235 , n57236 );
and ( n57238 , n57237 , n40163 );
or ( n57239 , n57232 , n57238 );
and ( n57240 , n57239 , n32498 );
nor ( n57241 , n42179 , n42246 , n40188 , n40194 , C0 );
not ( n57242 , n57241 );
not ( n57243 , n57233 );
and ( n57244 , n57243 , n31850 );
and ( n57245 , n42188 , n57233 );
or ( n57246 , n57244 , n57245 );
and ( n57247 , n57242 , n57246 );
and ( n57248 , n42188 , n57241 );
or ( n57249 , n57247 , n57248 );
and ( n57250 , n57249 , n32473 );
not ( n57251 , n32475 );
not ( n57252 , n57241 );
not ( n57253 , n57233 );
and ( n57254 , n57253 , n31850 );
and ( n57255 , n42188 , n57233 );
or ( n57256 , n57254 , n57255 );
and ( n57257 , n57252 , n57256 );
and ( n57258 , n42188 , n57241 );
or ( n57259 , n57257 , n57258 );
and ( n57260 , n57251 , n57259 );
nor ( n57261 , n42205 , n42272 , n40435 , n40445 , C0 );
not ( n57262 , n57261 );
nor ( n57263 , n42208 , n42275 , n40430 , n40440 , C0 );
not ( n57264 , n57263 );
and ( n57265 , n57264 , n57259 );
and ( n57266 , n42216 , n57263 );
or ( n57267 , n57265 , n57266 );
and ( n57268 , n57262 , n57267 );
and ( n57269 , n42224 , n57261 );
or ( n57270 , n57268 , n57269 );
and ( n57271 , n57270 , n32475 );
or ( n57272 , n57260 , n57271 );
and ( n57273 , n57272 , n32486 );
and ( n57274 , n31850 , n41278 );
or ( n57275 , C0 , n57240 , n57250 , n57273 , n57274 );
buf ( n57276 , n57275 );
buf ( n57277 , n57276 );
buf ( n57278 , n30987 );
buf ( n57279 , n31655 );
and ( n57280 , n42376 , n42402 );
xor ( n57281 , n52404 , n57280 );
and ( n57282 , n57281 , n48455 );
not ( n57283 , n48457 );
and ( n57284 , n57283 , n52404 );
and ( n57285 , n57281 , n48457 );
or ( n57286 , n57284 , n57285 );
and ( n57287 , n57286 , n31373 );
not ( n57288 , n44807 );
and ( n57289 , n57288 , n52404 );
and ( n57290 , n57281 , n44807 );
or ( n57291 , n57289 , n57290 );
and ( n57292 , n57291 , n31408 );
not ( n57293 , n48468 );
and ( n57294 , n57293 , n52404 );
and ( n57295 , n57281 , n48468 );
or ( n57296 , n57294 , n57295 );
and ( n57297 , n57296 , n31468 );
not ( n57298 , n44817 );
and ( n57299 , n57298 , n52404 );
and ( n57300 , n57281 , n44817 );
or ( n57301 , n57299 , n57300 );
and ( n57302 , n57301 , n31521 );
not ( n57303 , n39979 );
and ( n57304 , n57303 , n52404 );
and ( n57305 , n42376 , n42383 );
xor ( n57306 , n52404 , n57305 );
and ( n57307 , n57306 , n39979 );
or ( n57308 , n57304 , n57307 );
and ( n57309 , n57308 , n31538 );
not ( n57310 , n45059 );
and ( n57311 , n57310 , n52404 );
and ( n57312 , n57306 , n45059 );
or ( n57313 , n57311 , n57312 );
and ( n57314 , n57313 , n31536 );
not ( n57315 , n33419 );
and ( n57316 , n57315 , n52404 );
and ( n57317 , n42384 , n42391 );
xor ( n57318 , n57306 , n57317 );
and ( n57319 , n57318 , n33419 );
or ( n57320 , n57316 , n57319 );
and ( n57321 , n57320 , n31529 );
not ( n57322 , n33734 );
and ( n57323 , n57322 , n52404 );
not ( n57324 , n33533 );
and ( n57325 , n42403 , n42410 );
xor ( n57326 , n57281 , n57325 );
and ( n57327 , n57324 , n57326 );
and ( n57328 , n42376 , n42416 );
xor ( n57329 , n52404 , n57328 );
or ( n57330 , n42417 , n42424 );
xnor ( n57331 , n57329 , n57330 );
and ( n57332 , n57331 , n33533 );
or ( n57333 , n57327 , n57332 );
and ( n57334 , n57333 , n33734 );
or ( n57335 , n57323 , n57334 );
and ( n57336 , n57335 , n31527 );
and ( n57337 , n57329 , n48513 );
or ( n57338 , n57282 , n57287 , n57292 , n57297 , n57302 , n57309 , n57314 , n57321 , n57336 , n57337 );
and ( n57339 , n57338 , n31557 );
and ( n57340 , n35391 , n33973 );
and ( n57341 , n52404 , n48524 );
or ( n57342 , C0 , n57339 , n57340 , n57341 );
buf ( n57343 , n57342 );
buf ( n57344 , n57343 );
buf ( n57345 , n30987 );
buf ( n57346 , n31655 );
not ( n57347 , n38443 );
and ( n57348 , n57347 , n38303 );
xor ( n57349 , n53464 , n53505 );
and ( n57350 , n57349 , n38443 );
or ( n57351 , n57348 , n57350 );
and ( n57352 , n57351 , n38450 );
not ( n57353 , n39339 );
and ( n57354 , n57353 , n39203 );
xor ( n57355 , n53520 , n53561 );
and ( n57356 , n57355 , n39339 );
or ( n57357 , n57354 , n57356 );
and ( n57358 , n57357 , n39346 );
and ( n57359 , n40220 , n39359 );
or ( n57360 , n57352 , n57358 , n57359 );
buf ( n57361 , n57360 );
buf ( n57362 , n57361 );
not ( n57363 , n46356 );
and ( n57364 , n57363 , n31189 );
not ( n57365 , n55263 );
and ( n57366 , n57365 , n31189 );
and ( n57367 , n31205 , n55263 );
or ( n57368 , n57366 , n57367 );
and ( n57369 , n57368 , n46356 );
or ( n57370 , n57364 , n57369 );
and ( n57371 , n57370 , n31649 );
not ( n57372 , n55271 );
not ( n57373 , n55263 );
and ( n57374 , n57373 , n31189 );
and ( n57375 , n50125 , n55263 );
or ( n57376 , n57374 , n57375 );
and ( n57377 , n57372 , n57376 );
and ( n57378 , n50125 , n55271 );
or ( n57379 , n57377 , n57378 );
and ( n57380 , n57379 , n31643 );
not ( n57381 , n31452 );
not ( n57382 , n55271 );
not ( n57383 , n55263 );
and ( n57384 , n57383 , n31189 );
and ( n57385 , n50125 , n55263 );
or ( n57386 , n57384 , n57385 );
and ( n57387 , n57382 , n57386 );
and ( n57388 , n50125 , n55271 );
or ( n57389 , n57387 , n57388 );
and ( n57390 , n57381 , n57389 );
not ( n57391 , n55291 );
not ( n57392 , n55293 );
and ( n57393 , n57392 , n57389 );
and ( n57394 , n50151 , n55293 );
or ( n57395 , n57393 , n57394 );
and ( n57396 , n57391 , n57395 );
and ( n57397 , n50159 , n55291 );
or ( n57398 , n57396 , n57397 );
and ( n57399 , n57398 , n31452 );
or ( n57400 , n57390 , n57399 );
and ( n57401 , n57400 , n31638 );
and ( n57402 , n31189 , n47277 );
or ( n57403 , C0 , n57371 , n57380 , n57401 , n57402 );
buf ( n57404 , n57403 );
buf ( n57405 , n57404 );
xor ( n57406 , n46159 , n49991 );
and ( n57407 , n57406 , n32431 );
not ( n57408 , n50002 );
and ( n57409 , n57408 , n46159 );
and ( n57410 , n40341 , n50002 );
or ( n57411 , n57409 , n57410 );
and ( n57412 , n57411 , n32419 );
not ( n57413 , n50008 );
and ( n57414 , n57413 , n46159 );
not ( n57415 , n47910 );
buf ( n57416 , RI15b5f310_1113);
and ( n57417 , n57415 , n57416 );
not ( n57418 , n48101 );
and ( n57419 , n57418 , n47989 );
xor ( n57420 , n48105 , n48117 );
and ( n57421 , n57420 , n48101 );
or ( n57422 , n57419 , n57421 );
and ( n57423 , n57422 , n47910 );
or ( n57424 , n57417 , n57423 );
and ( n57425 , n57424 , n50008 );
or ( n57426 , n57414 , n57425 );
and ( n57427 , n57426 , n32415 );
not ( n57428 , n50067 );
and ( n57429 , n57428 , n46159 );
and ( n57430 , n31858 , n50067 );
or ( n57431 , n57429 , n57430 );
and ( n57432 , n57431 , n32411 );
and ( n57433 , n46159 , n50098 );
or ( n57434 , n57407 , n57412 , n57427 , n57432 , n57433 );
and ( n57435 , n57434 , n32456 );
and ( n57436 , n46159 , n47409 );
or ( n57437 , C0 , n57435 , n57436 );
buf ( n57438 , n57437 );
buf ( n57439 , n57438 );
buf ( n57440 , n30987 );
buf ( n57441 , n31655 );
buf ( n57442 , n31655 );
not ( n57443 , n38443 );
and ( n57444 , n57443 , n38252 );
xor ( n57445 , n53467 , n53502 );
and ( n57446 , n57445 , n38443 );
or ( n57447 , n57444 , n57446 );
and ( n57448 , n57447 , n38450 );
not ( n57449 , n39339 );
and ( n57450 , n57449 , n39152 );
xor ( n57451 , n53523 , n53558 );
and ( n57452 , n57451 , n39339 );
or ( n57453 , n57450 , n57452 );
and ( n57454 , n57453 , n39346 );
and ( n57455 , n40217 , n39359 );
or ( n57456 , n57448 , n57454 , n57455 );
buf ( n57457 , n57456 );
buf ( n57458 , n57457 );
buf ( n57459 , n30987 );
buf ( n57460 , n31655 );
and ( n57461 , n52404 , n57280 );
and ( n57462 , n52402 , n57461 );
and ( n57463 , n52400 , n57462 );
xor ( n57464 , n52398 , n57463 );
and ( n57465 , n57464 , n48455 );
not ( n57466 , n48457 );
and ( n57467 , n57466 , n52398 );
and ( n57468 , n57464 , n48457 );
or ( n57469 , n57467 , n57468 );
and ( n57470 , n57469 , n31373 );
not ( n57471 , n44807 );
and ( n57472 , n57471 , n52398 );
and ( n57473 , n57464 , n44807 );
or ( n57474 , n57472 , n57473 );
and ( n57475 , n57474 , n31408 );
not ( n57476 , n48468 );
and ( n57477 , n57476 , n52398 );
and ( n57478 , n57464 , n48468 );
or ( n57479 , n57477 , n57478 );
and ( n57480 , n57479 , n31468 );
not ( n57481 , n44817 );
and ( n57482 , n57481 , n52398 );
and ( n57483 , n57464 , n44817 );
or ( n57484 , n57482 , n57483 );
and ( n57485 , n57484 , n31521 );
not ( n57486 , n39979 );
and ( n57487 , n57486 , n52398 );
and ( n57488 , n52404 , n57305 );
and ( n57489 , n52402 , n57488 );
and ( n57490 , n52400 , n57489 );
xor ( n57491 , n52398 , n57490 );
and ( n57492 , n57491 , n39979 );
or ( n57493 , n57487 , n57492 );
and ( n57494 , n57493 , n31538 );
not ( n57495 , n45059 );
and ( n57496 , n57495 , n52398 );
and ( n57497 , n57491 , n45059 );
or ( n57498 , n57496 , n57497 );
and ( n57499 , n57498 , n31536 );
not ( n57500 , n33419 );
and ( n57501 , n57500 , n52398 );
xor ( n57502 , n52400 , n57489 );
xor ( n57503 , n52402 , n57488 );
and ( n57504 , n57306 , n57317 );
and ( n57505 , n57503 , n57504 );
and ( n57506 , n57502 , n57505 );
xor ( n57507 , n57491 , n57506 );
and ( n57508 , n57507 , n33419 );
or ( n57509 , n57501 , n57508 );
and ( n57510 , n57509 , n31529 );
not ( n57511 , n33734 );
and ( n57512 , n57511 , n52398 );
not ( n57513 , n33533 );
xor ( n57514 , n52400 , n57462 );
xor ( n57515 , n52402 , n57461 );
and ( n57516 , n57281 , n57325 );
and ( n57517 , n57515 , n57516 );
and ( n57518 , n57514 , n57517 );
xor ( n57519 , n57464 , n57518 );
and ( n57520 , n57513 , n57519 );
and ( n57521 , n52404 , n57328 );
and ( n57522 , n52402 , n57521 );
and ( n57523 , n52400 , n57522 );
xor ( n57524 , n52398 , n57523 );
xor ( n57525 , n52400 , n57522 );
xor ( n57526 , n52402 , n57521 );
or ( n57527 , n57329 , n57330 );
or ( n57528 , n57526 , n57527 );
or ( n57529 , n57525 , n57528 );
xnor ( n57530 , n57524 , n57529 );
and ( n57531 , n57530 , n33533 );
or ( n57532 , n57520 , n57531 );
and ( n57533 , n57532 , n33734 );
or ( n57534 , n57512 , n57533 );
and ( n57535 , n57534 , n31527 );
and ( n57536 , n57524 , n48513 );
or ( n57537 , n57465 , n57470 , n57475 , n57480 , n57485 , n57494 , n57499 , n57510 , n57535 , n57536 );
and ( n57538 , n57537 , n31557 );
and ( n57539 , n35388 , n33973 );
and ( n57540 , n52398 , n48524 );
or ( n57541 , C0 , n57538 , n57539 , n57540 );
buf ( n57542 , n57541 );
buf ( n57543 , n57542 );
buf ( n57544 , n30987 );
buf ( n57545 , n30987 );
buf ( n57546 , n31655 );
buf ( n57547 , n31655 );
not ( n57548 , n34150 );
and ( n57549 , n57548 , n33381 );
not ( n57550 , n56687 );
and ( n57551 , n57550 , n33379 );
not ( n57552 , n32967 );
and ( n57553 , n57552 , n32511 );
buf ( n57554 , n32967 );
or ( n57555 , n57553 , n57554 );
and ( n57556 , n57555 , n33377 );
not ( n57557 , n48642 );
and ( n57558 , n57557 , n32531 );
buf ( n57559 , n57558 );
and ( n57560 , n57559 , n32890 );
not ( n57561 , n48648 );
and ( n57562 , n57561 , n32531 );
and ( n57563 , n32535 , n52245 );
xor ( n57564 , n32531 , n57563 );
and ( n57565 , n57564 , n48648 );
or ( n57566 , n57562 , n57565 );
and ( n57567 , n57566 , n32924 );
not ( n57568 , n48654 );
and ( n57569 , n57568 , n32531 );
buf ( n57570 , n57569 );
and ( n57571 , n57570 , n33038 );
not ( n57572 , n48660 );
and ( n57573 , n57572 , n32531 );
buf ( n57574 , n57573 );
and ( n57575 , n57574 , n33172 );
not ( n57576 , n41576 );
and ( n57577 , n57576 , n32531 );
buf ( n57578 , n57577 );
and ( n57579 , n57578 , n33189 );
not ( n57580 , n48730 );
and ( n57581 , n57580 , n32531 );
buf ( n57582 , n57581 );
and ( n57583 , n57582 , n33187 );
or ( n57584 , n33178 , n33180 );
and ( n57585 , n32531 , n57584 );
or ( n57586 , C0 , n57560 , n57567 , n57571 , n57575 , n57579 , n57583 , n57585 , C0 );
not ( n57587 , n57586 );
and ( n57588 , n57587 , n32530 );
and ( n57589 , n52250 , n48639 );
not ( n57590 , n48642 );
and ( n57591 , n57590 , n32535 );
and ( n57592 , n52250 , n48642 );
or ( n57593 , n57591 , n57592 );
and ( n57594 , n57593 , n32890 );
not ( n57595 , n48648 );
and ( n57596 , n57595 , n32535 );
and ( n57597 , n52246 , n48648 );
or ( n57598 , n57596 , n57597 );
and ( n57599 , n57598 , n32924 );
not ( n57600 , n48654 );
and ( n57601 , n57600 , n32535 );
and ( n57602 , n52250 , n48654 );
or ( n57603 , n57601 , n57602 );
and ( n57604 , n57603 , n33038 );
not ( n57605 , n48660 );
and ( n57606 , n57605 , n32535 );
and ( n57607 , n52250 , n48660 );
or ( n57608 , n57606 , n57607 );
and ( n57609 , n57608 , n33172 );
not ( n57610 , n41576 );
and ( n57611 , n57610 , n32535 );
and ( n57612 , n32543 , n32547 );
or ( n57613 , n32539 , n57612 );
xor ( n57614 , n32535 , n57613 );
not ( n57615 , n57614 );
buf ( n57616 , n57615 );
buf ( n57617 , n57616 );
not ( n57618 , n57617 );
and ( n57619 , n57618 , n41576 );
or ( n57620 , n57611 , n57619 );
and ( n57621 , n57620 , n33189 );
not ( n57622 , n48730 );
and ( n57623 , n57622 , n32535 );
and ( n57624 , n57618 , n48730 );
or ( n57625 , n57623 , n57624 );
and ( n57626 , n57625 , n33187 );
and ( n57627 , n32535 , n57584 );
and ( n57628 , n48811 , n49275 );
or ( n57629 , n57589 , n57594 , n57599 , n57604 , n57609 , n57621 , n57626 , n57627 , n57628 );
not ( n57630 , n57629 );
and ( n57631 , n57630 , n32534 );
and ( n57632 , n52243 , n48639 );
not ( n57633 , n48642 );
and ( n57634 , n57633 , n32539 );
and ( n57635 , n52243 , n48642 );
or ( n57636 , n57634 , n57635 );
and ( n57637 , n57636 , n32890 );
not ( n57638 , n48648 );
and ( n57639 , n57638 , n32539 );
and ( n57640 , n52239 , n48648 );
or ( n57641 , n57639 , n57640 );
and ( n57642 , n57641 , n32924 );
not ( n57643 , n48654 );
and ( n57644 , n57643 , n32539 );
and ( n57645 , n52243 , n48654 );
or ( n57646 , n57644 , n57645 );
and ( n57647 , n57646 , n33038 );
not ( n57648 , n48660 );
and ( n57649 , n57648 , n32539 );
and ( n57650 , n52243 , n48660 );
or ( n57651 , n57649 , n57650 );
and ( n57652 , n57651 , n33172 );
not ( n57653 , n41576 );
and ( n57654 , n57653 , n32539 );
xnor ( n57655 , n32539 , n57612 );
not ( n57656 , n57655 );
buf ( n57657 , n57656 );
buf ( n57658 , n57657 );
not ( n57659 , n57658 );
and ( n57660 , n57659 , n41576 );
or ( n57661 , n57654 , n57660 );
and ( n57662 , n57661 , n33189 );
not ( n57663 , n48730 );
and ( n57664 , n57663 , n32539 );
and ( n57665 , n57659 , n48730 );
or ( n57666 , n57664 , n57665 );
and ( n57667 , n57666 , n33187 );
and ( n57668 , n32539 , n57584 );
and ( n57669 , n48805 , n49275 );
or ( n57670 , n57632 , n57637 , n57642 , n57647 , n57652 , n57662 , n57667 , n57668 , n57669 );
not ( n57671 , n57670 );
and ( n57672 , n57671 , n32538 );
and ( n57673 , n52237 , n48639 );
not ( n57674 , n48642 );
and ( n57675 , n57674 , n32543 );
and ( n57676 , n52237 , n48642 );
or ( n57677 , n57675 , n57676 );
and ( n57678 , n57677 , n32890 );
not ( n57679 , n48648 );
and ( n57680 , n57679 , n32543 );
and ( n57681 , n52233 , n48648 );
or ( n57682 , n57680 , n57681 );
and ( n57683 , n57682 , n32924 );
not ( n57684 , n48654 );
and ( n57685 , n57684 , n32543 );
and ( n57686 , n52237 , n48654 );
or ( n57687 , n57685 , n57686 );
and ( n57688 , n57687 , n33038 );
not ( n57689 , n48660 );
and ( n57690 , n57689 , n32543 );
and ( n57691 , n52237 , n48660 );
or ( n57692 , n57690 , n57691 );
and ( n57693 , n57692 , n33172 );
not ( n57694 , n41576 );
and ( n57695 , n57694 , n32543 );
xor ( n57696 , n32543 , n32547 );
not ( n57697 , n57696 );
buf ( n57698 , n57697 );
buf ( n57699 , n57698 );
not ( n57700 , n57699 );
and ( n57701 , n57700 , n41576 );
or ( n57702 , n57695 , n57701 );
and ( n57703 , n57702 , n33189 );
not ( n57704 , n48730 );
and ( n57705 , n57704 , n32543 );
and ( n57706 , n57700 , n48730 );
or ( n57707 , n57705 , n57706 );
and ( n57708 , n57707 , n33187 );
and ( n57709 , n32543 , n57584 );
and ( n57710 , n48799 , n49275 );
or ( n57711 , n57673 , n57678 , n57683 , n57688 , n57693 , n57703 , n57708 , n57709 , n57710 );
not ( n57712 , n57711 );
and ( n57713 , n57712 , n32542 );
and ( n57714 , n52231 , n48639 );
buf ( n57715 , n32547 );
and ( n57716 , n57715 , n32890 );
buf ( n57717 , n32547 );
and ( n57718 , n57717 , n32924 );
buf ( n57719 , n32547 );
and ( n57720 , n57719 , n33038 );
buf ( n57721 , n32547 );
and ( n57722 , n57721 , n33172 );
not ( n57723 , n41576 );
and ( n57724 , n57723 , n32547 );
not ( n57725 , n32547 );
not ( n57726 , n57725 );
buf ( n57727 , n57726 );
not ( n57728 , n57727 );
and ( n57729 , n57728 , n41576 );
or ( n57730 , n57724 , n57729 );
and ( n57731 , n57730 , n33189 );
not ( n57732 , n48730 );
and ( n57733 , n57732 , n32547 );
and ( n57734 , n57728 , n48730 );
or ( n57735 , n57733 , n57734 );
and ( n57736 , n57735 , n33187 );
and ( n57737 , n32547 , n57584 );
and ( n57738 , n48793 , n49275 );
or ( n57739 , n57714 , n57716 , n57718 , n57720 , n57722 , n57731 , n57736 , n57737 , n57738 );
not ( n57740 , n57739 );
and ( n57741 , n57740 , n32546 );
xnor ( n57742 , n57711 , n32542 );
and ( n57743 , n57741 , n57742 );
or ( n57744 , n57713 , n57743 );
xnor ( n57745 , n57670 , n32538 );
and ( n57746 , n57744 , n57745 );
or ( n57747 , n57672 , n57746 );
xnor ( n57748 , n57629 , n32534 );
and ( n57749 , n57747 , n57748 );
or ( n57750 , n57631 , n57749 );
xnor ( n57751 , n57586 , n32530 );
and ( n57752 , n57750 , n57751 );
or ( n57753 , n57588 , n57752 );
not ( n57754 , n57753 );
not ( n57755 , n57586 );
not ( n57756 , n57629 );
buf ( n57757 , n57586 );
buf ( n57758 , n57586 );
buf ( n57759 , n57586 );
buf ( n57760 , n57586 );
buf ( n57761 , n57586 );
buf ( n57762 , n57586 );
buf ( n57763 , n57586 );
buf ( n57764 , n57586 );
buf ( n57765 , n57586 );
buf ( n57766 , n57586 );
buf ( n57767 , n57586 );
buf ( n57768 , n57586 );
buf ( n57769 , n57586 );
buf ( n57770 , n57586 );
buf ( n57771 , n57586 );
buf ( n57772 , n57586 );
buf ( n57773 , n57586 );
buf ( n57774 , n57586 );
buf ( n57775 , n57586 );
buf ( n57776 , n57586 );
buf ( n57777 , n57586 );
buf ( n57778 , n57586 );
buf ( n57779 , n57586 );
buf ( n57780 , n57586 );
buf ( n57781 , n57586 );
buf ( n57782 , n57586 );
not ( n57783 , n57670 );
or ( n57784 , n57756 , n57586 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 );
nand ( n57785 , n57755 , n57784 );
not ( n57786 , n48641 );
and ( n57787 , n32598 , n57786 );
and ( n57788 , n56464 , n57787 );
and ( n57789 , n57788 , n32890 );
and ( n57790 , n32919 , n32966 );
and ( n57791 , n56464 , n57790 );
and ( n57792 , n57791 , n32924 );
and ( n57793 , n32953 , n57786 );
and ( n57794 , n56464 , n57793 );
and ( n57795 , n57794 , n33038 );
and ( n57796 , n33067 , n32966 );
and ( n57797 , n56464 , n57796 );
and ( n57798 , n57797 , n33172 );
and ( n57799 , n48765 , n33180 );
and ( n57800 , n49054 , n33178 );
or ( n57801 , n57789 , n57792 , n57795 , n57798 , n57799 , n57800 , C0 );
or ( n57802 , n57785 , n57801 );
not ( n57803 , n32598 );
buf ( n57804 , n57803 );
buf ( n57805 , RI15b44c40_211);
not ( n57806 , n48641 );
and ( n57807 , n57805 , n57806 );
and ( n57808 , n57807 , n32598 );
or ( n57809 , n57804 , n57808 );
and ( n57810 , n57809 , n32890 );
not ( n57811 , n32919 );
buf ( n57812 , n57811 );
not ( n57813 , n32967 );
and ( n57814 , n57805 , n57813 );
and ( n57815 , n57814 , n32919 );
or ( n57816 , n57812 , n57815 );
and ( n57817 , n57816 , n32924 );
not ( n57818 , n32953 );
buf ( n57819 , n57818 );
and ( n57820 , n57807 , n32953 );
or ( n57821 , n57819 , n57820 );
and ( n57822 , n57821 , n33038 );
not ( n57823 , n33067 );
buf ( n57824 , n57823 );
and ( n57825 , n57814 , n33067 );
or ( n57826 , n57824 , n57825 );
and ( n57827 , n57826 , n33172 );
not ( n57828 , n41576 );
and ( n57829 , n57828 , n33189 );
not ( n57830 , n48730 );
and ( n57831 , n57830 , n33187 );
not ( n57832 , n48765 );
and ( n57833 , n57832 , n33180 );
not ( n57834 , n49054 );
and ( n57835 , n57834 , n33178 );
or ( n57836 , n57810 , n57817 , n57822 , n57827 , n57829 , n57831 , n57833 , n57835 , C0 );
or ( n57837 , n57802 , n57836 );
or ( n57838 , n57754 , n57837 );
not ( n57839 , n57838 );
and ( n57840 , n32953 , n32971 );
not ( n57841 , n57840 );
and ( n57842 , n57841 , n32511 );
buf ( n57843 , n57842 );
and ( n57844 , n57843 , n33038 );
or ( n57845 , n48564 , n32890 );
or ( n57846 , n57845 , n33191 );
or ( n57847 , n57846 , n33193 );
or ( n57848 , n57847 , n33195 );
or ( n57849 , n57848 , n33197 );
or ( n57850 , n57849 , n33199 );
or ( n57851 , n57850 , n33201 );
or ( n57852 , n57851 , n33203 );
and ( n57853 , n32511 , n57852 );
or ( n57854 , n57844 , n57853 );
and ( n57855 , n57839 , n57854 );
buf ( n57856 , n57838 );
or ( n57857 , n57855 , n57856 );
and ( n57858 , n57857 , n33208 );
buf ( n57859 , n33375 );
not ( n57860 , n32967 );
and ( n57861 , n57860 , n33373 );
buf ( n57862 , n33370 );
and ( n57863 , n57860 , n33372 );
or ( n57864 , n35056 , n32528 );
buf ( n57865 , n57864 );
or ( n57866 , C0 , n57549 , n57551 , n57556 , n57858 , n57859 , n57861 , n57862 , n57863 , n57865 );
buf ( n57867 , n57866 );
buf ( n57868 , n57867 );
buf ( n57869 , n31655 );
not ( n57870 , n34150 );
and ( n57871 , n57870 , n32625 );
and ( n57872 , n32546 , n34153 , n41390 , n32534 , n41391 );
not ( n57873 , n57872 );
and ( n57874 , n57873 , n32625 );
and ( n57875 , n32655 , n57872 );
or ( n57876 , n57874 , n57875 );
and ( n57877 , n57876 , n34150 );
or ( n57878 , n57871 , n57877 );
and ( n57879 , n57878 , n33381 );
and ( n57880 , n34165 , n34171 , n41401 , n34183 , C1 );
not ( n57881 , n57880 );
not ( n57882 , n57872 );
and ( n57883 , n57882 , n32625 );
and ( n57884 , n56044 , n57872 );
or ( n57885 , n57883 , n57884 );
and ( n57886 , n57881 , n57885 );
and ( n57887 , n56044 , n57880 );
or ( n57888 , n57886 , n57887 );
and ( n57889 , n57888 , n33375 );
not ( n57890 , n32968 );
not ( n57891 , n57880 );
not ( n57892 , n57872 );
and ( n57893 , n57892 , n32625 );
and ( n57894 , n56044 , n57872 );
or ( n57895 , n57893 , n57894 );
and ( n57896 , n57891 , n57895 );
and ( n57897 , n56044 , n57880 );
or ( n57898 , n57896 , n57897 );
and ( n57899 , n57890 , n57898 );
and ( n57900 , n34325 , n34334 , n41423 , n34354 , C1 );
not ( n57901 , n57900 );
and ( n57902 , n34321 , n34357 , n41427 , n34349 , C1 );
not ( n57903 , n57902 );
and ( n57904 , n57903 , n57898 );
and ( n57905 , n56068 , n57902 );
or ( n57906 , n57904 , n57905 );
and ( n57907 , n57901 , n57906 );
and ( n57908 , n56076 , n57900 );
or ( n57909 , n57907 , n57908 );
and ( n57910 , n57909 , n32968 );
or ( n57911 , n57899 , n57910 );
and ( n57912 , n57911 , n33370 );
and ( n57913 , n32625 , n35062 );
or ( n57914 , C0 , n57879 , n57889 , n57912 , n57913 );
buf ( n57915 , n57914 );
buf ( n57916 , n57915 );
buf ( n57917 , n31655 );
buf ( n57918 , n30987 );
buf ( n57919 , n30987 );
buf ( n57920 , n31655 );
buf ( n57921 , n30987 );
not ( n57922 , n46356 );
and ( n57923 , n57922 , n31021 );
and ( n57924 , n46379 , n46356 );
or ( n57925 , n57923 , n57924 );
and ( n57926 , n57925 , n31649 );
not ( n57927 , n52614 );
not ( n57928 , n44702 );
and ( n57929 , n57928 , n31021 );
buf ( n57930 , n57929 );
and ( n57931 , n57927 , n57930 );
buf ( n57932 , n57931 );
and ( n57933 , n57932 , n31647 );
and ( n57934 , n46524 , n31643 );
not ( n57935 , n31452 );
and ( n57936 , n57935 , n46524 );
xor ( n57937 , n46528 , n46519 );
not ( n57938 , n57937 );
buf ( n57939 , n57938 );
not ( n57940 , n57939 );
and ( n57941 , n57940 , n31452 );
or ( n57942 , n57936 , n57941 );
and ( n57943 , n57942 , n31638 );
and ( n57944 , n31021 , n52626 );
or ( n57945 , C0 , n57926 , n57933 , n57934 , n57943 , n57944 );
buf ( n57946 , n57945 );
buf ( n57947 , n57946 );
buf ( n57948 , n30987 );
buf ( n57949 , n31655 );
not ( n57950 , n31728 );
and ( n57951 , n57950 , n32461 );
xor ( n57952 , n31895 , n31928 );
xor ( n57953 , n57952 , n32078 );
and ( n57954 , n57953 , n31728 );
or ( n57955 , n57951 , n57954 );
and ( n57956 , n57955 , n32253 );
not ( n57957 , n32283 );
and ( n57958 , n57957 , n32461 );
not ( n57959 , n31823 );
xor ( n57960 , n32300 , n31928 );
xor ( n57961 , n57960 , n32317 );
and ( n57962 , n57959 , n57961 );
xor ( n57963 , n32352 , n32354 );
xor ( n57964 , n57963 , n32380 );
and ( n57965 , n57964 , n31823 );
or ( n57966 , n57962 , n57965 );
and ( n57967 , n57966 , n32283 );
or ( n57968 , n57958 , n57967 );
and ( n57969 , n57968 , n32398 );
and ( n57970 , n32461 , n32436 );
or ( n57971 , n57956 , n57969 , n57970 );
and ( n57972 , n57971 , n32456 );
and ( n57973 , n49699 , n32473 );
not ( n57974 , n32475 );
and ( n57975 , n57974 , n49699 );
xor ( n57976 , n32461 , n32478 );
and ( n57977 , n57976 , n32475 );
or ( n57978 , n57975 , n57977 );
and ( n57979 , n57978 , n32486 );
and ( n57980 , n37581 , n32489 );
and ( n57981 , n32461 , n32501 );
or ( n57982 , C0 , n57972 , n57973 , n57979 , n57980 , n57981 );
buf ( n57983 , n57982 );
buf ( n57984 , n57983 );
buf ( n57985 , n30987 );
buf ( n57986 , n30987 );
buf ( n57987 , n31655 );
not ( n57988 , n32967 );
and ( n57989 , n57988 , n32514 );
buf ( n57990 , n57989 );
and ( n57991 , n57990 , n33377 );
not ( n57992 , n57838 );
not ( n57993 , n57840 );
and ( n57994 , n57993 , n32514 );
buf ( n57995 , n57840 );
or ( n57996 , n57994 , n57995 );
and ( n57997 , n57996 , n33038 );
and ( n57998 , n32514 , n57852 );
or ( n57999 , n57997 , n57998 );
and ( n58000 , n57992 , n57999 );
buf ( n58001 , n57838 );
or ( n58002 , n58000 , n58001 );
and ( n58003 , n58002 , n33208 );
and ( n58004 , n57860 , n33373 );
not ( n58005 , n32968 );
and ( n58006 , n58005 , n33370 );
not ( n58007 , n57860 );
and ( n58008 , n58007 , n33372 );
or ( n58009 , C0 , C0 , C0 , n57991 , n58003 , C0 , n58004 , n58006 , n58008 , C0 );
buf ( n58010 , n58009 );
buf ( n58011 , n58010 );
buf ( n58012 , n31655 );
buf ( n58013 , n30987 );
buf ( n58014 , n31655 );
buf ( n58015 , n31655 );
buf ( n58016 , n30987 );
not ( n58017 , n32953 );
buf ( n58018 , RI15b46a40_275);
and ( n58019 , n58017 , n58018 );
not ( n58020 , n39572 );
and ( n58021 , n58020 , n39451 );
xor ( n58022 , n42622 , n42631 );
and ( n58023 , n58022 , n39572 );
or ( n58024 , n58021 , n58023 );
and ( n58025 , n58024 , n32953 );
or ( n58026 , n58019 , n58025 );
and ( n58027 , n58026 , n33038 );
not ( n58028 , n39586 );
and ( n58029 , n58028 , n58018 );
not ( n58030 , n39775 );
and ( n58031 , n58030 , n39663 );
xor ( n58032 , n42658 , n42667 );
and ( n58033 , n58032 , n39775 );
or ( n58034 , n58031 , n58033 );
and ( n58035 , n58034 , n39586 );
or ( n58036 , n58029 , n58035 );
and ( n58037 , n58036 , n33172 );
and ( n58038 , n58018 , n39795 );
or ( n58039 , n58027 , n58037 , n58038 );
and ( n58040 , n58039 , n33208 );
and ( n58041 , n58018 , n39805 );
or ( n58042 , C0 , n58040 , n58041 );
buf ( n58043 , n58042 );
buf ( n58044 , n58043 );
not ( n58045 , n46356 );
and ( n58046 , n58045 , n31288 );
not ( n58047 , n48214 );
and ( n58048 , n58047 , n31288 );
and ( n58049 , n31306 , n48214 );
or ( n58050 , n58048 , n58049 );
and ( n58051 , n58050 , n46356 );
or ( n58052 , n58046 , n58051 );
and ( n58053 , n58052 , n31649 );
not ( n58054 , n48223 );
not ( n58055 , n48214 );
and ( n58056 , n58055 , n31288 );
not ( n58057 , n46487 );
and ( n58058 , n58057 , n46459 );
xor ( n58059 , n47438 , n47445 );
and ( n58060 , n58059 , n46487 );
or ( n58061 , n58058 , n58060 );
and ( n58062 , n58061 , n48214 );
or ( n58063 , n58056 , n58062 );
and ( n58064 , n58054 , n58063 );
and ( n58065 , n58061 , n48223 );
or ( n58066 , n58064 , n58065 );
and ( n58067 , n58066 , n31643 );
not ( n58068 , n31452 );
not ( n58069 , n48223 );
not ( n58070 , n48214 );
and ( n58071 , n58070 , n31288 );
and ( n58072 , n58061 , n48214 );
or ( n58073 , n58071 , n58072 );
and ( n58074 , n58069 , n58073 );
and ( n58075 , n58061 , n48223 );
or ( n58076 , n58074 , n58075 );
and ( n58077 , n58068 , n58076 );
not ( n58078 , n48244 );
not ( n58079 , n48247 );
and ( n58080 , n58079 , n58076 );
not ( n58081 , n46976 );
and ( n58082 , n58081 , n46938 );
xor ( n58083 , n47474 , n47481 );
and ( n58084 , n58083 , n46976 );
or ( n58085 , n58082 , n58084 );
and ( n58086 , n58085 , n48247 );
or ( n58087 , n58080 , n58086 );
and ( n58088 , n58078 , n58087 );
not ( n58089 , n47259 );
and ( n58090 , n58089 , n47225 );
xor ( n58091 , n47492 , n47499 );
and ( n58092 , n58091 , n47259 );
or ( n58093 , n58090 , n58092 );
and ( n58094 , n58093 , n48244 );
or ( n58095 , n58088 , n58094 );
and ( n58096 , n58095 , n31452 );
or ( n58097 , n58077 , n58096 );
and ( n58098 , n58097 , n31638 );
and ( n58099 , n31288 , n47277 );
or ( n58100 , C0 , n58053 , n58067 , n58098 , n58099 );
buf ( n58101 , n58100 );
buf ( n58102 , n58101 );
buf ( n58103 , n31655 );
buf ( n58104 , n30987 );
buf ( n58105 , n31655 );
not ( n58106 , n52719 );
not ( n58107 , n58106 );
not ( n58108 , n58107 );
and ( n58109 , n58108 , n52720 );
buf ( n58110 , RI15b60af8_1164);
and ( n58111 , n58110 , n52726 );
or ( n58112 , n58109 , C0 , n58111 );
buf ( n58113 , n58112 );
buf ( n58114 , n58113 );
buf ( n58115 , n31655 );
buf ( n58116 , n31655 );
buf ( n58117 , n30987 );
not ( n58118 , n34150 );
and ( n58119 , n58118 , n32712 );
not ( n58120 , n56192 );
and ( n58121 , n58120 , n32712 );
and ( n58122 , n32722 , n56192 );
or ( n58123 , n58121 , n58122 );
and ( n58124 , n58123 , n34150 );
or ( n58125 , n58119 , n58124 );
and ( n58126 , n58125 , n33381 );
not ( n58127 , n56200 );
not ( n58128 , n56192 );
and ( n58129 , n58128 , n32712 );
and ( n58130 , n42565 , n56192 );
or ( n58131 , n58129 , n58130 );
and ( n58132 , n58127 , n58131 );
and ( n58133 , n42565 , n56200 );
or ( n58134 , n58132 , n58133 );
and ( n58135 , n58134 , n33375 );
not ( n58136 , n32968 );
not ( n58137 , n56200 );
not ( n58138 , n56192 );
and ( n58139 , n58138 , n32712 );
and ( n58140 , n42565 , n56192 );
or ( n58141 , n58139 , n58140 );
and ( n58142 , n58137 , n58141 );
and ( n58143 , n42565 , n56200 );
or ( n58144 , n58142 , n58143 );
and ( n58145 , n58136 , n58144 );
not ( n58146 , n56220 );
not ( n58147 , n56222 );
and ( n58148 , n58147 , n58144 );
and ( n58149 , n42589 , n56222 );
or ( n58150 , n58148 , n58149 );
and ( n58151 , n58146 , n58150 );
and ( n58152 , n42597 , n56220 );
or ( n58153 , n58151 , n58152 );
and ( n58154 , n58153 , n32968 );
or ( n58155 , n58145 , n58154 );
and ( n58156 , n58155 , n33370 );
and ( n58157 , n32712 , n35062 );
or ( n58158 , C0 , n58126 , n58135 , n58156 , n58157 );
buf ( n58159 , n58158 );
buf ( n58160 , n58159 );
not ( n58161 , n34150 );
and ( n58162 , n58161 , n32821 );
not ( n58163 , n56239 );
and ( n58164 , n58163 , n32821 );
and ( n58165 , n32823 , n56239 );
or ( n58166 , n58164 , n58165 );
and ( n58167 , n58166 , n34150 );
or ( n58168 , n58162 , n58167 );
and ( n58169 , n58168 , n33381 );
not ( n58170 , n56247 );
not ( n58171 , n56239 );
and ( n58172 , n58171 , n32821 );
and ( n58173 , n41464 , n56239 );
or ( n58174 , n58172 , n58173 );
and ( n58175 , n58170 , n58174 );
and ( n58176 , n41464 , n56247 );
or ( n58177 , n58175 , n58176 );
and ( n58178 , n58177 , n33375 );
not ( n58179 , n32968 );
not ( n58180 , n56247 );
not ( n58181 , n56239 );
and ( n58182 , n58181 , n32821 );
and ( n58183 , n41464 , n56239 );
or ( n58184 , n58182 , n58183 );
and ( n58185 , n58180 , n58184 );
and ( n58186 , n41464 , n56247 );
or ( n58187 , n58185 , n58186 );
and ( n58188 , n58179 , n58187 );
not ( n58189 , n56267 );
not ( n58190 , n56269 );
and ( n58191 , n58190 , n58187 );
and ( n58192 , n41490 , n56269 );
or ( n58193 , n58191 , n58192 );
and ( n58194 , n58189 , n58193 );
and ( n58195 , n41500 , n56267 );
or ( n58196 , n58194 , n58195 );
and ( n58197 , n58196 , n32968 );
or ( n58198 , n58188 , n58197 );
and ( n58199 , n58198 , n33370 );
and ( n58200 , n32821 , n35062 );
or ( n58201 , C0 , n58169 , n58178 , n58199 , n58200 );
buf ( n58202 , n58201 );
buf ( n58203 , n58202 );
buf ( n58204 , n30987 );
buf ( n58205 , n30987 );
buf ( n58206 , RI15b47f58_320);
or ( n58207 , n44682 , n43774 );
and ( n58208 , n58206 , n58207 );
and ( n58209 , n54726 , n44695 );
or ( n58210 , n58208 , n58209 );
buf ( n58211 , n58210 );
buf ( n58212 , n58211 );
buf ( n58213 , n30987 );
buf ( n58214 , n31655 );
buf ( n58215 , n31655 );
not ( n58216 , n34150 );
and ( n58217 , n58216 , n32869 );
not ( n58218 , n57872 );
and ( n58219 , n58218 , n32869 );
and ( n58220 , n32889 , n57872 );
or ( n58221 , n58219 , n58220 );
and ( n58222 , n58221 , n34150 );
or ( n58223 , n58217 , n58222 );
and ( n58224 , n58223 , n33381 );
not ( n58225 , n57880 );
not ( n58226 , n57872 );
and ( n58227 , n58226 , n32869 );
and ( n58228 , n52819 , n57872 );
or ( n58229 , n58227 , n58228 );
and ( n58230 , n58225 , n58229 );
and ( n58231 , n52819 , n57880 );
or ( n58232 , n58230 , n58231 );
and ( n58233 , n58232 , n33375 );
not ( n58234 , n32968 );
not ( n58235 , n57880 );
not ( n58236 , n57872 );
and ( n58237 , n58236 , n32869 );
and ( n58238 , n52819 , n57872 );
or ( n58239 , n58237 , n58238 );
and ( n58240 , n58235 , n58239 );
and ( n58241 , n52819 , n57880 );
or ( n58242 , n58240 , n58241 );
and ( n58243 , n58234 , n58242 );
not ( n58244 , n57900 );
not ( n58245 , n57902 );
and ( n58246 , n58245 , n58242 );
and ( n58247 , n52845 , n57902 );
or ( n58248 , n58246 , n58247 );
and ( n58249 , n58244 , n58248 );
and ( n58250 , n52855 , n57900 );
or ( n58251 , n58249 , n58250 );
and ( n58252 , n58251 , n32968 );
or ( n58253 , n58243 , n58252 );
and ( n58254 , n58253 , n33370 );
and ( n58255 , n32869 , n35062 );
or ( n58256 , C0 , n58224 , n58233 , n58254 , n58255 );
buf ( n58257 , n58256 );
buf ( n58258 , n58257 );
buf ( n58259 , n30987 );
buf ( n58260 , n31655 );
buf ( n58261 , n31655 );
buf ( n58262 , n30987 );
buf ( n58263 , n31655 );
and ( n58264 , n33239 , n32528 );
not ( n58265 , n32598 );
and ( n58266 , n58265 , n33002 );
and ( n58267 , n48801 , n32598 );
or ( n58268 , n58266 , n58267 );
and ( n58269 , n58268 , n32890 );
not ( n58270 , n32919 );
and ( n58271 , n58270 , n33002 );
and ( n58272 , n48801 , n32919 );
or ( n58273 , n58271 , n58272 );
and ( n58274 , n58273 , n32924 );
not ( n58275 , n32953 );
and ( n58276 , n58275 , n33002 );
not ( n58277 , n32971 );
and ( n58278 , n58277 , n33129 );
xor ( n58279 , n33002 , n33003 );
and ( n58280 , n58279 , n32971 );
or ( n58281 , n58278 , n58280 );
and ( n58282 , n58281 , n32953 );
or ( n58283 , n58276 , n58282 );
and ( n58284 , n58283 , n33038 );
not ( n58285 , n33067 );
and ( n58286 , n58285 , n33002 );
not ( n58287 , n32970 );
not ( n58288 , n33071 );
and ( n58289 , n58288 , n33129 );
xor ( n58290 , n33130 , n33135 );
and ( n58291 , n58290 , n33071 );
or ( n58292 , n58289 , n58291 );
and ( n58293 , n58287 , n58292 );
and ( n58294 , n58279 , n32970 );
or ( n58295 , n58293 , n58294 );
and ( n58296 , n58295 , n33067 );
or ( n58297 , n58286 , n58296 );
and ( n58298 , n58297 , n33172 );
and ( n58299 , n33002 , n33204 );
or ( n58300 , n58269 , n58274 , n58284 , n58298 , n58299 );
and ( n58301 , n58300 , n33208 );
not ( n58302 , n32968 );
not ( n58303 , n33270 );
and ( n58304 , n58303 , n33329 );
xor ( n58305 , n33330 , n33335 );
and ( n58306 , n58305 , n33270 );
or ( n58307 , n58304 , n58306 );
and ( n58308 , n58302 , n58307 );
and ( n58309 , n33002 , n32968 );
or ( n58310 , n58308 , n58309 );
and ( n58311 , n58310 , n33370 );
and ( n58312 , n33002 , n33382 );
or ( n58313 , C0 , n58264 , n58301 , n58311 , C0 , n58312 );
buf ( n58314 , n58313 );
buf ( n58315 , n58314 );
buf ( n58316 , n30987 );
and ( n58317 , n32461 , n32500 );
not ( n58318 , n35211 );
and ( n58319 , n58318 , n37581 );
and ( n58320 , n31662 , n31769 );
xor ( n58321 , n31658 , n58320 );
and ( n58322 , n58321 , n35211 );
or ( n58323 , n58319 , n58322 );
and ( n58324 , n58323 , n32421 );
not ( n58325 , n35245 );
and ( n58326 , n58325 , n37581 );
and ( n58327 , n58321 , n35245 );
or ( n58328 , n58326 , n58327 );
and ( n58329 , n58328 , n32419 );
not ( n58330 , n35278 );
and ( n58331 , n58330 , n37581 );
not ( n58332 , n35295 );
and ( n58333 , n58332 , n47289 );
xor ( n58334 , n37581 , n49524 );
and ( n58335 , n58334 , n35295 );
or ( n58336 , n58333 , n58335 );
and ( n58337 , n58336 , n35278 );
or ( n58338 , n58331 , n58337 );
and ( n58339 , n58338 , n32417 );
not ( n58340 , n35331 );
and ( n58341 , n58340 , n37581 );
not ( n58342 , n35294 );
not ( n58343 , n45995 );
and ( n58344 , n58343 , n47289 );
xor ( n58345 , n49607 , n49610 );
and ( n58346 , n58345 , n45995 );
or ( n58347 , n58344 , n58346 );
and ( n58348 , n58342 , n58347 );
and ( n58349 , n58334 , n35294 );
or ( n58350 , n58348 , n58349 );
and ( n58351 , n58350 , n35331 );
or ( n58352 , n58341 , n58351 );
and ( n58353 , n58352 , n32415 );
and ( n58354 , n37581 , n35354 );
or ( n58355 , n58324 , n58329 , n58339 , n58353 , n58354 );
and ( n58356 , n58355 , n32456 );
not ( n58357 , n32475 );
not ( n58358 , n46060 );
and ( n58359 , n58358 , n49699 );
xor ( n58360 , n49700 , n49704 );
and ( n58361 , n58360 , n46060 );
or ( n58362 , n58359 , n58361 );
and ( n58363 , n58357 , n58362 );
and ( n58364 , n37581 , n32475 );
or ( n58365 , n58363 , n58364 );
and ( n58366 , n58365 , n32486 );
buf ( n58367 , n32489 );
and ( n58368 , n37581 , n35367 );
or ( n58369 , C0 , n58317 , n58356 , n58366 , n58367 , n58368 );
buf ( n58370 , n58369 );
buf ( n58371 , n58370 );
buf ( n58372 , n30987 );
buf ( n58373 , n31655 );
not ( n58374 , n35542 );
and ( n58375 , n58374 , n41841 );
and ( n58376 , n52795 , n35542 );
or ( n58377 , n58375 , n58376 );
buf ( n58378 , n58377 );
buf ( n58379 , n58378 );
buf ( n58380 , n31655 );
buf ( n58381 , n31655 );
buf ( n58382 , n30987 );
and ( n58383 , n33103 , n56362 );
and ( n58384 , n33101 , n58383 );
and ( n58385 , n33099 , n58384 );
and ( n58386 , n33097 , n58385 );
and ( n58387 , n33095 , n58386 );
and ( n58388 , n33093 , n58387 );
and ( n58389 , n33091 , n58388 );
and ( n58390 , n33089 , n58389 );
and ( n58391 , n33087 , n58390 );
and ( n58392 , n33085 , n58391 );
and ( n58393 , n33083 , n58392 );
and ( n58394 , n33081 , n58393 );
and ( n58395 , n33079 , n58394 );
and ( n58396 , n33077 , n58395 );
and ( n58397 , n33075 , n58396 );
xor ( n58398 , n32973 , n58397 );
and ( n58399 , n58398 , n33201 );
not ( n58400 , n41576 );
and ( n58401 , n58400 , n32973 );
not ( n58402 , n32547 );
buf ( n58403 , n58402 );
not ( n58404 , n58403 );
not ( n58405 , n58404 );
not ( n58406 , n32543 );
buf ( n58407 , n58406 );
buf ( n58408 , n58407 );
not ( n58409 , n58408 );
not ( n58410 , n58409 );
not ( n58411 , n32539 );
not ( n58412 , n58411 );
buf ( n58413 , n58412 );
buf ( n58414 , n58413 );
not ( n58415 , n58414 );
not ( n58416 , n58415 );
xor ( n58417 , n32535 , n32539 );
not ( n58418 , n58417 );
buf ( n58419 , n58418 );
buf ( n58420 , n58419 );
not ( n58421 , n58420 );
not ( n58422 , n58421 );
nor ( n58423 , n58405 , n58410 , n58416 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58424 , n32857 , n58423 );
nor ( n58425 , n58404 , n58410 , n58416 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58426 , n32859 , n58425 );
nor ( n58427 , n58405 , n58409 , n58416 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58428 , n32861 , n58427 );
nor ( n58429 , n58404 , n58409 , n58416 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58430 , n32863 , n58429 );
nor ( n58431 , n58405 , n58410 , n58415 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58432 , n32865 , n58431 );
nor ( n58433 , n58404 , n58410 , n58415 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58434 , n32867 , n58433 );
nor ( n58435 , n58405 , n58409 , n58415 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58436 , n32869 , n58435 );
nor ( n58437 , n58404 , n58409 , n58415 , n58422 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58438 , n32871 , n58437 );
nor ( n58439 , n58405 , n58410 , n58416 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58440 , n32873 , n58439 );
nor ( n58441 , n58404 , n58410 , n58416 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58442 , n32875 , n58441 );
nor ( n58443 , n58405 , n58409 , n58416 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58444 , n32877 , n58443 );
nor ( n58445 , n58404 , n58409 , n58416 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58446 , n32879 , n58445 );
nor ( n58447 , n58405 , n58410 , n58415 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58448 , n32881 , n58447 );
nor ( n58449 , n58404 , n58410 , n58415 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58450 , n32883 , n58449 );
nor ( n58451 , n58405 , n58409 , n58415 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58452 , n32885 , n58451 );
nor ( n58453 , n58404 , n58409 , n58415 , n58421 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n58454 , n32887 , n58453 );
or ( n58455 , n58424 , n58426 , n58428 , n58430 , n58432 , n58434 , n58436 , n58438 , n58440 , n58442 , n58444 , n58446 , n58448 , n58450 , n58452 , n58454 );
and ( n58456 , n32824 , n58423 );
and ( n58457 , n32826 , n58425 );
and ( n58458 , n32828 , n58427 );
and ( n58459 , n32830 , n58429 );
and ( n58460 , n32832 , n58431 );
and ( n58461 , n32834 , n58433 );
and ( n58462 , n32836 , n58435 );
and ( n58463 , n32838 , n58437 );
and ( n58464 , n32840 , n58439 );
and ( n58465 , n32842 , n58441 );
and ( n58466 , n32844 , n58443 );
and ( n58467 , n32846 , n58445 );
and ( n58468 , n32848 , n58447 );
and ( n58469 , n32850 , n58449 );
and ( n58470 , n32852 , n58451 );
and ( n58471 , n32854 , n58453 );
or ( n58472 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 );
and ( n58473 , n32791 , n58423 );
and ( n58474 , n32793 , n58425 );
and ( n58475 , n32795 , n58427 );
and ( n58476 , n32797 , n58429 );
and ( n58477 , n32799 , n58431 );
and ( n58478 , n32801 , n58433 );
and ( n58479 , n32803 , n58435 );
and ( n58480 , n32805 , n58437 );
and ( n58481 , n32807 , n58439 );
and ( n58482 , n32809 , n58441 );
and ( n58483 , n32811 , n58443 );
and ( n58484 , n32813 , n58445 );
and ( n58485 , n32815 , n58447 );
and ( n58486 , n32817 , n58449 );
and ( n58487 , n32819 , n58451 );
and ( n58488 , n32821 , n58453 );
or ( n58489 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 );
and ( n58490 , n32757 , n58423 );
and ( n58491 , n32759 , n58425 );
and ( n58492 , n32761 , n58427 );
and ( n58493 , n32763 , n58429 );
and ( n58494 , n32765 , n58431 );
and ( n58495 , n32767 , n58433 );
and ( n58496 , n32769 , n58435 );
and ( n58497 , n32771 , n58437 );
and ( n58498 , n32773 , n58439 );
and ( n58499 , n32775 , n58441 );
and ( n58500 , n32777 , n58443 );
and ( n58501 , n32779 , n58445 );
and ( n58502 , n32781 , n58447 );
and ( n58503 , n32783 , n58449 );
and ( n58504 , n32785 , n58451 );
and ( n58505 , n32787 , n58453 );
or ( n58506 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 );
and ( n58507 , n32723 , n58423 );
and ( n58508 , n32725 , n58425 );
and ( n58509 , n32727 , n58427 );
and ( n58510 , n32729 , n58429 );
and ( n58511 , n32731 , n58431 );
and ( n58512 , n32733 , n58433 );
and ( n58513 , n32735 , n58435 );
and ( n58514 , n32737 , n58437 );
and ( n58515 , n32739 , n58439 );
and ( n58516 , n32741 , n58441 );
and ( n58517 , n32743 , n58443 );
and ( n58518 , n32745 , n58445 );
and ( n58519 , n32747 , n58447 );
and ( n58520 , n32749 , n58449 );
and ( n58521 , n32751 , n58451 );
and ( n58522 , n32753 , n58453 );
or ( n58523 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 );
and ( n58524 , n32690 , n58423 );
and ( n58525 , n32692 , n58425 );
and ( n58526 , n32694 , n58427 );
and ( n58527 , n32696 , n58429 );
and ( n58528 , n32698 , n58431 );
and ( n58529 , n32700 , n58433 );
and ( n58530 , n32702 , n58435 );
and ( n58531 , n32704 , n58437 );
and ( n58532 , n32706 , n58439 );
and ( n58533 , n32708 , n58441 );
and ( n58534 , n32710 , n58443 );
and ( n58535 , n32712 , n58445 );
and ( n58536 , n32714 , n58447 );
and ( n58537 , n32716 , n58449 );
and ( n58538 , n32718 , n58451 );
and ( n58539 , n32720 , n58453 );
or ( n58540 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 );
and ( n58541 , n32657 , n58423 );
and ( n58542 , n32659 , n58425 );
and ( n58543 , n32661 , n58427 );
and ( n58544 , n32663 , n58429 );
and ( n58545 , n32665 , n58431 );
and ( n58546 , n32667 , n58433 );
and ( n58547 , n32669 , n58435 );
and ( n58548 , n32671 , n58437 );
and ( n58549 , n32673 , n58439 );
and ( n58550 , n32675 , n58441 );
and ( n58551 , n32677 , n58443 );
and ( n58552 , n32679 , n58445 );
and ( n58553 , n32681 , n58447 );
and ( n58554 , n32683 , n58449 );
and ( n58555 , n32685 , n58451 );
and ( n58556 , n32687 , n58453 );
or ( n58557 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 );
and ( n58558 , n32603 , n58423 );
and ( n58559 , n32607 , n58425 );
and ( n58560 , n32611 , n58427 );
and ( n58561 , n32615 , n58429 );
and ( n58562 , n32618 , n58431 );
and ( n58563 , n32622 , n58433 );
and ( n58564 , n32625 , n58435 );
and ( n58565 , n32628 , n58437 );
and ( n58566 , n32631 , n58439 );
and ( n58567 , n32634 , n58441 );
and ( n58568 , n32637 , n58443 );
and ( n58569 , n32640 , n58445 );
and ( n58570 , n32643 , n58447 );
and ( n58571 , n32646 , n58449 );
and ( n58572 , n32649 , n58451 );
and ( n58573 , n32652 , n58453 );
or ( n58574 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 );
and ( n58575 , n32857 , n55215 );
and ( n58576 , n32859 , n55217 );
and ( n58577 , n32861 , n55219 );
and ( n58578 , n32863 , n55221 );
and ( n58579 , n32865 , n55223 );
and ( n58580 , n32867 , n55225 );
and ( n58581 , n32869 , n55227 );
and ( n58582 , n32871 , n55229 );
and ( n58583 , n32873 , n55231 );
and ( n58584 , n32875 , n55233 );
and ( n58585 , n32877 , n55235 );
and ( n58586 , n32879 , n55237 );
and ( n58587 , n32881 , n55239 );
and ( n58588 , n32883 , n55241 );
and ( n58589 , n32885 , n55243 );
and ( n58590 , n32887 , n55245 );
or ( n58591 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 );
and ( n58592 , n58574 , n58591 );
and ( n58593 , n58557 , n58592 );
and ( n58594 , n58540 , n58593 );
and ( n58595 , n58523 , n58594 );
and ( n58596 , n58506 , n58595 );
and ( n58597 , n58489 , n58596 );
and ( n58598 , n58472 , n58597 );
xor ( n58599 , n58455 , n58598 );
and ( n58600 , n58599 , n41576 );
or ( n58601 , n58401 , n58600 );
and ( n58602 , n58601 , n33189 );
and ( n58603 , n32973 , n41592 );
or ( n58604 , n58399 , n58602 , n58603 );
and ( n58605 , n58604 , n33208 );
and ( n58606 , n32973 , n39805 );
or ( n58607 , C0 , n58605 , n58606 );
buf ( n58608 , n58607 );
buf ( n58609 , n58608 );
buf ( n58610 , n30987 );
not ( n58611 , n50828 );
not ( n58612 , n50834 );
and ( n58613 , n58612 , n40512 );
buf ( n58614 , RI15b53718_712);
and ( n58615 , n58614 , n50834 );
or ( n58616 , n58613 , n58615 );
and ( n58617 , n58611 , n58616 );
buf ( n58618 , RI15b5fb80_1131);
and ( n58619 , n58618 , n50828 );
or ( n58620 , n58617 , n58619 );
buf ( n58621 , n58620 );
buf ( n58622 , n58621 );
buf ( n58623 , n30987 );
xor ( n58624 , n41652 , n44779 );
and ( n58625 , n58624 , n31548 );
not ( n58626 , n44807 );
and ( n58627 , n58626 , n41652 );
and ( n58628 , n41934 , n44807 );
or ( n58629 , n58627 , n58628 );
and ( n58630 , n58629 , n31408 );
not ( n58631 , n44817 );
and ( n58632 , n58631 , n41652 );
not ( n58633 , n41835 );
buf ( n58634 , RI15b52db8_692);
and ( n58635 , n58633 , n58634 );
not ( n58636 , n42124 );
and ( n58637 , n58636 , n41944 );
xor ( n58638 , n42131 , n42139 );
and ( n58639 , n58638 , n42124 );
or ( n58640 , n58637 , n58639 );
and ( n58641 , n58640 , n41835 );
or ( n58642 , n58635 , n58641 );
and ( n58643 , n58642 , n44817 );
or ( n58644 , n58632 , n58643 );
and ( n58645 , n58644 , n31521 );
not ( n58646 , n45059 );
and ( n58647 , n58646 , n41652 );
and ( n58648 , n33590 , n45059 );
or ( n58649 , n58647 , n58648 );
and ( n58650 , n58649 , n31536 );
and ( n58651 , n41652 , n45148 );
or ( n58652 , n58625 , n58630 , n58645 , n58650 , n58651 );
and ( n58653 , n58652 , n31557 );
and ( n58654 , n41652 , n40154 );
or ( n58655 , C0 , n58653 , n58654 );
buf ( n58656 , n58655 );
buf ( n58657 , n58656 );
buf ( n58658 , n31655 );
not ( n58659 , n40163 );
and ( n58660 , n58659 , n31912 );
not ( n58661 , n50540 );
and ( n58662 , n58661 , n31912 );
and ( n58663 , n32200 , n50540 );
or ( n58664 , n58662 , n58663 );
and ( n58665 , n58664 , n40163 );
or ( n58666 , n58660 , n58665 );
and ( n58667 , n58666 , n32498 );
not ( n58668 , n50548 );
not ( n58669 , n50540 );
and ( n58670 , n58669 , n31912 );
and ( n58671 , n53243 , n50540 );
or ( n58672 , n58670 , n58671 );
and ( n58673 , n58668 , n58672 );
and ( n58674 , n53243 , n50548 );
or ( n58675 , n58673 , n58674 );
and ( n58676 , n58675 , n32473 );
not ( n58677 , n32475 );
not ( n58678 , n50548 );
not ( n58679 , n50540 );
and ( n58680 , n58679 , n31912 );
and ( n58681 , n53243 , n50540 );
or ( n58682 , n58680 , n58681 );
and ( n58683 , n58678 , n58682 );
and ( n58684 , n53243 , n50548 );
or ( n58685 , n58683 , n58684 );
and ( n58686 , n58677 , n58685 );
not ( n58687 , n50568 );
not ( n58688 , n50570 );
and ( n58689 , n58688 , n58685 );
and ( n58690 , n53269 , n50570 );
or ( n58691 , n58689 , n58690 );
and ( n58692 , n58687 , n58691 );
and ( n58693 , n53277 , n50568 );
or ( n58694 , n58692 , n58693 );
and ( n58695 , n58694 , n32475 );
or ( n58696 , n58686 , n58695 );
and ( n58697 , n58696 , n32486 );
and ( n58698 , n31912 , n41278 );
or ( n58699 , C0 , n58667 , n58676 , n58697 , n58698 );
buf ( n58700 , n58699 );
buf ( n58701 , n58700 );
buf ( n58702 , n30987 );
not ( n58703 , n35542 );
and ( n58704 , n58703 , n41866 );
buf ( n58705 , RI15b45d20_247);
and ( n58706 , n58705 , n35542 );
or ( n58707 , n58704 , n58706 );
buf ( n58708 , n58707 );
buf ( n58709 , n58708 );
not ( n58710 , n34150 );
and ( n58711 , n58710 , n32842 );
not ( n58712 , n56836 );
and ( n58713 , n58712 , n32842 );
and ( n58714 , n32856 , n56836 );
or ( n58715 , n58713 , n58714 );
and ( n58716 , n58715 , n34150 );
or ( n58717 , n58711 , n58716 );
and ( n58718 , n58717 , n33381 );
not ( n58719 , n56844 );
not ( n58720 , n56836 );
and ( n58721 , n58720 , n32842 );
and ( n58722 , n48160 , n56836 );
or ( n58723 , n58721 , n58722 );
and ( n58724 , n58719 , n58723 );
and ( n58725 , n48160 , n56844 );
or ( n58726 , n58724 , n58725 );
and ( n58727 , n58726 , n33375 );
not ( n58728 , n32968 );
not ( n58729 , n56844 );
not ( n58730 , n56836 );
and ( n58731 , n58730 , n32842 );
and ( n58732 , n48160 , n56836 );
or ( n58733 , n58731 , n58732 );
and ( n58734 , n58729 , n58733 );
and ( n58735 , n48160 , n56844 );
or ( n58736 , n58734 , n58735 );
and ( n58737 , n58728 , n58736 );
not ( n58738 , n56864 );
not ( n58739 , n56866 );
and ( n58740 , n58739 , n58736 );
and ( n58741 , n48186 , n56866 );
or ( n58742 , n58740 , n58741 );
and ( n58743 , n58738 , n58742 );
and ( n58744 , n48196 , n56864 );
or ( n58745 , n58743 , n58744 );
and ( n58746 , n58745 , n32968 );
or ( n58747 , n58737 , n58746 );
and ( n58748 , n58747 , n33370 );
and ( n58749 , n32842 , n35062 );
or ( n58750 , C0 , n58718 , n58727 , n58748 , n58749 );
buf ( n58751 , n58750 );
buf ( n58752 , n58751 );
buf ( n58753 , n30987 );
buf ( n58754 , n31655 );
buf ( n58755 , n31655 );
buf ( n58756 , n30987 );
buf ( n58757 , n30987 );
buf ( n58758 , n31655 );
buf ( n58759 , n31655 );
not ( n58760 , n34150 );
and ( n58761 , n58760 , n32834 );
and ( n58762 , n41389 , n32542 , n41390 , n32534 , n41391 );
not ( n58763 , n58762 );
and ( n58764 , n58763 , n32834 );
and ( n58765 , n32856 , n58762 );
or ( n58766 , n58764 , n58765 );
and ( n58767 , n58766 , n34150 );
or ( n58768 , n58761 , n58767 );
and ( n58769 , n58768 , n33381 );
and ( n58770 , n41400 , n34170 , n41401 , n34183 , C1 );
not ( n58771 , n58770 );
not ( n58772 , n58762 );
and ( n58773 , n58772 , n32834 );
and ( n58774 , n48160 , n58762 );
or ( n58775 , n58773 , n58774 );
and ( n58776 , n58771 , n58775 );
and ( n58777 , n48160 , n58770 );
or ( n58778 , n58776 , n58777 );
and ( n58779 , n58778 , n33375 );
not ( n58780 , n32968 );
not ( n58781 , n58770 );
not ( n58782 , n58762 );
and ( n58783 , n58782 , n32834 );
and ( n58784 , n48160 , n58762 );
or ( n58785 , n58783 , n58784 );
and ( n58786 , n58781 , n58785 );
and ( n58787 , n48160 , n58770 );
or ( n58788 , n58786 , n58787 );
and ( n58789 , n58780 , n58788 );
and ( n58790 , n41422 , n34333 , n41423 , n34354 , C1 );
not ( n58791 , n58790 );
and ( n58792 , n41426 , n34329 , n41427 , n34349 , C1 );
not ( n58793 , n58792 );
and ( n58794 , n58793 , n58788 );
and ( n58795 , n48186 , n58792 );
or ( n58796 , n58794 , n58795 );
and ( n58797 , n58791 , n58796 );
and ( n58798 , n48196 , n58790 );
or ( n58799 , n58797 , n58798 );
and ( n58800 , n58799 , n32968 );
or ( n58801 , n58789 , n58800 );
and ( n58802 , n58801 , n33370 );
and ( n58803 , n32834 , n35062 );
or ( n58804 , C0 , n58769 , n58779 , n58802 , n58803 );
buf ( n58805 , n58804 );
buf ( n58806 , n58805 );
buf ( n58807 , n30987 );
not ( n58808 , n31437 );
buf ( n58809 , RI15b52f20_695);
and ( n58810 , n58808 , n58809 );
not ( n58811 , n41809 );
and ( n58812 , n58811 , n41701 );
xor ( n58813 , n41813 , n41827 );
and ( n58814 , n58813 , n41809 );
or ( n58815 , n58812 , n58814 );
and ( n58816 , n58815 , n31437 );
or ( n58817 , n58810 , n58816 );
and ( n58818 , n58817 , n31468 );
not ( n58819 , n41837 );
and ( n58820 , n58819 , n58809 );
not ( n58821 , n42124 );
and ( n58822 , n58821 , n41992 );
xor ( n58823 , n42128 , n42142 );
and ( n58824 , n58823 , n42124 );
or ( n58825 , n58822 , n58824 );
and ( n58826 , n58825 , n41837 );
or ( n58827 , n58820 , n58826 );
and ( n58828 , n58827 , n31521 );
and ( n58829 , n58809 , n42158 );
or ( n58830 , n58818 , n58828 , n58829 );
and ( n58831 , n58830 , n31557 );
and ( n58832 , n58809 , n40154 );
or ( n58833 , C0 , n58831 , n58832 );
buf ( n58834 , n58833 );
buf ( n58835 , n58834 );
not ( n58836 , n40163 );
and ( n58837 , n58836 , n31778 );
not ( n58838 , n42171 );
and ( n58839 , n58838 , n31778 );
and ( n58840 , n32252 , n42171 );
or ( n58841 , n58839 , n58840 );
and ( n58842 , n58841 , n40163 );
or ( n58843 , n58837 , n58842 );
and ( n58844 , n58843 , n32498 );
not ( n58845 , n42180 );
not ( n58846 , n42171 );
and ( n58847 , n58846 , n31778 );
and ( n58848 , n40393 , n42171 );
or ( n58849 , n58847 , n58848 );
and ( n58850 , n58845 , n58849 );
and ( n58851 , n40393 , n42180 );
or ( n58852 , n58850 , n58851 );
and ( n58853 , n58852 , n32473 );
not ( n58854 , n32475 );
not ( n58855 , n42180 );
not ( n58856 , n42171 );
and ( n58857 , n58856 , n31778 );
and ( n58858 , n40393 , n42171 );
or ( n58859 , n58857 , n58858 );
and ( n58860 , n58855 , n58859 );
and ( n58861 , n40393 , n42180 );
or ( n58862 , n58860 , n58861 );
and ( n58863 , n58854 , n58862 );
not ( n58864 , n42206 );
not ( n58865 , n42209 );
and ( n58866 , n58865 , n58862 );
and ( n58867 , n40972 , n42209 );
or ( n58868 , n58866 , n58867 );
and ( n58869 , n58864 , n58868 );
and ( n58870 , n41267 , n42206 );
or ( n58871 , n58869 , n58870 );
and ( n58872 , n58871 , n32475 );
or ( n58873 , n58863 , n58872 );
and ( n58874 , n58873 , n32486 );
and ( n58875 , n31778 , n41278 );
or ( n58876 , C0 , n58844 , n58853 , n58874 , n58875 );
buf ( n58877 , n58876 );
buf ( n58878 , n58877 );
buf ( n58879 , n30987 );
buf ( n58880 , n31655 );
buf ( n58881 , n30987 );
buf ( n58882 , n31655 );
buf ( n58883 , RI15b47ee0_319);
not ( n58884 , n32598 );
and ( n58885 , n58883 , n58884 );
and ( n58886 , n58885 , n32890 );
not ( n58887 , n32919 );
and ( n58888 , n58887 , n58883 );
buf ( n58889 , n32919 );
or ( n58890 , n58888 , n58889 );
and ( n58891 , n58890 , n32924 );
not ( n58892 , n32953 );
and ( n58893 , n58883 , n58892 );
and ( n58894 , n58893 , n33038 );
not ( n58895 , n33067 );
and ( n58896 , n58895 , n58883 );
buf ( n58897 , n33067 );
or ( n58898 , n58896 , n58897 );
and ( n58899 , n58898 , n33172 );
and ( n58900 , n58883 , n33204 );
or ( n58901 , n58886 , n58891 , n58894 , n58899 , n58900 );
and ( n58902 , n58901 , n33208 );
or ( n58903 , n33370 , n33373 );
or ( n58904 , n58903 , n33375 );
or ( n58905 , n58904 , n33377 );
or ( n58906 , n58905 , n33379 );
or ( n58907 , n58906 , n33381 );
or ( n58908 , n58907 , n32528 );
and ( n58909 , n58883 , n58908 );
or ( n58910 , n35056 , n33372 );
buf ( n58911 , n58910 );
or ( n58912 , C0 , n58902 , n58909 , n58911 );
buf ( n58913 , n58912 );
buf ( n58914 , n58913 );
buf ( n58915 , n31655 );
buf ( n58916 , n30987 );
buf ( n58917 , n31655 );
buf ( n58918 , n30987 );
buf ( n58919 , RI15b543c0_739);
not ( n58920 , n58919 );
or ( n58921 , n37494 , n36596 );
and ( n58922 , n58920 , n58921 );
buf ( n58923 , n37497 );
or ( n58924 , n37496 , n37499 );
or ( n58925 , n58924 , n37501 );
or ( n58926 , n58925 , n37503 );
or ( n58927 , n58926 , n37505 );
and ( n58928 , n41522 , n58927 );
or ( n58929 , n58922 , n58923 , n58928 );
buf ( n58930 , n58929 );
buf ( n58931 , n58930 );
and ( n58932 , n47663 , n50275 );
not ( n58933 , n50278 );
and ( n58934 , n58933 , n47576 );
and ( n58935 , n47663 , n50278 );
or ( n58936 , n58934 , n58935 );
and ( n58937 , n58936 , n32421 );
not ( n58938 , n50002 );
and ( n58939 , n58938 , n47576 );
and ( n58940 , n47663 , n50002 );
or ( n58941 , n58939 , n58940 );
and ( n58942 , n58941 , n32419 );
not ( n58943 , n50289 );
and ( n58944 , n58943 , n47576 );
and ( n58945 , n47663 , n50289 );
or ( n58946 , n58944 , n58945 );
and ( n58947 , n58946 , n32417 );
not ( n58948 , n50008 );
and ( n58949 , n58948 , n47576 );
and ( n58950 , n47663 , n50008 );
or ( n58951 , n58949 , n58950 );
and ( n58952 , n58951 , n32415 );
not ( n58953 , n47331 );
and ( n58954 , n58953 , n47576 );
and ( n58955 , n47608 , n47331 );
or ( n58956 , n58954 , n58955 );
and ( n58957 , n58956 , n32413 );
not ( n58958 , n50067 );
and ( n58959 , n58958 , n47576 );
and ( n58960 , n47608 , n50067 );
or ( n58961 , n58959 , n58960 );
and ( n58962 , n58961 , n32411 );
not ( n58963 , n31728 );
and ( n58964 , n58963 , n47576 );
xor ( n58965 , n47608 , n47621 );
and ( n58966 , n58965 , n31728 );
or ( n58967 , n58964 , n58966 );
and ( n58968 , n58967 , n32253 );
not ( n58969 , n32283 );
and ( n58970 , n58969 , n47576 );
not ( n58971 , n31823 );
xor ( n58972 , n47663 , n47676 );
and ( n58973 , n58971 , n58972 );
xnor ( n58974 , n47713 , n47726 );
and ( n58975 , n58974 , n31823 );
or ( n58976 , n58973 , n58975 );
and ( n58977 , n58976 , n32283 );
or ( n58978 , n58970 , n58977 );
and ( n58979 , n58978 , n32398 );
and ( n58980 , n47713 , n50334 );
or ( n58981 , n58932 , n58937 , n58942 , n58947 , n58952 , n58957 , n58962 , n58968 , n58979 , n58980 );
and ( n58982 , n58981 , n32456 );
and ( n58983 , n37559 , n32489 );
and ( n58984 , n47576 , n50345 );
or ( n58985 , C0 , n58982 , n58983 , n58984 );
buf ( n58986 , n58985 );
buf ( n58987 , n58986 );
buf ( n58988 , n30987 );
not ( n58989 , n40163 );
and ( n58990 , n58989 , n31980 );
not ( n58991 , n52120 );
and ( n58992 , n58991 , n31980 );
and ( n58993 , n32165 , n52120 );
or ( n58994 , n58992 , n58993 );
and ( n58995 , n58994 , n40163 );
or ( n58996 , n58990 , n58995 );
and ( n58997 , n58996 , n32498 );
not ( n58998 , n52128 );
not ( n58999 , n52120 );
and ( n59000 , n58999 , n31980 );
not ( n59001 , n40373 );
and ( n59002 , n59001 , n40279 );
xor ( n59003 , n40381 , n40385 );
and ( n59004 , n59003 , n40373 );
or ( n59005 , n59002 , n59004 );
and ( n59006 , n59005 , n52120 );
or ( n59007 , n59000 , n59006 );
and ( n59008 , n58998 , n59007 );
and ( n59009 , n59005 , n52128 );
or ( n59010 , n59008 , n59009 );
and ( n59011 , n59010 , n32473 );
not ( n59012 , n32475 );
not ( n59013 , n52128 );
not ( n59014 , n52120 );
and ( n59015 , n59014 , n31980 );
and ( n59016 , n59005 , n52120 );
or ( n59017 , n59015 , n59016 );
and ( n59018 , n59013 , n59017 );
and ( n59019 , n59005 , n52128 );
or ( n59020 , n59018 , n59019 );
and ( n59021 , n59012 , n59020 );
not ( n59022 , n52148 );
not ( n59023 , n52150 );
and ( n59024 , n59023 , n59020 );
not ( n59025 , n40952 );
and ( n59026 , n59025 , n40863 );
xor ( n59027 , n40960 , n40964 );
and ( n59028 , n59027 , n40952 );
or ( n59029 , n59026 , n59028 );
and ( n59030 , n59029 , n52150 );
or ( n59031 , n59024 , n59030 );
and ( n59032 , n59022 , n59031 );
not ( n59033 , n41247 );
and ( n59034 , n59033 , n41162 );
xor ( n59035 , n41255 , n41259 );
and ( n59036 , n59035 , n41247 );
or ( n59037 , n59034 , n59036 );
and ( n59038 , n59037 , n52148 );
or ( n59039 , n59032 , n59038 );
and ( n59040 , n59039 , n32475 );
or ( n59041 , n59021 , n59040 );
and ( n59042 , n59041 , n32486 );
and ( n59043 , n31980 , n41278 );
or ( n59044 , C0 , n58997 , n59011 , n59042 , n59043 );
buf ( n59045 , n59044 );
buf ( n59046 , n59045 );
buf ( n59047 , n31655 );
not ( n59048 , n54795 );
not ( n59049 , n54797 );
not ( n59050 , n54800 );
and ( n59051 , n59050 , n54804 );
buf ( n59052 , n54800 );
or ( n59053 , n59051 , n59052 );
and ( n59054 , n59049 , n59053 );
buf ( n59055 , n59054 );
and ( n59056 , n59048 , n59055 );
buf ( n59057 , n54795 );
or ( n59058 , n59056 , n59057 );
and ( n59059 , n59058 , n37505 );
not ( n59060 , n31451 );
and ( n59061 , n59060 , n36596 );
and ( n59062 , n54815 , n37503 );
not ( n59063 , n54824 );
not ( n59064 , n54827 );
and ( n59065 , n59064 , n48294 );
buf ( n59066 , n54827 );
or ( n59067 , n59065 , n59066 );
and ( n59068 , n59063 , n59067 );
buf ( n59069 , n54824 );
or ( n59070 , n59068 , n59069 );
and ( n59071 , n59070 , n37501 );
not ( n59072 , n54800 );
not ( n59073 , n54838 );
not ( n59074 , n54842 );
not ( n59075 , n54845 );
not ( n59076 , n54847 );
not ( n59077 , n54849 );
and ( n59078 , n59076 , n59077 );
buf ( n59079 , n59078 );
and ( n59080 , n59075 , n59079 );
buf ( n59081 , n54845 );
or ( n59082 , n59080 , n59081 );
and ( n59083 , n59074 , n59082 );
buf ( n59084 , n54842 );
or ( n59085 , n59083 , n59084 );
and ( n59086 , n59073 , n59085 );
and ( n59087 , n31441 , n54838 );
or ( n59088 , n59086 , n59087 );
and ( n59089 , n59072 , n59088 );
buf ( n59090 , n54800 );
or ( n59091 , n59089 , n59090 );
and ( n59092 , n59091 , n37499 );
buf ( n59093 , n37494 );
and ( n59094 , n54792 , n37496 );
or ( n59095 , n59059 , n59061 , n59062 , n59071 , n59092 , n59093 , n59094 , C0 );
buf ( n59096 , n59095 );
buf ( n59097 , n59096 );
buf ( n59098 , n30987 );
buf ( n59099 , n30987 );
buf ( n59100 , n30987 );
buf ( n59101 , n31655 );
buf ( n59102 , n31655 );
not ( n59103 , n34150 );
and ( n59104 , n59103 , n32799 );
and ( n59105 , n32546 , n32542 , n41390 , n32534 , n41391 );
not ( n59106 , n59105 );
and ( n59107 , n59106 , n32799 );
and ( n59108 , n32823 , n59105 );
or ( n59109 , n59107 , n59108 );
and ( n59110 , n59109 , n34150 );
or ( n59111 , n59104 , n59110 );
and ( n59112 , n59111 , n33381 );
and ( n59113 , n34165 , n34170 , n41401 , n34183 , C1 );
not ( n59114 , n59113 );
not ( n59115 , n59105 );
and ( n59116 , n59115 , n32799 );
and ( n59117 , n41464 , n59105 );
or ( n59118 , n59116 , n59117 );
and ( n59119 , n59114 , n59118 );
and ( n59120 , n41464 , n59113 );
or ( n59121 , n59119 , n59120 );
and ( n59122 , n59121 , n33375 );
not ( n59123 , n32968 );
not ( n59124 , n59113 );
not ( n59125 , n59105 );
and ( n59126 , n59125 , n32799 );
and ( n59127 , n41464 , n59105 );
or ( n59128 , n59126 , n59127 );
and ( n59129 , n59124 , n59128 );
and ( n59130 , n41464 , n59113 );
or ( n59131 , n59129 , n59130 );
and ( n59132 , n59123 , n59131 );
and ( n59133 , n34325 , n34333 , n41423 , n34354 , C1 );
not ( n59134 , n59133 );
and ( n59135 , n34321 , n34329 , n41427 , n34349 , C1 );
not ( n59136 , n59135 );
and ( n59137 , n59136 , n59131 );
and ( n59138 , n41490 , n59135 );
or ( n59139 , n59137 , n59138 );
and ( n59140 , n59134 , n59139 );
and ( n59141 , n41500 , n59133 );
or ( n59142 , n59140 , n59141 );
and ( n59143 , n59142 , n32968 );
or ( n59144 , n59132 , n59143 );
and ( n59145 , n59144 , n33370 );
and ( n59146 , n32799 , n35062 );
or ( n59147 , C0 , n59112 , n59122 , n59145 , n59146 );
buf ( n59148 , n59147 );
buf ( n59149 , n59148 );
buf ( n59150 , n30987 );
buf ( n59151 , n30987 );
buf ( n59152 , n31655 );
and ( n59153 , n57836 , n33208 );
and ( n59154 , n57805 , n39805 );
or ( n59155 , C0 , n59153 , n59154 );
buf ( n59156 , n59155 );
buf ( n59157 , n59156 );
buf ( n59158 , n31655 );
buf ( n59159 , n31655 );
buf ( n59160 , n30987 );
and ( n59161 , n33443 , n48455 );
buf ( n59162 , n33443 );
and ( n59163 , n59162 , n31373 );
buf ( n59164 , n33443 );
and ( n59165 , n59164 , n31408 );
buf ( n59166 , n33443 );
and ( n59167 , n59166 , n31468 );
buf ( n59168 , n33443 );
and ( n59169 , n59168 , n31521 );
not ( n59170 , n39979 );
and ( n59171 , n59170 , n33443 );
and ( n59172 , n33649 , n39979 );
or ( n59173 , n59171 , n59172 );
and ( n59174 , n59173 , n31538 );
not ( n59175 , n45059 );
and ( n59176 , n59175 , n33443 );
and ( n59177 , n33649 , n45059 );
or ( n59178 , n59176 , n59177 );
and ( n59179 , n59178 , n31536 );
not ( n59180 , n33419 );
and ( n59181 , n59180 , n33443 );
xor ( n59182 , n33649 , n33666 );
and ( n59183 , n59182 , n33419 );
or ( n59184 , n59181 , n59183 );
and ( n59185 , n59184 , n31529 );
not ( n59186 , n33734 );
and ( n59187 , n59186 , n33443 );
not ( n59188 , n33533 );
xor ( n59189 , n33443 , n33666 );
and ( n59190 , n59188 , n59189 );
xor ( n59191 , n33884 , n33885 );
and ( n59192 , n59191 , n33533 );
or ( n59193 , n59190 , n59192 );
and ( n59194 , n59193 , n33734 );
or ( n59195 , n59187 , n59194 );
and ( n59196 , n59195 , n31527 );
and ( n59197 , n33884 , n48513 );
or ( n59198 , n59161 , n59163 , n59165 , n59167 , n59169 , n59174 , n59179 , n59185 , n59196 , n59197 );
and ( n59199 , n59198 , n31557 );
and ( n59200 , n35687 , n33973 );
and ( n59201 , n33443 , n48524 );
or ( n59202 , C0 , n59199 , n59200 , n59201 );
buf ( n59203 , n59202 );
buf ( n59204 , n59203 );
not ( n59205 , n35278 );
buf ( n59206 , RI15b5ef50_1105);
and ( n59207 , n59205 , n59206 );
not ( n59208 , n51396 );
and ( n59209 , n59208 , n51375 );
xor ( n59210 , n51375 , n51155 );
xor ( n59211 , n51358 , n51155 );
and ( n59212 , n53327 , n53336 );
and ( n59213 , n59211 , n59212 );
xor ( n59214 , n59210 , n59213 );
and ( n59215 , n59214 , n51396 );
or ( n59216 , n59209 , n59215 );
and ( n59217 , n59216 , n35278 );
or ( n59218 , n59207 , n59217 );
and ( n59219 , n59218 , n32417 );
not ( n59220 , n50008 );
and ( n59221 , n59220 , n59206 );
not ( n59222 , n51594 );
and ( n59223 , n59222 , n51578 );
xor ( n59224 , n51578 , n40244 );
xor ( n59225 , n51566 , n40244 );
xor ( n59226 , n51554 , n40244 );
xor ( n59227 , n51542 , n40244 );
xor ( n59228 , n51530 , n40244 );
xor ( n59229 , n51518 , n40244 );
xor ( n59230 , n51506 , n40244 );
and ( n59231 , n51597 , n51609 );
and ( n59232 , n59230 , n59231 );
and ( n59233 , n59229 , n59232 );
and ( n59234 , n59228 , n59233 );
and ( n59235 , n59227 , n59234 );
and ( n59236 , n59226 , n59235 );
and ( n59237 , n59225 , n59236 );
xor ( n59238 , n59224 , n59237 );
and ( n59239 , n59238 , n51594 );
or ( n59240 , n59223 , n59239 );
and ( n59241 , n59240 , n50008 );
or ( n59242 , n59221 , n59241 );
and ( n59243 , n59242 , n32415 );
and ( n59244 , n59206 , n48133 );
or ( n59245 , n59219 , n59243 , n59244 );
and ( n59246 , n59245 , n32456 );
and ( n59247 , n59206 , n47409 );
or ( n59248 , C0 , n59246 , n59247 );
buf ( n59249 , n59248 );
buf ( n59250 , n59249 );
buf ( n59251 , n30987 );
not ( n59252 , n35278 );
buf ( n59253 , RI15b5ec80_1099);
and ( n59254 , n59252 , n59253 );
not ( n59255 , n51396 );
and ( n59256 , n59255 , n51273 );
xor ( n59257 , n53331 , n53332 );
and ( n59258 , n59257 , n51396 );
or ( n59259 , n59256 , n59258 );
and ( n59260 , n59259 , n35278 );
or ( n59261 , n59254 , n59260 );
and ( n59262 , n59261 , n32417 );
not ( n59263 , n50008 );
and ( n59264 , n59263 , n59253 );
not ( n59265 , n51594 );
and ( n59266 , n59265 , n51506 );
xor ( n59267 , n59230 , n59231 );
and ( n59268 , n59267 , n51594 );
or ( n59269 , n59266 , n59268 );
and ( n59270 , n59269 , n50008 );
or ( n59271 , n59264 , n59270 );
and ( n59272 , n59271 , n32415 );
and ( n59273 , n59253 , n48133 );
or ( n59274 , n59262 , n59272 , n59273 );
and ( n59275 , n59274 , n32456 );
and ( n59276 , n59253 , n47409 );
or ( n59277 , C0 , n59275 , n59276 );
buf ( n59278 , n59277 );
buf ( n59279 , n59278 );
buf ( n59280 , n31655 );
and ( n59281 , n33773 , n48455 );
not ( n59282 , n48457 );
and ( n59283 , n59282 , n33437 );
and ( n59284 , n33773 , n48457 );
or ( n59285 , n59283 , n59284 );
and ( n59286 , n59285 , n31373 );
not ( n59287 , n44807 );
and ( n59288 , n59287 , n33437 );
and ( n59289 , n33773 , n44807 );
or ( n59290 , n59288 , n59289 );
and ( n59291 , n59290 , n31408 );
not ( n59292 , n48468 );
and ( n59293 , n59292 , n33437 );
and ( n59294 , n33773 , n48468 );
or ( n59295 , n59293 , n59294 );
and ( n59296 , n59295 , n31468 );
not ( n59297 , n44817 );
and ( n59298 , n59297 , n33437 );
and ( n59299 , n33773 , n44817 );
or ( n59300 , n59298 , n59299 );
and ( n59301 , n59300 , n31521 );
not ( n59302 , n39979 );
and ( n59303 , n59302 , n33437 );
and ( n59304 , n33535 , n39979 );
or ( n59305 , n59303 , n59304 );
and ( n59306 , n59305 , n31538 );
not ( n59307 , n45059 );
and ( n59308 , n59307 , n33437 );
and ( n59309 , n33535 , n45059 );
or ( n59310 , n59308 , n59309 );
and ( n59311 , n59310 , n31536 );
not ( n59312 , n33419 );
and ( n59313 , n59312 , n33437 );
xor ( n59314 , n33535 , n33552 );
xor ( n59315 , n59314 , n33682 );
and ( n59316 , n59315 , n33419 );
or ( n59317 , n59313 , n59316 );
and ( n59318 , n59317 , n31529 );
not ( n59319 , n33734 );
and ( n59320 , n59319 , n33437 );
not ( n59321 , n33533 );
xor ( n59322 , n33773 , n33552 );
xor ( n59323 , n59322 , n33800 );
and ( n59324 , n59321 , n59323 );
xor ( n59325 , n33860 , n33862 );
xor ( n59326 , n59325 , n33902 );
and ( n59327 , n59326 , n33533 );
or ( n59328 , n59324 , n59327 );
and ( n59329 , n59328 , n33734 );
or ( n59330 , n59320 , n59329 );
and ( n59331 , n59330 , n31527 );
and ( n59332 , n33860 , n48513 );
or ( n59333 , n59281 , n59286 , n59291 , n59296 , n59301 , n59306 , n59311 , n59318 , n59331 , n59332 );
and ( n59334 , n59333 , n31557 );
and ( n59335 , n34009 , n33973 );
and ( n59336 , n33437 , n48524 );
or ( n59337 , C0 , n59334 , n59335 , n59336 );
buf ( n59338 , n59337 );
buf ( n59339 , n59338 );
buf ( n59340 , n30987 );
and ( n59341 , n31584 , n31007 );
not ( n59342 , n31077 );
and ( n59343 , n59342 , n34008 );
buf ( n59344 , n59343 );
and ( n59345 , n59344 , n31373 );
not ( n59346 , n31402 );
and ( n59347 , n59346 , n34008 );
buf ( n59348 , n59347 );
and ( n59349 , n59348 , n31408 );
not ( n59350 , n31437 );
and ( n59351 , n59350 , n34008 );
not ( n59352 , n31455 );
and ( n59353 , n59352 , n34056 );
xor ( n59354 , n34008 , n34015 );
and ( n59355 , n59354 , n31455 );
or ( n59356 , n59353 , n59355 );
and ( n59357 , n59356 , n31437 );
or ( n59358 , n59351 , n59357 );
and ( n59359 , n59358 , n31468 );
not ( n59360 , n31497 );
and ( n59361 , n59360 , n34008 );
not ( n59362 , n31454 );
not ( n59363 , n31501 );
and ( n59364 , n59363 , n34056 );
xor ( n59365 , n34057 , n34067 );
and ( n59366 , n59365 , n31501 );
or ( n59367 , n59364 , n59366 );
and ( n59368 , n59362 , n59367 );
and ( n59369 , n59354 , n31454 );
or ( n59370 , n59368 , n59369 );
and ( n59371 , n59370 , n31497 );
or ( n59372 , n59361 , n59371 );
and ( n59373 , n59372 , n31521 );
and ( n59374 , n34008 , n31553 );
or ( n59375 , n59345 , n59349 , n59359 , n59373 , n59374 );
and ( n59376 , n59375 , n31557 );
not ( n59377 , n31452 );
not ( n59378 , n31619 );
and ( n59379 , n59378 , n34113 );
xor ( n59380 , n34114 , n34124 );
and ( n59381 , n59380 , n31619 );
or ( n59382 , n59379 , n59381 );
and ( n59383 , n59377 , n59382 );
and ( n59384 , n34008 , n31452 );
or ( n59385 , n59383 , n59384 );
and ( n59386 , n59385 , n31638 );
buf ( n59387 , n33973 );
and ( n59388 , n34008 , n31650 );
or ( n59389 , C0 , n59341 , n59376 , n59386 , n59387 , n59388 );
buf ( n59390 , n59389 );
buf ( n59391 , n59390 );
buf ( n59392 , n31655 );
buf ( n59393 , n31655 );
not ( n59394 , n33419 );
and ( n59395 , n59394 , n31560 );
and ( n59396 , n52398 , n57490 );
and ( n59397 , n52396 , n59396 );
xor ( n59398 , n52394 , n59397 );
xor ( n59399 , n52396 , n59396 );
and ( n59400 , n57491 , n57506 );
and ( n59401 , n59399 , n59400 );
xor ( n59402 , n59398 , n59401 );
and ( n59403 , n59402 , n33419 );
or ( n59404 , n59395 , n59403 );
and ( n59405 , n59404 , n31529 );
not ( n59406 , n33734 );
and ( n59407 , n59406 , n31560 );
not ( n59408 , n33533 );
and ( n59409 , n52398 , n57463 );
and ( n59410 , n52396 , n59409 );
xor ( n59411 , n52394 , n59410 );
xor ( n59412 , n52396 , n59409 );
and ( n59413 , n57464 , n57518 );
and ( n59414 , n59412 , n59413 );
xor ( n59415 , n59411 , n59414 );
and ( n59416 , n59408 , n59415 );
and ( n59417 , n52398 , n57523 );
and ( n59418 , n52396 , n59417 );
xor ( n59419 , n52394 , n59418 );
xor ( n59420 , n52396 , n59417 );
or ( n59421 , n57524 , n57529 );
or ( n59422 , n59420 , n59421 );
xnor ( n59423 , n59419 , n59422 );
and ( n59424 , n59423 , n33533 );
or ( n59425 , n59416 , n59424 );
and ( n59426 , n59425 , n33734 );
or ( n59427 , n59407 , n59426 );
and ( n59428 , n59427 , n31527 );
and ( n59429 , n31560 , n33942 );
or ( n59430 , n59405 , n59428 , n59429 );
and ( n59431 , n59430 , n31557 );
and ( n59432 , n31619 , n31643 );
not ( n59433 , n31452 );
and ( n59434 , n59433 , n31619 );
and ( n59435 , n31566 , n42440 );
and ( n59436 , n31565 , n59435 );
and ( n59437 , n31564 , n59436 );
and ( n59438 , n31563 , n59437 );
and ( n59439 , n31562 , n59438 );
and ( n59440 , n31561 , n59439 );
xor ( n59441 , n31560 , n59440 );
and ( n59442 , n59441 , n31452 );
or ( n59443 , n59434 , n59442 );
and ( n59444 , n59443 , n31638 );
and ( n59445 , n35375 , n33973 );
and ( n59446 , n31560 , n33978 );
or ( n59447 , C0 , n59431 , n59432 , n59444 , n59445 , n59446 );
buf ( n59448 , n59447 );
buf ( n59449 , n59448 );
buf ( n59450 , n30987 );
buf ( n59451 , n40222 );
buf ( n59452 , n31655 );
buf ( n59453 , n30987 );
not ( n59454 , n40163 );
and ( n59455 , n59454 , n31856 );
not ( n59456 , n40166 );
and ( n59457 , n59456 , n31856 );
and ( n59458 , n32235 , n40166 );
or ( n59459 , n59457 , n59458 );
and ( n59460 , n59459 , n40163 );
or ( n59461 , n59455 , n59460 );
and ( n59462 , n59461 , n32498 );
not ( n59463 , n40195 );
not ( n59464 , n40166 );
and ( n59465 , n59464 , n31856 );
and ( n59466 , n42188 , n40166 );
or ( n59467 , n59465 , n59466 );
and ( n59468 , n59463 , n59467 );
and ( n59469 , n42188 , n40195 );
or ( n59470 , n59468 , n59469 );
and ( n59471 , n59470 , n32473 );
not ( n59472 , n32475 );
not ( n59473 , n40195 );
not ( n59474 , n40166 );
and ( n59475 , n59474 , n31856 );
and ( n59476 , n42188 , n40166 );
or ( n59477 , n59475 , n59476 );
and ( n59478 , n59473 , n59477 );
and ( n59479 , n42188 , n40195 );
or ( n59480 , n59478 , n59479 );
and ( n59481 , n59472 , n59480 );
not ( n59482 , n40446 );
not ( n59483 , n40448 );
and ( n59484 , n59483 , n59480 );
and ( n59485 , n42216 , n40448 );
or ( n59486 , n59484 , n59485 );
and ( n59487 , n59482 , n59486 );
and ( n59488 , n42224 , n40446 );
or ( n59489 , n59487 , n59488 );
and ( n59490 , n59489 , n32475 );
or ( n59491 , n59481 , n59490 );
and ( n59492 , n59491 , n32486 );
and ( n59493 , n31856 , n41278 );
or ( n59494 , C0 , n59462 , n59471 , n59492 , n59493 );
buf ( n59495 , n59494 );
buf ( n59496 , n59495 );
and ( n59497 , n35433 , n39947 );
xor ( n59498 , n35431 , n59497 );
and ( n59499 , n59498 , n31550 );
not ( n59500 , n39979 );
and ( n59501 , n59500 , n35431 );
and ( n59502 , n40035 , n40129 );
xor ( n59503 , n45129 , n59502 );
and ( n59504 , n59503 , n39979 );
or ( n59505 , n59501 , n59504 );
and ( n59506 , n59505 , n31538 );
and ( n59507 , n35431 , n40143 );
or ( n59508 , n59499 , n59506 , n59507 );
and ( n59509 , n59508 , n31557 );
and ( n59510 , n35431 , n40154 );
or ( n59511 , C0 , n59509 , n59510 );
buf ( n59512 , n59511 );
buf ( n59513 , n59512 );
buf ( n59514 , n30987 );
buf ( n59515 , n31655 );
buf ( n59516 , n30987 );
xor ( n59517 , n33125 , n52216 );
and ( n59518 , n59517 , n33201 );
not ( n59519 , n41576 );
and ( n59520 , n59519 , n33125 );
buf ( n59521 , n32787 );
and ( n59522 , n59521 , n41576 );
or ( n59523 , n59520 , n59522 );
and ( n59524 , n59523 , n33189 );
and ( n59525 , n33125 , n41592 );
or ( n59526 , n59518 , n59524 , n59525 );
and ( n59527 , n59526 , n33208 );
and ( n59528 , n33125 , n39805 );
or ( n59529 , C0 , n59527 , n59528 );
buf ( n59530 , n59529 );
buf ( n59531 , n59530 );
buf ( n59532 , n30987 );
buf ( n59533 , n31655 );
not ( n59534 , n41532 );
and ( n59535 , n59534 , n34208 );
buf ( n59536 , RI15b53448_706);
and ( n59537 , n59536 , n41532 );
or ( n59538 , n59535 , n59537 );
buf ( n59539 , n59538 );
buf ( n59540 , n59539 );
buf ( n59541 , n30987 );
buf ( n59542 , n30987 );
buf ( n59543 , n31655 );
not ( n59544 , n32967 );
and ( n59545 , n59544 , n32515 );
buf ( n59546 , n32967 );
or ( n59547 , n59545 , n59546 );
and ( n59548 , n59547 , n33377 );
not ( n59549 , n57838 );
not ( n59550 , n57840 );
and ( n59551 , n59550 , n32515 );
buf ( n59552 , n57840 );
or ( n59553 , n59551 , n59552 );
and ( n59554 , n59553 , n33038 );
and ( n59555 , n32515 , n57852 );
or ( n59556 , n59554 , n59555 );
and ( n59557 , n59549 , n59556 );
buf ( n59558 , n57838 );
or ( n59559 , n59557 , n59558 );
and ( n59560 , n59559 , n33208 );
buf ( n59561 , n33375 );
not ( n59562 , n57860 );
and ( n59563 , n59562 , n33373 );
and ( n59564 , n32968 , n33370 );
or ( n59565 , C0 , C0 , C0 , n59548 , n59560 , n59561 , n59563 , n59564 , C0 , C0 );
buf ( n59566 , n59565 );
buf ( n59567 , n59566 );
buf ( n59568 , n31655 );
buf ( n59569 , n31655 );
buf ( n59570 , n31655 );
buf ( n59571 , n30987 );
not ( n59572 , n34150 );
and ( n59573 , n59572 , n32763 );
and ( n59574 , n41389 , n34153 , n32538 , n32534 , n41391 );
not ( n59575 , n59574 );
and ( n59576 , n59575 , n32763 );
and ( n59577 , n32789 , n59574 );
or ( n59578 , n59576 , n59577 );
and ( n59579 , n59578 , n34150 );
or ( n59580 , n59573 , n59579 );
and ( n59581 , n59580 , n33381 );
and ( n59582 , n41400 , n34171 , n34177 , n34183 , C1 );
not ( n59583 , n59582 );
not ( n59584 , n59574 );
and ( n59585 , n59584 , n32763 );
and ( n59586 , n34301 , n59574 );
or ( n59587 , n59585 , n59586 );
and ( n59588 , n59583 , n59587 );
and ( n59589 , n34301 , n59582 );
or ( n59590 , n59588 , n59589 );
and ( n59591 , n59590 , n33375 );
not ( n59592 , n32968 );
not ( n59593 , n59582 );
not ( n59594 , n59574 );
and ( n59595 , n59594 , n32763 );
and ( n59596 , n34301 , n59574 );
or ( n59597 , n59595 , n59596 );
and ( n59598 , n59593 , n59597 );
and ( n59599 , n34301 , n59582 );
or ( n59600 , n59598 , n59599 );
and ( n59601 , n59592 , n59600 );
and ( n59602 , n41422 , n34334 , n34344 , n34354 , C1 );
not ( n59603 , n59602 );
and ( n59604 , n41426 , n34357 , n34339 , n34349 , C1 );
not ( n59605 , n59604 );
and ( n59606 , n59605 , n59600 );
and ( n59607 , n34761 , n59604 );
or ( n59608 , n59606 , n59607 );
and ( n59609 , n59603 , n59608 );
and ( n59610 , n35050 , n59602 );
or ( n59611 , n59609 , n59610 );
and ( n59612 , n59611 , n32968 );
or ( n59613 , n59601 , n59612 );
and ( n59614 , n59613 , n33370 );
and ( n59615 , n32763 , n35062 );
or ( n59616 , C0 , n59581 , n59591 , n59614 , n59615 );
buf ( n59617 , n59616 );
buf ( n59618 , n59617 );
buf ( n59619 , n30987 );
buf ( n59620 , n40207 );
and ( n59621 , n46034 , n32500 );
not ( n59622 , n35211 );
and ( n59623 , n59622 , n37565 );
buf ( n59624 , n59623 );
and ( n59625 , n59624 , n32421 );
not ( n59626 , n35245 );
and ( n59627 , n59626 , n37565 );
buf ( n59628 , n59627 );
and ( n59629 , n59628 , n32419 );
not ( n59630 , n35278 );
and ( n59631 , n59630 , n37565 );
not ( n59632 , n35295 );
and ( n59633 , n59632 , n49595 );
xor ( n59634 , n37565 , n49533 );
and ( n59635 , n59634 , n35295 );
or ( n59636 , n59633 , n59635 );
and ( n59637 , n59636 , n35278 );
or ( n59638 , n59631 , n59637 );
and ( n59639 , n59638 , n32417 );
not ( n59640 , n35331 );
and ( n59641 , n59640 , n37565 );
not ( n59642 , n35294 );
not ( n59643 , n45995 );
and ( n59644 , n59643 , n49595 );
xor ( n59645 , n49596 , n49619 );
and ( n59646 , n59645 , n45995 );
or ( n59647 , n59644 , n59646 );
and ( n59648 , n59642 , n59647 );
and ( n59649 , n59634 , n35294 );
or ( n59650 , n59648 , n59649 );
and ( n59651 , n59650 , n35331 );
or ( n59652 , n59641 , n59651 );
and ( n59653 , n59652 , n32415 );
and ( n59654 , n37565 , n35354 );
or ( n59655 , n59625 , n59629 , n59639 , n59653 , n59654 );
and ( n59656 , n59655 , n32456 );
not ( n59657 , n32475 );
not ( n59658 , n46060 );
and ( n59659 , n59658 , n49685 );
xor ( n59660 , n49686 , n49713 );
and ( n59661 , n59660 , n46060 );
or ( n59662 , n59659 , n59661 );
and ( n59663 , n59657 , n59662 );
and ( n59664 , n37565 , n32475 );
or ( n59665 , n59663 , n59664 );
and ( n59666 , n59665 , n32486 );
buf ( n59667 , n32489 );
and ( n59668 , n37565 , n35367 );
or ( n59669 , C0 , n59621 , n59656 , n59666 , n59667 , n59668 );
buf ( n59670 , n59669 );
buf ( n59671 , n59670 );
buf ( n59672 , n31655 );
buf ( n59673 , n30987 );
not ( n59674 , n48765 );
and ( n59675 , n59674 , n33216 );
xor ( n59676 , n48771 , n49017 );
and ( n59677 , n59676 , n48765 );
or ( n59678 , n59675 , n59677 );
and ( n59679 , n59678 , n33180 );
not ( n59680 , n49054 );
and ( n59681 , n59680 , n33216 );
not ( n59682 , n48845 );
xor ( n59683 , n49061 , n49131 );
and ( n59684 , n59682 , n59683 );
xnor ( n59685 , n49170 , n49257 );
and ( n59686 , n59685 , n48845 );
or ( n59687 , n59684 , n59686 );
and ( n59688 , n59687 , n49054 );
or ( n59689 , n59681 , n59688 );
and ( n59690 , n59689 , n33178 );
and ( n59691 , n33216 , n49774 );
or ( n59692 , n59679 , n59690 , n59691 );
and ( n59693 , n59692 , n33208 );
and ( n59694 , n33283 , n33375 );
not ( n59695 , n32968 );
and ( n59696 , n59695 , n33283 );
and ( n59697 , n33222 , n53907 );
and ( n59698 , n33221 , n59697 );
and ( n59699 , n33220 , n59698 );
and ( n59700 , n33219 , n59699 );
and ( n59701 , n33218 , n59700 );
and ( n59702 , n33217 , n59701 );
xor ( n59703 , n33216 , n59702 );
and ( n59704 , n59703 , n32968 );
or ( n59705 , n59696 , n59704 );
and ( n59706 , n59705 , n33370 );
and ( n59707 , n32979 , n35056 );
and ( n59708 , n33216 , n49794 );
or ( n59709 , C0 , n59693 , n59694 , n59706 , n59707 , n59708 );
buf ( n59710 , n59709 );
buf ( n59711 , n59710 );
buf ( n59712 , n30987 );
buf ( n59713 , n31655 );
buf ( n59714 , n30987 );
buf ( n59715 , n30987 );
and ( n59716 , n46016 , n32500 );
not ( n59717 , n35211 );
and ( n59718 , n59717 , n37512 );
buf ( n59719 , n59718 );
and ( n59720 , n59719 , n32421 );
not ( n59721 , n35245 );
and ( n59722 , n59721 , n37512 );
buf ( n59723 , n59722 );
and ( n59724 , n59723 , n32419 );
not ( n59725 , n35278 );
and ( n59726 , n59725 , n37512 );
not ( n59727 , n35295 );
and ( n59728 , n59727 , n45995 );
and ( n59729 , n37531 , n49550 );
xor ( n59730 , n37512 , n59729 );
and ( n59731 , n59730 , n35295 );
or ( n59732 , n59728 , n59731 );
and ( n59733 , n59732 , n35278 );
or ( n59734 , n59726 , n59733 );
and ( n59735 , n59734 , n32417 );
not ( n59736 , n35331 );
and ( n59737 , n59736 , n37512 );
not ( n59738 , n35294 );
not ( n59739 , n45995 );
and ( n59740 , n49562 , n49636 );
xor ( n59741 , n59739 , n59740 );
buf ( n59742 , n45995 );
and ( n59743 , n59741 , n59742 );
buf ( n59744 , n59743 );
and ( n59745 , n59738 , n59744 );
and ( n59746 , n59730 , n35294 );
or ( n59747 , n59745 , n59746 );
and ( n59748 , n59747 , n35331 );
or ( n59749 , n59737 , n59748 );
and ( n59750 , n59749 , n32415 );
and ( n59751 , n37512 , n35354 );
or ( n59752 , n59720 , n59724 , n59735 , n59750 , n59751 );
and ( n59753 , n59752 , n32456 );
not ( n59754 , n32475 );
not ( n59755 , n46060 );
and ( n59756 , n49653 , n49730 );
xor ( n59757 , n59755 , n59756 );
buf ( n59758 , n46060 );
and ( n59759 , n59757 , n59758 );
buf ( n59760 , n59759 );
and ( n59761 , n59754 , n59760 );
and ( n59762 , n37512 , n32475 );
or ( n59763 , n59761 , n59762 );
and ( n59764 , n59763 , n32486 );
and ( n59765 , n37512 , n35367 );
or ( n59766 , C0 , n59716 , n59753 , n59764 , C0 , n59765 );
buf ( n59767 , n59766 );
buf ( n59768 , n59767 );
buf ( n59769 , n31655 );
not ( n59770 , n48765 );
and ( n59771 , n59770 , n33234 );
xor ( n59772 , n48789 , n48845 );
xor ( n59773 , n59772 , n48997 );
and ( n59774 , n59773 , n48765 );
or ( n59775 , n59771 , n59774 );
and ( n59776 , n59775 , n33180 );
not ( n59777 , n49054 );
and ( n59778 , n59777 , n33234 );
not ( n59779 , n48845 );
xor ( n59780 , n49079 , n48845 );
xor ( n59781 , n59780 , n49111 );
and ( n59782 , n59779 , n59781 );
xor ( n59783 , n49188 , n49190 );
xor ( n59784 , n59783 , n49237 );
and ( n59785 , n59784 , n48845 );
or ( n59786 , n59782 , n59785 );
and ( n59787 , n59786 , n49054 );
or ( n59788 , n59778 , n59787 );
and ( n59789 , n59788 , n33178 );
and ( n59790 , n33234 , n49774 );
or ( n59791 , n59776 , n59789 , n59790 );
and ( n59792 , n59791 , n33208 );
and ( n59793 , n33319 , n33375 );
not ( n59794 , n32968 );
and ( n59795 , n59794 , n33319 );
xor ( n59796 , n33234 , n49784 );
and ( n59797 , n59796 , n32968 );
or ( n59798 , n59795 , n59797 );
and ( n59799 , n59798 , n33370 );
and ( n59800 , n32997 , n35056 );
and ( n59801 , n33234 , n49794 );
or ( n59802 , C0 , n59792 , n59793 , n59799 , n59800 , n59801 );
buf ( n59803 , n59802 );
buf ( n59804 , n59803 );
buf ( n59805 , n31655 );
buf ( n59806 , n30987 );
buf ( n59807 , n30987 );
buf ( n59808 , n31655 );
not ( n59809 , n34150 );
and ( n59810 , n59809 , n32710 );
not ( n59811 , n56413 );
and ( n59812 , n59811 , n32710 );
and ( n59813 , n32722 , n56413 );
or ( n59814 , n59812 , n59813 );
and ( n59815 , n59814 , n34150 );
or ( n59816 , n59810 , n59815 );
and ( n59817 , n59816 , n33381 );
not ( n59818 , n56421 );
not ( n59819 , n56413 );
and ( n59820 , n59819 , n32710 );
and ( n59821 , n42565 , n56413 );
or ( n59822 , n59820 , n59821 );
and ( n59823 , n59818 , n59822 );
and ( n59824 , n42565 , n56421 );
or ( n59825 , n59823 , n59824 );
and ( n59826 , n59825 , n33375 );
not ( n59827 , n32968 );
not ( n59828 , n56421 );
not ( n59829 , n56413 );
and ( n59830 , n59829 , n32710 );
and ( n59831 , n42565 , n56413 );
or ( n59832 , n59830 , n59831 );
and ( n59833 , n59828 , n59832 );
and ( n59834 , n42565 , n56421 );
or ( n59835 , n59833 , n59834 );
and ( n59836 , n59827 , n59835 );
not ( n59837 , n56441 );
not ( n59838 , n56443 );
and ( n59839 , n59838 , n59835 );
and ( n59840 , n42589 , n56443 );
or ( n59841 , n59839 , n59840 );
and ( n59842 , n59837 , n59841 );
and ( n59843 , n42597 , n56441 );
or ( n59844 , n59842 , n59843 );
and ( n59845 , n59844 , n32968 );
or ( n59846 , n59836 , n59845 );
and ( n59847 , n59846 , n33370 );
and ( n59848 , n32710 , n35062 );
or ( n59849 , C0 , n59817 , n59826 , n59847 , n59848 );
buf ( n59850 , n59849 );
buf ( n59851 , n59850 );
not ( n59852 , n34150 );
and ( n59853 , n59852 , n32538 );
and ( n59854 , n34177 , n34150 );
or ( n59855 , n59853 , n59854 );
and ( n59856 , n59855 , n33381 );
not ( n59857 , n56687 );
not ( n59858 , n56464 );
and ( n59859 , n59858 , n32538 );
buf ( n59860 , n59859 );
and ( n59861 , n59857 , n59860 );
buf ( n59862 , n59861 );
and ( n59863 , n59862 , n33379 );
and ( n59864 , n34339 , n33375 );
not ( n59865 , n32968 );
and ( n59866 , n59865 , n34339 );
and ( n59867 , n34333 , n34325 );
xor ( n59868 , n34344 , n59867 );
not ( n59869 , n59868 );
buf ( n59870 , n59869 );
not ( n59871 , n59870 );
and ( n59872 , n59871 , n32968 );
or ( n59873 , n59866 , n59872 );
and ( n59874 , n59873 , n33370 );
and ( n59875 , n32538 , n56699 );
or ( n59876 , C0 , n59856 , n59863 , n59864 , n59874 , n59875 );
buf ( n59877 , n59876 );
buf ( n59878 , n59877 );
buf ( n59879 , n31655 );
buf ( n59880 , n30987 );
buf ( n59881 , n30987 );
not ( n59882 , n34150 );
and ( n59883 , n59882 , n32844 );
not ( n59884 , n56413 );
and ( n59885 , n59884 , n32844 );
and ( n59886 , n32856 , n56413 );
or ( n59887 , n59885 , n59886 );
and ( n59888 , n59887 , n34150 );
or ( n59889 , n59883 , n59888 );
and ( n59890 , n59889 , n33381 );
not ( n59891 , n56421 );
not ( n59892 , n56413 );
and ( n59893 , n59892 , n32844 );
and ( n59894 , n48160 , n56413 );
or ( n59895 , n59893 , n59894 );
and ( n59896 , n59891 , n59895 );
and ( n59897 , n48160 , n56421 );
or ( n59898 , n59896 , n59897 );
and ( n59899 , n59898 , n33375 );
not ( n59900 , n32968 );
not ( n59901 , n56421 );
not ( n59902 , n56413 );
and ( n59903 , n59902 , n32844 );
and ( n59904 , n48160 , n56413 );
or ( n59905 , n59903 , n59904 );
and ( n59906 , n59901 , n59905 );
and ( n59907 , n48160 , n56421 );
or ( n59908 , n59906 , n59907 );
and ( n59909 , n59900 , n59908 );
not ( n59910 , n56441 );
not ( n59911 , n56443 );
and ( n59912 , n59911 , n59908 );
and ( n59913 , n48186 , n56443 );
or ( n59914 , n59912 , n59913 );
and ( n59915 , n59910 , n59914 );
and ( n59916 , n48196 , n56441 );
or ( n59917 , n59915 , n59916 );
and ( n59918 , n59917 , n32968 );
or ( n59919 , n59909 , n59918 );
and ( n59920 , n59919 , n33370 );
and ( n59921 , n32844 , n35062 );
or ( n59922 , C0 , n59890 , n59899 , n59920 , n59921 );
buf ( n59923 , n59922 );
buf ( n59924 , n59923 );
buf ( n59925 , n31655 );
buf ( n59926 , n31655 );
buf ( n59927 , n54724 );
buf ( n59928 , n30987 );
buf ( n59929 , n31655 );
buf ( n59930 , n31655 );
buf ( n59931 , n30987 );
not ( n59932 , n34150 );
and ( n59933 , n59932 , n32733 );
not ( n59934 , n58762 );
and ( n59935 , n59934 , n32733 );
and ( n59936 , n32755 , n58762 );
or ( n59937 , n59935 , n59936 );
and ( n59938 , n59937 , n34150 );
or ( n59939 , n59933 , n59938 );
and ( n59940 , n59939 , n33381 );
not ( n59941 , n58770 );
not ( n59942 , n58762 );
and ( n59943 , n59942 , n32733 );
and ( n59944 , n35083 , n58762 );
or ( n59945 , n59943 , n59944 );
and ( n59946 , n59941 , n59945 );
and ( n59947 , n35083 , n58770 );
or ( n59948 , n59946 , n59947 );
and ( n59949 , n59948 , n33375 );
not ( n59950 , n32968 );
not ( n59951 , n58770 );
not ( n59952 , n58762 );
and ( n59953 , n59952 , n32733 );
and ( n59954 , n35083 , n58762 );
or ( n59955 , n59953 , n59954 );
and ( n59956 , n59951 , n59955 );
and ( n59957 , n35083 , n58770 );
or ( n59958 , n59956 , n59957 );
and ( n59959 , n59950 , n59958 );
not ( n59960 , n58790 );
not ( n59961 , n58792 );
and ( n59962 , n59961 , n59958 );
and ( n59963 , n35107 , n58792 );
or ( n59964 , n59962 , n59963 );
and ( n59965 , n59960 , n59964 );
and ( n59966 , n35115 , n58790 );
or ( n59967 , n59965 , n59966 );
and ( n59968 , n59967 , n32968 );
or ( n59969 , n59959 , n59968 );
and ( n59970 , n59969 , n33370 );
and ( n59971 , n32733 , n35062 );
or ( n59972 , C0 , n59940 , n59949 , n59970 , n59971 );
buf ( n59973 , n59972 );
buf ( n59974 , n59973 );
buf ( n59975 , RI15b529f8_684);
and ( n59976 , n59975 , n31645 );
not ( n59977 , n45274 );
buf ( n59978 , RI15b54000_731);
and ( n59979 , n59977 , n59978 );
buf ( n59980 , n59979 );
and ( n59981 , n59980 , n31373 );
not ( n59982 , n45280 );
and ( n59983 , n59982 , n59978 );
not ( n59984 , n45766 );
and ( n59985 , n59984 , n45711 );
xor ( n59986 , n45888 , n45891 );
and ( n59987 , n59986 , n45766 );
or ( n59988 , n59985 , n59987 );
and ( n59989 , n59988 , n45280 );
or ( n59990 , n59983 , n59989 );
and ( n59991 , n59990 , n31468 );
and ( n59992 , n59978 , n45802 );
or ( n59993 , n59981 , n59991 , n59992 );
and ( n59994 , n59993 , n31557 );
and ( n59995 , n59978 , n45808 );
or ( n59996 , C0 , n59976 , n59994 , n59995 );
buf ( n59997 , n59996 );
buf ( n59998 , n59997 );
buf ( n59999 , n31655 );
buf ( n60000 , n30987 );
buf ( n60001 , n30987 );
not ( n60002 , n40163 );
and ( n60003 , n60002 , n31941 );
not ( n60004 , n45227 );
and ( n60005 , n60004 , n31941 );
and ( n60006 , n32183 , n45227 );
or ( n60007 , n60005 , n60006 );
and ( n60008 , n60007 , n40163 );
or ( n60009 , n60003 , n60008 );
and ( n60010 , n60009 , n32498 );
not ( n60011 , n45235 );
not ( n60012 , n45227 );
and ( n60013 , n60012 , n31941 );
and ( n60014 , n45178 , n45227 );
or ( n60015 , n60013 , n60014 );
and ( n60016 , n60011 , n60015 );
and ( n60017 , n45178 , n45235 );
or ( n60018 , n60016 , n60017 );
and ( n60019 , n60018 , n32473 );
not ( n60020 , n32475 );
not ( n60021 , n45235 );
not ( n60022 , n45227 );
and ( n60023 , n60022 , n31941 );
and ( n60024 , n45178 , n45227 );
or ( n60025 , n60023 , n60024 );
and ( n60026 , n60021 , n60025 );
and ( n60027 , n45178 , n45235 );
or ( n60028 , n60026 , n60027 );
and ( n60029 , n60020 , n60028 );
not ( n60030 , n45255 );
not ( n60031 , n45257 );
and ( n60032 , n60031 , n60028 );
and ( n60033 , n45206 , n45257 );
or ( n60034 , n60032 , n60033 );
and ( n60035 , n60030 , n60034 );
and ( n60036 , n45214 , n45255 );
or ( n60037 , n60035 , n60036 );
and ( n60038 , n60037 , n32475 );
or ( n60039 , n60029 , n60038 );
and ( n60040 , n60039 , n32486 );
and ( n60041 , n31941 , n41278 );
or ( n60042 , C0 , n60010 , n60019 , n60040 , n60041 );
buf ( n60043 , n60042 );
buf ( n60044 , n60043 );
buf ( n60045 , n31655 );
buf ( n60046 , n30987 );
xor ( n60047 , n34050 , n39932 );
and ( n60048 , n60047 , n31550 );
not ( n60049 , n39979 );
and ( n60050 , n60049 , n34050 );
and ( n60051 , n31173 , n42330 );
and ( n60052 , n31175 , n42332 );
and ( n60053 , n31177 , n42334 );
and ( n60054 , n31179 , n42336 );
and ( n60055 , n31181 , n42338 );
and ( n60056 , n31183 , n42340 );
and ( n60057 , n31185 , n42342 );
and ( n60058 , n31187 , n42344 );
and ( n60059 , n31189 , n42346 );
and ( n60060 , n31191 , n42348 );
and ( n60061 , n31193 , n42350 );
and ( n60062 , n31195 , n42352 );
and ( n60063 , n31197 , n42354 );
and ( n60064 , n31199 , n42356 );
and ( n60065 , n31201 , n42358 );
and ( n60066 , n31203 , n42360 );
or ( n60067 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 );
and ( n60068 , n60067 , n39979 );
or ( n60069 , n60050 , n60068 );
and ( n60070 , n60069 , n31538 );
and ( n60071 , n34050 , n40143 );
or ( n60072 , n60048 , n60070 , n60071 );
and ( n60073 , n60072 , n31557 );
and ( n60074 , n34050 , n40154 );
or ( n60075 , C0 , n60073 , n60074 );
buf ( n60076 , n60075 );
buf ( n60077 , n60076 );
not ( n60078 , n40163 );
and ( n60079 , n60078 , n31852 );
not ( n60080 , n42238 );
and ( n60081 , n60080 , n31852 );
and ( n60082 , n32235 , n42238 );
or ( n60083 , n60081 , n60082 );
and ( n60084 , n60083 , n40163 );
or ( n60085 , n60079 , n60084 );
and ( n60086 , n60085 , n32498 );
not ( n60087 , n42247 );
not ( n60088 , n42238 );
and ( n60089 , n60088 , n31852 );
and ( n60090 , n42188 , n42238 );
or ( n60091 , n60089 , n60090 );
and ( n60092 , n60087 , n60091 );
and ( n60093 , n42188 , n42247 );
or ( n60094 , n60092 , n60093 );
and ( n60095 , n60094 , n32473 );
not ( n60096 , n32475 );
not ( n60097 , n42247 );
not ( n60098 , n42238 );
and ( n60099 , n60098 , n31852 );
and ( n60100 , n42188 , n42238 );
or ( n60101 , n60099 , n60100 );
and ( n60102 , n60097 , n60101 );
and ( n60103 , n42188 , n42247 );
or ( n60104 , n60102 , n60103 );
and ( n60105 , n60096 , n60104 );
not ( n60106 , n42273 );
not ( n60107 , n42276 );
and ( n60108 , n60107 , n60104 );
and ( n60109 , n42216 , n42276 );
or ( n60110 , n60108 , n60109 );
and ( n60111 , n60106 , n60110 );
and ( n60112 , n42224 , n42273 );
or ( n60113 , n60111 , n60112 );
and ( n60114 , n60113 , n32475 );
or ( n60115 , n60105 , n60114 );
and ( n60116 , n60115 , n32486 );
and ( n60117 , n31852 , n41278 );
or ( n60118 , C0 , n60086 , n60095 , n60116 , n60117 );
buf ( n60119 , n60118 );
buf ( n60120 , n60119 );
buf ( n60121 , n30987 );
buf ( n60122 , n31655 );
buf ( n60123 , n30987 );
not ( n60124 , n34150 );
and ( n60125 , n60124 , n32727 );
and ( n60126 , n32546 , n34153 , n32538 , n32534 , n41391 );
not ( n60127 , n60126 );
and ( n60128 , n60127 , n32727 );
and ( n60129 , n32755 , n60126 );
or ( n60130 , n60128 , n60129 );
and ( n60131 , n60130 , n34150 );
or ( n60132 , n60125 , n60131 );
and ( n60133 , n60132 , n33381 );
and ( n60134 , n34165 , n34171 , n34177 , n34183 , C1 );
not ( n60135 , n60134 );
not ( n60136 , n60126 );
and ( n60137 , n60136 , n32727 );
and ( n60138 , n35083 , n60126 );
or ( n60139 , n60137 , n60138 );
and ( n60140 , n60135 , n60139 );
and ( n60141 , n35083 , n60134 );
or ( n60142 , n60140 , n60141 );
and ( n60143 , n60142 , n33375 );
not ( n60144 , n32968 );
not ( n60145 , n60134 );
not ( n60146 , n60126 );
and ( n60147 , n60146 , n32727 );
and ( n60148 , n35083 , n60126 );
or ( n60149 , n60147 , n60148 );
and ( n60150 , n60145 , n60149 );
and ( n60151 , n35083 , n60134 );
or ( n60152 , n60150 , n60151 );
and ( n60153 , n60144 , n60152 );
and ( n60154 , n34325 , n34334 , n34344 , n34354 , C1 );
not ( n60155 , n60154 );
and ( n60156 , n34321 , n34357 , n34339 , n34349 , C1 );
not ( n60157 , n60156 );
and ( n60158 , n60157 , n60152 );
and ( n60159 , n35107 , n60156 );
or ( n60160 , n60158 , n60159 );
and ( n60161 , n60155 , n60160 );
and ( n60162 , n35115 , n60154 );
or ( n60163 , n60161 , n60162 );
and ( n60164 , n60163 , n32968 );
or ( n60165 , n60153 , n60164 );
and ( n60166 , n60165 , n33370 );
and ( n60167 , n32727 , n35062 );
or ( n60168 , C0 , n60133 , n60143 , n60166 , n60167 );
buf ( n60169 , n60168 );
buf ( n60170 , n60169 );
buf ( n60171 , n30987 );
buf ( n60172 , n31655 );
not ( n60173 , n46356 );
and ( n60174 , n60173 , n31278 );
not ( n60175 , n55473 );
and ( n60176 , n60175 , n31278 );
and ( n60177 , n31306 , n55473 );
or ( n60178 , n60176 , n60177 );
and ( n60179 , n60178 , n46356 );
or ( n60180 , n60174 , n60179 );
and ( n60181 , n60180 , n31649 );
not ( n60182 , n55481 );
not ( n60183 , n55473 );
and ( n60184 , n60183 , n31278 );
and ( n60185 , n58061 , n55473 );
or ( n60186 , n60184 , n60185 );
and ( n60187 , n60182 , n60186 );
and ( n60188 , n58061 , n55481 );
or ( n60189 , n60187 , n60188 );
and ( n60190 , n60189 , n31643 );
not ( n60191 , n31452 );
not ( n60192 , n55481 );
not ( n60193 , n55473 );
and ( n60194 , n60193 , n31278 );
and ( n60195 , n58061 , n55473 );
or ( n60196 , n60194 , n60195 );
and ( n60197 , n60192 , n60196 );
and ( n60198 , n58061 , n55481 );
or ( n60199 , n60197 , n60198 );
and ( n60200 , n60191 , n60199 );
not ( n60201 , n55501 );
not ( n60202 , n55503 );
and ( n60203 , n60202 , n60199 );
and ( n60204 , n58085 , n55503 );
or ( n60205 , n60203 , n60204 );
and ( n60206 , n60201 , n60205 );
and ( n60207 , n58093 , n55501 );
or ( n60208 , n60206 , n60207 );
and ( n60209 , n60208 , n31452 );
or ( n60210 , n60200 , n60209 );
and ( n60211 , n60210 , n31638 );
and ( n60212 , n31278 , n47277 );
or ( n60213 , C0 , n60181 , n60190 , n60211 , n60212 );
buf ( n60214 , n60213 );
buf ( n60215 , n60214 );
and ( n60216 , n55319 , n32494 );
not ( n60217 , n46083 );
buf ( n60218 , RI15b5f838_1124);
and ( n60219 , n60217 , n60218 );
not ( n60220 , n46290 );
and ( n60221 , n60220 , n46104 );
xor ( n60222 , n46305 , n46307 );
and ( n60223 , n60222 , n46290 );
or ( n60224 , n60221 , n60223 );
and ( n60225 , n60224 , n46083 );
or ( n60226 , n60219 , n60225 );
and ( n60227 , n60226 , n32421 );
not ( n60228 , n46326 );
and ( n60229 , n60228 , n60218 );
and ( n60230 , n60224 , n46326 );
or ( n60231 , n60229 , n60230 );
and ( n60232 , n60231 , n32417 );
and ( n60233 , n60218 , n46340 );
or ( n60234 , n60227 , n60232 , n60233 );
and ( n60235 , n60234 , n32456 );
and ( n60236 , n60218 , n46349 );
or ( n60237 , C0 , n60216 , n60235 , n60236 );
buf ( n60238 , n60237 );
buf ( n60239 , n60238 );
buf ( n60240 , n31655 );
buf ( n60241 , n31655 );
buf ( n60242 , n30987 );
buf ( n60243 , n31655 );
buf ( n60244 , n31655 );
buf ( n60245 , n30987 );
not ( n60246 , n50828 );
not ( n60247 , n50834 );
and ( n60248 , n60247 , n40491 );
buf ( n60249 , RI15b53880_715);
and ( n60250 , n60249 , n50834 );
or ( n60251 , n60248 , n60250 );
and ( n60252 , n60246 , n60251 );
buf ( n60253 , RI15b5fce8_1134);
and ( n60254 , n60253 , n50828 );
or ( n60255 , n60252 , n60254 );
buf ( n60256 , n60255 );
buf ( n60257 , n60256 );
buf ( n60258 , n30987 );
xor ( n60259 , n33079 , n58394 );
and ( n60260 , n60259 , n33201 );
not ( n60261 , n41576 );
and ( n60262 , n60261 , n33079 );
xor ( n60263 , n58506 , n58595 );
and ( n60264 , n60263 , n41576 );
or ( n60265 , n60262 , n60264 );
and ( n60266 , n60265 , n33189 );
and ( n60267 , n33079 , n41592 );
or ( n60268 , n60260 , n60266 , n60267 );
and ( n60269 , n60268 , n33208 );
and ( n60270 , n33079 , n39805 );
or ( n60271 , C0 , n60269 , n60270 );
buf ( n60272 , n60271 );
buf ( n60273 , n60272 );
buf ( n60274 , n30987 );
buf ( n60275 , n30987 );
buf ( n60276 , n31655 );
buf ( n60277 , n31655 );
xor ( n60278 , n39376 , n39369 );
and ( n60279 , n60278 , n33199 );
not ( n60280 , n48648 );
and ( n60281 , n60280 , n39376 );
and ( n60282 , n34195 , n48648 );
or ( n60283 , n60281 , n60282 );
and ( n60284 , n60283 , n32924 );
not ( n60285 , n48660 );
and ( n60286 , n60285 , n39376 );
not ( n60287 , n39584 );
and ( n60288 , n60287 , n39367 );
and ( n60289 , n39783 , n39584 );
or ( n60290 , n60288 , n60289 );
and ( n60291 , n60290 , n48660 );
or ( n60292 , n60286 , n60291 );
and ( n60293 , n60292 , n33172 );
not ( n60294 , n48730 );
and ( n60295 , n60294 , n39376 );
and ( n60296 , n48959 , n48730 );
or ( n60297 , n60295 , n60296 );
and ( n60298 , n60297 , n33187 );
and ( n60299 , n39376 , n54713 );
or ( n60300 , n60279 , n60284 , n60293 , n60298 , n60299 );
and ( n60301 , n60300 , n33208 );
and ( n60302 , n39376 , n39805 );
or ( n60303 , C0 , n60301 , n60302 );
buf ( n60304 , n60303 );
buf ( n60305 , n60304 );
and ( n60306 , n47283 , n47299 );
and ( n60307 , n49599 , n60306 );
and ( n60308 , n49597 , n60307 );
and ( n60309 , n49595 , n60308 );
and ( n60310 , n49593 , n60309 );
and ( n60311 , n49591 , n60310 );
and ( n60312 , n49589 , n60311 );
and ( n60313 , n49587 , n60312 );
and ( n60314 , n49585 , n60313 );
and ( n60315 , n49583 , n60314 );
and ( n60316 , n49581 , n60315 );
and ( n60317 , n49579 , n60316 );
and ( n60318 , n49577 , n60317 );
and ( n60319 , n49575 , n60318 );
and ( n60320 , n49573 , n60319 );
and ( n60321 , n49571 , n60320 );
and ( n60322 , n49569 , n60321 );
and ( n60323 , n49567 , n60322 );
and ( n60324 , n49565 , n60323 );
xor ( n60325 , n49563 , n60324 );
and ( n60326 , n60325 , n32433 );
not ( n60327 , n47331 );
and ( n60328 , n60327 , n49563 );
not ( n60329 , n31674 );
buf ( n60330 , n60329 );
not ( n60331 , n60330 );
not ( n60332 , n60331 );
not ( n60333 , n31670 );
buf ( n60334 , n60333 );
buf ( n60335 , n60334 );
not ( n60336 , n60335 );
not ( n60337 , n60336 );
not ( n60338 , n31666 );
not ( n60339 , n60338 );
buf ( n60340 , n60339 );
buf ( n60341 , n60340 );
not ( n60342 , n60341 );
not ( n60343 , n60342 );
xor ( n60344 , n31662 , n31666 );
not ( n60345 , n60344 );
buf ( n60346 , n60345 );
buf ( n60347 , n60346 );
not ( n60348 , n60347 );
not ( n60349 , n60348 );
nor ( n60350 , n60332 , n60337 , n60343 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60351 , n31826 , n60350 );
nor ( n60352 , n60331 , n60337 , n60343 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60353 , n31828 , n60352 );
nor ( n60354 , n60332 , n60336 , n60343 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60355 , n31830 , n60354 );
nor ( n60356 , n60331 , n60336 , n60343 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60357 , n31832 , n60356 );
nor ( n60358 , n60332 , n60337 , n60342 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60359 , n31834 , n60358 );
nor ( n60360 , n60331 , n60337 , n60342 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60361 , n31836 , n60360 );
nor ( n60362 , n60332 , n60336 , n60342 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60363 , n31838 , n60362 );
nor ( n60364 , n60331 , n60336 , n60342 , n60349 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60365 , n31840 , n60364 );
nor ( n60366 , n60332 , n60337 , n60343 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60367 , n31842 , n60366 );
nor ( n60368 , n60331 , n60337 , n60343 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60369 , n31844 , n60368 );
nor ( n60370 , n60332 , n60336 , n60343 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60371 , n31846 , n60370 );
nor ( n60372 , n60331 , n60336 , n60343 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60373 , n31848 , n60372 );
nor ( n60374 , n60332 , n60337 , n60342 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60375 , n31850 , n60374 );
nor ( n60376 , n60331 , n60337 , n60342 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60377 , n31852 , n60376 );
nor ( n60378 , n60332 , n60336 , n60342 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60379 , n31854 , n60378 );
nor ( n60380 , n60331 , n60336 , n60342 , n60348 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60381 , n31856 , n60380 );
or ( n60382 , n60351 , n60353 , n60355 , n60357 , n60359 , n60361 , n60363 , n60365 , n60367 , n60369 , n60371 , n60373 , n60375 , n60377 , n60379 , n60381 );
and ( n60383 , n31861 , n60350 );
and ( n60384 , n31863 , n60352 );
and ( n60385 , n31865 , n60354 );
and ( n60386 , n31867 , n60356 );
and ( n60387 , n31869 , n60358 );
and ( n60388 , n31871 , n60360 );
and ( n60389 , n31873 , n60362 );
and ( n60390 , n31875 , n60364 );
and ( n60391 , n31877 , n60366 );
and ( n60392 , n31879 , n60368 );
and ( n60393 , n31881 , n60370 );
and ( n60394 , n31883 , n60372 );
and ( n60395 , n31885 , n60374 );
and ( n60396 , n31887 , n60376 );
and ( n60397 , n31889 , n60378 );
and ( n60398 , n31891 , n60380 );
or ( n60399 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 );
and ( n60400 , n31896 , n60350 );
and ( n60401 , n31898 , n60352 );
and ( n60402 , n31900 , n60354 );
and ( n60403 , n31902 , n60356 );
and ( n60404 , n31904 , n60358 );
and ( n60405 , n31906 , n60360 );
and ( n60406 , n31908 , n60362 );
and ( n60407 , n31910 , n60364 );
and ( n60408 , n31912 , n60366 );
and ( n60409 , n31914 , n60368 );
and ( n60410 , n31916 , n60370 );
and ( n60411 , n31918 , n60372 );
and ( n60412 , n31920 , n60374 );
and ( n60413 , n31922 , n60376 );
and ( n60414 , n31924 , n60378 );
and ( n60415 , n31926 , n60380 );
or ( n60416 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 );
and ( n60417 , n31931 , n60350 );
and ( n60418 , n31933 , n60352 );
and ( n60419 , n31935 , n60354 );
and ( n60420 , n31937 , n60356 );
and ( n60421 , n31939 , n60358 );
and ( n60422 , n31941 , n60360 );
and ( n60423 , n31943 , n60362 );
and ( n60424 , n31945 , n60364 );
and ( n60425 , n31947 , n60366 );
and ( n60426 , n31949 , n60368 );
and ( n60427 , n31951 , n60370 );
and ( n60428 , n31953 , n60372 );
and ( n60429 , n31955 , n60374 );
and ( n60430 , n31957 , n60376 );
and ( n60431 , n31959 , n60378 );
and ( n60432 , n31961 , n60380 );
or ( n60433 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 );
and ( n60434 , n31966 , n60350 );
and ( n60435 , n31968 , n60352 );
and ( n60436 , n31970 , n60354 );
and ( n60437 , n31972 , n60356 );
and ( n60438 , n31974 , n60358 );
and ( n60439 , n31976 , n60360 );
and ( n60440 , n31978 , n60362 );
and ( n60441 , n31980 , n60364 );
and ( n60442 , n31982 , n60366 );
and ( n60443 , n31984 , n60368 );
and ( n60444 , n31986 , n60370 );
and ( n60445 , n31988 , n60372 );
and ( n60446 , n31990 , n60374 );
and ( n60447 , n31992 , n60376 );
and ( n60448 , n31994 , n60378 );
and ( n60449 , n31996 , n60380 );
or ( n60450 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 );
and ( n60451 , n32001 , n60350 );
and ( n60452 , n32003 , n60352 );
and ( n60453 , n32005 , n60354 );
and ( n60454 , n32007 , n60356 );
and ( n60455 , n32009 , n60358 );
and ( n60456 , n32011 , n60360 );
and ( n60457 , n32013 , n60362 );
and ( n60458 , n32015 , n60364 );
and ( n60459 , n32017 , n60366 );
and ( n60460 , n32019 , n60368 );
and ( n60461 , n32021 , n60370 );
and ( n60462 , n32023 , n60372 );
and ( n60463 , n32025 , n60374 );
and ( n60464 , n32027 , n60376 );
and ( n60465 , n32029 , n60378 );
and ( n60466 , n32031 , n60380 );
or ( n60467 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 );
and ( n60468 , n32036 , n60350 );
and ( n60469 , n32038 , n60352 );
and ( n60470 , n32040 , n60354 );
and ( n60471 , n32042 , n60356 );
and ( n60472 , n32044 , n60358 );
and ( n60473 , n32046 , n60360 );
and ( n60474 , n32048 , n60362 );
and ( n60475 , n32050 , n60364 );
and ( n60476 , n32052 , n60366 );
and ( n60477 , n32054 , n60368 );
and ( n60478 , n32056 , n60370 );
and ( n60479 , n32058 , n60372 );
and ( n60480 , n32060 , n60374 );
and ( n60481 , n32062 , n60376 );
and ( n60482 , n32064 , n60378 );
and ( n60483 , n32066 , n60380 );
or ( n60484 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 );
not ( n60485 , n31674 );
not ( n60486 , n60485 );
buf ( n60487 , n60486 );
not ( n60488 , n60487 );
not ( n60489 , n60488 );
xnor ( n60490 , n31670 , n31674 );
not ( n60491 , n60490 );
buf ( n60492 , n60491 );
buf ( n60493 , n60492 );
not ( n60494 , n60493 );
not ( n60495 , n60494 );
or ( n60496 , n31670 , n31674 );
xor ( n60497 , n31666 , n60496 );
not ( n60498 , n60497 );
buf ( n60499 , n60498 );
buf ( n60500 , n60499 );
not ( n60501 , n60500 );
not ( n60502 , n60501 );
and ( n60503 , n31666 , n60496 );
xor ( n60504 , n31662 , n60503 );
not ( n60505 , n60504 );
buf ( n60506 , n60505 );
buf ( n60507 , n60506 );
not ( n60508 , n60507 );
not ( n60509 , n60508 );
nor ( n60510 , n60489 , n60495 , n60502 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60511 , n31750 , n60510 );
nor ( n60512 , n60488 , n60495 , n60502 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60513 , n31778 , n60512 );
nor ( n60514 , n60489 , n60494 , n60502 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60515 , n31781 , n60514 );
nor ( n60516 , n60488 , n60494 , n60502 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60517 , n31784 , n60516 );
nor ( n60518 , n60489 , n60495 , n60501 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60519 , n31787 , n60518 );
nor ( n60520 , n60488 , n60495 , n60501 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60521 , n31790 , n60520 );
nor ( n60522 , n60489 , n60494 , n60501 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60523 , n31793 , n60522 );
nor ( n60524 , n60488 , n60494 , n60501 , n60509 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60525 , n31796 , n60524 );
nor ( n60526 , n60489 , n60495 , n60502 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60527 , n31799 , n60526 );
nor ( n60528 , n60488 , n60495 , n60502 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60529 , n31802 , n60528 );
nor ( n60530 , n60489 , n60494 , n60502 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60531 , n31805 , n60530 );
nor ( n60532 , n60488 , n60494 , n60502 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60533 , n31808 , n60532 );
nor ( n60534 , n60489 , n60495 , n60501 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60535 , n31811 , n60534 );
nor ( n60536 , n60488 , n60495 , n60501 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60537 , n31814 , n60536 );
nor ( n60538 , n60489 , n60494 , n60501 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60539 , n31817 , n60538 );
nor ( n60540 , n60488 , n60494 , n60501 , n60508 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n60541 , n31820 , n60540 );
or ( n60542 , n60511 , n60513 , n60515 , n60517 , n60519 , n60521 , n60523 , n60525 , n60527 , n60529 , n60531 , n60533 , n60535 , n60537 , n60539 , n60541 );
and ( n60543 , n60484 , n60542 );
and ( n60544 , n60467 , n60543 );
and ( n60545 , n60450 , n60544 );
and ( n60546 , n60433 , n60545 );
and ( n60547 , n60416 , n60546 );
and ( n60548 , n60399 , n60547 );
xor ( n60549 , n60382 , n60548 );
and ( n60550 , n60549 , n47331 );
or ( n60551 , n60328 , n60550 );
and ( n60552 , n60551 , n32413 );
and ( n60553 , n49563 , n47402 );
or ( n60554 , n60326 , n60552 , n60553 );
and ( n60555 , n60554 , n32456 );
and ( n60556 , n49563 , n47409 );
or ( n60557 , C0 , n60555 , n60556 );
buf ( n60558 , n60557 );
buf ( n60559 , n60558 );
buf ( n60560 , n31655 );
buf ( n60561 , n30987 );
not ( n60562 , n46356 );
and ( n60563 , n60562 , n31236 );
nor ( n60564 , n31025 , n31021 , n31017 , n31013 , n31009 );
not ( n60565 , n60564 );
and ( n60566 , n60565 , n31236 );
and ( n60567 , n31238 , n60564 );
or ( n60568 , n60566 , n60567 );
and ( n60569 , n60568 , n46356 );
or ( n60570 , n60563 , n60569 );
and ( n60571 , n60570 , n31649 );
nor ( n60572 , n46373 , n46379 , n46386 , n46392 , C0 );
not ( n60573 , n60572 );
not ( n60574 , n60564 );
and ( n60575 , n60574 , n31236 );
and ( n60576 , n49901 , n60564 );
or ( n60577 , n60575 , n60576 );
and ( n60578 , n60573 , n60577 );
and ( n60579 , n49901 , n60572 );
or ( n60580 , n60578 , n60579 );
and ( n60581 , n60580 , n31643 );
not ( n60582 , n31452 );
not ( n60583 , n60572 );
not ( n60584 , n60564 );
and ( n60585 , n60584 , n31236 );
and ( n60586 , n49901 , n60564 );
or ( n60587 , n60585 , n60586 );
and ( n60588 , n60583 , n60587 );
and ( n60589 , n49901 , n60572 );
or ( n60590 , n60588 , n60589 );
and ( n60591 , n60582 , n60590 );
nor ( n60592 , n46519 , n46528 , n46539 , n46549 , C0 );
not ( n60593 , n60592 );
nor ( n60594 , n46515 , n46524 , n46534 , n46544 , C0 );
not ( n60595 , n60594 );
and ( n60596 , n60595 , n60590 );
and ( n60597 , n49925 , n60594 );
or ( n60598 , n60596 , n60597 );
and ( n60599 , n60593 , n60598 );
and ( n60600 , n49933 , n60592 );
or ( n60601 , n60599 , n60600 );
and ( n60602 , n60601 , n31452 );
or ( n60603 , n60591 , n60602 );
and ( n60604 , n60603 , n31638 );
and ( n60605 , n31236 , n47277 );
or ( n60606 , C0 , n60571 , n60581 , n60604 , n60605 );
buf ( n60607 , n60606 );
buf ( n60608 , n60607 );
buf ( n60609 , n30987 );
buf ( n60610 , n31655 );
buf ( n60611 , n31655 );
buf ( n60612 , n30987 );
buf ( n60613 , n30987 );
buf ( n60614 , n31655 );
not ( n60615 , n32953 );
buf ( n60616 , RI15b46d10_281);
and ( n60617 , n60615 , n60616 );
not ( n60618 , n39572 );
and ( n60619 , n60618 , n39529 );
xor ( n60620 , n42616 , n42637 );
and ( n60621 , n60620 , n39572 );
or ( n60622 , n60619 , n60621 );
and ( n60623 , n60622 , n32953 );
or ( n60624 , n60617 , n60623 );
and ( n60625 , n60624 , n33038 );
not ( n60626 , n39586 );
and ( n60627 , n60626 , n60616 );
not ( n60628 , n39775 );
and ( n60629 , n60628 , n39735 );
xor ( n60630 , n42652 , n42673 );
and ( n60631 , n60630 , n39775 );
or ( n60632 , n60629 , n60631 );
and ( n60633 , n60632 , n39586 );
or ( n60634 , n60627 , n60633 );
and ( n60635 , n60634 , n33172 );
and ( n60636 , n60616 , n39795 );
or ( n60637 , n60625 , n60635 , n60636 );
and ( n60638 , n60637 , n33208 );
and ( n60639 , n60616 , n39805 );
or ( n60640 , C0 , n60638 , n60639 );
buf ( n60641 , n60640 );
buf ( n60642 , n60641 );
buf ( n60643 , n31655 );
buf ( n60644 , n30987 );
not ( n60645 , n34150 );
and ( n60646 , n60645 , n32692 );
not ( n60647 , n50731 );
and ( n60648 , n60647 , n32692 );
and ( n60649 , n32722 , n50731 );
or ( n60650 , n60648 , n60649 );
and ( n60651 , n60650 , n34150 );
or ( n60652 , n60646 , n60651 );
and ( n60653 , n60652 , n33381 );
not ( n60654 , n50739 );
not ( n60655 , n50731 );
and ( n60656 , n60655 , n32692 );
and ( n60657 , n42565 , n50731 );
or ( n60658 , n60656 , n60657 );
and ( n60659 , n60654 , n60658 );
and ( n60660 , n42565 , n50739 );
or ( n60661 , n60659 , n60660 );
and ( n60662 , n60661 , n33375 );
not ( n60663 , n32968 );
not ( n60664 , n50739 );
not ( n60665 , n50731 );
and ( n60666 , n60665 , n32692 );
and ( n60667 , n42565 , n50731 );
or ( n60668 , n60666 , n60667 );
and ( n60669 , n60664 , n60668 );
and ( n60670 , n42565 , n50739 );
or ( n60671 , n60669 , n60670 );
and ( n60672 , n60663 , n60671 );
not ( n60673 , n50759 );
not ( n60674 , n50761 );
and ( n60675 , n60674 , n60671 );
and ( n60676 , n42589 , n50761 );
or ( n60677 , n60675 , n60676 );
and ( n60678 , n60673 , n60677 );
and ( n60679 , n42597 , n50759 );
or ( n60680 , n60678 , n60679 );
and ( n60681 , n60680 , n32968 );
or ( n60682 , n60672 , n60681 );
and ( n60683 , n60682 , n33370 );
and ( n60684 , n32692 , n35062 );
or ( n60685 , C0 , n60653 , n60662 , n60683 , n60684 );
buf ( n60686 , n60685 );
buf ( n60687 , n60686 );
buf ( n60688 , n30987 );
buf ( n60689 , n31655 );
and ( n60690 , n32298 , n50275 );
not ( n60691 , n50278 );
and ( n60692 , n60691 , n31735 );
and ( n60693 , n32298 , n50278 );
or ( n60694 , n60692 , n60693 );
and ( n60695 , n60694 , n32421 );
not ( n60696 , n50002 );
and ( n60697 , n60696 , n31735 );
and ( n60698 , n32298 , n50002 );
or ( n60699 , n60697 , n60698 );
and ( n60700 , n60699 , n32419 );
not ( n60701 , n50289 );
and ( n60702 , n60701 , n31735 );
and ( n60703 , n32298 , n50289 );
or ( n60704 , n60702 , n60703 );
and ( n60705 , n60704 , n32417 );
not ( n60706 , n50008 );
and ( n60707 , n60706 , n31735 );
and ( n60708 , n32298 , n50008 );
or ( n60709 , n60707 , n60708 );
and ( n60710 , n60709 , n32415 );
not ( n60711 , n47331 );
and ( n60712 , n60711 , n31735 );
and ( n60713 , n31860 , n47331 );
or ( n60714 , n60712 , n60713 );
and ( n60715 , n60714 , n32413 );
not ( n60716 , n50067 );
and ( n60717 , n60716 , n31735 );
and ( n60718 , n31860 , n50067 );
or ( n60719 , n60717 , n60718 );
and ( n60720 , n60719 , n32411 );
not ( n60721 , n31728 );
and ( n60722 , n60721 , n31735 );
and ( n60723 , n52636 , n31728 );
or ( n60724 , n60722 , n60723 );
and ( n60725 , n60724 , n32253 );
not ( n60726 , n32283 );
and ( n60727 , n60726 , n31735 );
and ( n60728 , n52649 , n32283 );
or ( n60729 , n60727 , n60728 );
and ( n60730 , n60729 , n32398 );
and ( n60731 , n32348 , n50334 );
or ( n60732 , n60690 , n60695 , n60700 , n60705 , n60710 , n60715 , n60720 , n60725 , n60730 , n60731 );
and ( n60733 , n60732 , n32456 );
and ( n60734 , n37579 , n32489 );
and ( n60735 , n31735 , n50345 );
or ( n60736 , C0 , n60733 , n60734 , n60735 );
buf ( n60737 , n60736 );
buf ( n60738 , n60737 );
buf ( n60739 , n30987 );
not ( n60740 , n31437 );
buf ( n60741 , RI15b52890_681);
and ( n60742 , n60740 , n60741 );
not ( n60743 , n45766 );
and ( n60744 , n60743 , n45660 );
xor ( n60745 , n45770 , n45786 );
and ( n60746 , n60745 , n45766 );
or ( n60747 , n60744 , n60746 );
and ( n60748 , n60747 , n31437 );
or ( n60749 , n60742 , n60748 );
and ( n60750 , n60749 , n31468 );
not ( n60751 , n44817 );
and ( n60752 , n60751 , n60741 );
not ( n60753 , n44994 );
and ( n60754 , n60753 , n44918 );
xor ( n60755 , n45002 , n45018 );
and ( n60756 , n60755 , n44994 );
or ( n60757 , n60754 , n60756 );
and ( n60758 , n60757 , n44817 );
or ( n60759 , n60752 , n60758 );
and ( n60760 , n60759 , n31521 );
and ( n60761 , n60741 , n42158 );
or ( n60762 , n60750 , n60760 , n60761 );
and ( n60763 , n60762 , n31557 );
and ( n60764 , n60741 , n40154 );
or ( n60765 , C0 , n60763 , n60764 );
buf ( n60766 , n60765 );
buf ( n60767 , n60766 );
buf ( n60768 , n31655 );
not ( n60769 , n31728 );
and ( n60770 , n60769 , n46035 );
xor ( n60771 , n47612 , n47617 );
and ( n60772 , n60771 , n31728 );
or ( n60773 , n60770 , n60772 );
and ( n60774 , n60773 , n32253 );
not ( n60775 , n32283 );
and ( n60776 , n60775 , n46035 );
not ( n60777 , n31823 );
xor ( n60778 , n47667 , n47672 );
and ( n60779 , n60777 , n60778 );
xnor ( n60780 , n47717 , n47722 );
and ( n60781 , n60780 , n31823 );
or ( n60782 , n60779 , n60781 );
and ( n60783 , n60782 , n32283 );
or ( n60784 , n60776 , n60783 );
and ( n60785 , n60784 , n32398 );
and ( n60786 , n46035 , n32436 );
or ( n60787 , n60774 , n60785 , n60786 );
and ( n60788 , n60787 , n32456 );
and ( n60789 , n49687 , n32473 );
not ( n60790 , n32475 );
and ( n60791 , n60790 , n49687 );
xor ( n60792 , n46035 , n47751 );
and ( n60793 , n60792 , n32475 );
or ( n60794 , n60791 , n60793 );
and ( n60795 , n60794 , n32486 );
and ( n60796 , n37567 , n32489 );
and ( n60797 , n46035 , n32501 );
or ( n60798 , C0 , n60788 , n60789 , n60795 , n60796 , n60797 );
buf ( n60799 , n60798 );
buf ( n60800 , n60799 );
buf ( n60801 , n31655 );
buf ( n60802 , n30987 );
and ( n60803 , n33215 , n32528 );
not ( n60804 , n32598 );
and ( n60805 , n60804 , n32978 );
buf ( n60806 , n60805 );
and ( n60807 , n60806 , n32890 );
not ( n60808 , n32919 );
and ( n60809 , n60808 , n32978 );
buf ( n60810 , n60809 );
and ( n60811 , n60810 , n32924 );
not ( n60812 , n32953 );
and ( n60813 , n60812 , n32978 );
not ( n60814 , n32971 );
and ( n60815 , n60814 , n33081 );
xor ( n60816 , n32978 , n33027 );
and ( n60817 , n60816 , n32971 );
or ( n60818 , n60815 , n60817 );
and ( n60819 , n60818 , n32953 );
or ( n60820 , n60813 , n60819 );
and ( n60821 , n60820 , n33038 );
not ( n60822 , n33067 );
and ( n60823 , n60822 , n32978 );
not ( n60824 , n32970 );
not ( n60825 , n33071 );
and ( n60826 , n60825 , n33081 );
xor ( n60827 , n33082 , n33159 );
and ( n60828 , n60827 , n33071 );
or ( n60829 , n60826 , n60828 );
and ( n60830 , n60824 , n60829 );
and ( n60831 , n60816 , n32970 );
or ( n60832 , n60830 , n60831 );
and ( n60833 , n60832 , n33067 );
or ( n60834 , n60823 , n60833 );
and ( n60835 , n60834 , n33172 );
and ( n60836 , n32978 , n33204 );
or ( n60837 , n60807 , n60811 , n60821 , n60835 , n60836 );
and ( n60838 , n60837 , n33208 );
not ( n60839 , n32968 );
not ( n60840 , n33270 );
and ( n60841 , n60840 , n33281 );
xor ( n60842 , n33282 , n33359 );
and ( n60843 , n60842 , n33270 );
or ( n60844 , n60841 , n60843 );
and ( n60845 , n60839 , n60844 );
and ( n60846 , n32978 , n32968 );
or ( n60847 , n60845 , n60846 );
and ( n60848 , n60847 , n33370 );
and ( n60849 , n32978 , n33382 );
or ( n60850 , C0 , n60803 , n60838 , n60848 , C0 , n60849 );
buf ( n60851 , n60850 );
buf ( n60852 , n60851 );
buf ( n60853 , n30987 );
buf ( n60854 , n31655 );
buf ( n60855 , n31655 );
buf ( n60856 , n30987 );
not ( n60857 , n46356 );
and ( n60858 , n60857 , n31179 );
not ( n60859 , n46362 );
and ( n60860 , n60859 , n31179 );
and ( n60861 , n31205 , n46362 );
or ( n60862 , n60860 , n60861 );
and ( n60863 , n60862 , n46356 );
or ( n60864 , n60858 , n60863 );
and ( n60865 , n60864 , n31649 );
not ( n60866 , n46393 );
not ( n60867 , n46362 );
and ( n60868 , n60867 , n31179 );
and ( n60869 , n50125 , n46362 );
or ( n60870 , n60868 , n60869 );
and ( n60871 , n60866 , n60870 );
and ( n60872 , n50125 , n46393 );
or ( n60873 , n60871 , n60872 );
and ( n60874 , n60873 , n31643 );
not ( n60875 , n31452 );
not ( n60876 , n46393 );
not ( n60877 , n46362 );
and ( n60878 , n60877 , n31179 );
and ( n60879 , n50125 , n46362 );
or ( n60880 , n60878 , n60879 );
and ( n60881 , n60876 , n60880 );
and ( n60882 , n50125 , n46393 );
or ( n60883 , n60881 , n60882 );
and ( n60884 , n60875 , n60883 );
not ( n60885 , n46550 );
not ( n60886 , n46554 );
and ( n60887 , n60886 , n60883 );
and ( n60888 , n50151 , n46554 );
or ( n60889 , n60887 , n60888 );
and ( n60890 , n60885 , n60889 );
and ( n60891 , n50159 , n46550 );
or ( n60892 , n60890 , n60891 );
and ( n60893 , n60892 , n31452 );
or ( n60894 , n60884 , n60893 );
and ( n60895 , n60894 , n31638 );
and ( n60896 , n31179 , n47277 );
or ( n60897 , C0 , n60865 , n60874 , n60895 , n60896 );
buf ( n60898 , n60897 );
buf ( n60899 , n60898 );
buf ( n60900 , n31655 );
buf ( n60901 , RI15b5f5e0_1119);
and ( n60902 , n60901 , n32494 );
not ( n60903 , n46083 );
buf ( n60904 , RI15b5fd60_1135);
and ( n60905 , n60903 , n60904 );
not ( n60906 , n46290 );
and ( n60907 , n60906 , n46247 );
xor ( n60908 , n46294 , n46318 );
and ( n60909 , n60908 , n46290 );
or ( n60910 , n60907 , n60909 );
and ( n60911 , n60910 , n46083 );
or ( n60912 , n60905 , n60911 );
and ( n60913 , n60912 , n32421 );
not ( n60914 , n46326 );
and ( n60915 , n60914 , n60904 );
and ( n60916 , n60910 , n46326 );
or ( n60917 , n60915 , n60916 );
and ( n60918 , n60917 , n32417 );
and ( n60919 , n60904 , n46340 );
or ( n60920 , n60913 , n60918 , n60919 );
and ( n60921 , n60920 , n32456 );
and ( n60922 , n60904 , n46349 );
or ( n60923 , C0 , n60902 , n60921 , n60922 );
buf ( n60924 , n60923 );
buf ( n60925 , n60924 );
and ( n60926 , n33231 , n32528 );
not ( n60927 , n32598 );
and ( n60928 , n60927 , n32994 );
buf ( n60929 , n60928 );
and ( n60930 , n60929 , n32890 );
not ( n60931 , n32919 );
and ( n60932 , n60931 , n32994 );
buf ( n60933 , n60932 );
and ( n60934 , n60933 , n32924 );
not ( n60935 , n32953 );
and ( n60936 , n60935 , n32994 );
not ( n60937 , n32971 );
and ( n60938 , n60937 , n33113 );
xor ( n60939 , n32994 , n33011 );
and ( n60940 , n60939 , n32971 );
or ( n60941 , n60938 , n60940 );
and ( n60942 , n60941 , n32953 );
or ( n60943 , n60936 , n60942 );
and ( n60944 , n60943 , n33038 );
not ( n60945 , n33067 );
and ( n60946 , n60945 , n32994 );
not ( n60947 , n32970 );
not ( n60948 , n33071 );
and ( n60949 , n60948 , n33113 );
xor ( n60950 , n33114 , n33143 );
and ( n60951 , n60950 , n33071 );
or ( n60952 , n60949 , n60951 );
and ( n60953 , n60947 , n60952 );
and ( n60954 , n60939 , n32970 );
or ( n60955 , n60953 , n60954 );
and ( n60956 , n60955 , n33067 );
or ( n60957 , n60946 , n60956 );
and ( n60958 , n60957 , n33172 );
and ( n60959 , n32994 , n33204 );
or ( n60960 , n60930 , n60934 , n60944 , n60958 , n60959 );
and ( n60961 , n60960 , n33208 );
not ( n60962 , n32968 );
not ( n60963 , n33270 );
and ( n60964 , n60963 , n33313 );
xor ( n60965 , n33314 , n33343 );
and ( n60966 , n60965 , n33270 );
or ( n60967 , n60964 , n60966 );
and ( n60968 , n60962 , n60967 );
and ( n60969 , n32994 , n32968 );
or ( n60970 , n60968 , n60969 );
and ( n60971 , n60970 , n33370 );
buf ( n60972 , n35056 );
and ( n60973 , n32994 , n33382 );
or ( n60974 , C0 , n60926 , n60961 , n60971 , n60972 , n60973 );
buf ( n60975 , n60974 );
buf ( n60976 , n60975 );
buf ( n60977 , n31655 );
buf ( n60978 , n30987 );
buf ( n60979 , n30987 );
buf ( n60980 , n31655 );
not ( n60981 , n31728 );
and ( n60982 , n60981 , n46019 );
xor ( n60983 , n50419 , n50424 );
and ( n60984 , n60983 , n31728 );
or ( n60985 , n60982 , n60984 );
and ( n60986 , n60985 , n32253 );
not ( n60987 , n32283 );
and ( n60988 , n60987 , n46019 );
not ( n60989 , n31823 );
xor ( n60990 , n50441 , n50446 );
and ( n60991 , n60989 , n60990 );
xnor ( n60992 , n50458 , n50463 );
and ( n60993 , n60992 , n31823 );
or ( n60994 , n60991 , n60993 );
and ( n60995 , n60994 , n32283 );
or ( n60996 , n60988 , n60995 );
and ( n60997 , n60996 , n32398 );
and ( n60998 , n46019 , n32436 );
or ( n60999 , n60986 , n60997 , n60998 );
and ( n61000 , n60999 , n32456 );
and ( n61001 , n49656 , n32473 );
not ( n61002 , n32475 );
and ( n61003 , n61002 , n49656 );
xor ( n61004 , n46019 , n50480 );
and ( n61005 , n61004 , n32475 );
or ( n61006 , n61003 , n61005 );
and ( n61007 , n61006 , n32486 );
and ( n61008 , n37535 , n32489 );
and ( n61009 , n46019 , n32501 );
or ( n61010 , C0 , n61000 , n61001 , n61007 , n61008 , n61009 );
buf ( n61011 , n61010 );
buf ( n61012 , n61011 );
buf ( n61013 , n31655 );
buf ( n61014 , n30987 );
not ( n61015 , n33419 );
and ( n61016 , n61015 , n31586 );
xor ( n61017 , n33554 , n33571 );
xor ( n61018 , n61017 , n33679 );
and ( n61019 , n61018 , n33419 );
or ( n61020 , n61016 , n61019 );
and ( n61021 , n61020 , n31529 );
not ( n61022 , n33734 );
and ( n61023 , n61022 , n31586 );
not ( n61024 , n33533 );
xor ( n61025 , n33775 , n33571 );
xor ( n61026 , n61025 , n33797 );
and ( n61027 , n61024 , n61026 );
xor ( n61028 , n33864 , n33866 );
xor ( n61029 , n61028 , n33899 );
and ( n61030 , n61029 , n33533 );
or ( n61031 , n61027 , n61030 );
and ( n61032 , n61031 , n33734 );
or ( n61033 , n61023 , n61032 );
and ( n61034 , n61033 , n31527 );
and ( n61035 , n31586 , n33942 );
or ( n61036 , n61021 , n61034 , n61035 );
and ( n61037 , n61036 , n31557 );
and ( n61038 , n34117 , n31643 );
not ( n61039 , n31452 );
and ( n61040 , n61039 , n34117 );
xor ( n61041 , n31586 , n33951 );
and ( n61042 , n61041 , n31452 );
or ( n61043 , n61040 , n61042 );
and ( n61044 , n61043 , n31638 );
and ( n61045 , n34010 , n33973 );
and ( n61046 , n31586 , n33978 );
or ( n61047 , C0 , n61037 , n61038 , n61044 , n61045 , n61046 );
buf ( n61048 , n61047 );
buf ( n61049 , n61048 );
not ( n61050 , n40163 );
and ( n61051 , n61050 , n31673 );
and ( n61052 , n40177 , n40163 );
or ( n61053 , n61051 , n61052 );
and ( n61054 , n61053 , n32498 );
not ( n61055 , n55780 );
not ( n61056 , n55558 );
and ( n61057 , n61056 , n31673 );
buf ( n61058 , n55558 );
or ( n61059 , n61057 , n61058 );
and ( n61060 , n61055 , n61059 );
buf ( n61061 , n61060 );
and ( n61062 , n61061 , n32496 );
and ( n61063 , n40413 , n32473 );
buf ( n61064 , n40413 );
and ( n61065 , n61064 , n32486 );
and ( n61066 , n31673 , n55800 );
or ( n61067 , C0 , n61054 , n61062 , n61063 , n61065 , n61066 );
buf ( n61068 , n61067 );
buf ( n61069 , n61068 );
buf ( n61070 , n30987 );
not ( n61071 , n35542 );
and ( n61072 , n61071 , n41848 );
buf ( n61073 , RI15b454b0_229);
and ( n61074 , n61073 , n35542 );
or ( n61075 , n61072 , n61074 );
buf ( n61076 , n61075 );
buf ( n61077 , n61076 );
buf ( n61078 , n31655 );
buf ( n61079 , n30987 );
not ( n61080 , n34150 );
and ( n61081 , n61080 , n32863 );
not ( n61082 , n59574 );
and ( n61083 , n61082 , n32863 );
and ( n61084 , n32889 , n59574 );
or ( n61085 , n61083 , n61084 );
and ( n61086 , n61085 , n34150 );
or ( n61087 , n61081 , n61086 );
and ( n61088 , n61087 , n33381 );
not ( n61089 , n59582 );
not ( n61090 , n59574 );
and ( n61091 , n61090 , n32863 );
and ( n61092 , n52819 , n59574 );
or ( n61093 , n61091 , n61092 );
and ( n61094 , n61089 , n61093 );
and ( n61095 , n52819 , n59582 );
or ( n61096 , n61094 , n61095 );
and ( n61097 , n61096 , n33375 );
not ( n61098 , n32968 );
not ( n61099 , n59582 );
not ( n61100 , n59574 );
and ( n61101 , n61100 , n32863 );
and ( n61102 , n52819 , n59574 );
or ( n61103 , n61101 , n61102 );
and ( n61104 , n61099 , n61103 );
and ( n61105 , n52819 , n59582 );
or ( n61106 , n61104 , n61105 );
and ( n61107 , n61098 , n61106 );
not ( n61108 , n59602 );
not ( n61109 , n59604 );
and ( n61110 , n61109 , n61106 );
and ( n61111 , n52845 , n59604 );
or ( n61112 , n61110 , n61111 );
and ( n61113 , n61108 , n61112 );
and ( n61114 , n52855 , n59602 );
or ( n61115 , n61113 , n61114 );
and ( n61116 , n61115 , n32968 );
or ( n61117 , n61107 , n61116 );
and ( n61118 , n61117 , n33370 );
and ( n61119 , n32863 , n35062 );
or ( n61120 , C0 , n61088 , n61097 , n61118 , n61119 );
buf ( n61121 , n61120 );
buf ( n61122 , n61121 );
buf ( n61123 , n30987 );
buf ( n61124 , n31655 );
buf ( n61125 , n31655 );
buf ( n61126 , n30987 );
not ( n61127 , n34150 );
and ( n61128 , n61127 , n32657 );
not ( n61129 , n56708 );
and ( n61130 , n61129 , n32657 );
and ( n61131 , n32689 , n56708 );
or ( n61132 , n61130 , n61131 );
and ( n61133 , n61132 , n34150 );
or ( n61134 , n61128 , n61133 );
and ( n61135 , n61134 , n33381 );
not ( n61136 , n56716 );
not ( n61137 , n56708 );
and ( n61138 , n61137 , n32657 );
and ( n61139 , n50682 , n56708 );
or ( n61140 , n61138 , n61139 );
and ( n61141 , n61136 , n61140 );
and ( n61142 , n50682 , n56716 );
or ( n61143 , n61141 , n61142 );
and ( n61144 , n61143 , n33375 );
not ( n61145 , n32968 );
not ( n61146 , n56716 );
not ( n61147 , n56708 );
and ( n61148 , n61147 , n32657 );
and ( n61149 , n50682 , n56708 );
or ( n61150 , n61148 , n61149 );
and ( n61151 , n61146 , n61150 );
and ( n61152 , n50682 , n56716 );
or ( n61153 , n61151 , n61152 );
and ( n61154 , n61145 , n61153 );
not ( n61155 , n56736 );
not ( n61156 , n56738 );
and ( n61157 , n61156 , n61153 );
and ( n61158 , n50706 , n56738 );
or ( n61159 , n61157 , n61158 );
and ( n61160 , n61155 , n61159 );
and ( n61161 , n50714 , n56736 );
or ( n61162 , n61160 , n61161 );
and ( n61163 , n61162 , n32968 );
or ( n61164 , n61154 , n61163 );
and ( n61165 , n61164 , n33370 );
and ( n61166 , n32657 , n35062 );
or ( n61167 , C0 , n61135 , n61144 , n61165 , n61166 );
buf ( n61168 , n61167 );
buf ( n61169 , n61168 );
buf ( n61170 , n30987 );
buf ( n61171 , n31655 );
not ( n61172 , n38443 );
and ( n61173 , n61172 , n38133 );
xor ( n61174 , n53474 , n53495 );
and ( n61175 , n61174 , n38443 );
or ( n61176 , n61173 , n61175 );
and ( n61177 , n61176 , n38450 );
not ( n61178 , n39339 );
and ( n61179 , n61178 , n39033 );
xor ( n61180 , n53530 , n53551 );
and ( n61181 , n61180 , n39339 );
or ( n61182 , n61179 , n61181 );
and ( n61183 , n61182 , n39346 );
and ( n61184 , n40210 , n39359 );
or ( n61185 , n61177 , n61183 , n61184 );
buf ( n61186 , n61185 );
buf ( n61187 , n61186 );
and ( n61188 , n52390 , n31647 );
not ( n61189 , n48457 );
and ( n61190 , n61189 , n31010 );
buf ( n61191 , n61190 );
and ( n61192 , n61191 , n31373 );
not ( n61193 , n44807 );
and ( n61194 , n61193 , n31010 );
and ( n61195 , n31014 , n42323 );
xor ( n61196 , n31010 , n61195 );
and ( n61197 , n61196 , n44807 );
or ( n61198 , n61194 , n61197 );
and ( n61199 , n61198 , n31408 );
not ( n61200 , n48468 );
and ( n61201 , n61200 , n31010 );
buf ( n61202 , n61201 );
and ( n61203 , n61202 , n31468 );
not ( n61204 , n44817 );
and ( n61205 , n61204 , n31010 );
buf ( n61206 , n61205 );
and ( n61207 , n61206 , n31521 );
not ( n61208 , n39979 );
and ( n61209 , n61208 , n31010 );
buf ( n61210 , n61209 );
and ( n61211 , n61210 , n31538 );
not ( n61212 , n45059 );
and ( n61213 , n61212 , n31010 );
buf ( n61214 , n61213 );
and ( n61215 , n61214 , n31536 );
or ( n61216 , n31527 , n31529 );
and ( n61217 , n31010 , n61216 );
or ( n61218 , C0 , n61192 , n61199 , n61203 , n61207 , n61211 , n61215 , n61217 , C0 );
and ( n61219 , n61218 , n31557 );
or ( n61220 , n40151 , n31007 );
and ( n61221 , n31010 , n61220 );
or ( n61222 , C0 , C0 , n61188 , n61219 , n61221 );
buf ( n61223 , n61222 );
buf ( n61224 , n61223 );
buf ( n61225 , n31655 );
buf ( n61226 , n30987 );
buf ( n61227 , n30987 );
buf ( n61228 , n31655 );
buf ( n61229 , n31655 );
buf ( n61230 , n30987 );
not ( n61231 , n32953 );
buf ( n61232 , RI15b46860_271);
and ( n61233 , n61231 , n61232 );
not ( n61234 , n39572 );
and ( n61235 , n61234 , n39399 );
xor ( n61236 , n42626 , n42627 );
and ( n61237 , n61236 , n39572 );
or ( n61238 , n61235 , n61237 );
and ( n61239 , n61238 , n32953 );
or ( n61240 , n61233 , n61239 );
and ( n61241 , n61240 , n33038 );
not ( n61242 , n39586 );
and ( n61243 , n61242 , n61232 );
not ( n61244 , n39775 );
and ( n61245 , n61244 , n39615 );
xor ( n61246 , n42662 , n42663 );
and ( n61247 , n61246 , n39775 );
or ( n61248 , n61245 , n61247 );
and ( n61249 , n61248 , n39586 );
or ( n61250 , n61243 , n61249 );
and ( n61251 , n61250 , n33172 );
and ( n61252 , n61232 , n39795 );
or ( n61253 , n61241 , n61251 , n61252 );
and ( n61254 , n61253 , n33208 );
and ( n61255 , n61232 , n39805 );
or ( n61256 , C0 , n61254 , n61255 );
buf ( n61257 , n61256 );
buf ( n61258 , n61257 );
buf ( n61259 , n30987 );
buf ( n61260 , n31655 );
buf ( n61261 , n31655 );
not ( n61262 , n34150 );
and ( n61263 , n61262 , n32731 );
not ( n61264 , n59105 );
and ( n61265 , n61264 , n32731 );
and ( n61266 , n32755 , n59105 );
or ( n61267 , n61265 , n61266 );
and ( n61268 , n61267 , n34150 );
or ( n61269 , n61263 , n61268 );
and ( n61270 , n61269 , n33381 );
not ( n61271 , n59113 );
not ( n61272 , n59105 );
and ( n61273 , n61272 , n32731 );
and ( n61274 , n35083 , n59105 );
or ( n61275 , n61273 , n61274 );
and ( n61276 , n61271 , n61275 );
and ( n61277 , n35083 , n59113 );
or ( n61278 , n61276 , n61277 );
and ( n61279 , n61278 , n33375 );
not ( n61280 , n32968 );
not ( n61281 , n59113 );
not ( n61282 , n59105 );
and ( n61283 , n61282 , n32731 );
and ( n61284 , n35083 , n59105 );
or ( n61285 , n61283 , n61284 );
and ( n61286 , n61281 , n61285 );
and ( n61287 , n35083 , n59113 );
or ( n61288 , n61286 , n61287 );
and ( n61289 , n61280 , n61288 );
not ( n61290 , n59133 );
not ( n61291 , n59135 );
and ( n61292 , n61291 , n61288 );
and ( n61293 , n35107 , n59135 );
or ( n61294 , n61292 , n61293 );
and ( n61295 , n61290 , n61294 );
and ( n61296 , n35115 , n59133 );
or ( n61297 , n61295 , n61296 );
and ( n61298 , n61297 , n32968 );
or ( n61299 , n61289 , n61298 );
and ( n61300 , n61299 , n33370 );
and ( n61301 , n32731 , n35062 );
or ( n61302 , C0 , n61270 , n61279 , n61300 , n61301 );
buf ( n61303 , n61302 );
buf ( n61304 , n61303 );
buf ( n61305 , n30987 );
buf ( n61306 , n30987 );
buf ( n61307 , n30987 );
buf ( n61308 , n31655 );
and ( n61309 , n56467 , n33379 );
and ( n61310 , n57586 , n33208 );
or ( n61311 , n39802 , n32528 );
and ( n61312 , n32531 , n61311 );
or ( n61313 , C0 , C0 , n61309 , n61310 , n61312 );
buf ( n61314 , n61313 );
buf ( n61315 , n61314 );
buf ( n61316 , n31655 );
buf ( n61317 , n30987 );
buf ( n61318 , n30987 );
buf ( n61319 , n31655 );
not ( n61320 , n41532 );
and ( n61321 , n61320 , n34193 );
and ( n61322 , n35534 , n41532 );
or ( n61323 , n61321 , n61322 );
buf ( n61324 , n61323 );
buf ( n61325 , n61324 );
xor ( n61326 , n39454 , n54970 );
and ( n61327 , n61326 , n33199 );
not ( n61328 , n48648 );
and ( n61329 , n61328 , n39454 );
and ( n61330 , n34273 , n48648 );
or ( n61331 , n61329 , n61330 );
and ( n61332 , n61331 , n32924 );
not ( n61333 , n48660 );
and ( n61334 , n61333 , n39454 );
not ( n61335 , n39584 );
buf ( n61336 , RI15b46ab8_276);
and ( n61337 , n61335 , n61336 );
not ( n61338 , n39775 );
and ( n61339 , n61338 , n39675 );
xor ( n61340 , n42657 , n42668 );
and ( n61341 , n61340 , n39775 );
or ( n61342 , n61339 , n61341 );
and ( n61343 , n61342 , n39584 );
or ( n61344 , n61337 , n61343 );
and ( n61345 , n61344 , n48660 );
or ( n61346 , n61334 , n61345 );
and ( n61347 , n61346 , n33172 );
not ( n61348 , n48730 );
and ( n61349 , n61348 , n39454 );
and ( n61350 , n48845 , n48730 );
or ( n61351 , n61349 , n61350 );
and ( n61352 , n61351 , n33187 );
and ( n61353 , n39454 , n54713 );
or ( n61354 , n61327 , n61332 , n61347 , n61352 , n61353 );
and ( n61355 , n61354 , n33208 );
and ( n61356 , n39454 , n39805 );
or ( n61357 , C0 , n61355 , n61356 );
buf ( n61358 , n61357 );
buf ( n61359 , n61358 );
buf ( n61360 , n31655 );
buf ( n61361 , n31655 );
buf ( n61362 , n30987 );
and ( n61363 , n48668 , n48639 );
buf ( n61364 , n48668 );
and ( n61365 , n61364 , n32890 );
buf ( n61366 , n48668 );
and ( n61367 , n61366 , n32924 );
buf ( n61368 , n48668 );
and ( n61369 , n61368 , n33038 );
buf ( n61370 , n48668 );
and ( n61371 , n61370 , n33172 );
not ( n61372 , n41576 );
and ( n61373 , n61372 , n48668 );
and ( n61374 , n48961 , n41576 );
or ( n61375 , n61373 , n61374 );
and ( n61376 , n61375 , n33189 );
not ( n61377 , n48730 );
and ( n61378 , n61377 , n48668 );
and ( n61379 , n48961 , n48730 );
or ( n61380 , n61378 , n61379 );
and ( n61381 , n61380 , n33187 );
not ( n61382 , n48765 );
and ( n61383 , n61382 , n48668 );
xor ( n61384 , n48961 , n48978 );
and ( n61385 , n61384 , n48765 );
or ( n61386 , n61383 , n61385 );
and ( n61387 , n61386 , n33180 );
not ( n61388 , n49054 );
and ( n61389 , n61388 , n48668 );
not ( n61390 , n48845 );
xor ( n61391 , n48668 , n48978 );
and ( n61392 , n61390 , n61391 );
xor ( n61393 , n49216 , n49217 );
and ( n61394 , n61393 , n48845 );
or ( n61395 , n61392 , n61394 );
and ( n61396 , n61395 , n49054 );
or ( n61397 , n61389 , n61396 );
and ( n61398 , n61397 , n33178 );
and ( n61399 , n49216 , n49275 );
or ( n61400 , n61363 , n61365 , n61367 , n61369 , n61371 , n61376 , n61381 , n61387 , n61398 , n61399 );
and ( n61401 , n61400 , n33208 );
and ( n61402 , n42695 , n35056 );
and ( n61403 , n48668 , n49286 );
or ( n61404 , C0 , n61401 , n61402 , n61403 );
buf ( n61405 , n61404 );
buf ( n61406 , n61405 );
buf ( n61407 , n30987 );
buf ( n61408 , n31655 );
buf ( n61409 , n30987 );
buf ( n61410 , n31655 );
not ( n61411 , n34150 );
and ( n61412 , n61411 , n32865 );
not ( n61413 , n59105 );
and ( n61414 , n61413 , n32865 );
and ( n61415 , n32889 , n59105 );
or ( n61416 , n61414 , n61415 );
and ( n61417 , n61416 , n34150 );
or ( n61418 , n61412 , n61417 );
and ( n61419 , n61418 , n33381 );
not ( n61420 , n59113 );
not ( n61421 , n59105 );
and ( n61422 , n61421 , n32865 );
and ( n61423 , n52819 , n59105 );
or ( n61424 , n61422 , n61423 );
and ( n61425 , n61420 , n61424 );
and ( n61426 , n52819 , n59113 );
or ( n61427 , n61425 , n61426 );
and ( n61428 , n61427 , n33375 );
not ( n61429 , n32968 );
not ( n61430 , n59113 );
not ( n61431 , n59105 );
and ( n61432 , n61431 , n32865 );
and ( n61433 , n52819 , n59105 );
or ( n61434 , n61432 , n61433 );
and ( n61435 , n61430 , n61434 );
and ( n61436 , n52819 , n59113 );
or ( n61437 , n61435 , n61436 );
and ( n61438 , n61429 , n61437 );
not ( n61439 , n59133 );
not ( n61440 , n59135 );
and ( n61441 , n61440 , n61437 );
and ( n61442 , n52845 , n59135 );
or ( n61443 , n61441 , n61442 );
and ( n61444 , n61439 , n61443 );
and ( n61445 , n52855 , n59133 );
or ( n61446 , n61444 , n61445 );
and ( n61447 , n61446 , n32968 );
or ( n61448 , n61438 , n61447 );
and ( n61449 , n61448 , n33370 );
and ( n61450 , n32865 , n35062 );
or ( n61451 , C0 , n61419 , n61428 , n61449 , n61450 );
buf ( n61452 , n61451 );
buf ( n61453 , n61452 );
buf ( n61454 , n31655 );
buf ( n61455 , n30987 );
xor ( n61456 , n46198 , n49994 );
and ( n61457 , n61456 , n32431 );
not ( n61458 , n50002 );
and ( n61459 , n61458 , n46198 );
and ( n61460 , n40507 , n50002 );
or ( n61461 , n61459 , n61460 );
and ( n61462 , n61461 , n32419 );
not ( n61463 , n50008 );
and ( n61464 , n61463 , n46198 );
not ( n61465 , n47910 );
buf ( n61466 , RI15b5f478_1116);
and ( n61467 , n61465 , n61466 );
not ( n61468 , n48101 );
and ( n61469 , n61468 , n48025 );
xor ( n61470 , n50021 , n50024 );
and ( n61471 , n61470 , n48101 );
or ( n61472 , n61469 , n61471 );
and ( n61473 , n61472 , n47910 );
or ( n61474 , n61467 , n61473 );
and ( n61475 , n61474 , n50008 );
or ( n61476 , n61464 , n61475 );
and ( n61477 , n61476 , n32415 );
not ( n61478 , n50067 );
and ( n61479 , n61478 , n46198 );
and ( n61480 , n32001 , n47357 );
and ( n61481 , n32003 , n47359 );
and ( n61482 , n32005 , n47361 );
and ( n61483 , n32007 , n47363 );
and ( n61484 , n32009 , n47365 );
and ( n61485 , n32011 , n47367 );
and ( n61486 , n32013 , n47369 );
and ( n61487 , n32015 , n47371 );
and ( n61488 , n32017 , n47373 );
and ( n61489 , n32019 , n47375 );
and ( n61490 , n32021 , n47377 );
and ( n61491 , n32023 , n47379 );
and ( n61492 , n32025 , n47381 );
and ( n61493 , n32027 , n47383 );
and ( n61494 , n32029 , n47385 );
and ( n61495 , n32031 , n47387 );
or ( n61496 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 );
and ( n61497 , n61496 , n50067 );
or ( n61498 , n61479 , n61497 );
and ( n61499 , n61498 , n32411 );
and ( n61500 , n46198 , n50098 );
or ( n61501 , n61457 , n61462 , n61477 , n61499 , n61500 );
and ( n61502 , n61501 , n32456 );
and ( n61503 , n46198 , n47409 );
or ( n61504 , C0 , n61502 , n61503 );
buf ( n61505 , n61504 );
buf ( n61506 , n61505 );
not ( n61507 , n46356 );
and ( n61508 , n61507 , n31358 );
not ( n61509 , n50109 );
and ( n61510 , n61509 , n31358 );
and ( n61511 , n31372 , n50109 );
or ( n61512 , n61510 , n61511 );
and ( n61513 , n61512 , n46356 );
or ( n61514 , n61508 , n61513 );
and ( n61515 , n61514 , n31649 );
not ( n61516 , n50117 );
not ( n61517 , n50109 );
and ( n61518 , n61517 , n31358 );
and ( n61519 , n47849 , n50109 );
or ( n61520 , n61518 , n61519 );
and ( n61521 , n61516 , n61520 );
and ( n61522 , n47849 , n50117 );
or ( n61523 , n61521 , n61522 );
and ( n61524 , n61523 , n31643 );
not ( n61525 , n31452 );
not ( n61526 , n50117 );
not ( n61527 , n50109 );
and ( n61528 , n61527 , n31358 );
and ( n61529 , n47849 , n50109 );
or ( n61530 , n61528 , n61529 );
and ( n61531 , n61526 , n61530 );
and ( n61532 , n47849 , n50117 );
or ( n61533 , n61531 , n61532 );
and ( n61534 , n61525 , n61533 );
not ( n61535 , n50142 );
not ( n61536 , n50144 );
and ( n61537 , n61536 , n61533 );
and ( n61538 , n47877 , n50144 );
or ( n61539 , n61537 , n61538 );
and ( n61540 , n61535 , n61539 );
and ( n61541 , n47887 , n50142 );
or ( n61542 , n61540 , n61541 );
and ( n61543 , n61542 , n31452 );
or ( n61544 , n61534 , n61543 );
and ( n61545 , n61544 , n31638 );
and ( n61546 , n31358 , n47277 );
or ( n61547 , C0 , n61515 , n61524 , n61545 , n61546 );
buf ( n61548 , n61547 );
buf ( n61549 , n61548 );
buf ( n61550 , n30987 );
buf ( n61551 , n31655 );
buf ( n61552 , n31655 );
buf ( n61553 , n30987 );
xor ( n61554 , n33115 , n52221 );
and ( n61555 , n61554 , n33201 );
not ( n61556 , n41576 );
and ( n61557 , n61556 , n33115 );
and ( n61558 , n32657 , n52252 );
and ( n61559 , n32659 , n52254 );
and ( n61560 , n32661 , n52256 );
and ( n61561 , n32663 , n52258 );
and ( n61562 , n32665 , n52260 );
and ( n61563 , n32667 , n52262 );
and ( n61564 , n32669 , n52264 );
and ( n61565 , n32671 , n52266 );
and ( n61566 , n32673 , n52268 );
and ( n61567 , n32675 , n52270 );
and ( n61568 , n32677 , n52272 );
and ( n61569 , n32679 , n52274 );
and ( n61570 , n32681 , n52276 );
and ( n61571 , n32683 , n52278 );
and ( n61572 , n32685 , n52280 );
and ( n61573 , n32687 , n52282 );
or ( n61574 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 );
and ( n61575 , n61574 , n41576 );
or ( n61576 , n61557 , n61575 );
and ( n61577 , n61576 , n33189 );
and ( n61578 , n33115 , n41592 );
or ( n61579 , n61555 , n61577 , n61578 );
and ( n61580 , n61579 , n33208 );
and ( n61581 , n33115 , n39805 );
or ( n61582 , C0 , n61580 , n61581 );
buf ( n61583 , n61582 );
buf ( n61584 , n61583 );
buf ( n61585 , n30987 );
buf ( n61586 , n31655 );
buf ( n61587 , n31655 );
not ( n61588 , n50828 );
not ( n61589 , n50834 );
and ( n61590 , n61589 , n40562 );
buf ( n61591 , RI15b540f0_733);
and ( n61592 , n61591 , n50834 );
or ( n61593 , n61590 , n61592 );
and ( n61594 , n61588 , n61593 );
buf ( n61595 , RI15b60558_1152);
and ( n61596 , n61595 , n50828 );
or ( n61597 , n61594 , n61596 );
buf ( n61598 , n61597 );
buf ( n61599 , n61598 );
buf ( n61600 , n31655 );
buf ( n61601 , n30987 );
not ( n61602 , n34150 );
and ( n61603 , n61602 , n32643 );
not ( n61604 , n56093 );
and ( n61605 , n61604 , n32643 );
and ( n61606 , n32655 , n56093 );
or ( n61607 , n61605 , n61606 );
and ( n61608 , n61607 , n34150 );
or ( n61609 , n61603 , n61608 );
and ( n61610 , n61609 , n33381 );
not ( n61611 , n56101 );
not ( n61612 , n56093 );
and ( n61613 , n61612 , n32643 );
and ( n61614 , n56044 , n56093 );
or ( n61615 , n61613 , n61614 );
and ( n61616 , n61611 , n61615 );
and ( n61617 , n56044 , n56101 );
or ( n61618 , n61616 , n61617 );
and ( n61619 , n61618 , n33375 );
not ( n61620 , n32968 );
not ( n61621 , n56101 );
not ( n61622 , n56093 );
and ( n61623 , n61622 , n32643 );
and ( n61624 , n56044 , n56093 );
or ( n61625 , n61623 , n61624 );
and ( n61626 , n61621 , n61625 );
and ( n61627 , n56044 , n56101 );
or ( n61628 , n61626 , n61627 );
and ( n61629 , n61620 , n61628 );
not ( n61630 , n56121 );
not ( n61631 , n56123 );
and ( n61632 , n61631 , n61628 );
and ( n61633 , n56068 , n56123 );
or ( n61634 , n61632 , n61633 );
and ( n61635 , n61630 , n61634 );
and ( n61636 , n56076 , n56121 );
or ( n61637 , n61635 , n61636 );
and ( n61638 , n61637 , n32968 );
or ( n61639 , n61629 , n61638 );
and ( n61640 , n61639 , n33370 );
and ( n61641 , n32643 , n35062 );
or ( n61642 , C0 , n61610 , n61619 , n61640 , n61641 );
buf ( n61643 , n61642 );
buf ( n61644 , n61643 );
not ( n61645 , n34150 );
and ( n61646 , n61645 , n32885 );
not ( n61647 , n56140 );
and ( n61648 , n61647 , n32885 );
and ( n61649 , n32889 , n56140 );
or ( n61650 , n61648 , n61649 );
and ( n61651 , n61650 , n34150 );
or ( n61652 , n61646 , n61651 );
and ( n61653 , n61652 , n33381 );
not ( n61654 , n56148 );
not ( n61655 , n56140 );
and ( n61656 , n61655 , n32885 );
and ( n61657 , n52819 , n56140 );
or ( n61658 , n61656 , n61657 );
and ( n61659 , n61654 , n61658 );
and ( n61660 , n52819 , n56148 );
or ( n61661 , n61659 , n61660 );
and ( n61662 , n61661 , n33375 );
not ( n61663 , n32968 );
not ( n61664 , n56148 );
not ( n61665 , n56140 );
and ( n61666 , n61665 , n32885 );
and ( n61667 , n52819 , n56140 );
or ( n61668 , n61666 , n61667 );
and ( n61669 , n61664 , n61668 );
and ( n61670 , n52819 , n56148 );
or ( n61671 , n61669 , n61670 );
and ( n61672 , n61663 , n61671 );
not ( n61673 , n56168 );
not ( n61674 , n56170 );
and ( n61675 , n61674 , n61671 );
and ( n61676 , n52845 , n56170 );
or ( n61677 , n61675 , n61676 );
and ( n61678 , n61673 , n61677 );
and ( n61679 , n52855 , n56168 );
or ( n61680 , n61678 , n61679 );
and ( n61681 , n61680 , n32968 );
or ( n61682 , n61672 , n61681 );
and ( n61683 , n61682 , n33370 );
and ( n61684 , n32885 , n35062 );
or ( n61685 , C0 , n61653 , n61662 , n61683 , n61684 );
buf ( n61686 , n61685 );
buf ( n61687 , n61686 );
buf ( n61688 , n30987 );
buf ( n61689 , n31655 );
buf ( n61690 , n30987 );
and ( n61691 , n60616 , n33377 );
not ( n61692 , n48545 );
buf ( n61693 , RI15b47490_297);
and ( n61694 , n61692 , n61693 );
and ( n61695 , n60622 , n48545 );
or ( n61696 , n61694 , n61695 );
and ( n61697 , n61696 , n32890 );
not ( n61698 , n48557 );
and ( n61699 , n61698 , n61693 );
and ( n61700 , n60622 , n48557 );
or ( n61701 , n61699 , n61700 );
and ( n61702 , n61701 , n33038 );
and ( n61703 , n61693 , n48571 );
or ( n61704 , n61697 , n61702 , n61703 );
and ( n61705 , n61704 , n33208 );
and ( n61706 , n61693 , n48577 );
or ( n61707 , C0 , n61691 , n61705 , n61706 );
buf ( n61708 , n61707 );
buf ( n61709 , n61708 );
buf ( n61710 , n30987 );
buf ( n61711 , n31655 );
buf ( n61712 , n31655 );
buf ( n61713 , n30987 );
buf ( n61714 , n30987 );
buf ( n61715 , n31655 );
buf ( n61716 , n33381 );
buf ( n61717 , n33379 );
not ( n61718 , n57838 );
not ( n61719 , n57840 );
and ( n61720 , n61719 , n32513 );
buf ( n61721 , n61720 );
and ( n61722 , n61721 , n33038 );
and ( n61723 , n32513 , n57852 );
or ( n61724 , n61722 , n61723 );
and ( n61725 , n61718 , n61724 );
buf ( n61726 , n61725 );
and ( n61727 , n61726 , n33208 );
or ( n61728 , C0 , n61716 , n61717 , C0 , n61727 , C0 , C0 , C0 , C0 , C0 );
buf ( n61729 , n61728 );
buf ( n61730 , n61729 );
buf ( n61731 , n31655 );
buf ( n61732 , n30987 );
buf ( n61733 , n30987 );
and ( n61734 , n58018 , n33377 );
not ( n61735 , n48545 );
buf ( n61736 , RI15b471c0_291);
and ( n61737 , n61735 , n61736 );
and ( n61738 , n58024 , n48545 );
or ( n61739 , n61737 , n61738 );
and ( n61740 , n61739 , n32890 );
not ( n61741 , n48557 );
and ( n61742 , n61741 , n61736 );
and ( n61743 , n58024 , n48557 );
or ( n61744 , n61742 , n61743 );
and ( n61745 , n61744 , n33038 );
and ( n61746 , n61736 , n48571 );
or ( n61747 , n61740 , n61745 , n61746 );
and ( n61748 , n61747 , n33208 );
and ( n61749 , n61736 , n48577 );
or ( n61750 , C0 , n61734 , n61748 , n61749 );
buf ( n61751 , n61750 );
buf ( n61752 , n61751 );
buf ( n61753 , n31655 );
buf ( n61754 , n31655 );
buf ( n61755 , n30987 );
and ( n61756 , n49079 , n48639 );
not ( n61757 , n48642 );
and ( n61758 , n61757 , n48604 );
and ( n61759 , n49079 , n48642 );
or ( n61760 , n61758 , n61759 );
and ( n61761 , n61760 , n32890 );
not ( n61762 , n48648 );
and ( n61763 , n61762 , n48604 );
and ( n61764 , n49079 , n48648 );
or ( n61765 , n61763 , n61764 );
and ( n61766 , n61765 , n32924 );
not ( n61767 , n48654 );
and ( n61768 , n61767 , n48604 );
and ( n61769 , n49079 , n48654 );
or ( n61770 , n61768 , n61769 );
and ( n61771 , n61770 , n33038 );
not ( n61772 , n48660 );
and ( n61773 , n61772 , n48604 );
and ( n61774 , n49079 , n48660 );
or ( n61775 , n61773 , n61774 );
and ( n61776 , n61775 , n33172 );
not ( n61777 , n41576 );
and ( n61778 , n61777 , n48604 );
and ( n61779 , n48789 , n41576 );
or ( n61780 , n61778 , n61779 );
and ( n61781 , n61780 , n33189 );
not ( n61782 , n48730 );
and ( n61783 , n61782 , n48604 );
and ( n61784 , n48789 , n48730 );
or ( n61785 , n61783 , n61784 );
and ( n61786 , n61785 , n33187 );
not ( n61787 , n48765 );
and ( n61788 , n61787 , n48604 );
and ( n61789 , n59773 , n48765 );
or ( n61790 , n61788 , n61789 );
and ( n61791 , n61790 , n33180 );
not ( n61792 , n49054 );
and ( n61793 , n61792 , n48604 );
and ( n61794 , n59786 , n49054 );
or ( n61795 , n61793 , n61794 );
and ( n61796 , n61795 , n33178 );
and ( n61797 , n49188 , n49275 );
or ( n61798 , n61756 , n61761 , n61766 , n61771 , n61776 , n61781 , n61786 , n61791 , n61796 , n61797 );
and ( n61799 , n61798 , n33208 );
and ( n61800 , n32997 , n35056 );
and ( n61801 , n48604 , n49286 );
or ( n61802 , C0 , n61799 , n61800 , n61801 );
buf ( n61803 , n61802 );
buf ( n61804 , n61803 );
buf ( n61805 , n30987 );
buf ( n61806 , n31655 );
buf ( n61807 , n31655 );
buf ( n61808 , n30987 );
not ( n61809 , n40163 );
and ( n61810 , n61809 , n32023 );
not ( n61811 , n45161 );
and ( n61812 , n61811 , n32023 );
and ( n61813 , n32147 , n45161 );
or ( n61814 , n61812 , n61813 );
and ( n61815 , n61814 , n40163 );
or ( n61816 , n61810 , n61815 );
and ( n61817 , n61816 , n32498 );
not ( n61818 , n45170 );
not ( n61819 , n45161 );
and ( n61820 , n61819 , n32023 );
and ( n61821 , n49314 , n45161 );
or ( n61822 , n61820 , n61821 );
and ( n61823 , n61818 , n61822 );
and ( n61824 , n49314 , n45170 );
or ( n61825 , n61823 , n61824 );
and ( n61826 , n61825 , n32473 );
not ( n61827 , n32475 );
not ( n61828 , n45170 );
not ( n61829 , n45161 );
and ( n61830 , n61829 , n32023 );
and ( n61831 , n49314 , n45161 );
or ( n61832 , n61830 , n61831 );
and ( n61833 , n61828 , n61832 );
and ( n61834 , n49314 , n45170 );
or ( n61835 , n61833 , n61834 );
and ( n61836 , n61827 , n61835 );
not ( n61837 , n45196 );
not ( n61838 , n45199 );
and ( n61839 , n61838 , n61835 );
and ( n61840 , n49340 , n45199 );
or ( n61841 , n61839 , n61840 );
and ( n61842 , n61837 , n61841 );
and ( n61843 , n49348 , n45196 );
or ( n61844 , n61842 , n61843 );
and ( n61845 , n61844 , n32475 );
or ( n61846 , n61836 , n61845 );
and ( n61847 , n61846 , n32486 );
and ( n61848 , n32023 , n41278 );
or ( n61849 , C0 , n61817 , n61826 , n61847 , n61848 );
buf ( n61850 , n61849 );
buf ( n61851 , n61850 );
and ( n61852 , n44763 , n44804 );
and ( n61853 , n45330 , n61852 );
xor ( n61854 , n41611 , n61853 );
and ( n61855 , n61854 , n31548 );
not ( n61856 , n44807 );
and ( n61857 , n61856 , n41611 );
and ( n61858 , n41881 , n44807 );
or ( n61859 , n61857 , n61858 );
and ( n61860 , n61859 , n31408 );
not ( n61861 , n44817 );
and ( n61862 , n61861 , n41611 );
buf ( n61863 , n61862 );
and ( n61864 , n61863 , n31521 );
not ( n61865 , n45059 );
and ( n61866 , n61865 , n41611 );
buf ( n61867 , n61866 );
and ( n61868 , n61867 , n31536 );
and ( n61869 , n41611 , n45148 );
or ( n61870 , n61855 , n61860 , n61864 , n61868 , n61869 );
and ( n61871 , n61870 , n31557 );
and ( n61872 , n41611 , n40154 );
or ( n61873 , C0 , n61871 , n61872 );
buf ( n61874 , n61873 );
buf ( n61875 , n61874 );
buf ( n61876 , n30987 );
buf ( n61877 , n31655 );
buf ( n61878 , n31655 );
and ( n61879 , n47660 , n50275 );
not ( n61880 , n50278 );
and ( n61881 , n61880 , n47573 );
and ( n61882 , n47660 , n50278 );
or ( n61883 , n61881 , n61882 );
and ( n61884 , n61883 , n32421 );
not ( n61885 , n50002 );
and ( n61886 , n61885 , n47573 );
and ( n61887 , n47660 , n50002 );
or ( n61888 , n61886 , n61887 );
and ( n61889 , n61888 , n32419 );
not ( n61890 , n50289 );
and ( n61891 , n61890 , n47573 );
and ( n61892 , n47660 , n50289 );
or ( n61893 , n61891 , n61892 );
and ( n61894 , n61893 , n32417 );
not ( n61895 , n50008 );
and ( n61896 , n61895 , n47573 );
and ( n61897 , n47660 , n50008 );
or ( n61898 , n61896 , n61897 );
and ( n61899 , n61898 , n32415 );
not ( n61900 , n47331 );
and ( n61901 , n61900 , n47573 );
and ( n61902 , n47605 , n47331 );
or ( n61903 , n61901 , n61902 );
and ( n61904 , n61903 , n32413 );
not ( n61905 , n50067 );
and ( n61906 , n61905 , n47573 );
and ( n61907 , n47605 , n50067 );
or ( n61908 , n61906 , n61907 );
and ( n61909 , n61908 , n32411 );
not ( n61910 , n31728 );
and ( n61911 , n61910 , n47573 );
xor ( n61912 , n47605 , n47624 );
and ( n61913 , n61912 , n31728 );
or ( n61914 , n61911 , n61913 );
and ( n61915 , n61914 , n32253 );
not ( n61916 , n32283 );
and ( n61917 , n61916 , n47573 );
not ( n61918 , n31823 );
xor ( n61919 , n47660 , n47679 );
and ( n61920 , n61918 , n61919 );
xnor ( n61921 , n47710 , n47729 );
and ( n61922 , n61921 , n31823 );
or ( n61923 , n61920 , n61922 );
and ( n61924 , n61923 , n32283 );
or ( n61925 , n61917 , n61924 );
and ( n61926 , n61925 , n32398 );
and ( n61927 , n47710 , n50334 );
or ( n61928 , n61879 , n61884 , n61889 , n61894 , n61899 , n61904 , n61909 , n61915 , n61926 , n61927 );
and ( n61929 , n61928 , n32456 );
and ( n61930 , n37553 , n32489 );
and ( n61931 , n47573 , n50345 );
or ( n61932 , C0 , n61929 , n61930 , n61931 );
buf ( n61933 , n61932 );
buf ( n61934 , n61933 );
buf ( n61935 , n30987 );
not ( n61936 , n36587 );
and ( n61937 , n61936 , n36566 );
xor ( n61938 , n36566 , n36091 );
xor ( n61939 , n36549 , n36091 );
xor ( n61940 , n36532 , n36091 );
xor ( n61941 , n36515 , n36091 );
xor ( n61942 , n36498 , n36091 );
and ( n61943 , n50172 , n50215 );
and ( n61944 , n61942 , n61943 );
and ( n61945 , n61941 , n61944 );
and ( n61946 , n61940 , n61945 );
and ( n61947 , n61939 , n61946 );
xor ( n61948 , n61938 , n61947 );
and ( n61949 , n61948 , n36587 );
or ( n61950 , n61937 , n61949 );
and ( n61951 , n61950 , n36596 );
not ( n61952 , n37485 );
and ( n61953 , n61952 , n37468 );
xor ( n61954 , n37468 , n36993 );
xor ( n61955 , n37451 , n36993 );
xor ( n61956 , n37434 , n36993 );
xor ( n61957 , n37417 , n36993 );
xor ( n61958 , n37400 , n36993 );
and ( n61959 , n50222 , n50265 );
and ( n61960 , n61958 , n61959 );
and ( n61961 , n61957 , n61960 );
and ( n61962 , n61956 , n61961 );
and ( n61963 , n61955 , n61962 );
xor ( n61964 , n61954 , n61963 );
and ( n61965 , n61964 , n37485 );
or ( n61966 , n61953 , n61965 );
and ( n61967 , n61966 , n37494 );
and ( n61968 , n41867 , n37506 );
or ( n61969 , n61951 , n61967 , n61968 );
buf ( n61970 , n61969 );
buf ( n61971 , n61970 );
buf ( n61972 , n30987 );
not ( n61973 , n46356 );
and ( n61974 , n61973 , n31201 );
nor ( n61975 , n46359 , n31021 , n31017 , n31013 , n31009 );
not ( n61976 , n61975 );
and ( n61977 , n61976 , n31201 );
and ( n61978 , n31205 , n61975 );
or ( n61979 , n61977 , n61978 );
and ( n61980 , n61979 , n46356 );
or ( n61981 , n61974 , n61980 );
and ( n61982 , n61981 , n31649 );
nor ( n61983 , n46374 , n46379 , n46386 , n46392 , C0 );
not ( n61984 , n61983 );
not ( n61985 , n61975 );
and ( n61986 , n61985 , n31201 );
and ( n61987 , n50125 , n61975 );
or ( n61988 , n61986 , n61987 );
and ( n61989 , n61984 , n61988 );
and ( n61990 , n50125 , n61983 );
or ( n61991 , n61989 , n61990 );
and ( n61992 , n61991 , n31643 );
not ( n61993 , n31452 );
not ( n61994 , n61983 );
not ( n61995 , n61975 );
and ( n61996 , n61995 , n31201 );
and ( n61997 , n50125 , n61975 );
or ( n61998 , n61996 , n61997 );
and ( n61999 , n61994 , n61998 );
and ( n62000 , n50125 , n61983 );
or ( n62001 , n61999 , n62000 );
and ( n62002 , n61993 , n62001 );
nor ( n62003 , n46520 , n46528 , n46539 , n46549 , C0 );
not ( n62004 , n62003 );
nor ( n62005 , n46552 , n46524 , n46534 , n46544 , C0 );
not ( n62006 , n62005 );
and ( n62007 , n62006 , n62001 );
and ( n62008 , n50151 , n62005 );
or ( n62009 , n62007 , n62008 );
and ( n62010 , n62004 , n62009 );
and ( n62011 , n50159 , n62003 );
or ( n62012 , n62010 , n62011 );
and ( n62013 , n62012 , n31452 );
or ( n62014 , n62002 , n62013 );
and ( n62015 , n62014 , n31638 );
and ( n62016 , n31201 , n47277 );
or ( n62017 , C0 , n61982 , n61992 , n62015 , n62016 );
buf ( n62018 , n62017 );
buf ( n62019 , n62018 );
xor ( n62020 , n49577 , n60317 );
and ( n62021 , n62020 , n32433 );
not ( n62022 , n47331 );
and ( n62023 , n62022 , n49577 );
and ( n62024 , n31826 , n60510 );
and ( n62025 , n31828 , n60512 );
and ( n62026 , n31830 , n60514 );
and ( n62027 , n31832 , n60516 );
and ( n62028 , n31834 , n60518 );
and ( n62029 , n31836 , n60520 );
and ( n62030 , n31838 , n60522 );
and ( n62031 , n31840 , n60524 );
and ( n62032 , n31842 , n60526 );
and ( n62033 , n31844 , n60528 );
and ( n62034 , n31846 , n60530 );
and ( n62035 , n31848 , n60532 );
and ( n62036 , n31850 , n60534 );
and ( n62037 , n31852 , n60536 );
and ( n62038 , n31854 , n60538 );
and ( n62039 , n31856 , n60540 );
or ( n62040 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 );
and ( n62041 , n62040 , n47331 );
or ( n62042 , n62023 , n62041 );
and ( n62043 , n62042 , n32413 );
and ( n62044 , n49577 , n47402 );
or ( n62045 , n62021 , n62043 , n62044 );
and ( n62046 , n62045 , n32456 );
and ( n62047 , n49577 , n47409 );
or ( n62048 , C0 , n62046 , n62047 );
buf ( n62049 , n62048 );
buf ( n62050 , n62049 );
buf ( n62051 , n30987 );
buf ( n62052 , n31655 );
buf ( n62053 , n31655 );
not ( n62054 , n38443 );
and ( n62055 , n62054 , n38167 );
xor ( n62056 , n53472 , n53497 );
and ( n62057 , n62056 , n38443 );
or ( n62058 , n62055 , n62057 );
and ( n62059 , n62058 , n38450 );
not ( n62060 , n39339 );
and ( n62061 , n62060 , n39067 );
xor ( n62062 , n53528 , n53553 );
and ( n62063 , n62062 , n39339 );
or ( n62064 , n62061 , n62063 );
and ( n62065 , n62064 , n39346 );
and ( n62066 , n40212 , n39359 );
or ( n62067 , n62059 , n62065 , n62066 );
buf ( n62068 , n62067 );
buf ( n62069 , n62068 );
buf ( n62070 , n31655 );
and ( n62071 , n33494 , n46356 );
buf ( n62072 , n62071 );
and ( n62073 , n62072 , n31649 );
and ( n62074 , n52536 , n31647 );
and ( n62075 , n42321 , n48455 );
not ( n62076 , n48457 );
and ( n62077 , n62076 , n31018 );
and ( n62078 , n42321 , n48457 );
or ( n62079 , n62077 , n62078 );
and ( n62080 , n62079 , n31373 );
not ( n62081 , n44807 );
and ( n62082 , n62081 , n31018 );
and ( n62083 , n42317 , n44807 );
or ( n62084 , n62082 , n62083 );
and ( n62085 , n62084 , n31408 );
not ( n62086 , n48468 );
and ( n62087 , n62086 , n31018 );
and ( n62088 , n42321 , n48468 );
or ( n62089 , n62087 , n62088 );
and ( n62090 , n62089 , n31468 );
not ( n62091 , n44817 );
and ( n62092 , n62091 , n31018 );
and ( n62093 , n42321 , n44817 );
or ( n62094 , n62092 , n62093 );
and ( n62095 , n62094 , n31521 );
not ( n62096 , n39979 );
and ( n62097 , n62096 , n31018 );
and ( n62098 , n31022 , n31026 );
xnor ( n62099 , n31018 , n62098 );
not ( n62100 , n62099 );
buf ( n62101 , n62100 );
buf ( n62102 , n62101 );
not ( n62103 , n62102 );
and ( n62104 , n62103 , n39979 );
or ( n62105 , n62097 , n62104 );
and ( n62106 , n62105 , n31538 );
not ( n62107 , n45059 );
and ( n62108 , n62107 , n31018 );
and ( n62109 , n62103 , n45059 );
or ( n62110 , n62108 , n62109 );
and ( n62111 , n62110 , n31536 );
and ( n62112 , n31018 , n61216 );
and ( n62113 , n33494 , n48513 );
or ( n62114 , n62075 , n62080 , n62085 , n62090 , n62095 , n62106 , n62111 , n62112 , n62113 );
and ( n62115 , n62114 , n31557 );
and ( n62116 , n31018 , n61220 );
or ( n62117 , C0 , n62073 , n62074 , n62115 , n62116 );
buf ( n62118 , n62117 );
buf ( n62119 , n62118 );
buf ( n62120 , n30987 );
not ( n62121 , n34150 );
and ( n62122 , n62121 , n32628 );
not ( n62123 , n41392 );
and ( n62124 , n62123 , n32628 );
and ( n62125 , n32655 , n41392 );
or ( n62126 , n62124 , n62125 );
and ( n62127 , n62126 , n34150 );
or ( n62128 , n62122 , n62127 );
and ( n62129 , n62128 , n33381 );
not ( n62130 , n41402 );
not ( n62131 , n41392 );
and ( n62132 , n62131 , n32628 );
and ( n62133 , n56044 , n41392 );
or ( n62134 , n62132 , n62133 );
and ( n62135 , n62130 , n62134 );
and ( n62136 , n56044 , n41402 );
or ( n62137 , n62135 , n62136 );
and ( n62138 , n62137 , n33375 );
not ( n62139 , n32968 );
not ( n62140 , n41402 );
not ( n62141 , n41392 );
and ( n62142 , n62141 , n32628 );
and ( n62143 , n56044 , n41392 );
or ( n62144 , n62142 , n62143 );
and ( n62145 , n62140 , n62144 );
and ( n62146 , n56044 , n41402 );
or ( n62147 , n62145 , n62146 );
and ( n62148 , n62139 , n62147 );
not ( n62149 , n41424 );
not ( n62150 , n41428 );
and ( n62151 , n62150 , n62147 );
and ( n62152 , n56068 , n41428 );
or ( n62153 , n62151 , n62152 );
and ( n62154 , n62149 , n62153 );
and ( n62155 , n56076 , n41424 );
or ( n62156 , n62154 , n62155 );
and ( n62157 , n62156 , n32968 );
or ( n62158 , n62148 , n62157 );
and ( n62159 , n62158 , n33370 );
and ( n62160 , n32628 , n35062 );
or ( n62161 , C0 , n62129 , n62138 , n62159 , n62160 );
buf ( n62162 , n62161 );
buf ( n62163 , n62162 );
buf ( n62164 , n31655 );
buf ( n62165 , n30987 );
buf ( n62166 , n30987 );
buf ( n62167 , n31655 );
buf ( n62168 , RI15b47238_292);
buf ( n62169 , n62168 );
buf ( n62170 , n30987 );
xor ( n62171 , n41665 , n44780 );
and ( n62172 , n62171 , n31548 );
not ( n62173 , n44807 );
and ( n62174 , n62173 , n41665 );
and ( n62175 , n41950 , n44807 );
or ( n62176 , n62174 , n62175 );
and ( n62177 , n62176 , n31408 );
not ( n62178 , n44817 );
and ( n62179 , n62178 , n41665 );
not ( n62180 , n41835 );
and ( n62181 , n62180 , n56333 );
not ( n62182 , n42124 );
and ( n62183 , n62182 , n41960 );
xor ( n62184 , n42130 , n42140 );
and ( n62185 , n62184 , n42124 );
or ( n62186 , n62183 , n62185 );
and ( n62187 , n62186 , n41835 );
or ( n62188 , n62181 , n62187 );
and ( n62189 , n62188 , n44817 );
or ( n62190 , n62179 , n62189 );
and ( n62191 , n62190 , n31521 );
not ( n62192 , n45059 );
and ( n62193 , n62192 , n41665 );
and ( n62194 , n33571 , n45059 );
or ( n62195 , n62193 , n62194 );
and ( n62196 , n62195 , n31536 );
and ( n62197 , n41665 , n45148 );
or ( n62198 , n62172 , n62177 , n62191 , n62196 , n62197 );
and ( n62199 , n62198 , n31557 );
and ( n62200 , n41665 , n40154 );
or ( n62201 , C0 , n62199 , n62200 );
buf ( n62202 , n62201 );
buf ( n62203 , n62202 );
buf ( n62204 , n31655 );
not ( n62205 , n40163 );
and ( n62206 , n62205 , n31947 );
not ( n62207 , n50540 );
and ( n62208 , n62207 , n31947 );
and ( n62209 , n32183 , n50540 );
or ( n62210 , n62208 , n62209 );
and ( n62211 , n62210 , n40163 );
or ( n62212 , n62206 , n62211 );
and ( n62213 , n62212 , n32498 );
not ( n62214 , n50548 );
not ( n62215 , n50540 );
and ( n62216 , n62215 , n31947 );
and ( n62217 , n45178 , n50540 );
or ( n62218 , n62216 , n62217 );
and ( n62219 , n62214 , n62218 );
and ( n62220 , n45178 , n50548 );
or ( n62221 , n62219 , n62220 );
and ( n62222 , n62221 , n32473 );
not ( n62223 , n32475 );
not ( n62224 , n50548 );
not ( n62225 , n50540 );
and ( n62226 , n62225 , n31947 );
and ( n62227 , n45178 , n50540 );
or ( n62228 , n62226 , n62227 );
and ( n62229 , n62224 , n62228 );
and ( n62230 , n45178 , n50548 );
or ( n62231 , n62229 , n62230 );
and ( n62232 , n62223 , n62231 );
not ( n62233 , n50568 );
not ( n62234 , n50570 );
and ( n62235 , n62234 , n62231 );
and ( n62236 , n45206 , n50570 );
or ( n62237 , n62235 , n62236 );
and ( n62238 , n62233 , n62237 );
and ( n62239 , n45214 , n50568 );
or ( n62240 , n62238 , n62239 );
and ( n62241 , n62240 , n32475 );
or ( n62242 , n62232 , n62241 );
and ( n62243 , n62242 , n32486 );
and ( n62244 , n31947 , n41278 );
or ( n62245 , C0 , n62213 , n62222 , n62243 , n62244 );
buf ( n62246 , n62245 );
buf ( n62247 , n62246 );
buf ( n62248 , n30987 );
buf ( n62249 , n30987 );
xor ( n62250 , n49571 , n60320 );
and ( n62251 , n62250 , n32433 );
not ( n62252 , n47331 );
and ( n62253 , n62252 , n49571 );
xor ( n62254 , n60450 , n60544 );
and ( n62255 , n62254 , n47331 );
or ( n62256 , n62253 , n62255 );
and ( n62257 , n62256 , n32413 );
and ( n62258 , n49571 , n47402 );
or ( n62259 , n62251 , n62257 , n62258 );
and ( n62260 , n62259 , n32456 );
and ( n62261 , n49571 , n47409 );
or ( n62262 , C0 , n62260 , n62261 );
buf ( n62263 , n62262 );
buf ( n62264 , n62263 );
not ( n62265 , n46356 );
and ( n62266 , n62265 , n31370 );
not ( n62267 , n60564 );
and ( n62268 , n62267 , n31370 );
and ( n62269 , n31372 , n60564 );
or ( n62270 , n62268 , n62269 );
and ( n62271 , n62270 , n46356 );
or ( n62272 , n62266 , n62271 );
and ( n62273 , n62272 , n31649 );
not ( n62274 , n60572 );
not ( n62275 , n60564 );
and ( n62276 , n62275 , n31370 );
and ( n62277 , n47849 , n60564 );
or ( n62278 , n62276 , n62277 );
and ( n62279 , n62274 , n62278 );
and ( n62280 , n47849 , n60572 );
or ( n62281 , n62279 , n62280 );
and ( n62282 , n62281 , n31643 );
not ( n62283 , n31452 );
not ( n62284 , n60572 );
not ( n62285 , n60564 );
and ( n62286 , n62285 , n31370 );
and ( n62287 , n47849 , n60564 );
or ( n62288 , n62286 , n62287 );
and ( n62289 , n62284 , n62288 );
and ( n62290 , n47849 , n60572 );
or ( n62291 , n62289 , n62290 );
and ( n62292 , n62283 , n62291 );
not ( n62293 , n60592 );
not ( n62294 , n60594 );
and ( n62295 , n62294 , n62291 );
and ( n62296 , n47877 , n60594 );
or ( n62297 , n62295 , n62296 );
and ( n62298 , n62293 , n62297 );
and ( n62299 , n47887 , n60592 );
or ( n62300 , n62298 , n62299 );
and ( n62301 , n62300 , n31452 );
or ( n62302 , n62292 , n62301 );
and ( n62303 , n62302 , n31638 );
and ( n62304 , n31370 , n47277 );
or ( n62305 , C0 , n62273 , n62282 , n62303 , n62304 );
buf ( n62306 , n62305 );
buf ( n62307 , n62306 );
buf ( n62308 , n30987 );
buf ( n62309 , n31655 );
buf ( n62310 , n31655 );
buf ( n62311 , n31655 );
and ( n62312 , n49072 , n48639 );
not ( n62313 , n48642 );
and ( n62314 , n62313 , n48597 );
and ( n62315 , n49072 , n48642 );
or ( n62316 , n62314 , n62315 );
and ( n62317 , n62316 , n32890 );
not ( n62318 , n48648 );
and ( n62319 , n62318 , n48597 );
and ( n62320 , n49072 , n48648 );
or ( n62321 , n62319 , n62320 );
and ( n62322 , n62321 , n32924 );
not ( n62323 , n48654 );
and ( n62324 , n62323 , n48597 );
and ( n62325 , n49072 , n48654 );
or ( n62326 , n62324 , n62325 );
and ( n62327 , n62326 , n33038 );
not ( n62328 , n48660 );
and ( n62329 , n62328 , n48597 );
and ( n62330 , n49072 , n48660 );
or ( n62331 , n62329 , n62330 );
and ( n62332 , n62331 , n33172 );
not ( n62333 , n41576 );
and ( n62334 , n62333 , n48597 );
and ( n62335 , n48782 , n41576 );
or ( n62336 , n62334 , n62335 );
and ( n62337 , n62336 , n33189 );
not ( n62338 , n48730 );
and ( n62339 , n62338 , n48597 );
and ( n62340 , n48782 , n48730 );
or ( n62341 , n62339 , n62340 );
and ( n62342 , n62341 , n33187 );
not ( n62343 , n48765 );
and ( n62344 , n62343 , n48597 );
xor ( n62345 , n48782 , n49006 );
and ( n62346 , n62345 , n48765 );
or ( n62347 , n62344 , n62346 );
and ( n62348 , n62347 , n33180 );
not ( n62349 , n49054 );
and ( n62350 , n62349 , n48597 );
not ( n62351 , n48845 );
xor ( n62352 , n49072 , n49120 );
and ( n62353 , n62351 , n62352 );
xnor ( n62354 , n49181 , n49246 );
and ( n62355 , n62354 , n48845 );
or ( n62356 , n62353 , n62355 );
and ( n62357 , n62356 , n49054 );
or ( n62358 , n62350 , n62357 );
and ( n62359 , n62358 , n33178 );
and ( n62360 , n49181 , n49275 );
or ( n62361 , n62312 , n62317 , n62322 , n62327 , n62332 , n62337 , n62342 , n62348 , n62359 , n62360 );
and ( n62362 , n62361 , n33208 );
and ( n62363 , n32990 , n35056 );
and ( n62364 , n48597 , n49286 );
or ( n62365 , C0 , n62362 , n62363 , n62364 );
buf ( n62366 , n62365 );
buf ( n62367 , n62366 );
buf ( n62368 , n31655 );
buf ( n62369 , n30987 );
buf ( n62370 , n30987 );
buf ( n62371 , n30987 );
buf ( n62372 , n31655 );
buf ( n62373 , n31655 );
or ( n62374 , n44685 , n44682 );
or ( n62375 , n62374 , n44692 );
or ( n62376 , n62375 , n43774 );
or ( n62377 , n62376 , n44694 );
and ( n62378 , n42741 , n62377 );
buf ( n62379 , n62378 );
buf ( n62380 , n62379 );
buf ( n62381 , n30987 );
not ( n62382 , n40163 );
and ( n62383 , n62382 , n32042 );
not ( n62384 , n53227 );
and ( n62385 , n62384 , n32042 );
and ( n62386 , n32130 , n53227 );
or ( n62387 , n62385 , n62386 );
and ( n62388 , n62387 , n40163 );
or ( n62389 , n62383 , n62388 );
and ( n62390 , n62389 , n32498 );
not ( n62391 , n53235 );
not ( n62392 , n53227 );
and ( n62393 , n62392 , n32042 );
and ( n62394 , n45833 , n53227 );
or ( n62395 , n62393 , n62394 );
and ( n62396 , n62391 , n62395 );
and ( n62397 , n45833 , n53235 );
or ( n62398 , n62396 , n62397 );
and ( n62399 , n62398 , n32473 );
not ( n62400 , n32475 );
not ( n62401 , n53235 );
not ( n62402 , n53227 );
and ( n62403 , n62402 , n32042 );
and ( n62404 , n45833 , n53227 );
or ( n62405 , n62403 , n62404 );
and ( n62406 , n62401 , n62405 );
and ( n62407 , n45833 , n53235 );
or ( n62408 , n62406 , n62407 );
and ( n62409 , n62400 , n62408 );
not ( n62410 , n53260 );
not ( n62411 , n53262 );
and ( n62412 , n62411 , n62408 );
and ( n62413 , n45857 , n53262 );
or ( n62414 , n62412 , n62413 );
and ( n62415 , n62410 , n62414 );
and ( n62416 , n45865 , n53260 );
or ( n62417 , n62415 , n62416 );
and ( n62418 , n62417 , n32475 );
or ( n62419 , n62409 , n62418 );
and ( n62420 , n62419 , n32486 );
and ( n62421 , n32042 , n41278 );
or ( n62422 , C0 , n62390 , n62399 , n62420 , n62421 );
buf ( n62423 , n62422 );
buf ( n62424 , n62423 );
buf ( n62425 , RI15b53268_702);
and ( n62426 , n62425 , n31645 );
not ( n62427 , n45274 );
buf ( n62428 , RI15b539e8_718);
and ( n62429 , n62427 , n62428 );
not ( n62430 , n41809 );
and ( n62431 , n62430 , n41792 );
xor ( n62432 , n41792 , n41611 );
xor ( n62433 , n41779 , n41611 );
xor ( n62434 , n41766 , n41611 );
xor ( n62435 , n41753 , n41611 );
and ( n62436 , n53294 , n53297 );
and ( n62437 , n62435 , n62436 );
and ( n62438 , n62434 , n62437 );
and ( n62439 , n62433 , n62438 );
xor ( n62440 , n62432 , n62439 );
and ( n62441 , n62440 , n41809 );
or ( n62442 , n62431 , n62441 );
and ( n62443 , n62442 , n45274 );
or ( n62444 , n62429 , n62443 );
and ( n62445 , n62444 , n31373 );
not ( n62446 , n45280 );
and ( n62447 , n62446 , n62428 );
and ( n62448 , n62442 , n45280 );
or ( n62449 , n62447 , n62448 );
and ( n62450 , n62449 , n31468 );
and ( n62451 , n62428 , n45802 );
or ( n62452 , n62445 , n62450 , n62451 );
and ( n62453 , n62452 , n31557 );
and ( n62454 , n62428 , n45808 );
or ( n62455 , C0 , n62426 , n62453 , n62454 );
buf ( n62456 , n62455 );
buf ( n62457 , n62456 );
buf ( n62458 , n30987 );
buf ( n62459 , n31655 );
buf ( n62460 , n31655 );
buf ( n62461 , n30987 );
buf ( n62462 , n30987 );
buf ( n62463 , n31655 );
not ( n62464 , n34150 );
and ( n62465 , n62464 , n32669 );
not ( n62466 , n57872 );
and ( n62467 , n62466 , n32669 );
and ( n62468 , n32689 , n57872 );
or ( n62469 , n62467 , n62468 );
and ( n62470 , n62469 , n34150 );
or ( n62471 , n62465 , n62470 );
and ( n62472 , n62471 , n33381 );
not ( n62473 , n57880 );
not ( n62474 , n57872 );
and ( n62475 , n62474 , n32669 );
and ( n62476 , n50682 , n57872 );
or ( n62477 , n62475 , n62476 );
and ( n62478 , n62473 , n62477 );
and ( n62479 , n50682 , n57880 );
or ( n62480 , n62478 , n62479 );
and ( n62481 , n62480 , n33375 );
not ( n62482 , n32968 );
not ( n62483 , n57880 );
not ( n62484 , n57872 );
and ( n62485 , n62484 , n32669 );
and ( n62486 , n50682 , n57872 );
or ( n62487 , n62485 , n62486 );
and ( n62488 , n62483 , n62487 );
and ( n62489 , n50682 , n57880 );
or ( n62490 , n62488 , n62489 );
and ( n62491 , n62482 , n62490 );
not ( n62492 , n57900 );
not ( n62493 , n57902 );
and ( n62494 , n62493 , n62490 );
and ( n62495 , n50706 , n57902 );
or ( n62496 , n62494 , n62495 );
and ( n62497 , n62492 , n62496 );
and ( n62498 , n50714 , n57900 );
or ( n62499 , n62497 , n62498 );
and ( n62500 , n62499 , n32968 );
or ( n62501 , n62491 , n62500 );
and ( n62502 , n62501 , n33370 );
and ( n62503 , n32669 , n35062 );
or ( n62504 , C0 , n62472 , n62481 , n62502 , n62503 );
buf ( n62505 , n62504 );
buf ( n62506 , n62505 );
buf ( n62507 , n30987 );
buf ( n62508 , n31655 );
not ( n62509 , n48765 );
and ( n62510 , n62509 , n33221 );
xor ( n62511 , n48776 , n49012 );
and ( n62512 , n62511 , n48765 );
or ( n62513 , n62510 , n62512 );
and ( n62514 , n62513 , n33180 );
not ( n62515 , n49054 );
and ( n62516 , n62515 , n33221 );
not ( n62517 , n48845 );
xor ( n62518 , n49066 , n49126 );
and ( n62519 , n62517 , n62518 );
xnor ( n62520 , n49175 , n49252 );
and ( n62521 , n62520 , n48845 );
or ( n62522 , n62519 , n62521 );
and ( n62523 , n62522 , n49054 );
or ( n62524 , n62516 , n62523 );
and ( n62525 , n62524 , n33178 );
and ( n62526 , n33221 , n49774 );
or ( n62527 , n62514 , n62525 , n62526 );
and ( n62528 , n62527 , n33208 );
and ( n62529 , n33293 , n33375 );
not ( n62530 , n32968 );
and ( n62531 , n62530 , n33293 );
xor ( n62532 , n33221 , n59697 );
and ( n62533 , n62532 , n32968 );
or ( n62534 , n62531 , n62533 );
and ( n62535 , n62534 , n33370 );
and ( n62536 , n32984 , n35056 );
and ( n62537 , n33221 , n49794 );
or ( n62538 , C0 , n62528 , n62529 , n62535 , n62536 , n62537 );
buf ( n62539 , n62538 );
buf ( n62540 , n62539 );
buf ( n62541 , n31655 );
and ( n62542 , n46029 , n32500 );
not ( n62543 , n35211 );
and ( n62544 , n62543 , n37555 );
buf ( n62545 , n62544 );
and ( n62546 , n62545 , n32421 );
not ( n62547 , n35245 );
and ( n62548 , n62547 , n37555 );
buf ( n62549 , n62548 );
and ( n62550 , n62549 , n32419 );
not ( n62551 , n35278 );
and ( n62552 , n62551 , n37555 );
not ( n62553 , n35295 );
and ( n62554 , n62553 , n49585 );
xor ( n62555 , n37555 , n49538 );
and ( n62556 , n62555 , n35295 );
or ( n62557 , n62554 , n62556 );
and ( n62558 , n62557 , n35278 );
or ( n62559 , n62552 , n62558 );
and ( n62560 , n62559 , n32417 );
not ( n62561 , n35331 );
and ( n62562 , n62561 , n37555 );
not ( n62563 , n35294 );
not ( n62564 , n45995 );
and ( n62565 , n62564 , n49585 );
xor ( n62566 , n49586 , n49624 );
and ( n62567 , n62566 , n45995 );
or ( n62568 , n62565 , n62567 );
and ( n62569 , n62563 , n62568 );
and ( n62570 , n62555 , n35294 );
or ( n62571 , n62569 , n62570 );
and ( n62572 , n62571 , n35331 );
or ( n62573 , n62562 , n62572 );
and ( n62574 , n62573 , n32415 );
and ( n62575 , n37555 , n35354 );
or ( n62576 , n62546 , n62550 , n62560 , n62574 , n62575 );
and ( n62577 , n62576 , n32456 );
not ( n62578 , n32475 );
not ( n62579 , n46060 );
and ( n62580 , n62579 , n49675 );
xor ( n62581 , n49676 , n49718 );
and ( n62582 , n62581 , n46060 );
or ( n62583 , n62580 , n62582 );
and ( n62584 , n62578 , n62583 );
and ( n62585 , n37555 , n32475 );
or ( n62586 , n62584 , n62585 );
and ( n62587 , n62586 , n32486 );
buf ( n62588 , n32489 );
and ( n62589 , n37555 , n35367 );
or ( n62590 , C0 , n62542 , n62577 , n62587 , n62588 , n62589 );
buf ( n62591 , n62590 );
buf ( n62592 , n62591 );
buf ( n62593 , n30987 );
buf ( n62594 , n40226 );
buf ( n62595 , n30987 );
and ( n62596 , n49085 , n48639 );
not ( n62597 , n48642 );
and ( n62598 , n62597 , n48607 );
and ( n62599 , n49085 , n48642 );
or ( n62600 , n62598 , n62599 );
and ( n62601 , n62600 , n32890 );
not ( n62602 , n48648 );
and ( n62603 , n62602 , n48607 );
and ( n62604 , n49085 , n48648 );
or ( n62605 , n62603 , n62604 );
and ( n62606 , n62605 , n32924 );
not ( n62607 , n48654 );
and ( n62608 , n62607 , n48607 );
and ( n62609 , n49085 , n48654 );
or ( n62610 , n62608 , n62609 );
and ( n62611 , n62610 , n33038 );
not ( n62612 , n48660 );
and ( n62613 , n62612 , n48607 );
and ( n62614 , n49085 , n48660 );
or ( n62615 , n62613 , n62614 );
and ( n62616 , n62615 , n33172 );
not ( n62617 , n41576 );
and ( n62618 , n62617 , n48607 );
and ( n62619 , n48885 , n41576 );
or ( n62620 , n62618 , n62619 );
and ( n62621 , n62620 , n33189 );
not ( n62622 , n48730 );
and ( n62623 , n62622 , n48607 );
and ( n62624 , n48885 , n48730 );
or ( n62625 , n62623 , n62624 );
and ( n62626 , n62625 , n33187 );
not ( n62627 , n48765 );
and ( n62628 , n62627 , n48607 );
xor ( n62629 , n48885 , n48902 );
xor ( n62630 , n62629 , n48988 );
and ( n62631 , n62630 , n48765 );
or ( n62632 , n62628 , n62631 );
and ( n62633 , n62632 , n33180 );
not ( n62634 , n49054 );
and ( n62635 , n62634 , n48607 );
not ( n62636 , n48845 );
xor ( n62637 , n49085 , n48902 );
xor ( n62638 , n62637 , n49102 );
and ( n62639 , n62636 , n62638 );
xor ( n62640 , n49200 , n49202 );
xor ( n62641 , n62640 , n49228 );
and ( n62642 , n62641 , n48845 );
or ( n62643 , n62639 , n62642 );
and ( n62644 , n62643 , n49054 );
or ( n62645 , n62635 , n62644 );
and ( n62646 , n62645 , n33178 );
and ( n62647 , n49200 , n49275 );
or ( n62648 , n62596 , n62601 , n62606 , n62611 , n62616 , n62621 , n62626 , n62633 , n62646 , n62647 );
and ( n62649 , n62648 , n33208 );
and ( n62650 , n33000 , n35056 );
and ( n62651 , n48607 , n49286 );
or ( n62652 , C0 , n62649 , n62650 , n62651 );
buf ( n62653 , n62652 );
buf ( n62654 , n62653 );
buf ( n62655 , n30987 );
buf ( n62656 , n31655 );
buf ( n62657 , n31655 );
buf ( n62658 , n31655 );
buf ( n62659 , n30987 );
not ( n62660 , n46356 );
and ( n62661 , n62660 , n31017 );
and ( n62662 , n46386 , n46356 );
or ( n62663 , n62661 , n62662 );
and ( n62664 , n62663 , n31649 );
not ( n62665 , n52614 );
not ( n62666 , n44702 );
and ( n62667 , n62666 , n31017 );
buf ( n62668 , n62667 );
and ( n62669 , n62665 , n62668 );
buf ( n62670 , n62669 );
and ( n62671 , n62670 , n31647 );
and ( n62672 , n46534 , n31643 );
not ( n62673 , n31452 );
and ( n62674 , n62673 , n46534 );
and ( n62675 , n46528 , n46519 );
xor ( n62676 , n46539 , n62675 );
not ( n62677 , n62676 );
buf ( n62678 , n62677 );
not ( n62679 , n62678 );
and ( n62680 , n62679 , n31452 );
or ( n62681 , n62674 , n62680 );
and ( n62682 , n62681 , n31638 );
and ( n62683 , n31017 , n52626 );
or ( n62684 , C0 , n62664 , n62671 , n62672 , n62682 , n62683 );
buf ( n62685 , n62684 );
buf ( n62686 , n62685 );
buf ( n62687 , n30987 );
buf ( n62688 , n31655 );
not ( n62689 , n31728 );
and ( n62690 , n62689 , n32462 );
xor ( n62691 , n31930 , n31963 );
xor ( n62692 , n62691 , n32075 );
and ( n62693 , n62692 , n31728 );
or ( n62694 , n62690 , n62693 );
and ( n62695 , n62694 , n32253 );
not ( n62696 , n32283 );
and ( n62697 , n62696 , n32462 );
not ( n62698 , n31823 );
xor ( n62699 , n32302 , n31963 );
xor ( n62700 , n62699 , n32314 );
and ( n62701 , n62698 , n62700 );
xor ( n62702 , n32356 , n32358 );
xor ( n62703 , n62702 , n32377 );
and ( n62704 , n62703 , n31823 );
or ( n62705 , n62701 , n62704 );
and ( n62706 , n62705 , n32283 );
or ( n62707 , n62697 , n62706 );
and ( n62708 , n62707 , n32398 );
and ( n62709 , n32462 , n32436 );
or ( n62710 , n62695 , n62708 , n62709 );
and ( n62711 , n62710 , n32456 );
and ( n62712 , n49701 , n32473 );
not ( n62713 , n32475 );
and ( n62714 , n62713 , n49701 );
xor ( n62715 , n32462 , n32463 );
and ( n62716 , n62715 , n32475 );
or ( n62717 , n62714 , n62716 );
and ( n62718 , n62717 , n32486 );
and ( n62719 , n37583 , n32489 );
and ( n62720 , n32462 , n32501 );
or ( n62721 , C0 , n62711 , n62712 , n62718 , n62719 , n62720 );
buf ( n62722 , n62721 );
buf ( n62723 , n62722 );
buf ( n62724 , n30987 );
not ( n62725 , n40163 );
and ( n62726 , n62725 , n31945 );
not ( n62727 , n52120 );
and ( n62728 , n62727 , n31945 );
and ( n62729 , n32183 , n52120 );
or ( n62730 , n62728 , n62729 );
and ( n62731 , n62730 , n40163 );
or ( n62732 , n62726 , n62731 );
and ( n62733 , n62732 , n32498 );
not ( n62734 , n52128 );
not ( n62735 , n52120 );
and ( n62736 , n62735 , n31945 );
and ( n62737 , n45178 , n52120 );
or ( n62738 , n62736 , n62737 );
and ( n62739 , n62734 , n62738 );
and ( n62740 , n45178 , n52128 );
or ( n62741 , n62739 , n62740 );
and ( n62742 , n62741 , n32473 );
not ( n62743 , n32475 );
not ( n62744 , n52128 );
not ( n62745 , n52120 );
and ( n62746 , n62745 , n31945 );
and ( n62747 , n45178 , n52120 );
or ( n62748 , n62746 , n62747 );
and ( n62749 , n62744 , n62748 );
and ( n62750 , n45178 , n52128 );
or ( n62751 , n62749 , n62750 );
and ( n62752 , n62743 , n62751 );
not ( n62753 , n52148 );
not ( n62754 , n52150 );
and ( n62755 , n62754 , n62751 );
and ( n62756 , n45206 , n52150 );
or ( n62757 , n62755 , n62756 );
and ( n62758 , n62753 , n62757 );
and ( n62759 , n45214 , n52148 );
or ( n62760 , n62758 , n62759 );
and ( n62761 , n62760 , n32475 );
or ( n62762 , n62752 , n62761 );
and ( n62763 , n62762 , n32486 );
and ( n62764 , n31945 , n41278 );
or ( n62765 , C0 , n62733 , n62742 , n62763 , n62764 );
buf ( n62766 , n62765 );
buf ( n62767 , n62766 );
buf ( n62768 , n31655 );
not ( n62769 , n54795 );
not ( n62770 , n54797 );
not ( n62771 , n54800 );
and ( n62772 , n62770 , n62771 );
buf ( n62773 , n54797 );
or ( n62774 , n62772 , n62773 );
and ( n62775 , n62769 , n62774 );
buf ( n62776 , n62775 );
and ( n62777 , n62776 , n37505 );
not ( n62778 , n54815 );
and ( n62779 , n62778 , n37503 );
not ( n62780 , n54824 );
not ( n62781 , n54827 );
and ( n62782 , n62781 , n48294 );
buf ( n62783 , n54827 );
or ( n62784 , n62782 , n62783 );
and ( n62785 , n62780 , n62784 );
buf ( n62786 , n62785 );
and ( n62787 , n62786 , n37501 );
not ( n62788 , n54800 );
not ( n62789 , n54838 );
not ( n62790 , n54842 );
not ( n62791 , n54845 );
and ( n62792 , n62790 , n62791 );
buf ( n62793 , n54842 );
or ( n62794 , n62792 , n62793 );
and ( n62795 , n62789 , n62794 );
and ( n62796 , n31440 , n54838 );
or ( n62797 , n62795 , n62796 );
and ( n62798 , n62788 , n62797 );
buf ( n62799 , n62798 );
and ( n62800 , n62799 , n37499 );
buf ( n62801 , n37494 );
not ( n62802 , n54792 );
and ( n62803 , n62802 , n37496 );
buf ( n62804 , n37497 );
or ( n62805 , n62777 , C0 , n62779 , n62787 , n62800 , n62801 , n62803 , n62804 );
buf ( n62806 , n62805 );
buf ( n62807 , n62806 );
buf ( n62808 , n30987 );
buf ( n62809 , n30987 );
buf ( n62810 , n31655 );
not ( n62811 , n40163 );
and ( n62812 , n62811 , n32031 );
not ( n62813 , n40166 );
and ( n62814 , n62813 , n32031 );
and ( n62815 , n32147 , n40166 );
or ( n62816 , n62814 , n62815 );
and ( n62817 , n62816 , n40163 );
or ( n62818 , n62812 , n62817 );
and ( n62819 , n62818 , n32498 );
not ( n62820 , n40195 );
not ( n62821 , n40166 );
and ( n62822 , n62821 , n32031 );
and ( n62823 , n49314 , n40166 );
or ( n62824 , n62822 , n62823 );
and ( n62825 , n62820 , n62824 );
and ( n62826 , n49314 , n40195 );
or ( n62827 , n62825 , n62826 );
and ( n62828 , n62827 , n32473 );
not ( n62829 , n32475 );
not ( n62830 , n40195 );
not ( n62831 , n40166 );
and ( n62832 , n62831 , n32031 );
and ( n62833 , n49314 , n40166 );
or ( n62834 , n62832 , n62833 );
and ( n62835 , n62830 , n62834 );
and ( n62836 , n49314 , n40195 );
or ( n62837 , n62835 , n62836 );
and ( n62838 , n62829 , n62837 );
not ( n62839 , n40446 );
not ( n62840 , n40448 );
and ( n62841 , n62840 , n62837 );
and ( n62842 , n49340 , n40448 );
or ( n62843 , n62841 , n62842 );
and ( n62844 , n62839 , n62843 );
and ( n62845 , n49348 , n40446 );
or ( n62846 , n62844 , n62845 );
and ( n62847 , n62846 , n32475 );
or ( n62848 , n62838 , n62847 );
and ( n62849 , n62848 , n32486 );
and ( n62850 , n32031 , n41278 );
or ( n62851 , C0 , n62819 , n62828 , n62849 , n62850 );
buf ( n62852 , n62851 );
buf ( n62853 , n62852 );
and ( n62854 , n35431 , n59497 );
and ( n62855 , n35429 , n62854 );
and ( n62856 , n35427 , n62855 );
and ( n62857 , n35425 , n62856 );
and ( n62858 , n35423 , n62857 );
xor ( n62859 , n31501 , n62858 );
and ( n62860 , n62859 , n31550 );
not ( n62861 , n39979 );
and ( n62862 , n62861 , n31501 );
buf ( n62863 , n62862 );
and ( n62864 , n62863 , n31538 );
and ( n62865 , n31501 , n40143 );
or ( n62866 , n62860 , n62864 , n62865 );
and ( n62867 , n62866 , n31557 );
and ( n62868 , n31501 , n40154 );
or ( n62869 , C0 , n62867 , n62868 );
buf ( n62870 , n62869 );
buf ( n62871 , n62870 );
buf ( n62872 , n40202 );
buf ( n62873 , n30987 );
buf ( n62874 , n31655 );
buf ( n62875 , n31655 );
buf ( n62876 , n30987 );
buf ( n62877 , n30987 );
and ( n62878 , n49065 , n48639 );
not ( n62879 , n48642 );
and ( n62880 , n62879 , n48590 );
and ( n62881 , n49065 , n48642 );
or ( n62882 , n62880 , n62881 );
and ( n62883 , n62882 , n32890 );
not ( n62884 , n48648 );
and ( n62885 , n62884 , n48590 );
and ( n62886 , n49065 , n48648 );
or ( n62887 , n62885 , n62886 );
and ( n62888 , n62887 , n32924 );
not ( n62889 , n48654 );
and ( n62890 , n62889 , n48590 );
and ( n62891 , n49065 , n48654 );
or ( n62892 , n62890 , n62891 );
and ( n62893 , n62892 , n33038 );
not ( n62894 , n48660 );
and ( n62895 , n62894 , n48590 );
and ( n62896 , n49065 , n48660 );
or ( n62897 , n62895 , n62896 );
and ( n62898 , n62897 , n33172 );
not ( n62899 , n41576 );
and ( n62900 , n62899 , n48590 );
and ( n62901 , n48775 , n41576 );
or ( n62902 , n62900 , n62901 );
and ( n62903 , n62902 , n33189 );
not ( n62904 , n48730 );
and ( n62905 , n62904 , n48590 );
and ( n62906 , n48775 , n48730 );
or ( n62907 , n62905 , n62906 );
and ( n62908 , n62907 , n33187 );
not ( n62909 , n48765 );
and ( n62910 , n62909 , n48590 );
xor ( n62911 , n48775 , n49013 );
and ( n62912 , n62911 , n48765 );
or ( n62913 , n62910 , n62912 );
and ( n62914 , n62913 , n33180 );
not ( n62915 , n49054 );
and ( n62916 , n62915 , n48590 );
not ( n62917 , n48845 );
xor ( n62918 , n49065 , n49127 );
and ( n62919 , n62917 , n62918 );
xnor ( n62920 , n49174 , n49253 );
and ( n62921 , n62920 , n48845 );
or ( n62922 , n62919 , n62921 );
and ( n62923 , n62922 , n49054 );
or ( n62924 , n62916 , n62923 );
and ( n62925 , n62924 , n33178 );
and ( n62926 , n49174 , n49275 );
or ( n62927 , n62878 , n62883 , n62888 , n62893 , n62898 , n62903 , n62908 , n62914 , n62925 , n62926 );
and ( n62928 , n62927 , n33208 );
and ( n62929 , n32983 , n35056 );
and ( n62930 , n48590 , n49286 );
or ( n62931 , C0 , n62928 , n62929 , n62930 );
buf ( n62932 , n62931 );
buf ( n62933 , n62932 );
buf ( n62934 , n30987 );
and ( n62935 , n31577 , n31007 );
not ( n62936 , n31077 );
and ( n62937 , n62936 , n34001 );
buf ( n62938 , n62937 );
and ( n62939 , n62938 , n31373 );
not ( n62940 , n31402 );
and ( n62941 , n62940 , n34001 );
buf ( n62942 , n62941 );
and ( n62943 , n62942 , n31408 );
not ( n62944 , n31437 );
and ( n62945 , n62944 , n34001 );
not ( n62946 , n31455 );
and ( n62947 , n62946 , n34042 );
xor ( n62948 , n34001 , n34022 );
and ( n62949 , n62948 , n31455 );
or ( n62950 , n62947 , n62949 );
and ( n62951 , n62950 , n31437 );
or ( n62952 , n62945 , n62951 );
and ( n62953 , n62952 , n31468 );
not ( n62954 , n31497 );
and ( n62955 , n62954 , n34001 );
not ( n62956 , n31454 );
not ( n62957 , n31501 );
and ( n62958 , n62957 , n34042 );
xor ( n62959 , n34043 , n34074 );
and ( n62960 , n62959 , n31501 );
or ( n62961 , n62958 , n62960 );
and ( n62962 , n62956 , n62961 );
and ( n62963 , n62948 , n31454 );
or ( n62964 , n62962 , n62963 );
and ( n62965 , n62964 , n31497 );
or ( n62966 , n62955 , n62965 );
and ( n62967 , n62966 , n31521 );
and ( n62968 , n34001 , n31553 );
or ( n62969 , n62939 , n62943 , n62953 , n62967 , n62968 );
and ( n62970 , n62969 , n31557 );
not ( n62971 , n31452 );
not ( n62972 , n31619 );
and ( n62973 , n62972 , n34099 );
xor ( n62974 , n34100 , n34131 );
and ( n62975 , n62974 , n31619 );
or ( n62976 , n62973 , n62975 );
and ( n62977 , n62971 , n62976 );
and ( n62978 , n34001 , n31452 );
or ( n62979 , n62977 , n62978 );
and ( n62980 , n62979 , n31638 );
buf ( n62981 , n33973 );
and ( n62982 , n34001 , n31650 );
or ( n62983 , C0 , n62935 , n62970 , n62980 , n62981 , n62982 );
buf ( n62984 , n62983 );
buf ( n62985 , n62984 );
buf ( n62986 , n31655 );
buf ( n62987 , n31655 );
not ( n62988 , n33419 );
and ( n62989 , n62988 , n31567 );
xor ( n62990 , n42385 , n42390 );
and ( n62991 , n62990 , n33419 );
or ( n62992 , n62989 , n62991 );
and ( n62993 , n62992 , n31529 );
not ( n62994 , n33734 );
and ( n62995 , n62994 , n31567 );
not ( n62996 , n33533 );
xor ( n62997 , n42404 , n42409 );
and ( n62998 , n62996 , n62997 );
xnor ( n62999 , n42418 , n42423 );
and ( n63000 , n62999 , n33533 );
or ( n63001 , n62998 , n63000 );
and ( n63002 , n63001 , n33734 );
or ( n63003 , n62995 , n63002 );
and ( n63004 , n63003 , n31527 );
and ( n63005 , n31567 , n33942 );
or ( n63006 , n62993 , n63004 , n63005 );
and ( n63007 , n63006 , n31557 );
and ( n63008 , n35490 , n31643 );
not ( n63009 , n31452 );
and ( n63010 , n63009 , n35490 );
xor ( n63011 , n31567 , n42439 );
and ( n63012 , n63011 , n31452 );
or ( n63013 , n63010 , n63012 );
and ( n63014 , n63013 , n31638 );
and ( n63015 , n35393 , n33973 );
and ( n63016 , n31567 , n33978 );
or ( n63017 , C0 , n63007 , n63008 , n63014 , n63015 , n63016 );
buf ( n63018 , n63017 );
buf ( n63019 , n63018 );
buf ( n63020 , n30987 );
buf ( n63021 , n30987 );
not ( n63022 , n46356 );
and ( n63023 , n63022 , n31240 );
and ( n63024 , n31025 , n31021 , n31017 , n31013 , n46361 );
not ( n63025 , n63024 );
and ( n63026 , n63025 , n31240 );
and ( n63027 , n31272 , n63024 );
or ( n63028 , n63026 , n63027 );
and ( n63029 , n63028 , n46356 );
or ( n63030 , n63023 , n63029 );
and ( n63031 , n63030 , n31649 );
and ( n63032 , n46373 , n46379 , n46386 , n46392 , C1 );
not ( n63033 , n63032 );
not ( n63034 , n63024 );
and ( n63035 , n63034 , n31240 );
and ( n63036 , n49443 , n63024 );
or ( n63037 , n63035 , n63036 );
and ( n63038 , n63033 , n63037 );
and ( n63039 , n49443 , n63032 );
or ( n63040 , n63038 , n63039 );
and ( n63041 , n63040 , n31643 );
not ( n63042 , n31452 );
not ( n63043 , n63032 );
not ( n63044 , n63024 );
and ( n63045 , n63044 , n31240 );
and ( n63046 , n49443 , n63024 );
or ( n63047 , n63045 , n63046 );
and ( n63048 , n63043 , n63047 );
and ( n63049 , n49443 , n63032 );
or ( n63050 , n63048 , n63049 );
and ( n63051 , n63042 , n63050 );
and ( n63052 , n46519 , n46528 , n46539 , n46549 , C1 );
not ( n63053 , n63052 );
and ( n63054 , n46515 , n46524 , n46534 , n46544 , C1 );
not ( n63055 , n63054 );
and ( n63056 , n63055 , n63050 );
and ( n63057 , n49469 , n63054 );
or ( n63058 , n63056 , n63057 );
and ( n63059 , n63053 , n63058 );
and ( n63060 , n49477 , n63052 );
or ( n63061 , n63059 , n63060 );
and ( n63062 , n63061 , n31452 );
or ( n63063 , n63051 , n63062 );
and ( n63064 , n63063 , n31638 );
and ( n63065 , n31240 , n47277 );
or ( n63066 , C0 , n63031 , n63041 , n63064 , n63065 );
buf ( n63067 , n63066 );
buf ( n63068 , n63067 );
not ( n63069 , n35278 );
buf ( n63070 , RI15b5f130_1109);
and ( n63071 , n63069 , n63070 );
not ( n63072 , n46290 );
and ( n63073 , n63072 , n46117 );
xor ( n63074 , n46304 , n46308 );
and ( n63075 , n63074 , n46290 );
or ( n63076 , n63073 , n63075 );
and ( n63077 , n63076 , n35278 );
or ( n63078 , n63071 , n63077 );
and ( n63079 , n63078 , n32417 );
not ( n63080 , n47912 );
and ( n63081 , n63080 , n63070 );
not ( n63082 , n48101 );
and ( n63083 , n63082 , n47941 );
xor ( n63084 , n48109 , n48113 );
and ( n63085 , n63084 , n48101 );
or ( n63086 , n63083 , n63085 );
and ( n63087 , n63086 , n47912 );
or ( n63088 , n63081 , n63087 );
and ( n63089 , n63088 , n32415 );
and ( n63090 , n63070 , n48133 );
or ( n63091 , n63079 , n63089 , n63090 );
and ( n63092 , n63091 , n32456 );
and ( n63093 , n63070 , n47409 );
or ( n63094 , C0 , n63092 , n63093 );
buf ( n63095 , n63094 );
buf ( n63096 , n63095 );
buf ( n63097 , n31655 );
buf ( n63098 , n31655 );
buf ( n63099 , n31655 );
not ( n63100 , n35211 );
and ( n63101 , n56812 , n63100 );
and ( n63102 , n63101 , n32421 );
not ( n63103 , n35245 );
and ( n63104 , n56812 , n63103 );
and ( n63105 , n63104 , n32419 );
not ( n63106 , n35278 );
and ( n63107 , n56812 , n63106 );
and ( n63108 , n63107 , n32417 );
not ( n63109 , n35331 );
and ( n63110 , n56812 , n63109 );
and ( n63111 , n63110 , n32415 );
and ( n63112 , n56812 , n35354 );
or ( n63113 , n63102 , n63105 , n63108 , n63111 , n63112 );
and ( n63114 , n63113 , n32456 );
buf ( n63115 , n32491 );
or ( n63116 , n32489 , n32486 );
or ( n63117 , n63116 , n32492 );
or ( n63118 , n63117 , n32473 );
or ( n63119 , n63118 , n32494 );
or ( n63120 , n63119 , n32496 );
or ( n63121 , n63120 , n32498 );
or ( n63122 , n63121 , n32500 );
and ( n63123 , n56812 , n63122 );
or ( n63124 , C0 , n63114 , n63115 , n63123 );
buf ( n63125 , n63124 );
buf ( n63126 , n63125 );
not ( n63127 , n46356 );
and ( n63128 , n63127 , n31185 );
not ( n63129 , n52734 );
and ( n63130 , n63129 , n31185 );
and ( n63131 , n31205 , n52734 );
or ( n63132 , n63130 , n63131 );
and ( n63133 , n63132 , n46356 );
or ( n63134 , n63128 , n63133 );
and ( n63135 , n63134 , n31649 );
not ( n63136 , n52742 );
not ( n63137 , n52734 );
and ( n63138 , n63137 , n31185 );
and ( n63139 , n50125 , n52734 );
or ( n63140 , n63138 , n63139 );
and ( n63141 , n63136 , n63140 );
and ( n63142 , n50125 , n52742 );
or ( n63143 , n63141 , n63142 );
and ( n63144 , n63143 , n31643 );
not ( n63145 , n31452 );
not ( n63146 , n52742 );
not ( n63147 , n52734 );
and ( n63148 , n63147 , n31185 );
and ( n63149 , n50125 , n52734 );
or ( n63150 , n63148 , n63149 );
and ( n63151 , n63146 , n63150 );
and ( n63152 , n50125 , n52742 );
or ( n63153 , n63151 , n63152 );
and ( n63154 , n63145 , n63153 );
not ( n63155 , n52762 );
not ( n63156 , n52764 );
and ( n63157 , n63156 , n63153 );
and ( n63158 , n50151 , n52764 );
or ( n63159 , n63157 , n63158 );
and ( n63160 , n63155 , n63159 );
and ( n63161 , n50159 , n52762 );
or ( n63162 , n63160 , n63161 );
and ( n63163 , n63162 , n31452 );
or ( n63164 , n63154 , n63163 );
and ( n63165 , n63164 , n31638 );
and ( n63166 , n31185 , n47277 );
or ( n63167 , C0 , n63135 , n63144 , n63165 , n63166 );
buf ( n63168 , n63167 );
buf ( n63169 , n63168 );
buf ( n63170 , n30987 );
not ( n63171 , n46356 );
and ( n63172 , n63171 , n31346 );
not ( n63173 , n46362 );
and ( n63174 , n63173 , n31346 );
and ( n63175 , n31372 , n46362 );
or ( n63176 , n63174 , n63175 );
and ( n63177 , n63176 , n46356 );
or ( n63178 , n63172 , n63177 );
and ( n63179 , n63178 , n31649 );
not ( n63180 , n46393 );
not ( n63181 , n46362 );
and ( n63182 , n63181 , n31346 );
and ( n63183 , n47849 , n46362 );
or ( n63184 , n63182 , n63183 );
and ( n63185 , n63180 , n63184 );
and ( n63186 , n47849 , n46393 );
or ( n63187 , n63185 , n63186 );
and ( n63188 , n63187 , n31643 );
not ( n63189 , n31452 );
not ( n63190 , n46393 );
not ( n63191 , n46362 );
and ( n63192 , n63191 , n31346 );
and ( n63193 , n47849 , n46362 );
or ( n63194 , n63192 , n63193 );
and ( n63195 , n63190 , n63194 );
and ( n63196 , n47849 , n46393 );
or ( n63197 , n63195 , n63196 );
and ( n63198 , n63189 , n63197 );
not ( n63199 , n46550 );
not ( n63200 , n46554 );
and ( n63201 , n63200 , n63197 );
and ( n63202 , n47877 , n46554 );
or ( n63203 , n63201 , n63202 );
and ( n63204 , n63199 , n63203 );
and ( n63205 , n47887 , n46550 );
or ( n63206 , n63204 , n63205 );
and ( n63207 , n63206 , n31452 );
or ( n63208 , n63198 , n63207 );
and ( n63209 , n63208 , n31638 );
and ( n63210 , n31346 , n47277 );
or ( n63211 , C0 , n63179 , n63188 , n63209 , n63210 );
buf ( n63212 , n63211 );
buf ( n63213 , n63212 );
buf ( n63214 , n31655 );
buf ( n63215 , n31655 );
and ( n63216 , n47900 , n32494 );
not ( n63217 , n46083 );
buf ( n63218 , RI15b5fb08_1130);
and ( n63219 , n63217 , n63218 );
and ( n63220 , n47906 , n46083 );
or ( n63221 , n63219 , n63220 );
and ( n63222 , n63221 , n32421 );
not ( n63223 , n46326 );
and ( n63224 , n63223 , n63218 );
and ( n63225 , n47906 , n46326 );
or ( n63226 , n63224 , n63225 );
and ( n63227 , n63226 , n32417 );
and ( n63228 , n63218 , n46340 );
or ( n63229 , n63222 , n63227 , n63228 );
and ( n63230 , n63229 , n32456 );
and ( n63231 , n63218 , n46349 );
or ( n63232 , C0 , n63216 , n63230 , n63231 );
buf ( n63233 , n63232 );
buf ( n63234 , n63233 );
buf ( n63235 , n30987 );
and ( n63236 , n33761 , n48455 );
not ( n63237 , n48457 );
and ( n63238 , n63237 , n33426 );
and ( n63239 , n33761 , n48457 );
or ( n63240 , n63238 , n63239 );
and ( n63241 , n63240 , n31373 );
not ( n63242 , n44807 );
and ( n63243 , n63242 , n33426 );
and ( n63244 , n33761 , n44807 );
or ( n63245 , n63243 , n63244 );
and ( n63246 , n63245 , n31408 );
not ( n63247 , n48468 );
and ( n63248 , n63247 , n33426 );
and ( n63249 , n33761 , n48468 );
or ( n63250 , n63248 , n63249 );
and ( n63251 , n63250 , n31468 );
not ( n63252 , n44817 );
and ( n63253 , n63252 , n33426 );
and ( n63254 , n33761 , n44817 );
or ( n63255 , n63253 , n63254 );
and ( n63256 , n63255 , n31521 );
not ( n63257 , n39979 );
and ( n63258 , n63257 , n33426 );
and ( n63259 , n33468 , n39979 );
or ( n63260 , n63258 , n63259 );
and ( n63261 , n63260 , n31538 );
not ( n63262 , n45059 );
and ( n63263 , n63262 , n33426 );
and ( n63264 , n33468 , n45059 );
or ( n63265 , n63263 , n63264 );
and ( n63266 , n63265 , n31536 );
not ( n63267 , n33419 );
and ( n63268 , n63267 , n33426 );
xor ( n63269 , n33468 , n33697 );
and ( n63270 , n63269 , n33419 );
or ( n63271 , n63268 , n63270 );
and ( n63272 , n63271 , n31529 );
not ( n63273 , n33734 );
and ( n63274 , n63273 , n33426 );
not ( n63275 , n33533 );
xor ( n63276 , n33761 , n33815 );
and ( n63277 , n63275 , n63276 );
xnor ( n63278 , n33846 , n33917 );
and ( n63279 , n63278 , n33533 );
or ( n63280 , n63277 , n63279 );
and ( n63281 , n63280 , n33734 );
or ( n63282 , n63274 , n63281 );
and ( n63283 , n63282 , n31527 );
and ( n63284 , n33846 , n48513 );
or ( n63285 , n63236 , n63241 , n63246 , n63251 , n63256 , n63261 , n63266 , n63272 , n63283 , n63284 );
and ( n63286 , n63285 , n31557 );
and ( n63287 , n33986 , n33973 );
and ( n63288 , n33426 , n48524 );
or ( n63289 , C0 , n63286 , n63287 , n63288 );
buf ( n63290 , n63289 );
buf ( n63291 , n63290 );
buf ( n63292 , n31655 );
buf ( n63293 , RI15b607b0_1157);
not ( n63294 , n63293 );
and ( n63295 , n63294 , n48531 );
and ( n63296 , n50821 , n39359 );
or ( n63297 , n63295 , n63296 );
buf ( n63298 , n63297 );
buf ( n63299 , n63298 );
buf ( n63300 , n30987 );
buf ( n63301 , n31655 );
not ( n63302 , n46356 );
and ( n63303 , n63302 , n31224 );
not ( n63304 , n50109 );
and ( n63305 , n63304 , n31224 );
and ( n63306 , n31238 , n50109 );
or ( n63307 , n63305 , n63306 );
and ( n63308 , n63307 , n46356 );
or ( n63309 , n63303 , n63308 );
and ( n63310 , n63309 , n31649 );
not ( n63311 , n50117 );
not ( n63312 , n50109 );
and ( n63313 , n63312 , n31224 );
and ( n63314 , n49901 , n50109 );
or ( n63315 , n63313 , n63314 );
and ( n63316 , n63311 , n63315 );
and ( n63317 , n49901 , n50117 );
or ( n63318 , n63316 , n63317 );
and ( n63319 , n63318 , n31643 );
not ( n63320 , n31452 );
not ( n63321 , n50117 );
not ( n63322 , n50109 );
and ( n63323 , n63322 , n31224 );
and ( n63324 , n49901 , n50109 );
or ( n63325 , n63323 , n63324 );
and ( n63326 , n63321 , n63325 );
and ( n63327 , n49901 , n50117 );
or ( n63328 , n63326 , n63327 );
and ( n63329 , n63320 , n63328 );
not ( n63330 , n50142 );
not ( n63331 , n50144 );
and ( n63332 , n63331 , n63328 );
and ( n63333 , n49925 , n50144 );
or ( n63334 , n63332 , n63333 );
and ( n63335 , n63330 , n63334 );
and ( n63336 , n49933 , n50142 );
or ( n63337 , n63335 , n63336 );
and ( n63338 , n63337 , n31452 );
or ( n63339 , n63329 , n63338 );
and ( n63340 , n63339 , n31638 );
and ( n63341 , n31224 , n47277 );
or ( n63342 , C0 , n63310 , n63319 , n63340 , n63341 );
buf ( n63343 , n63342 );
buf ( n63344 , n63343 );
buf ( n63345 , n30987 );
buf ( n63346 , n31655 );
xor ( n63347 , n46250 , n49998 );
and ( n63348 , n63347 , n32431 );
not ( n63349 , n50002 );
and ( n63350 , n63349 , n46250 );
and ( n63351 , n40479 , n50002 );
or ( n63352 , n63350 , n63351 );
and ( n63353 , n63352 , n32419 );
not ( n63354 , n50008 );
and ( n63355 , n63354 , n46250 );
not ( n63356 , n47910 );
and ( n63357 , n63356 , n46081 );
not ( n63358 , n48101 );
and ( n63359 , n63358 , n48073 );
xor ( n63360 , n50017 , n50028 );
and ( n63361 , n63360 , n48101 );
or ( n63362 , n63359 , n63361 );
and ( n63363 , n63362 , n47910 );
or ( n63364 , n63357 , n63363 );
and ( n63365 , n63364 , n50008 );
or ( n63366 , n63355 , n63365 );
and ( n63367 , n63366 , n32415 );
not ( n63368 , n50067 );
and ( n63369 , n63368 , n46250 );
and ( n63370 , n31861 , n47357 );
and ( n63371 , n31863 , n47359 );
and ( n63372 , n31865 , n47361 );
and ( n63373 , n31867 , n47363 );
and ( n63374 , n31869 , n47365 );
and ( n63375 , n31871 , n47367 );
and ( n63376 , n31873 , n47369 );
and ( n63377 , n31875 , n47371 );
and ( n63378 , n31877 , n47373 );
and ( n63379 , n31879 , n47375 );
and ( n63380 , n31881 , n47377 );
and ( n63381 , n31883 , n47379 );
and ( n63382 , n31885 , n47381 );
and ( n63383 , n31887 , n47383 );
and ( n63384 , n31889 , n47385 );
and ( n63385 , n31891 , n47387 );
or ( n63386 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 );
and ( n63387 , n63386 , n50067 );
or ( n63388 , n63369 , n63387 );
and ( n63389 , n63388 , n32411 );
and ( n63390 , n46250 , n50098 );
or ( n63391 , n63348 , n63353 , n63367 , n63389 , n63390 );
and ( n63392 , n63391 , n32456 );
and ( n63393 , n46250 , n47409 );
or ( n63394 , C0 , n63392 , n63393 );
buf ( n63395 , n63394 );
buf ( n63396 , n63395 );
not ( n63397 , n38443 );
and ( n63398 , n63397 , n38014 );
xor ( n63399 , n53481 , n53488 );
and ( n63400 , n63399 , n38443 );
or ( n63401 , n63398 , n63400 );
and ( n63402 , n63401 , n38450 );
not ( n63403 , n39339 );
and ( n63404 , n63403 , n38914 );
xor ( n63405 , n53537 , n53544 );
and ( n63406 , n63405 , n39339 );
or ( n63407 , n63404 , n63406 );
and ( n63408 , n63407 , n39346 );
and ( n63409 , n40203 , n39359 );
or ( n63410 , n63402 , n63408 , n63409 );
buf ( n63411 , n63410 );
buf ( n63412 , n63411 );
buf ( n63413 , RI15b544b0_741);
and ( n63414 , n63413 , n58921 );
and ( n63415 , n41528 , n37506 );
or ( n63416 , n63414 , n63415 );
buf ( n63417 , n63416 );
buf ( n63418 , n63417 );
buf ( n63419 , n30987 );
buf ( n63420 , n31655 );
buf ( n63421 , n31655 );
and ( n63422 , n47656 , n50275 );
not ( n63423 , n50278 );
and ( n63424 , n63423 , n47569 );
and ( n63425 , n47656 , n50278 );
or ( n63426 , n63424 , n63425 );
and ( n63427 , n63426 , n32421 );
not ( n63428 , n50002 );
and ( n63429 , n63428 , n47569 );
and ( n63430 , n47656 , n50002 );
or ( n63431 , n63429 , n63430 );
and ( n63432 , n63431 , n32419 );
not ( n63433 , n50289 );
and ( n63434 , n63433 , n47569 );
and ( n63435 , n47656 , n50289 );
or ( n63436 , n63434 , n63435 );
and ( n63437 , n63436 , n32417 );
not ( n63438 , n50008 );
and ( n63439 , n63438 , n47569 );
and ( n63440 , n47656 , n50008 );
or ( n63441 , n63439 , n63440 );
and ( n63442 , n63441 , n32415 );
not ( n63443 , n47331 );
and ( n63444 , n63443 , n47569 );
and ( n63445 , n47601 , n47331 );
or ( n63446 , n63444 , n63445 );
and ( n63447 , n63446 , n32413 );
not ( n63448 , n50067 );
and ( n63449 , n63448 , n47569 );
and ( n63450 , n47601 , n50067 );
or ( n63451 , n63449 , n63450 );
and ( n63452 , n63451 , n32411 );
not ( n63453 , n31728 );
and ( n63454 , n63453 , n47569 );
xor ( n63455 , n47601 , n47628 );
and ( n63456 , n63455 , n31728 );
or ( n63457 , n63454 , n63456 );
and ( n63458 , n63457 , n32253 );
not ( n63459 , n32283 );
and ( n63460 , n63459 , n47569 );
not ( n63461 , n31823 );
xor ( n63462 , n47656 , n47683 );
and ( n63463 , n63461 , n63462 );
xnor ( n63464 , n47706 , n47733 );
and ( n63465 , n63464 , n31823 );
or ( n63466 , n63463 , n63465 );
and ( n63467 , n63466 , n32283 );
or ( n63468 , n63460 , n63467 );
and ( n63469 , n63468 , n32398 );
and ( n63470 , n47706 , n50334 );
or ( n63471 , n63422 , n63427 , n63432 , n63437 , n63442 , n63447 , n63452 , n63458 , n63469 , n63470 );
and ( n63472 , n63471 , n32456 );
and ( n63473 , n37545 , n32489 );
and ( n63474 , n47569 , n50345 );
or ( n63475 , C0 , n63472 , n63473 , n63474 );
buf ( n63476 , n63475 );
buf ( n63477 , n63476 );
buf ( n63478 , n30987 );
not ( n63479 , n36587 );
and ( n63480 , n63479 , n36498 );
xor ( n63481 , n61942 , n61943 );
and ( n63482 , n63481 , n36587 );
or ( n63483 , n63480 , n63482 );
and ( n63484 , n63483 , n36596 );
not ( n63485 , n37485 );
and ( n63486 , n63485 , n37400 );
xor ( n63487 , n61958 , n61959 );
and ( n63488 , n63487 , n37485 );
or ( n63489 , n63486 , n63488 );
and ( n63490 , n63489 , n37494 );
and ( n63491 , n41863 , n37506 );
or ( n63492 , n63484 , n63490 , n63491 );
buf ( n63493 , n63492 );
buf ( n63494 , n63493 );
buf ( n63495 , n30987 );
buf ( n63496 , n31655 );
buf ( n63497 , n31655 );
buf ( n63498 , n30987 );
and ( n63499 , n49058 , n48639 );
not ( n63500 , n48642 );
and ( n63501 , n63500 , n48583 );
and ( n63502 , n49058 , n48642 );
or ( n63503 , n63501 , n63502 );
and ( n63504 , n63503 , n32890 );
not ( n63505 , n48648 );
and ( n63506 , n63505 , n48583 );
and ( n63507 , n49058 , n48648 );
or ( n63508 , n63506 , n63507 );
and ( n63509 , n63508 , n32924 );
not ( n63510 , n48654 );
and ( n63511 , n63510 , n48583 );
and ( n63512 , n49058 , n48654 );
or ( n63513 , n63511 , n63512 );
and ( n63514 , n63513 , n33038 );
not ( n63515 , n48660 );
and ( n63516 , n63515 , n48583 );
and ( n63517 , n49058 , n48660 );
or ( n63518 , n63516 , n63517 );
and ( n63519 , n63518 , n33172 );
not ( n63520 , n41576 );
and ( n63521 , n63520 , n48583 );
and ( n63522 , n48768 , n41576 );
or ( n63523 , n63521 , n63522 );
and ( n63524 , n63523 , n33189 );
not ( n63525 , n48730 );
and ( n63526 , n63525 , n48583 );
and ( n63527 , n48768 , n48730 );
or ( n63528 , n63526 , n63527 );
and ( n63529 , n63528 , n33187 );
not ( n63530 , n48765 );
and ( n63531 , n63530 , n48583 );
xor ( n63532 , n48768 , n49020 );
and ( n63533 , n63532 , n48765 );
or ( n63534 , n63531 , n63533 );
and ( n63535 , n63534 , n33180 );
not ( n63536 , n49054 );
and ( n63537 , n63536 , n48583 );
not ( n63538 , n48845 );
xor ( n63539 , n49058 , n49134 );
and ( n63540 , n63538 , n63539 );
xnor ( n63541 , n49167 , n49260 );
and ( n63542 , n63541 , n48845 );
or ( n63543 , n63540 , n63542 );
and ( n63544 , n63543 , n49054 );
or ( n63545 , n63537 , n63544 );
and ( n63546 , n63545 , n33178 );
and ( n63547 , n49167 , n49275 );
or ( n63548 , n63499 , n63504 , n63509 , n63514 , n63519 , n63524 , n63529 , n63535 , n63546 , n63547 );
and ( n63549 , n63548 , n33208 );
and ( n63550 , n32976 , n35056 );
and ( n63551 , n48583 , n49286 );
or ( n63552 , C0 , n63549 , n63550 , n63551 );
buf ( n63553 , n63552 );
buf ( n63554 , n63553 );
buf ( n63555 , RI15b5eed8_1104);
and ( n63556 , n63555 , n32494 );
not ( n63557 , n46083 );
buf ( n63558 , RI15b604e0_1151);
and ( n63559 , n63557 , n63558 );
buf ( n63560 , n63559 );
and ( n63561 , n63560 , n32421 );
not ( n63562 , n46326 );
and ( n63563 , n63562 , n63558 );
not ( n63564 , n51396 );
and ( n63565 , n63564 , n51358 );
xor ( n63566 , n59211 , n59212 );
and ( n63567 , n63566 , n51396 );
or ( n63568 , n63565 , n63567 );
and ( n63569 , n63568 , n46326 );
or ( n63570 , n63563 , n63569 );
and ( n63571 , n63570 , n32417 );
and ( n63572 , n63558 , n46340 );
or ( n63573 , n63561 , n63571 , n63572 );
and ( n63574 , n63573 , n32456 );
and ( n63575 , n63558 , n46349 );
or ( n63576 , C0 , n63556 , n63574 , n63575 );
buf ( n63577 , n63576 );
buf ( n63578 , n63577 );
buf ( n63579 , n31655 );
not ( n63580 , n46356 );
and ( n63581 , n63580 , n31183 );
not ( n63582 , n53353 );
and ( n63583 , n63582 , n31183 );
and ( n63584 , n31205 , n53353 );
or ( n63585 , n63583 , n63584 );
and ( n63586 , n63585 , n46356 );
or ( n63587 , n63581 , n63586 );
and ( n63588 , n63587 , n31649 );
not ( n63589 , n53361 );
not ( n63590 , n53353 );
and ( n63591 , n63590 , n31183 );
and ( n63592 , n50125 , n53353 );
or ( n63593 , n63591 , n63592 );
and ( n63594 , n63589 , n63593 );
and ( n63595 , n50125 , n53361 );
or ( n63596 , n63594 , n63595 );
and ( n63597 , n63596 , n31643 );
not ( n63598 , n31452 );
not ( n63599 , n53361 );
not ( n63600 , n53353 );
and ( n63601 , n63600 , n31183 );
and ( n63602 , n50125 , n53353 );
or ( n63603 , n63601 , n63602 );
and ( n63604 , n63599 , n63603 );
and ( n63605 , n50125 , n53361 );
or ( n63606 , n63604 , n63605 );
and ( n63607 , n63598 , n63606 );
not ( n63608 , n53381 );
not ( n63609 , n53383 );
and ( n63610 , n63609 , n63606 );
and ( n63611 , n50151 , n53383 );
or ( n63612 , n63610 , n63611 );
and ( n63613 , n63608 , n63612 );
and ( n63614 , n50159 , n53381 );
or ( n63615 , n63613 , n63614 );
and ( n63616 , n63615 , n31452 );
or ( n63617 , n63607 , n63616 );
and ( n63618 , n63617 , n31638 );
and ( n63619 , n31183 , n47277 );
or ( n63620 , C0 , n63588 , n63597 , n63618 , n63619 );
buf ( n63621 , n63620 );
buf ( n63622 , n63621 );
buf ( n63623 , n30987 );
buf ( n63624 , n31655 );
not ( n63625 , n38443 );
and ( n63626 , n63625 , n38099 );
xor ( n63627 , n53476 , n53493 );
and ( n63628 , n63627 , n38443 );
or ( n63629 , n63626 , n63628 );
and ( n63630 , n63629 , n38450 );
not ( n63631 , n39339 );
and ( n63632 , n63631 , n38999 );
xor ( n63633 , n53532 , n53549 );
and ( n63634 , n63633 , n39339 );
or ( n63635 , n63632 , n63634 );
and ( n63636 , n63635 , n39346 );
and ( n63637 , n40208 , n39359 );
or ( n63638 , n63630 , n63636 , n63637 );
buf ( n63639 , n63638 );
buf ( n63640 , n63639 );
not ( n63641 , n46356 );
and ( n63642 , n63641 , n31649 );
not ( n63643 , n52614 );
and ( n63644 , n63643 , n31647 );
not ( n63645 , n31451 );
and ( n63646 , n63645 , n30990 );
buf ( n63647 , n31451 );
or ( n63648 , n63646 , n63647 );
and ( n63649 , n63648 , n31645 );
not ( n63650 , n61218 );
and ( n63651 , n63650 , n31009 );
and ( n63652 , n42328 , n48455 );
not ( n63653 , n48457 );
and ( n63654 , n63653 , n31014 );
and ( n63655 , n42328 , n48457 );
or ( n63656 , n63654 , n63655 );
and ( n63657 , n63656 , n31373 );
not ( n63658 , n44807 );
and ( n63659 , n63658 , n31014 );
and ( n63660 , n42324 , n44807 );
or ( n63661 , n63659 , n63660 );
and ( n63662 , n63661 , n31408 );
not ( n63663 , n48468 );
and ( n63664 , n63663 , n31014 );
and ( n63665 , n42328 , n48468 );
or ( n63666 , n63664 , n63665 );
and ( n63667 , n63666 , n31468 );
not ( n63668 , n44817 );
and ( n63669 , n63668 , n31014 );
and ( n63670 , n42328 , n44817 );
or ( n63671 , n63669 , n63670 );
and ( n63672 , n63671 , n31521 );
not ( n63673 , n39979 );
and ( n63674 , n63673 , n31014 );
or ( n63675 , n31018 , n62098 );
xor ( n63676 , n31014 , n63675 );
not ( n63677 , n63676 );
buf ( n63678 , n63677 );
buf ( n63679 , n63678 );
not ( n63680 , n63679 );
and ( n63681 , n63680 , n39979 );
or ( n63682 , n63674 , n63681 );
and ( n63683 , n63682 , n31538 );
not ( n63684 , n45059 );
and ( n63685 , n63684 , n31014 );
and ( n63686 , n63680 , n45059 );
or ( n63687 , n63685 , n63686 );
and ( n63688 , n63687 , n31536 );
and ( n63689 , n31014 , n61216 );
and ( n63690 , n33499 , n48513 );
or ( n63691 , n63652 , n63657 , n63662 , n63667 , n63672 , n63683 , n63688 , n63689 , n63690 );
not ( n63692 , n63691 );
and ( n63693 , n63692 , n31013 );
not ( n63694 , n62114 );
and ( n63695 , n63694 , n31017 );
and ( n63696 , n42315 , n48455 );
not ( n63697 , n48457 );
and ( n63698 , n63697 , n31022 );
and ( n63699 , n42315 , n48457 );
or ( n63700 , n63698 , n63699 );
and ( n63701 , n63700 , n31373 );
not ( n63702 , n44807 );
and ( n63703 , n63702 , n31022 );
and ( n63704 , n42311 , n44807 );
or ( n63705 , n63703 , n63704 );
and ( n63706 , n63705 , n31408 );
not ( n63707 , n48468 );
and ( n63708 , n63707 , n31022 );
and ( n63709 , n42315 , n48468 );
or ( n63710 , n63708 , n63709 );
and ( n63711 , n63710 , n31468 );
not ( n63712 , n44817 );
and ( n63713 , n63712 , n31022 );
and ( n63714 , n42315 , n44817 );
or ( n63715 , n63713 , n63714 );
and ( n63716 , n63715 , n31521 );
not ( n63717 , n39979 );
and ( n63718 , n63717 , n31022 );
xor ( n63719 , n31022 , n31026 );
not ( n63720 , n63719 );
buf ( n63721 , n63720 );
buf ( n63722 , n63721 );
not ( n63723 , n63722 );
and ( n63724 , n63723 , n39979 );
or ( n63725 , n63718 , n63724 );
and ( n63726 , n63725 , n31538 );
not ( n63727 , n45059 );
and ( n63728 , n63727 , n31022 );
and ( n63729 , n63723 , n45059 );
or ( n63730 , n63728 , n63729 );
and ( n63731 , n63730 , n31536 );
and ( n63732 , n31022 , n61216 );
and ( n63733 , n33488 , n48513 );
or ( n63734 , n63696 , n63701 , n63706 , n63711 , n63716 , n63726 , n63731 , n63732 , n63733 );
not ( n63735 , n63734 );
and ( n63736 , n63735 , n31021 );
and ( n63737 , n42309 , n48455 );
buf ( n63738 , n31026 );
and ( n63739 , n63738 , n31373 );
buf ( n63740 , n31026 );
and ( n63741 , n63740 , n31408 );
buf ( n63742 , n31026 );
and ( n63743 , n63742 , n31468 );
buf ( n63744 , n31026 );
and ( n63745 , n63744 , n31521 );
not ( n63746 , n39979 );
and ( n63747 , n63746 , n31026 );
not ( n63748 , n31026 );
not ( n63749 , n63748 );
buf ( n63750 , n63749 );
not ( n63751 , n63750 );
and ( n63752 , n63751 , n39979 );
or ( n63753 , n63747 , n63752 );
and ( n63754 , n63753 , n31538 );
not ( n63755 , n45059 );
and ( n63756 , n63755 , n31026 );
and ( n63757 , n63751 , n45059 );
or ( n63758 , n63756 , n63757 );
and ( n63759 , n63758 , n31536 );
and ( n63760 , n31026 , n61216 );
and ( n63761 , n33482 , n48513 );
or ( n63762 , n63737 , n63739 , n63741 , n63743 , n63745 , n63754 , n63759 , n63760 , n63761 );
not ( n63763 , n63762 );
and ( n63764 , n63763 , n31025 );
xnor ( n63765 , n63734 , n31021 );
and ( n63766 , n63764 , n63765 );
or ( n63767 , n63736 , n63766 );
xnor ( n63768 , n62114 , n31017 );
and ( n63769 , n63767 , n63768 );
or ( n63770 , n63695 , n63769 );
xnor ( n63771 , n63691 , n31013 );
and ( n63772 , n63770 , n63771 );
or ( n63773 , n63693 , n63772 );
xnor ( n63774 , n61218 , n31009 );
and ( n63775 , n63773 , n63774 );
or ( n63776 , n63651 , n63775 );
not ( n63777 , n63776 );
not ( n63778 , n61218 );
not ( n63779 , n63691 );
buf ( n63780 , n61218 );
buf ( n63781 , n61218 );
buf ( n63782 , n61218 );
buf ( n63783 , n61218 );
buf ( n63784 , n61218 );
buf ( n63785 , n61218 );
buf ( n63786 , n61218 );
buf ( n63787 , n61218 );
buf ( n63788 , n61218 );
buf ( n63789 , n61218 );
buf ( n63790 , n61218 );
buf ( n63791 , n61218 );
buf ( n63792 , n61218 );
buf ( n63793 , n61218 );
buf ( n63794 , n61218 );
buf ( n63795 , n61218 );
buf ( n63796 , n61218 );
buf ( n63797 , n61218 );
buf ( n63798 , n61218 );
buf ( n63799 , n61218 );
buf ( n63800 , n61218 );
buf ( n63801 , n61218 );
buf ( n63802 , n61218 );
buf ( n63803 , n61218 );
buf ( n63804 , n61218 );
buf ( n63805 , n61218 );
not ( n63806 , n62114 );
or ( n63807 , n63779 , n61218 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 );
nand ( n63808 , n63778 , n63807 );
or ( n63809 , n63808 , n44719 );
not ( n63810 , n31077 );
buf ( n63811 , n63810 );
buf ( n63812 , RI15b510a8_630);
not ( n63813 , n44703 );
and ( n63814 , n63812 , n63813 );
and ( n63815 , n63814 , n31077 );
or ( n63816 , n63811 , n63815 );
and ( n63817 , n63816 , n31373 );
not ( n63818 , n31402 );
buf ( n63819 , n63818 );
not ( n63820 , n31451 );
and ( n63821 , n63812 , n63820 );
and ( n63822 , n63821 , n31402 );
or ( n63823 , n63819 , n63822 );
and ( n63824 , n63823 , n31408 );
not ( n63825 , n31437 );
buf ( n63826 , n63825 );
and ( n63827 , n63814 , n31437 );
or ( n63828 , n63826 , n63827 );
and ( n63829 , n63828 , n31468 );
not ( n63830 , n31497 );
buf ( n63831 , n63830 );
and ( n63832 , n63821 , n31497 );
or ( n63833 , n63831 , n63832 );
and ( n63834 , n63833 , n31521 );
not ( n63835 , n39979 );
and ( n63836 , n63835 , n31538 );
not ( n63837 , n45059 );
and ( n63838 , n63837 , n31536 );
not ( n63839 , n33419 );
and ( n63840 , n63839 , n31529 );
not ( n63841 , n33734 );
and ( n63842 , n63841 , n31527 );
or ( n63843 , n63817 , n63824 , n63829 , n63834 , n63836 , n63838 , n63840 , n63842 , C0 );
or ( n63844 , n63809 , n63843 );
or ( n63845 , n63777 , n63844 );
not ( n63846 , n63845 );
and ( n63847 , n31437 , n31455 );
not ( n63848 , n63847 );
and ( n63849 , n63848 , n30990 );
buf ( n63850 , n63849 );
and ( n63851 , n63850 , n31468 );
or ( n63852 , n45795 , n31373 );
or ( n63853 , n63852 , n31540 );
or ( n63854 , n63853 , n31542 );
or ( n63855 , n63854 , n31544 );
or ( n63856 , n63855 , n31546 );
or ( n63857 , n63856 , n31548 );
or ( n63858 , n63857 , n31550 );
or ( n63859 , n63858 , n31552 );
and ( n63860 , n30990 , n63859 );
or ( n63861 , n63851 , n63860 );
and ( n63862 , n63846 , n63861 );
buf ( n63863 , n63845 );
or ( n63864 , n63862 , n63863 );
and ( n63865 , n63864 , n31557 );
buf ( n63866 , n31643 );
and ( n63867 , n59060 , n31641 );
buf ( n63868 , n31638 );
and ( n63869 , n59060 , n31640 );
or ( n63870 , n33973 , n31007 );
buf ( n63871 , n63870 );
or ( n63872 , C0 , n63642 , n63644 , n63649 , n63865 , n63866 , n63867 , n63868 , n63869 , n63871 );
buf ( n63873 , n63872 );
buf ( n63874 , n63873 );
buf ( n63875 , n31655 );
buf ( n63876 , n30987 );
xor ( n63877 , n34060 , n39927 );
and ( n63878 , n63877 , n31550 );
not ( n63879 , n39979 );
and ( n63880 , n63879 , n34060 );
buf ( n63881 , n31304 );
and ( n63882 , n63881 , n39979 );
or ( n63883 , n63880 , n63882 );
and ( n63884 , n63883 , n31538 );
and ( n63885 , n34060 , n40143 );
or ( n63886 , n63878 , n63884 , n63885 );
and ( n63887 , n63886 , n31557 );
and ( n63888 , n34060 , n40154 );
or ( n63889 , C0 , n63887 , n63888 );
buf ( n63890 , n63889 );
buf ( n63891 , n63890 );
not ( n63892 , n40163 );
and ( n63893 , n63892 , n31955 );
not ( n63894 , n57233 );
and ( n63895 , n63894 , n31955 );
and ( n63896 , n32183 , n57233 );
or ( n63897 , n63895 , n63896 );
and ( n63898 , n63897 , n40163 );
or ( n63899 , n63893 , n63898 );
and ( n63900 , n63899 , n32498 );
not ( n63901 , n57241 );
not ( n63902 , n57233 );
and ( n63903 , n63902 , n31955 );
and ( n63904 , n45178 , n57233 );
or ( n63905 , n63903 , n63904 );
and ( n63906 , n63901 , n63905 );
and ( n63907 , n45178 , n57241 );
or ( n63908 , n63906 , n63907 );
and ( n63909 , n63908 , n32473 );
not ( n63910 , n32475 );
not ( n63911 , n57241 );
not ( n63912 , n57233 );
and ( n63913 , n63912 , n31955 );
and ( n63914 , n45178 , n57233 );
or ( n63915 , n63913 , n63914 );
and ( n63916 , n63911 , n63915 );
and ( n63917 , n45178 , n57241 );
or ( n63918 , n63916 , n63917 );
and ( n63919 , n63910 , n63918 );
not ( n63920 , n57261 );
not ( n63921 , n57263 );
and ( n63922 , n63921 , n63918 );
and ( n63923 , n45206 , n57263 );
or ( n63924 , n63922 , n63923 );
and ( n63925 , n63920 , n63924 );
and ( n63926 , n45214 , n57261 );
or ( n63927 , n63925 , n63926 );
and ( n63928 , n63927 , n32475 );
or ( n63929 , n63919 , n63928 );
and ( n63930 , n63929 , n32486 );
and ( n63931 , n31955 , n41278 );
or ( n63932 , C0 , n63900 , n63909 , n63930 , n63931 );
buf ( n63933 , n63932 );
buf ( n63934 , n63933 );
buf ( n63935 , n31655 );
buf ( n63936 , n30987 );
buf ( n63937 , n30987 );
and ( n63938 , n31760 , n40163 );
buf ( n63939 , n63938 );
and ( n63940 , n63939 , n32498 );
and ( n63941 , n55776 , n32496 );
and ( n63942 , n47342 , n50275 );
not ( n63943 , n50278 );
and ( n63944 , n63943 , n31670 );
and ( n63945 , n47342 , n50278 );
or ( n63946 , n63944 , n63945 );
and ( n63947 , n63946 , n32421 );
not ( n63948 , n50002 );
and ( n63949 , n63948 , n31670 );
and ( n63950 , n47338 , n50002 );
or ( n63951 , n63949 , n63950 );
and ( n63952 , n63951 , n32419 );
not ( n63953 , n50289 );
and ( n63954 , n63953 , n31670 );
and ( n63955 , n47342 , n50289 );
or ( n63956 , n63954 , n63955 );
and ( n63957 , n63956 , n32417 );
not ( n63958 , n50008 );
and ( n63959 , n63958 , n31670 );
and ( n63960 , n47342 , n50008 );
or ( n63961 , n63959 , n63960 );
and ( n63962 , n63961 , n32415 );
not ( n63963 , n47331 );
and ( n63964 , n63963 , n31670 );
xor ( n63965 , n31670 , n31674 );
not ( n63966 , n63965 );
buf ( n63967 , n63966 );
buf ( n63968 , n63967 );
not ( n63969 , n63968 );
and ( n63970 , n63969 , n47331 );
or ( n63971 , n63964 , n63970 );
and ( n63972 , n63971 , n32413 );
not ( n63973 , n50067 );
and ( n63974 , n63973 , n31670 );
and ( n63975 , n63969 , n50067 );
or ( n63976 , n63974 , n63975 );
and ( n63977 , n63976 , n32411 );
or ( n63978 , n32398 , n32253 );
and ( n63979 , n31670 , n63978 );
and ( n63980 , n31760 , n50334 );
or ( n63981 , n63942 , n63947 , n63952 , n63957 , n63962 , n63972 , n63977 , n63979 , n63980 );
and ( n63982 , n63981 , n32456 );
or ( n63983 , n47406 , n32500 );
and ( n63984 , n31670 , n63983 );
or ( n63985 , C0 , n63940 , n63941 , n63982 , n63984 );
buf ( n63986 , n63985 );
buf ( n63987 , n63986 );
buf ( n63988 , n30987 );
buf ( n63989 , n31655 );
not ( n63990 , n36587 );
and ( n63991 , n63990 , n36328 );
xor ( n63992 , n50181 , n50206 );
and ( n63993 , n63992 , n36587 );
or ( n63994 , n63991 , n63993 );
and ( n63995 , n63994 , n36596 );
not ( n63996 , n37485 );
and ( n63997 , n63996 , n37230 );
xor ( n63998 , n50231 , n50256 );
and ( n63999 , n63998 , n37485 );
or ( n64000 , n63997 , n63999 );
and ( n64001 , n64000 , n37494 );
and ( n64002 , n41853 , n37506 );
or ( n64003 , n63995 , n64001 , n64002 );
buf ( n64004 , n64003 );
buf ( n64005 , n64004 );
buf ( n64006 , n31655 );
buf ( n64007 , n30987 );
buf ( n64008 , n31655 );
buf ( n64009 , n30987 );
not ( n64010 , n32953 );
buf ( n64011 , RI15b463b0_261);
and ( n64012 , n64010 , n64011 );
not ( n64013 , n54581 );
and ( n64014 , n64013 , n54458 );
xor ( n64015 , n54458 , n54340 );
xor ( n64016 , n54441 , n54340 );
xor ( n64017 , n54424 , n54340 );
xor ( n64018 , n54407 , n54340 );
xor ( n64019 , n54390 , n54340 );
xor ( n64020 , n54373 , n54340 );
and ( n64021 , n54584 , n54586 );
and ( n64022 , n64020 , n64021 );
and ( n64023 , n64019 , n64022 );
and ( n64024 , n64018 , n64023 );
and ( n64025 , n64017 , n64024 );
and ( n64026 , n64016 , n64025 );
xor ( n64027 , n64015 , n64026 );
and ( n64028 , n64027 , n54581 );
or ( n64029 , n64014 , n64028 );
and ( n64030 , n64029 , n32953 );
or ( n64031 , n64012 , n64030 );
and ( n64032 , n64031 , n33038 );
not ( n64033 , n48660 );
and ( n64034 , n64033 , n64011 );
not ( n64035 , n55168 );
and ( n64036 , n64035 , n55080 );
xor ( n64037 , n55080 , n34193 );
xor ( n64038 , n55068 , n34193 );
and ( n64039 , n55171 , n55181 );
and ( n64040 , n64038 , n64039 );
xor ( n64041 , n64037 , n64040 );
and ( n64042 , n64041 , n55168 );
or ( n64043 , n64036 , n64042 );
and ( n64044 , n64043 , n48660 );
or ( n64045 , n64034 , n64044 );
and ( n64046 , n64045 , n33172 );
and ( n64047 , n64011 , n39795 );
or ( n64048 , n64032 , n64046 , n64047 );
and ( n64049 , n64048 , n33208 );
and ( n64050 , n64011 , n39805 );
or ( n64051 , C0 , n64049 , n64050 );
buf ( n64052 , n64051 );
buf ( n64053 , n64052 );
buf ( n64054 , n31655 );
buf ( n64055 , n30987 );
not ( n64056 , n32953 );
buf ( n64057 , RI15b46428_262);
and ( n64058 , n64056 , n64057 );
not ( n64059 , n54581 );
and ( n64060 , n64059 , n54475 );
xor ( n64061 , n54475 , n54340 );
and ( n64062 , n64015 , n64026 );
xor ( n64063 , n64061 , n64062 );
and ( n64064 , n64063 , n54581 );
or ( n64065 , n64060 , n64064 );
and ( n64066 , n64065 , n32953 );
or ( n64067 , n64058 , n64066 );
and ( n64068 , n64067 , n33038 );
not ( n64069 , n48660 );
and ( n64070 , n64069 , n64057 );
not ( n64071 , n55168 );
and ( n64072 , n64071 , n55092 );
xor ( n64073 , n55092 , n34193 );
and ( n64074 , n64037 , n64040 );
xor ( n64075 , n64073 , n64074 );
and ( n64076 , n64075 , n55168 );
or ( n64077 , n64072 , n64076 );
and ( n64078 , n64077 , n48660 );
or ( n64079 , n64070 , n64078 );
and ( n64080 , n64079 , n33172 );
and ( n64081 , n64057 , n39795 );
or ( n64082 , n64068 , n64080 , n64081 );
and ( n64083 , n64082 , n33208 );
and ( n64084 , n64057 , n39805 );
or ( n64085 , C0 , n64083 , n64084 );
buf ( n64086 , n64085 );
buf ( n64087 , n64086 );
buf ( n64088 , n30987 );
buf ( n64089 , n31655 );
buf ( n64090 , n31655 );
xor ( n64091 , n49591 , n60310 );
and ( n64092 , n64091 , n32433 );
not ( n64093 , n47331 );
and ( n64094 , n64093 , n49591 );
and ( n64095 , n31750 , n47357 );
and ( n64096 , n31778 , n47359 );
and ( n64097 , n31781 , n47361 );
and ( n64098 , n31784 , n47363 );
and ( n64099 , n31787 , n47365 );
and ( n64100 , n31790 , n47367 );
and ( n64101 , n31793 , n47369 );
and ( n64102 , n31796 , n47371 );
and ( n64103 , n31799 , n47373 );
and ( n64104 , n31802 , n47375 );
and ( n64105 , n31805 , n47377 );
and ( n64106 , n31808 , n47379 );
and ( n64107 , n31811 , n47381 );
and ( n64108 , n31814 , n47383 );
and ( n64109 , n31817 , n47385 );
and ( n64110 , n31820 , n47387 );
or ( n64111 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 );
and ( n64112 , n64111 , n47331 );
or ( n64113 , n64094 , n64112 );
and ( n64114 , n64113 , n32413 );
and ( n64115 , n49591 , n47402 );
or ( n64116 , n64092 , n64114 , n64115 );
and ( n64117 , n64116 , n32456 );
and ( n64118 , n49591 , n47409 );
or ( n64119 , C0 , n64117 , n64118 );
buf ( n64120 , n64119 );
buf ( n64121 , n64120 );
buf ( n64122 , n30987 );
buf ( n64123 , n30987 );
not ( n64124 , n46356 );
and ( n64125 , n64124 , n31166 );
not ( n64126 , n47423 );
and ( n64127 , n64126 , n31166 );
and ( n64128 , n31172 , n47423 );
or ( n64129 , n64127 , n64128 );
and ( n64130 , n64129 , n46356 );
or ( n64131 , n64125 , n64130 );
and ( n64132 , n64131 , n31649 );
not ( n64133 , n47431 );
not ( n64134 , n47423 );
and ( n64135 , n64134 , n31166 );
and ( n64136 , n46495 , n47423 );
or ( n64137 , n64135 , n64136 );
and ( n64138 , n64133 , n64137 );
and ( n64139 , n46495 , n47431 );
or ( n64140 , n64138 , n64139 );
and ( n64141 , n64140 , n31643 );
not ( n64142 , n31452 );
not ( n64143 , n47431 );
not ( n64144 , n47423 );
and ( n64145 , n64144 , n31166 );
and ( n64146 , n46495 , n47423 );
or ( n64147 , n64145 , n64146 );
and ( n64148 , n64143 , n64147 );
and ( n64149 , n46495 , n47431 );
or ( n64150 , n64148 , n64149 );
and ( n64151 , n64142 , n64150 );
not ( n64152 , n47466 );
not ( n64153 , n47468 );
and ( n64154 , n64153 , n64150 );
and ( n64155 , n46984 , n47468 );
or ( n64156 , n64154 , n64155 );
and ( n64157 , n64152 , n64156 );
and ( n64158 , n47267 , n47466 );
or ( n64159 , n64157 , n64158 );
and ( n64160 , n64159 , n31452 );
or ( n64161 , n64151 , n64160 );
and ( n64162 , n64161 , n31638 );
and ( n64163 , n31166 , n47277 );
or ( n64164 , C0 , n64132 , n64141 , n64162 , n64163 );
buf ( n64165 , n64164 );
buf ( n64166 , n64165 );
buf ( n64167 , n31655 );
buf ( n64168 , n30987 );
and ( n64169 , n31583 , n31007 );
not ( n64170 , n31077 );
and ( n64171 , n64170 , n34007 );
buf ( n64172 , n64171 );
and ( n64173 , n64172 , n31373 );
not ( n64174 , n31402 );
and ( n64175 , n64174 , n34007 );
buf ( n64176 , n64175 );
and ( n64177 , n64176 , n31408 );
not ( n64178 , n31437 );
and ( n64179 , n64178 , n34007 );
not ( n64180 , n31455 );
and ( n64181 , n64180 , n34054 );
xor ( n64182 , n34007 , n34016 );
and ( n64183 , n64182 , n31455 );
or ( n64184 , n64181 , n64183 );
and ( n64185 , n64184 , n31437 );
or ( n64186 , n64179 , n64185 );
and ( n64187 , n64186 , n31468 );
not ( n64188 , n31497 );
and ( n64189 , n64188 , n34007 );
not ( n64190 , n31454 );
not ( n64191 , n31501 );
and ( n64192 , n64191 , n34054 );
xor ( n64193 , n34055 , n34068 );
and ( n64194 , n64193 , n31501 );
or ( n64195 , n64192 , n64194 );
and ( n64196 , n64190 , n64195 );
and ( n64197 , n64182 , n31454 );
or ( n64198 , n64196 , n64197 );
and ( n64199 , n64198 , n31497 );
or ( n64200 , n64189 , n64199 );
and ( n64201 , n64200 , n31521 );
and ( n64202 , n34007 , n31553 );
or ( n64203 , n64173 , n64177 , n64187 , n64201 , n64202 );
and ( n64204 , n64203 , n31557 );
not ( n64205 , n31452 );
not ( n64206 , n31619 );
and ( n64207 , n64206 , n34111 );
xor ( n64208 , n34112 , n34125 );
and ( n64209 , n64208 , n31619 );
or ( n64210 , n64207 , n64209 );
and ( n64211 , n64205 , n64210 );
and ( n64212 , n34007 , n31452 );
or ( n64213 , n64211 , n64212 );
and ( n64214 , n64213 , n31638 );
buf ( n64215 , n33973 );
and ( n64216 , n34007 , n31650 );
or ( n64217 , C0 , n64169 , n64204 , n64214 , n64215 , n64216 );
buf ( n64218 , n64217 );
buf ( n64219 , n64218 );
buf ( n64220 , n31655 );
buf ( n64221 , n31655 );
not ( n64222 , n33419 );
and ( n64223 , n64222 , n31561 );
xor ( n64224 , n59399 , n59400 );
and ( n64225 , n64224 , n33419 );
or ( n64226 , n64223 , n64225 );
and ( n64227 , n64226 , n31529 );
not ( n64228 , n33734 );
and ( n64229 , n64228 , n31561 );
not ( n64230 , n33533 );
xor ( n64231 , n59412 , n59413 );
and ( n64232 , n64230 , n64231 );
xnor ( n64233 , n59420 , n59421 );
and ( n64234 , n64233 , n33533 );
or ( n64235 , n64232 , n64234 );
and ( n64236 , n64235 , n33734 );
or ( n64237 , n64229 , n64236 );
and ( n64238 , n64237 , n31527 );
and ( n64239 , n31561 , n33942 );
or ( n64240 , n64227 , n64238 , n64239 );
and ( n64241 , n64240 , n31557 );
and ( n64242 , n35478 , n31643 );
not ( n64243 , n31452 );
and ( n64244 , n64243 , n35478 );
xor ( n64245 , n31561 , n59439 );
and ( n64246 , n64245 , n31452 );
or ( n64247 , n64244 , n64246 );
and ( n64248 , n64247 , n31638 );
and ( n64249 , n35387 , n33973 );
and ( n64250 , n31561 , n33978 );
or ( n64251 , C0 , n64241 , n64242 , n64248 , n64249 , n64250 );
buf ( n64252 , n64251 );
buf ( n64253 , n64252 );
buf ( n64254 , n30987 );
buf ( n64255 , n30987 );
not ( n64256 , n35278 );
buf ( n64257 , RI15b5f298_1112);
and ( n64258 , n64256 , n64257 );
not ( n64259 , n46290 );
and ( n64260 , n64259 , n46156 );
xor ( n64261 , n46301 , n46311 );
and ( n64262 , n64261 , n46290 );
or ( n64263 , n64260 , n64262 );
and ( n64264 , n64263 , n35278 );
or ( n64265 , n64258 , n64264 );
and ( n64266 , n64265 , n32417 );
not ( n64267 , n47912 );
and ( n64268 , n64267 , n64257 );
not ( n64269 , n48101 );
and ( n64270 , n64269 , n47977 );
xor ( n64271 , n48106 , n48116 );
and ( n64272 , n64271 , n48101 );
or ( n64273 , n64270 , n64272 );
and ( n64274 , n64273 , n47912 );
or ( n64275 , n64268 , n64274 );
and ( n64276 , n64275 , n32415 );
and ( n64277 , n64257 , n48133 );
or ( n64278 , n64266 , n64276 , n64277 );
and ( n64279 , n64278 , n32456 );
and ( n64280 , n64257 , n47409 );
or ( n64281 , C0 , n64279 , n64280 );
buf ( n64282 , n64281 );
buf ( n64283 , n64282 );
not ( n64284 , n46356 );
and ( n64285 , n64284 , n31140 );
not ( n64286 , n63024 );
and ( n64287 , n64286 , n31140 );
and ( n64288 , n31172 , n63024 );
or ( n64289 , n64287 , n64288 );
and ( n64290 , n64289 , n46356 );
or ( n64291 , n64285 , n64290 );
and ( n64292 , n64291 , n31649 );
not ( n64293 , n63032 );
not ( n64294 , n63024 );
and ( n64295 , n64294 , n31140 );
and ( n64296 , n46495 , n63024 );
or ( n64297 , n64295 , n64296 );
and ( n64298 , n64293 , n64297 );
and ( n64299 , n46495 , n63032 );
or ( n64300 , n64298 , n64299 );
and ( n64301 , n64300 , n31643 );
not ( n64302 , n31452 );
not ( n64303 , n63032 );
not ( n64304 , n63024 );
and ( n64305 , n64304 , n31140 );
and ( n64306 , n46495 , n63024 );
or ( n64307 , n64305 , n64306 );
and ( n64308 , n64303 , n64307 );
and ( n64309 , n46495 , n63032 );
or ( n64310 , n64308 , n64309 );
and ( n64311 , n64302 , n64310 );
not ( n64312 , n63052 );
not ( n64313 , n63054 );
and ( n64314 , n64313 , n64310 );
and ( n64315 , n46984 , n63054 );
or ( n64316 , n64314 , n64315 );
and ( n64317 , n64312 , n64316 );
and ( n64318 , n47267 , n63052 );
or ( n64319 , n64317 , n64318 );
and ( n64320 , n64319 , n31452 );
or ( n64321 , n64311 , n64320 );
and ( n64322 , n64321 , n31638 );
and ( n64323 , n31140 , n47277 );
or ( n64324 , C0 , n64292 , n64301 , n64322 , n64323 );
buf ( n64325 , n64324 );
buf ( n64326 , n64325 );
buf ( n64327 , n31655 );
buf ( n64328 , n30987 );
not ( n64329 , n36587 );
and ( n64330 , n64329 , n36345 );
xor ( n64331 , n50180 , n50207 );
and ( n64332 , n64331 , n36587 );
or ( n64333 , n64330 , n64332 );
and ( n64334 , n64333 , n36596 );
not ( n64335 , n37485 );
and ( n64336 , n64335 , n37247 );
xor ( n64337 , n50230 , n50257 );
and ( n64338 , n64337 , n37485 );
or ( n64339 , n64336 , n64338 );
and ( n64340 , n64339 , n37494 );
and ( n64341 , n41854 , n37506 );
or ( n64342 , n64334 , n64340 , n64341 );
buf ( n64343 , n64342 );
buf ( n64344 , n64343 );
buf ( n64345 , n31655 );
and ( n64346 , n31754 , n40163 );
buf ( n64347 , n64346 );
and ( n64348 , n64347 , n32498 );
and ( n64349 , n55760 , n32496 );
and ( n64350 , n47336 , n50275 );
buf ( n64351 , n31674 );
and ( n64352 , n64351 , n32421 );
buf ( n64353 , n31674 );
and ( n64354 , n64353 , n32419 );
buf ( n64355 , n31674 );
and ( n64356 , n64355 , n32417 );
buf ( n64357 , n31674 );
and ( n64358 , n64357 , n32415 );
not ( n64359 , n47331 );
and ( n64360 , n64359 , n31674 );
not ( n64361 , n31674 );
not ( n64362 , n64361 );
buf ( n64363 , n64362 );
not ( n64364 , n64363 );
and ( n64365 , n64364 , n47331 );
or ( n64366 , n64360 , n64365 );
and ( n64367 , n64366 , n32413 );
not ( n64368 , n50067 );
and ( n64369 , n64368 , n31674 );
and ( n64370 , n64364 , n50067 );
or ( n64371 , n64369 , n64370 );
and ( n64372 , n64371 , n32411 );
and ( n64373 , n31674 , n63978 );
and ( n64374 , n31754 , n50334 );
or ( n64375 , n64350 , n64352 , n64354 , n64356 , n64358 , n64367 , n64372 , n64373 , n64374 );
and ( n64376 , n64375 , n32456 );
and ( n64377 , n31674 , n63983 );
or ( n64378 , C0 , n64348 , n64349 , n64376 , n64377 );
buf ( n64379 , n64378 );
buf ( n64380 , n64379 );
buf ( n64381 , n30987 );
buf ( n64382 , n30987 );
buf ( n64383 , n31655 );
and ( n64384 , n48811 , n34150 );
buf ( n64385 , n64384 );
and ( n64386 , n64385 , n33381 );
and ( n64387 , n56625 , n33379 );
and ( n64388 , n57629 , n33208 );
and ( n64389 , n32535 , n61311 );
or ( n64390 , C0 , n64386 , n64387 , n64388 , n64389 );
buf ( n64391 , n64390 );
buf ( n64392 , n64391 );
buf ( n64393 , n31655 );
buf ( n64394 , n31655 );
buf ( n64395 , n31655 );
buf ( n64396 , n30987 );
and ( n64397 , n49062 , n48639 );
not ( n64398 , n48642 );
and ( n64399 , n64398 , n48587 );
and ( n64400 , n49062 , n48642 );
or ( n64401 , n64399 , n64400 );
and ( n64402 , n64401 , n32890 );
not ( n64403 , n48648 );
and ( n64404 , n64403 , n48587 );
and ( n64405 , n49062 , n48648 );
or ( n64406 , n64404 , n64405 );
and ( n64407 , n64406 , n32924 );
not ( n64408 , n48654 );
and ( n64409 , n64408 , n48587 );
and ( n64410 , n49062 , n48654 );
or ( n64411 , n64409 , n64410 );
and ( n64412 , n64411 , n33038 );
not ( n64413 , n48660 );
and ( n64414 , n64413 , n48587 );
and ( n64415 , n49062 , n48660 );
or ( n64416 , n64414 , n64415 );
and ( n64417 , n64416 , n33172 );
not ( n64418 , n41576 );
and ( n64419 , n64418 , n48587 );
and ( n64420 , n48772 , n41576 );
or ( n64421 , n64419 , n64420 );
and ( n64422 , n64421 , n33189 );
not ( n64423 , n48730 );
and ( n64424 , n64423 , n48587 );
and ( n64425 , n48772 , n48730 );
or ( n64426 , n64424 , n64425 );
and ( n64427 , n64426 , n33187 );
not ( n64428 , n48765 );
and ( n64429 , n64428 , n48587 );
xor ( n64430 , n48772 , n49016 );
and ( n64431 , n64430 , n48765 );
or ( n64432 , n64429 , n64431 );
and ( n64433 , n64432 , n33180 );
not ( n64434 , n49054 );
and ( n64435 , n64434 , n48587 );
not ( n64436 , n48845 );
xor ( n64437 , n49062 , n49130 );
and ( n64438 , n64436 , n64437 );
xnor ( n64439 , n49171 , n49256 );
and ( n64440 , n64439 , n48845 );
or ( n64441 , n64438 , n64440 );
and ( n64442 , n64441 , n49054 );
or ( n64443 , n64435 , n64442 );
and ( n64444 , n64443 , n33178 );
and ( n64445 , n49171 , n49275 );
or ( n64446 , n64397 , n64402 , n64407 , n64412 , n64417 , n64422 , n64427 , n64433 , n64444 , n64445 );
and ( n64447 , n64446 , n33208 );
and ( n64448 , n32980 , n35056 );
and ( n64449 , n48587 , n49286 );
or ( n64450 , C0 , n64447 , n64448 , n64449 );
buf ( n64451 , n64450 );
buf ( n64452 , n64451 );
buf ( n64453 , n30987 );
and ( n64454 , n49074 , n48639 );
not ( n64455 , n48642 );
and ( n64456 , n64455 , n48599 );
and ( n64457 , n49074 , n48642 );
or ( n64458 , n64456 , n64457 );
and ( n64459 , n64458 , n32890 );
not ( n64460 , n48648 );
and ( n64461 , n64460 , n48599 );
and ( n64462 , n49074 , n48648 );
or ( n64463 , n64461 , n64462 );
and ( n64464 , n64463 , n32924 );
not ( n64465 , n48654 );
and ( n64466 , n64465 , n48599 );
and ( n64467 , n49074 , n48654 );
or ( n64468 , n64466 , n64467 );
and ( n64469 , n64468 , n33038 );
not ( n64470 , n48660 );
and ( n64471 , n64470 , n48599 );
and ( n64472 , n49074 , n48660 );
or ( n64473 , n64471 , n64472 );
and ( n64474 , n64473 , n33172 );
not ( n64475 , n41576 );
and ( n64476 , n64475 , n48599 );
and ( n64477 , n48784 , n41576 );
or ( n64478 , n64476 , n64477 );
and ( n64479 , n64478 , n33189 );
not ( n64480 , n48730 );
and ( n64481 , n64480 , n48599 );
and ( n64482 , n48784 , n48730 );
or ( n64483 , n64481 , n64482 );
and ( n64484 , n64483 , n33187 );
not ( n64485 , n48765 );
and ( n64486 , n64485 , n48599 );
xor ( n64487 , n48784 , n49004 );
and ( n64488 , n64487 , n48765 );
or ( n64489 , n64486 , n64488 );
and ( n64490 , n64489 , n33180 );
not ( n64491 , n49054 );
and ( n64492 , n64491 , n48599 );
not ( n64493 , n48845 );
xor ( n64494 , n49074 , n49118 );
and ( n64495 , n64493 , n64494 );
xnor ( n64496 , n49183 , n49244 );
and ( n64497 , n64496 , n48845 );
or ( n64498 , n64495 , n64497 );
and ( n64499 , n64498 , n49054 );
or ( n64500 , n64492 , n64499 );
and ( n64501 , n64500 , n33178 );
and ( n64502 , n49183 , n49275 );
or ( n64503 , n64454 , n64459 , n64464 , n64469 , n64474 , n64479 , n64484 , n64490 , n64501 , n64502 );
and ( n64504 , n64503 , n33208 );
and ( n64505 , n32992 , n35056 );
and ( n64506 , n48599 , n49286 );
or ( n64507 , C0 , n64504 , n64505 , n64506 );
buf ( n64508 , n64507 );
buf ( n64509 , n64508 );
buf ( n64510 , n31655 );
buf ( n64511 , n30987 );
buf ( n64512 , n30987 );
buf ( n64513 , n31655 );
not ( n64514 , n46356 );
and ( n64515 , n64514 , n31290 );
not ( n64516 , n55263 );
and ( n64517 , n64516 , n31290 );
and ( n64518 , n31306 , n55263 );
or ( n64519 , n64517 , n64518 );
and ( n64520 , n64519 , n46356 );
or ( n64521 , n64515 , n64520 );
and ( n64522 , n64521 , n31649 );
not ( n64523 , n55271 );
not ( n64524 , n55263 );
and ( n64525 , n64524 , n31290 );
and ( n64526 , n58061 , n55263 );
or ( n64527 , n64525 , n64526 );
and ( n64528 , n64523 , n64527 );
and ( n64529 , n58061 , n55271 );
or ( n64530 , n64528 , n64529 );
and ( n64531 , n64530 , n31643 );
not ( n64532 , n31452 );
not ( n64533 , n55271 );
not ( n64534 , n55263 );
and ( n64535 , n64534 , n31290 );
and ( n64536 , n58061 , n55263 );
or ( n64537 , n64535 , n64536 );
and ( n64538 , n64533 , n64537 );
and ( n64539 , n58061 , n55271 );
or ( n64540 , n64538 , n64539 );
and ( n64541 , n64532 , n64540 );
not ( n64542 , n55291 );
not ( n64543 , n55293 );
and ( n64544 , n64543 , n64540 );
and ( n64545 , n58085 , n55293 );
or ( n64546 , n64544 , n64545 );
and ( n64547 , n64542 , n64546 );
and ( n64548 , n58093 , n55291 );
or ( n64549 , n64547 , n64548 );
and ( n64550 , n64549 , n31452 );
or ( n64551 , n64541 , n64550 );
and ( n64552 , n64551 , n31638 );
and ( n64553 , n31290 , n47277 );
or ( n64554 , C0 , n64522 , n64531 , n64552 , n64553 );
buf ( n64555 , n64554 );
buf ( n64556 , n64555 );
xor ( n64557 , n46120 , n49988 );
and ( n64558 , n64557 , n32431 );
not ( n64559 , n50002 );
and ( n64560 , n64559 , n46120 );
and ( n64561 , n40287 , n50002 );
or ( n64562 , n64560 , n64561 );
and ( n64563 , n64562 , n32419 );
not ( n64564 , n50008 );
and ( n64565 , n64564 , n46120 );
not ( n64566 , n47910 );
buf ( n64567 , RI15b5f1a8_1110);
and ( n64568 , n64566 , n64567 );
not ( n64569 , n48101 );
and ( n64570 , n64569 , n47953 );
xor ( n64571 , n48108 , n48114 );
and ( n64572 , n64571 , n48101 );
or ( n64573 , n64570 , n64572 );
and ( n64574 , n64573 , n47910 );
or ( n64575 , n64568 , n64574 );
and ( n64576 , n64575 , n50008 );
or ( n64577 , n64565 , n64576 );
and ( n64578 , n64577 , n32415 );
not ( n64579 , n50067 );
and ( n64580 , n64579 , n46120 );
and ( n64581 , n31963 , n50067 );
or ( n64582 , n64580 , n64581 );
and ( n64583 , n64582 , n32411 );
and ( n64584 , n46120 , n50098 );
or ( n64585 , n64558 , n64563 , n64578 , n64583 , n64584 );
and ( n64586 , n64585 , n32456 );
and ( n64587 , n46120 , n47409 );
or ( n64588 , C0 , n64586 , n64587 );
buf ( n64589 , n64588 );
buf ( n64590 , n64589 );
buf ( n64591 , n30987 );
buf ( n64592 , n31655 );
buf ( n64593 , n31655 );
and ( n64594 , n31767 , n40163 );
buf ( n64595 , n64594 );
and ( n64596 , n64595 , n32498 );
and ( n64597 , n55702 , n32496 );
and ( n64598 , n47348 , n50275 );
not ( n64599 , n50278 );
and ( n64600 , n64599 , n31666 );
and ( n64601 , n47348 , n50278 );
or ( n64602 , n64600 , n64601 );
and ( n64603 , n64602 , n32421 );
not ( n64604 , n50002 );
and ( n64605 , n64604 , n31666 );
and ( n64606 , n47344 , n50002 );
or ( n64607 , n64605 , n64606 );
and ( n64608 , n64607 , n32419 );
not ( n64609 , n50289 );
and ( n64610 , n64609 , n31666 );
and ( n64611 , n47348 , n50289 );
or ( n64612 , n64610 , n64611 );
and ( n64613 , n64612 , n32417 );
not ( n64614 , n50008 );
and ( n64615 , n64614 , n31666 );
and ( n64616 , n47348 , n50008 );
or ( n64617 , n64615 , n64616 );
and ( n64618 , n64617 , n32415 );
not ( n64619 , n47331 );
and ( n64620 , n64619 , n31666 );
and ( n64621 , n31670 , n31674 );
xnor ( n64622 , n31666 , n64621 );
not ( n64623 , n64622 );
buf ( n64624 , n64623 );
buf ( n64625 , n64624 );
not ( n64626 , n64625 );
and ( n64627 , n64626 , n47331 );
or ( n64628 , n64620 , n64627 );
and ( n64629 , n64628 , n32413 );
not ( n64630 , n50067 );
and ( n64631 , n64630 , n31666 );
and ( n64632 , n64626 , n50067 );
or ( n64633 , n64631 , n64632 );
and ( n64634 , n64633 , n32411 );
and ( n64635 , n31666 , n63978 );
and ( n64636 , n31767 , n50334 );
or ( n64637 , n64598 , n64603 , n64608 , n64613 , n64618 , n64629 , n64634 , n64635 , n64636 );
and ( n64638 , n64637 , n32456 );
and ( n64639 , n31666 , n63983 );
or ( n64640 , C0 , n64596 , n64597 , n64638 , n64639 );
buf ( n64641 , n64640 );
buf ( n64642 , n64641 );
buf ( n64643 , n31655 );
not ( n64644 , n36587 );
and ( n64645 , n64644 , n36311 );
xor ( n64646 , n50182 , n50205 );
and ( n64647 , n64646 , n36587 );
or ( n64648 , n64645 , n64647 );
and ( n64649 , n64648 , n36596 );
not ( n64650 , n37485 );
and ( n64651 , n64650 , n37213 );
xor ( n64652 , n50232 , n50255 );
and ( n64653 , n64652 , n37485 );
or ( n64654 , n64651 , n64653 );
and ( n64655 , n64654 , n37494 );
and ( n64656 , n41852 , n37506 );
or ( n64657 , n64649 , n64655 , n64656 );
buf ( n64658 , n64657 );
buf ( n64659 , n64658 );
buf ( n64660 , n30987 );
buf ( n64661 , n31655 );
buf ( n64662 , n30987 );
not ( n64663 , n34150 );
and ( n64664 , n64663 , n32659 );
not ( n64665 , n50731 );
and ( n64666 , n64665 , n32659 );
and ( n64667 , n32689 , n50731 );
or ( n64668 , n64666 , n64667 );
and ( n64669 , n64668 , n34150 );
or ( n64670 , n64664 , n64669 );
and ( n64671 , n64670 , n33381 );
not ( n64672 , n50739 );
not ( n64673 , n50731 );
and ( n64674 , n64673 , n32659 );
and ( n64675 , n50682 , n50731 );
or ( n64676 , n64674 , n64675 );
and ( n64677 , n64672 , n64676 );
and ( n64678 , n50682 , n50739 );
or ( n64679 , n64677 , n64678 );
and ( n64680 , n64679 , n33375 );
not ( n64681 , n32968 );
not ( n64682 , n50739 );
not ( n64683 , n50731 );
and ( n64684 , n64683 , n32659 );
and ( n64685 , n50682 , n50731 );
or ( n64686 , n64684 , n64685 );
and ( n64687 , n64682 , n64686 );
and ( n64688 , n50682 , n50739 );
or ( n64689 , n64687 , n64688 );
and ( n64690 , n64681 , n64689 );
not ( n64691 , n50759 );
not ( n64692 , n50761 );
and ( n64693 , n64692 , n64689 );
and ( n64694 , n50706 , n50761 );
or ( n64695 , n64693 , n64694 );
and ( n64696 , n64691 , n64695 );
and ( n64697 , n50714 , n50759 );
or ( n64698 , n64696 , n64697 );
and ( n64699 , n64698 , n32968 );
or ( n64700 , n64690 , n64699 );
and ( n64701 , n64700 , n33370 );
and ( n64702 , n32659 , n35062 );
or ( n64703 , C0 , n64671 , n64680 , n64701 , n64702 );
buf ( n64704 , n64703 );
buf ( n64705 , n64704 );
buf ( n64706 , n30987 );
buf ( n64707 , n31655 );
and ( n64708 , n46263 , n49999 );
and ( n64709 , n46276 , n64708 );
and ( n64710 , n50900 , n64709 );
and ( n64711 , n50973 , n64710 );
and ( n64712 , n50971 , n64711 );
and ( n64713 , n50969 , n64712 );
and ( n64714 , n50967 , n64713 );
and ( n64715 , n50965 , n64714 );
and ( n64716 , n50963 , n64715 );
xor ( n64717 , n50961 , n64716 );
and ( n64718 , n64717 , n32431 );
not ( n64719 , n50002 );
and ( n64720 , n64719 , n50961 );
and ( n64721 , n40606 , n50002 );
or ( n64722 , n64720 , n64721 );
and ( n64723 , n64722 , n32419 );
not ( n64724 , n50008 );
and ( n64725 , n64724 , n50961 );
and ( n64726 , n59269 , n50008 );
or ( n64727 , n64725 , n64726 );
and ( n64728 , n64727 , n32415 );
not ( n64729 , n50067 );
and ( n64730 , n64729 , n50961 );
xor ( n64731 , n60484 , n60542 );
and ( n64732 , n64731 , n50067 );
or ( n64733 , n64730 , n64732 );
and ( n64734 , n64733 , n32411 );
and ( n64735 , n50961 , n50098 );
or ( n64736 , n64718 , n64723 , n64728 , n64734 , n64735 );
and ( n64737 , n64736 , n32456 );
and ( n64738 , n50961 , n47409 );
or ( n64739 , C0 , n64737 , n64738 );
buf ( n64740 , n64739 );
buf ( n64741 , n64740 );
buf ( n64742 , n31655 );
buf ( n64743 , n31655 );
not ( n64744 , n46356 );
and ( n64745 , n64744 , n31160 );
nor ( n64746 , n46359 , n31021 , n48213 , n31013 , n31009 );
not ( n64747 , n64746 );
and ( n64748 , n64747 , n31160 );
and ( n64749 , n31172 , n64746 );
or ( n64750 , n64748 , n64749 );
and ( n64751 , n64750 , n46356 );
or ( n64752 , n64745 , n64751 );
and ( n64753 , n64752 , n31649 );
nor ( n64754 , n46374 , n46379 , n48222 , n46392 , C0 );
not ( n64755 , n64754 );
not ( n64756 , n64746 );
and ( n64757 , n64756 , n31160 );
and ( n64758 , n46495 , n64746 );
or ( n64759 , n64757 , n64758 );
and ( n64760 , n64755 , n64759 );
and ( n64761 , n46495 , n64754 );
or ( n64762 , n64760 , n64761 );
and ( n64763 , n64762 , n31643 );
not ( n64764 , n31452 );
not ( n64765 , n64754 );
not ( n64766 , n64746 );
and ( n64767 , n64766 , n31160 );
and ( n64768 , n46495 , n64746 );
or ( n64769 , n64767 , n64768 );
and ( n64770 , n64765 , n64769 );
and ( n64771 , n46495 , n64754 );
or ( n64772 , n64770 , n64771 );
and ( n64773 , n64764 , n64772 );
nor ( n64774 , n46520 , n46528 , n48243 , n46549 , C0 );
not ( n64775 , n64774 );
nor ( n64776 , n46552 , n46524 , n48246 , n46544 , C0 );
not ( n64777 , n64776 );
and ( n64778 , n64777 , n64772 );
and ( n64779 , n46984 , n64776 );
or ( n64780 , n64778 , n64779 );
and ( n64781 , n64775 , n64780 );
and ( n64782 , n47267 , n64774 );
or ( n64783 , n64781 , n64782 );
and ( n64784 , n64783 , n31452 );
or ( n64785 , n64773 , n64784 );
and ( n64786 , n64785 , n31638 );
and ( n64787 , n31160 , n47277 );
or ( n64788 , C0 , n64753 , n64763 , n64786 , n64787 );
buf ( n64789 , n64788 );
buf ( n64790 , n64789 );
buf ( n64791 , n30987 );
buf ( n64792 , RI15b47a30_309);
buf ( n64793 , n64792 );
buf ( n64794 , n31655 );
buf ( n64795 , n31655 );
buf ( n64796 , n30987 );
buf ( n64797 , n30987 );
and ( n64798 , n49070 , n48639 );
not ( n64799 , n48642 );
and ( n64800 , n64799 , n48595 );
and ( n64801 , n49070 , n48642 );
or ( n64802 , n64800 , n64801 );
and ( n64803 , n64802 , n32890 );
not ( n64804 , n48648 );
and ( n64805 , n64804 , n48595 );
and ( n64806 , n49070 , n48648 );
or ( n64807 , n64805 , n64806 );
and ( n64808 , n64807 , n32924 );
not ( n64809 , n48654 );
and ( n64810 , n64809 , n48595 );
and ( n64811 , n49070 , n48654 );
or ( n64812 , n64810 , n64811 );
and ( n64813 , n64812 , n33038 );
not ( n64814 , n48660 );
and ( n64815 , n64814 , n48595 );
and ( n64816 , n49070 , n48660 );
or ( n64817 , n64815 , n64816 );
and ( n64818 , n64817 , n33172 );
not ( n64819 , n41576 );
and ( n64820 , n64819 , n48595 );
and ( n64821 , n48780 , n41576 );
or ( n64822 , n64820 , n64821 );
and ( n64823 , n64822 , n33189 );
not ( n64824 , n48730 );
and ( n64825 , n64824 , n48595 );
and ( n64826 , n48780 , n48730 );
or ( n64827 , n64825 , n64826 );
and ( n64828 , n64827 , n33187 );
not ( n64829 , n48765 );
and ( n64830 , n64829 , n48595 );
xor ( n64831 , n48780 , n49008 );
and ( n64832 , n64831 , n48765 );
or ( n64833 , n64830 , n64832 );
and ( n64834 , n64833 , n33180 );
not ( n64835 , n49054 );
and ( n64836 , n64835 , n48595 );
not ( n64837 , n48845 );
xor ( n64838 , n49070 , n49122 );
and ( n64839 , n64837 , n64838 );
xnor ( n64840 , n49179 , n49248 );
and ( n64841 , n64840 , n48845 );
or ( n64842 , n64839 , n64841 );
and ( n64843 , n64842 , n49054 );
or ( n64844 , n64836 , n64843 );
and ( n64845 , n64844 , n33178 );
and ( n64846 , n49179 , n49275 );
or ( n64847 , n64798 , n64803 , n64808 , n64813 , n64818 , n64823 , n64828 , n64834 , n64845 , n64846 );
and ( n64848 , n64847 , n33208 );
and ( n64849 , n32988 , n35056 );
and ( n64850 , n48595 , n49286 );
or ( n64851 , C0 , n64848 , n64849 , n64850 );
buf ( n64852 , n64851 );
buf ( n64853 , n64852 );
buf ( n64854 , n31655 );
buf ( n64855 , n30987 );
xor ( n64856 , n54152 , n54983 );
and ( n64857 , n64856 , n33199 );
not ( n64858 , n48648 );
and ( n64859 , n64858 , n54152 );
and ( n64860 , n34437 , n48648 );
or ( n64861 , n64859 , n64860 );
and ( n64862 , n64861 , n32924 );
not ( n64863 , n48660 );
and ( n64864 , n64863 , n54152 );
not ( n64865 , n55168 );
and ( n64866 , n64865 , n55044 );
xor ( n64867 , n55172 , n55180 );
and ( n64868 , n64867 , n55168 );
or ( n64869 , n64866 , n64868 );
and ( n64870 , n64869 , n48660 );
or ( n64871 , n64864 , n64870 );
and ( n64872 , n64871 , n33172 );
not ( n64873 , n48730 );
and ( n64874 , n64873 , n54152 );
and ( n64875 , n32757 , n55215 );
and ( n64876 , n32759 , n55217 );
and ( n64877 , n32761 , n55219 );
and ( n64878 , n32763 , n55221 );
and ( n64879 , n32765 , n55223 );
and ( n64880 , n32767 , n55225 );
and ( n64881 , n32769 , n55227 );
and ( n64882 , n32771 , n55229 );
and ( n64883 , n32773 , n55231 );
and ( n64884 , n32775 , n55233 );
and ( n64885 , n32777 , n55235 );
and ( n64886 , n32779 , n55237 );
and ( n64887 , n32781 , n55239 );
and ( n64888 , n32783 , n55241 );
and ( n64889 , n32785 , n55243 );
and ( n64890 , n32787 , n55245 );
or ( n64891 , n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , n64889 , n64890 );
and ( n64892 , n64891 , n48730 );
or ( n64893 , n64874 , n64892 );
and ( n64894 , n64893 , n33187 );
and ( n64895 , n54152 , n54713 );
or ( n64896 , n64857 , n64862 , n64872 , n64894 , n64895 );
and ( n64897 , n64896 , n33208 );
and ( n64898 , n54152 , n39805 );
or ( n64899 , C0 , n64897 , n64898 );
buf ( n64900 , n64899 );
buf ( n64901 , n64900 );
buf ( n64902 , n30987 );
buf ( n64903 , n31655 );
not ( n64904 , n41532 );
and ( n64905 , n64904 , n34441 );
buf ( n64906 , RI15b53bc8_722);
and ( n64907 , n64906 , n41532 );
or ( n64908 , n64905 , n64907 );
buf ( n64909 , n64908 );
buf ( n64910 , n64909 );
buf ( n64911 , n31655 );
buf ( n64912 , n30987 );
not ( n64913 , n32953 );
buf ( n64914 , RI15b46338_260);
and ( n64915 , n64913 , n64914 );
not ( n64916 , n54581 );
and ( n64917 , n64916 , n54441 );
xor ( n64918 , n64016 , n64025 );
and ( n64919 , n64918 , n54581 );
or ( n64920 , n64917 , n64919 );
and ( n64921 , n64920 , n32953 );
or ( n64922 , n64915 , n64921 );
and ( n64923 , n64922 , n33038 );
not ( n64924 , n48660 );
and ( n64925 , n64924 , n64914 );
not ( n64926 , n55168 );
and ( n64927 , n64926 , n55068 );
xor ( n64928 , n64038 , n64039 );
and ( n64929 , n64928 , n55168 );
or ( n64930 , n64927 , n64929 );
and ( n64931 , n64930 , n48660 );
or ( n64932 , n64925 , n64931 );
and ( n64933 , n64932 , n33172 );
and ( n64934 , n64914 , n39795 );
or ( n64935 , n64923 , n64933 , n64934 );
and ( n64936 , n64935 , n33208 );
and ( n64937 , n64914 , n39805 );
or ( n64938 , C0 , n64936 , n64937 );
buf ( n64939 , n64938 );
buf ( n64940 , n64939 );
buf ( n64941 , n30987 );
buf ( n64942 , n31655 );
buf ( n64943 , n31655 );
not ( n64944 , n46356 );
and ( n64945 , n64944 , n31193 );
not ( n64946 , n64746 );
and ( n64947 , n64946 , n31193 );
and ( n64948 , n31205 , n64746 );
or ( n64949 , n64947 , n64948 );
and ( n64950 , n64949 , n46356 );
or ( n64951 , n64945 , n64950 );
and ( n64952 , n64951 , n31649 );
not ( n64953 , n64754 );
not ( n64954 , n64746 );
and ( n64955 , n64954 , n31193 );
and ( n64956 , n50125 , n64746 );
or ( n64957 , n64955 , n64956 );
and ( n64958 , n64953 , n64957 );
and ( n64959 , n50125 , n64754 );
or ( n64960 , n64958 , n64959 );
and ( n64961 , n64960 , n31643 );
not ( n64962 , n31452 );
not ( n64963 , n64754 );
not ( n64964 , n64746 );
and ( n64965 , n64964 , n31193 );
and ( n64966 , n50125 , n64746 );
or ( n64967 , n64965 , n64966 );
and ( n64968 , n64963 , n64967 );
and ( n64969 , n50125 , n64754 );
or ( n64970 , n64968 , n64969 );
and ( n64971 , n64962 , n64970 );
not ( n64972 , n64774 );
not ( n64973 , n64776 );
and ( n64974 , n64973 , n64970 );
and ( n64975 , n50151 , n64776 );
or ( n64976 , n64974 , n64975 );
and ( n64977 , n64972 , n64976 );
and ( n64978 , n50159 , n64774 );
or ( n64979 , n64977 , n64978 );
and ( n64980 , n64979 , n31452 );
or ( n64981 , n64971 , n64980 );
and ( n64982 , n64981 , n31638 );
and ( n64983 , n31193 , n47277 );
or ( n64984 , C0 , n64952 , n64961 , n64982 , n64983 );
buf ( n64985 , n64984 );
buf ( n64986 , n64985 );
buf ( n64987 , n31655 );
xor ( n64988 , n50963 , n64715 );
and ( n64989 , n64988 , n32431 );
not ( n64990 , n50002 );
and ( n64991 , n64990 , n50963 );
and ( n64992 , n40613 , n50002 );
or ( n64993 , n64991 , n64992 );
and ( n64994 , n64993 , n32419 );
not ( n64995 , n50008 );
and ( n64996 , n64995 , n50963 );
and ( n64997 , n51612 , n50008 );
or ( n64998 , n64996 , n64997 );
and ( n64999 , n64998 , n32415 );
not ( n65000 , n50067 );
and ( n65001 , n65000 , n50963 );
and ( n65002 , n62040 , n50067 );
or ( n65003 , n65001 , n65002 );
and ( n65004 , n65003 , n32411 );
and ( n65005 , n50963 , n50098 );
or ( n65006 , n64989 , n64994 , n64999 , n65004 , n65005 );
and ( n65007 , n65006 , n32456 );
and ( n65008 , n50963 , n47409 );
or ( n65009 , C0 , n65007 , n65008 );
buf ( n65010 , n65009 );
buf ( n65011 , n65010 );
buf ( n65012 , n30987 );
buf ( n65013 , RI15b47c10_313);
buf ( n65014 , n65013 );
buf ( n65015 , n30987 );
buf ( n65016 , n30987 );
buf ( n65017 , n31655 );
buf ( n65018 , RI15b48048_322);
and ( n65019 , n65018 , n58207 );
and ( n65020 , n54734 , n44695 );
or ( n65021 , n65019 , n65020 );
buf ( n65022 , n65021 );
buf ( n65023 , n65022 );
buf ( n65024 , n31655 );
buf ( n65025 , n31655 );
buf ( n65026 , n30987 );
not ( n65027 , n34150 );
and ( n65028 , n65027 , n32690 );
not ( n65029 , n56708 );
and ( n65030 , n65029 , n32690 );
and ( n65031 , n32722 , n56708 );
or ( n65032 , n65030 , n65031 );
and ( n65033 , n65032 , n34150 );
or ( n65034 , n65028 , n65033 );
and ( n65035 , n65034 , n33381 );
not ( n65036 , n56716 );
not ( n65037 , n56708 );
and ( n65038 , n65037 , n32690 );
and ( n65039 , n42565 , n56708 );
or ( n65040 , n65038 , n65039 );
and ( n65041 , n65036 , n65040 );
and ( n65042 , n42565 , n56716 );
or ( n65043 , n65041 , n65042 );
and ( n65044 , n65043 , n33375 );
not ( n65045 , n32968 );
not ( n65046 , n56716 );
not ( n65047 , n56708 );
and ( n65048 , n65047 , n32690 );
and ( n65049 , n42565 , n56708 );
or ( n65050 , n65048 , n65049 );
and ( n65051 , n65046 , n65050 );
and ( n65052 , n42565 , n56716 );
or ( n65053 , n65051 , n65052 );
and ( n65054 , n65045 , n65053 );
not ( n65055 , n56736 );
not ( n65056 , n56738 );
and ( n65057 , n65056 , n65053 );
and ( n65058 , n42589 , n56738 );
or ( n65059 , n65057 , n65058 );
and ( n65060 , n65055 , n65059 );
and ( n65061 , n42597 , n56736 );
or ( n65062 , n65060 , n65061 );
and ( n65063 , n65062 , n32968 );
or ( n65064 , n65054 , n65063 );
and ( n65065 , n65064 , n33370 );
and ( n65066 , n32690 , n35062 );
or ( n65067 , C0 , n65035 , n65044 , n65065 , n65066 );
buf ( n65068 , n65067 );
buf ( n65069 , n65068 );
buf ( n65070 , n30987 );
buf ( n65071 , n31655 );
buf ( n65072 , n31655 );
buf ( n65073 , n30987 );
not ( n65074 , n32953 );
buf ( n65075 , RI15b464a0_263);
and ( n65076 , n65074 , n65075 );
not ( n65077 , n54581 );
and ( n65078 , n65077 , n54492 );
xor ( n65079 , n54492 , n54340 );
and ( n65080 , n64061 , n64062 );
xor ( n65081 , n65079 , n65080 );
and ( n65082 , n65081 , n54581 );
or ( n65083 , n65078 , n65082 );
and ( n65084 , n65083 , n32953 );
or ( n65085 , n65076 , n65084 );
and ( n65086 , n65085 , n33038 );
not ( n65087 , n48660 );
and ( n65088 , n65087 , n65075 );
not ( n65089 , n55168 );
and ( n65090 , n65089 , n55104 );
xor ( n65091 , n55104 , n34193 );
and ( n65092 , n64073 , n64074 );
xor ( n65093 , n65091 , n65092 );
and ( n65094 , n65093 , n55168 );
or ( n65095 , n65090 , n65094 );
and ( n65096 , n65095 , n48660 );
or ( n65097 , n65088 , n65096 );
and ( n65098 , n65097 , n33172 );
and ( n65099 , n65075 , n39795 );
or ( n65100 , n65086 , n65098 , n65099 );
and ( n65101 , n65100 , n33208 );
and ( n65102 , n65075 , n39805 );
or ( n65103 , C0 , n65101 , n65102 );
buf ( n65104 , n65103 );
buf ( n65105 , n65104 );
buf ( n65106 , n30987 );
buf ( n65107 , n31655 );
buf ( n65108 , n31655 );
and ( n65109 , n33775 , n48455 );
not ( n65110 , n48457 );
and ( n65111 , n65110 , n33438 );
and ( n65112 , n33775 , n48457 );
or ( n65113 , n65111 , n65112 );
and ( n65114 , n65113 , n31373 );
not ( n65115 , n44807 );
and ( n65116 , n65115 , n33438 );
and ( n65117 , n33775 , n44807 );
or ( n65118 , n65116 , n65117 );
and ( n65119 , n65118 , n31408 );
not ( n65120 , n48468 );
and ( n65121 , n65120 , n33438 );
and ( n65122 , n33775 , n48468 );
or ( n65123 , n65121 , n65122 );
and ( n65124 , n65123 , n31468 );
not ( n65125 , n44817 );
and ( n65126 , n65125 , n33438 );
and ( n65127 , n33775 , n44817 );
or ( n65128 , n65126 , n65127 );
and ( n65129 , n65128 , n31521 );
not ( n65130 , n39979 );
and ( n65131 , n65130 , n33438 );
and ( n65132 , n33554 , n39979 );
or ( n65133 , n65131 , n65132 );
and ( n65134 , n65133 , n31538 );
not ( n65135 , n45059 );
and ( n65136 , n65135 , n33438 );
and ( n65137 , n33554 , n45059 );
or ( n65138 , n65136 , n65137 );
and ( n65139 , n65138 , n31536 );
not ( n65140 , n33419 );
and ( n65141 , n65140 , n33438 );
and ( n65142 , n61018 , n33419 );
or ( n65143 , n65141 , n65142 );
and ( n65144 , n65143 , n31529 );
not ( n65145 , n33734 );
and ( n65146 , n65145 , n33438 );
and ( n65147 , n61031 , n33734 );
or ( n65148 , n65146 , n65147 );
and ( n65149 , n65148 , n31527 );
and ( n65150 , n33864 , n48513 );
or ( n65151 , n65109 , n65114 , n65119 , n65124 , n65129 , n65134 , n65139 , n65144 , n65149 , n65150 );
and ( n65152 , n65151 , n31557 );
and ( n65153 , n34010 , n33973 );
and ( n65154 , n33438 , n48524 );
or ( n65155 , C0 , n65152 , n65153 , n65154 );
buf ( n65156 , n65155 );
buf ( n65157 , n65156 );
buf ( n65158 , n30987 );
not ( n65159 , n35278 );
buf ( n65160 , RI15b5ecf8_1100);
and ( n65161 , n65159 , n65160 );
not ( n65162 , n51396 );
and ( n65163 , n65162 , n51290 );
xor ( n65164 , n53330 , n53333 );
and ( n65165 , n65164 , n51396 );
or ( n65166 , n65163 , n65165 );
and ( n65167 , n65166 , n35278 );
or ( n65168 , n65161 , n65167 );
and ( n65169 , n65168 , n32417 );
not ( n65170 , n50008 );
and ( n65171 , n65170 , n65160 );
not ( n65172 , n51594 );
and ( n65173 , n65172 , n51518 );
xor ( n65174 , n59229 , n59232 );
and ( n65175 , n65174 , n51594 );
or ( n65176 , n65173 , n65175 );
and ( n65177 , n65176 , n50008 );
or ( n65178 , n65171 , n65177 );
and ( n65179 , n65178 , n32415 );
and ( n65180 , n65160 , n48133 );
or ( n65181 , n65169 , n65179 , n65180 );
and ( n65182 , n65181 , n32456 );
and ( n65183 , n65160 , n47409 );
or ( n65184 , C0 , n65182 , n65183 );
buf ( n65185 , n65184 );
buf ( n65186 , n65185 );
buf ( n65187 , RI15b52ea8_694);
and ( n65188 , n65187 , n31645 );
not ( n65189 , n45274 );
buf ( n65190 , RI15b53628_710);
and ( n65191 , n65189 , n65190 );
not ( n65192 , n41809 );
and ( n65193 , n65192 , n41688 );
xor ( n65194 , n41814 , n41826 );
and ( n65195 , n65194 , n41809 );
or ( n65196 , n65193 , n65195 );
and ( n65197 , n65196 , n45274 );
or ( n65198 , n65191 , n65197 );
and ( n65199 , n65198 , n31373 );
not ( n65200 , n45280 );
and ( n65201 , n65200 , n65190 );
and ( n65202 , n65196 , n45280 );
or ( n65203 , n65201 , n65202 );
and ( n65204 , n65203 , n31468 );
and ( n65205 , n65190 , n45802 );
or ( n65206 , n65199 , n65204 , n65205 );
and ( n65207 , n65206 , n31557 );
and ( n65208 , n65190 , n45808 );
or ( n65209 , C0 , n65188 , n65207 , n65208 );
buf ( n65210 , n65209 );
buf ( n65211 , n65210 );
buf ( n65212 , n31655 );
buf ( n65213 , n30987 );
not ( n65214 , n40163 );
and ( n65215 , n65214 , n32040 );
not ( n65216 , n56287 );
and ( n65217 , n65216 , n32040 );
and ( n65218 , n32130 , n56287 );
or ( n65219 , n65217 , n65218 );
and ( n65220 , n65219 , n40163 );
or ( n65221 , n65215 , n65220 );
and ( n65222 , n65221 , n32498 );
not ( n65223 , n56295 );
not ( n65224 , n56287 );
and ( n65225 , n65224 , n32040 );
and ( n65226 , n45833 , n56287 );
or ( n65227 , n65225 , n65226 );
and ( n65228 , n65223 , n65227 );
and ( n65229 , n45833 , n56295 );
or ( n65230 , n65228 , n65229 );
and ( n65231 , n65230 , n32473 );
not ( n65232 , n32475 );
not ( n65233 , n56295 );
not ( n65234 , n56287 );
and ( n65235 , n65234 , n32040 );
and ( n65236 , n45833 , n56287 );
or ( n65237 , n65235 , n65236 );
and ( n65238 , n65233 , n65237 );
and ( n65239 , n45833 , n56295 );
or ( n65240 , n65238 , n65239 );
and ( n65241 , n65232 , n65240 );
not ( n65242 , n56315 );
not ( n65243 , n56317 );
and ( n65244 , n65243 , n65240 );
and ( n65245 , n45857 , n56317 );
or ( n65246 , n65244 , n65245 );
and ( n65247 , n65242 , n65246 );
and ( n65248 , n45865 , n56315 );
or ( n65249 , n65247 , n65248 );
and ( n65250 , n65249 , n32475 );
or ( n65251 , n65241 , n65250 );
and ( n65252 , n65251 , n32486 );
and ( n65253 , n32040 , n41278 );
or ( n65254 , C0 , n65222 , n65231 , n65252 , n65253 );
buf ( n65255 , n65254 );
buf ( n65256 , n65255 );
buf ( n65257 , n30987 );
not ( n65258 , n41532 );
and ( n65259 , n65258 , n34425 );
and ( n65260 , n52207 , n41532 );
or ( n65261 , n65259 , n65260 );
buf ( n65262 , n65261 );
buf ( n65263 , n65262 );
xor ( n65264 , n39519 , n54975 );
and ( n65265 , n65264 , n33199 );
not ( n65266 , n48648 );
and ( n65267 , n65266 , n39519 );
and ( n65268 , n34371 , n48648 );
or ( n65269 , n65267 , n65268 );
and ( n65270 , n65269 , n32924 );
not ( n65271 , n48660 );
and ( n65272 , n65271 , n39519 );
not ( n65273 , n39584 );
and ( n65274 , n65273 , n60616 );
and ( n65275 , n60632 , n39584 );
or ( n65276 , n65274 , n65275 );
and ( n65277 , n65276 , n48660 );
or ( n65278 , n65272 , n65277 );
and ( n65279 , n65278 , n33172 );
not ( n65280 , n48730 );
and ( n65281 , n65280 , n39519 );
and ( n65282 , n52284 , n48730 );
or ( n65283 , n65281 , n65282 );
and ( n65284 , n65283 , n33187 );
and ( n65285 , n39519 , n54713 );
or ( n65286 , n65265 , n65270 , n65279 , n65284 , n65285 );
and ( n65287 , n65286 , n33208 );
and ( n65288 , n39519 , n39805 );
or ( n65289 , C0 , n65287 , n65288 );
buf ( n65290 , n65289 );
buf ( n65291 , n65290 );
buf ( n65292 , n30987 );
buf ( n65293 , n31655 );
buf ( n65294 , n31655 );
and ( n65295 , n50961 , n64716 );
xor ( n65296 , n50959 , n65295 );
and ( n65297 , n65296 , n32431 );
not ( n65298 , n50002 );
and ( n65299 , n65298 , n50959 );
and ( n65300 , n40599 , n50002 );
or ( n65301 , n65299 , n65300 );
and ( n65302 , n65301 , n32419 );
not ( n65303 , n50008 );
and ( n65304 , n65303 , n50959 );
and ( n65305 , n65176 , n50008 );
or ( n65306 , n65304 , n65305 );
and ( n65307 , n65306 , n32415 );
not ( n65308 , n50067 );
and ( n65309 , n65308 , n50959 );
and ( n65310 , n60484 , n60542 );
xor ( n65311 , n60467 , n65310 );
and ( n65312 , n65311 , n50067 );
or ( n65313 , n65309 , n65312 );
and ( n65314 , n65313 , n32411 );
and ( n65315 , n50959 , n50098 );
or ( n65316 , n65297 , n65302 , n65307 , n65314 , n65315 );
and ( n65317 , n65316 , n32456 );
and ( n65318 , n50959 , n47409 );
or ( n65319 , C0 , n65317 , n65318 );
buf ( n65320 , n65319 );
buf ( n65321 , n65320 );
buf ( n65322 , n31655 );
not ( n65323 , n46356 );
and ( n65324 , n65323 , n31120 );
not ( n65325 , n64746 );
and ( n65326 , n65325 , n31120 );
and ( n65327 , n31138 , n64746 );
or ( n65328 , n65326 , n65327 );
and ( n65329 , n65328 , n46356 );
or ( n65330 , n65324 , n65329 );
and ( n65331 , n65330 , n31649 );
not ( n65332 , n64754 );
not ( n65333 , n64746 );
and ( n65334 , n65333 , n31120 );
and ( n65335 , n56920 , n64746 );
or ( n65336 , n65334 , n65335 );
and ( n65337 , n65332 , n65336 );
and ( n65338 , n56920 , n64754 );
or ( n65339 , n65337 , n65338 );
and ( n65340 , n65339 , n31643 );
not ( n65341 , n31452 );
not ( n65342 , n64754 );
not ( n65343 , n64746 );
and ( n65344 , n65343 , n31120 );
and ( n65345 , n56920 , n64746 );
or ( n65346 , n65344 , n65345 );
and ( n65347 , n65342 , n65346 );
and ( n65348 , n56920 , n64754 );
or ( n65349 , n65347 , n65348 );
and ( n65350 , n65341 , n65349 );
not ( n65351 , n64774 );
not ( n65352 , n64776 );
and ( n65353 , n65352 , n65349 );
and ( n65354 , n56946 , n64776 );
or ( n65355 , n65353 , n65354 );
and ( n65356 , n65351 , n65355 );
and ( n65357 , n56954 , n64774 );
or ( n65358 , n65356 , n65357 );
and ( n65359 , n65358 , n31452 );
or ( n65360 , n65350 , n65359 );
and ( n65361 , n65360 , n31638 );
and ( n65362 , n31120 , n47277 );
or ( n65363 , C0 , n65331 , n65340 , n65361 , n65362 );
buf ( n65364 , n65363 );
buf ( n65365 , n65364 );
buf ( n65366 , n31655 );
buf ( n65367 , RI15b47850_305);
buf ( n65368 , n65367 );
buf ( n65369 , n30987 );
not ( n65370 , n31728 );
and ( n65371 , n65370 , n46034 );
xor ( n65372 , n47611 , n47618 );
and ( n65373 , n65372 , n31728 );
or ( n65374 , n65371 , n65373 );
and ( n65375 , n65374 , n32253 );
not ( n65376 , n32283 );
and ( n65377 , n65376 , n46034 );
not ( n65378 , n31823 );
xor ( n65379 , n47666 , n47673 );
and ( n65380 , n65378 , n65379 );
xnor ( n65381 , n47716 , n47723 );
and ( n65382 , n65381 , n31823 );
or ( n65383 , n65380 , n65382 );
and ( n65384 , n65383 , n32283 );
or ( n65385 , n65377 , n65384 );
and ( n65386 , n65385 , n32398 );
and ( n65387 , n46034 , n32436 );
or ( n65388 , n65375 , n65386 , n65387 );
and ( n65389 , n65388 , n32456 );
and ( n65390 , n49685 , n32473 );
not ( n65391 , n32475 );
and ( n65392 , n65391 , n49685 );
xor ( n65393 , n46034 , n47752 );
and ( n65394 , n65393 , n32475 );
or ( n65395 , n65392 , n65394 );
and ( n65396 , n65395 , n32486 );
and ( n65397 , n37565 , n32489 );
and ( n65398 , n46034 , n32501 );
or ( n65399 , C0 , n65389 , n65390 , n65396 , n65397 , n65398 );
buf ( n65400 , n65399 );
buf ( n65401 , n65400 );
buf ( n65402 , n31655 );
buf ( n65403 , n30987 );
and ( n65404 , n33216 , n32528 );
not ( n65405 , n32598 );
and ( n65406 , n65405 , n32979 );
buf ( n65407 , n65406 );
and ( n65408 , n65407 , n32890 );
not ( n65409 , n32919 );
and ( n65410 , n65409 , n32979 );
buf ( n65411 , n65410 );
and ( n65412 , n65411 , n32924 );
not ( n65413 , n32953 );
and ( n65414 , n65413 , n32979 );
not ( n65415 , n32971 );
and ( n65416 , n65415 , n33083 );
xor ( n65417 , n32979 , n33026 );
and ( n65418 , n65417 , n32971 );
or ( n65419 , n65416 , n65418 );
and ( n65420 , n65419 , n32953 );
or ( n65421 , n65414 , n65420 );
and ( n65422 , n65421 , n33038 );
not ( n65423 , n33067 );
and ( n65424 , n65423 , n32979 );
not ( n65425 , n32970 );
not ( n65426 , n33071 );
and ( n65427 , n65426 , n33083 );
xor ( n65428 , n33084 , n33158 );
and ( n65429 , n65428 , n33071 );
or ( n65430 , n65427 , n65429 );
and ( n65431 , n65425 , n65430 );
and ( n65432 , n65417 , n32970 );
or ( n65433 , n65431 , n65432 );
and ( n65434 , n65433 , n33067 );
or ( n65435 , n65424 , n65434 );
and ( n65436 , n65435 , n33172 );
and ( n65437 , n32979 , n33204 );
or ( n65438 , n65408 , n65412 , n65422 , n65436 , n65437 );
and ( n65439 , n65438 , n33208 );
not ( n65440 , n32968 );
not ( n65441 , n33270 );
and ( n65442 , n65441 , n33283 );
xor ( n65443 , n33284 , n33358 );
and ( n65444 , n65443 , n33270 );
or ( n65445 , n65442 , n65444 );
and ( n65446 , n65440 , n65445 );
and ( n65447 , n32979 , n32968 );
or ( n65448 , n65446 , n65447 );
and ( n65449 , n65448 , n33370 );
and ( n65450 , n32979 , n33382 );
or ( n65451 , C0 , n65404 , n65439 , n65449 , C0 , n65450 );
buf ( n65452 , n65451 );
buf ( n65453 , n65452 );
buf ( n65454 , n30987 );
buf ( n65455 , n31655 );
buf ( n65456 , RI15b46068_254);
and ( n65457 , n65456 , n33377 );
not ( n65458 , n48545 );
buf ( n65459 , RI15b47670_301);
and ( n65460 , n65458 , n65459 );
xor ( n65461 , n39568 , n39374 );
and ( n65462 , n42614 , n42639 );
and ( n65463 , n65461 , n65462 );
buf ( n65464 , n65463 );
and ( n65465 , n65464 , n39572 );
buf ( n65466 , n65465 );
and ( n65467 , n65466 , n48545 );
or ( n65468 , n65460 , n65467 );
and ( n65469 , n65468 , n32890 );
not ( n65470 , n48557 );
and ( n65471 , n65470 , n65459 );
not ( n65472 , n54581 );
and ( n65473 , n65472 , n54130 );
xor ( n65474 , n54585 , n54340 );
and ( n65475 , n65474 , n54581 );
or ( n65476 , n65473 , n65475 );
and ( n65477 , n65476 , n48557 );
or ( n65478 , n65471 , n65477 );
and ( n65479 , n65478 , n33038 );
and ( n65480 , n65459 , n48571 );
or ( n65481 , n65469 , n65479 , n65480 );
and ( n65482 , n65481 , n33208 );
and ( n65483 , n65459 , n48577 );
or ( n65484 , C0 , n65457 , n65482 , n65483 );
buf ( n65485 , n65484 );
buf ( n65486 , n65485 );
buf ( n65487 , n31655 );
buf ( n65488 , n30987 );
buf ( n65489 , n30987 );
buf ( n65490 , n31655 );
buf ( n65491 , n30987 );
buf ( n65492 , n31655 );
not ( n65493 , n31437 );
buf ( n65494 , RI15b524d0_673);
and ( n65495 , n65493 , n65494 );
not ( n65496 , n45766 );
and ( n65497 , n65496 , n45328 );
xor ( n65498 , n45778 , n45525 );
and ( n65499 , n65498 , n45766 );
or ( n65500 , n65497 , n65499 );
and ( n65501 , n65500 , n31437 );
or ( n65502 , n65495 , n65501 );
and ( n65503 , n65502 , n31468 );
not ( n65504 , n44817 );
and ( n65505 , n65504 , n65494 );
not ( n65506 , n44994 );
and ( n65507 , n65506 , n44823 );
xor ( n65508 , n45010 , n41881 );
and ( n65509 , n65508 , n44994 );
or ( n65510 , n65507 , n65509 );
and ( n65511 , n65510 , n44817 );
or ( n65512 , n65505 , n65511 );
and ( n65513 , n65512 , n31521 );
and ( n65514 , n65494 , n42158 );
or ( n65515 , n65503 , n65513 , n65514 );
and ( n65516 , n65515 , n31557 );
and ( n65517 , n65494 , n40154 );
or ( n65518 , C0 , n65516 , n65517 );
buf ( n65519 , n65518 );
buf ( n65520 , n65519 );
and ( n65521 , n47666 , n50275 );
not ( n65522 , n50278 );
and ( n65523 , n65522 , n47579 );
and ( n65524 , n47666 , n50278 );
or ( n65525 , n65523 , n65524 );
and ( n65526 , n65525 , n32421 );
not ( n65527 , n50002 );
and ( n65528 , n65527 , n47579 );
and ( n65529 , n47666 , n50002 );
or ( n65530 , n65528 , n65529 );
and ( n65531 , n65530 , n32419 );
not ( n65532 , n50289 );
and ( n65533 , n65532 , n47579 );
and ( n65534 , n47666 , n50289 );
or ( n65535 , n65533 , n65534 );
and ( n65536 , n65535 , n32417 );
not ( n65537 , n50008 );
and ( n65538 , n65537 , n47579 );
and ( n65539 , n47666 , n50008 );
or ( n65540 , n65538 , n65539 );
and ( n65541 , n65540 , n32415 );
not ( n65542 , n47331 );
and ( n65543 , n65542 , n47579 );
and ( n65544 , n47611 , n47331 );
or ( n65545 , n65543 , n65544 );
and ( n65546 , n65545 , n32413 );
not ( n65547 , n50067 );
and ( n65548 , n65547 , n47579 );
and ( n65549 , n47611 , n50067 );
or ( n65550 , n65548 , n65549 );
and ( n65551 , n65550 , n32411 );
not ( n65552 , n31728 );
and ( n65553 , n65552 , n47579 );
and ( n65554 , n65372 , n31728 );
or ( n65555 , n65553 , n65554 );
and ( n65556 , n65555 , n32253 );
not ( n65557 , n32283 );
and ( n65558 , n65557 , n47579 );
and ( n65559 , n65383 , n32283 );
or ( n65560 , n65558 , n65559 );
and ( n65561 , n65560 , n32398 );
and ( n65562 , n47716 , n50334 );
or ( n65563 , n65521 , n65526 , n65531 , n65536 , n65541 , n65546 , n65551 , n65556 , n65561 , n65562 );
and ( n65564 , n65563 , n32456 );
and ( n65565 , n37565 , n32489 );
and ( n65566 , n47579 , n50345 );
or ( n65567 , C0 , n65564 , n65565 , n65566 );
buf ( n65568 , n65567 );
buf ( n65569 , n65568 );
buf ( n65570 , n31655 );
not ( n65571 , n40163 );
and ( n65572 , n65571 , n31914 );
not ( n65573 , n49298 );
and ( n65574 , n65573 , n31914 );
and ( n65575 , n32200 , n49298 );
or ( n65576 , n65574 , n65575 );
and ( n65577 , n65576 , n40163 );
or ( n65578 , n65572 , n65577 );
and ( n65579 , n65578 , n32498 );
not ( n65580 , n49306 );
not ( n65581 , n49298 );
and ( n65582 , n65581 , n31914 );
and ( n65583 , n53243 , n49298 );
or ( n65584 , n65582 , n65583 );
and ( n65585 , n65580 , n65584 );
and ( n65586 , n53243 , n49306 );
or ( n65587 , n65585 , n65586 );
and ( n65588 , n65587 , n32473 );
not ( n65589 , n32475 );
not ( n65590 , n49306 );
not ( n65591 , n49298 );
and ( n65592 , n65591 , n31914 );
and ( n65593 , n53243 , n49298 );
or ( n65594 , n65592 , n65593 );
and ( n65595 , n65590 , n65594 );
and ( n65596 , n53243 , n49306 );
or ( n65597 , n65595 , n65596 );
and ( n65598 , n65589 , n65597 );
not ( n65599 , n49331 );
not ( n65600 , n49333 );
and ( n65601 , n65600 , n65597 );
and ( n65602 , n53269 , n49333 );
or ( n65603 , n65601 , n65602 );
and ( n65604 , n65599 , n65603 );
and ( n65605 , n53277 , n49331 );
or ( n65606 , n65604 , n65605 );
and ( n65607 , n65606 , n32475 );
or ( n65608 , n65598 , n65607 );
and ( n65609 , n65608 , n32486 );
and ( n65610 , n31914 , n41278 );
or ( n65611 , C0 , n65579 , n65588 , n65609 , n65610 );
buf ( n65612 , n65611 );
buf ( n65613 , n65612 );
buf ( n65614 , n30987 );
buf ( n65615 , n30987 );
xor ( n65616 , n41756 , n44787 );
and ( n65617 , n65616 , n31548 );
not ( n65618 , n44807 );
and ( n65619 , n65618 , n41756 );
and ( n65620 , n42062 , n44807 );
or ( n65621 , n65619 , n65620 );
and ( n65622 , n65621 , n31408 );
not ( n65623 , n44817 );
and ( n65624 , n65623 , n41756 );
not ( n65625 , n41835 );
buf ( n65626 , RI15b53178_700);
and ( n65627 , n65625 , n65626 );
not ( n65628 , n42124 );
and ( n65629 , n65628 , n42072 );
xor ( n65630 , n49376 , n49383 );
and ( n65631 , n65630 , n42124 );
or ( n65632 , n65629 , n65631 );
and ( n65633 , n65632 , n41835 );
or ( n65634 , n65627 , n65633 );
and ( n65635 , n65634 , n44817 );
or ( n65636 , n65624 , n65635 );
and ( n65637 , n65636 , n31521 );
not ( n65638 , n45059 );
and ( n65639 , n65638 , n41756 );
and ( n65640 , n31240 , n42330 );
and ( n65641 , n31242 , n42332 );
and ( n65642 , n31244 , n42334 );
and ( n65643 , n31246 , n42336 );
and ( n65644 , n31248 , n42338 );
and ( n65645 , n31250 , n42340 );
and ( n65646 , n31252 , n42342 );
and ( n65647 , n31254 , n42344 );
and ( n65648 , n31256 , n42346 );
and ( n65649 , n31258 , n42348 );
and ( n65650 , n31260 , n42350 );
and ( n65651 , n31262 , n42352 );
and ( n65652 , n31264 , n42354 );
and ( n65653 , n31266 , n42356 );
and ( n65654 , n31268 , n42358 );
and ( n65655 , n31270 , n42360 );
or ( n65656 , n65640 , n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , n65655 );
and ( n65657 , n65656 , n45059 );
or ( n65658 , n65639 , n65657 );
and ( n65659 , n65658 , n31536 );
and ( n65660 , n41756 , n45148 );
or ( n65661 , n65617 , n65622 , n65637 , n65659 , n65660 );
and ( n65662 , n65661 , n31557 );
and ( n65663 , n41756 , n40154 );
or ( n65664 , C0 , n65662 , n65663 );
buf ( n65665 , n65664 );
buf ( n65666 , n65665 );
xor ( n65667 , n49587 , n60312 );
and ( n65668 , n65667 , n32433 );
not ( n65669 , n47331 );
and ( n65670 , n65669 , n49587 );
and ( n65671 , n32001 , n60510 );
and ( n65672 , n32003 , n60512 );
and ( n65673 , n32005 , n60514 );
and ( n65674 , n32007 , n60516 );
and ( n65675 , n32009 , n60518 );
and ( n65676 , n32011 , n60520 );
and ( n65677 , n32013 , n60522 );
and ( n65678 , n32015 , n60524 );
and ( n65679 , n32017 , n60526 );
and ( n65680 , n32019 , n60528 );
and ( n65681 , n32021 , n60530 );
and ( n65682 , n32023 , n60532 );
and ( n65683 , n32025 , n60534 );
and ( n65684 , n32027 , n60536 );
and ( n65685 , n32029 , n60538 );
and ( n65686 , n32031 , n60540 );
or ( n65687 , n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , n65685 , n65686 );
and ( n65688 , n65687 , n47331 );
or ( n65689 , n65670 , n65688 );
and ( n65690 , n65689 , n32413 );
and ( n65691 , n49587 , n47402 );
or ( n65692 , n65668 , n65690 , n65691 );
and ( n65693 , n65692 , n32456 );
and ( n65694 , n49587 , n47409 );
or ( n65695 , C0 , n65693 , n65694 );
buf ( n65696 , n65695 );
buf ( n65697 , n65696 );
buf ( n65698 , n31655 );
buf ( n65699 , n30987 );
buf ( n65700 , n30987 );
buf ( n65701 , n31655 );
not ( n65702 , n46356 );
and ( n65703 , n65702 , n31368 );
not ( n65704 , n61975 );
and ( n65705 , n65704 , n31368 );
and ( n65706 , n31372 , n61975 );
or ( n65707 , n65705 , n65706 );
and ( n65708 , n65707 , n46356 );
or ( n65709 , n65703 , n65708 );
and ( n65710 , n65709 , n31649 );
not ( n65711 , n61983 );
not ( n65712 , n61975 );
and ( n65713 , n65712 , n31368 );
and ( n65714 , n47849 , n61975 );
or ( n65715 , n65713 , n65714 );
and ( n65716 , n65711 , n65715 );
and ( n65717 , n47849 , n61983 );
or ( n65718 , n65716 , n65717 );
and ( n65719 , n65718 , n31643 );
not ( n65720 , n31452 );
not ( n65721 , n61983 );
not ( n65722 , n61975 );
and ( n65723 , n65722 , n31368 );
and ( n65724 , n47849 , n61975 );
or ( n65725 , n65723 , n65724 );
and ( n65726 , n65721 , n65725 );
and ( n65727 , n47849 , n61983 );
or ( n65728 , n65726 , n65727 );
and ( n65729 , n65720 , n65728 );
not ( n65730 , n62003 );
not ( n65731 , n62005 );
and ( n65732 , n65731 , n65728 );
and ( n65733 , n47877 , n62005 );
or ( n65734 , n65732 , n65733 );
and ( n65735 , n65730 , n65734 );
and ( n65736 , n47887 , n62003 );
or ( n65737 , n65735 , n65736 );
and ( n65738 , n65737 , n31452 );
or ( n65739 , n65729 , n65738 );
and ( n65740 , n65739 , n31638 );
and ( n65741 , n31368 , n47277 );
or ( n65742 , C0 , n65710 , n65719 , n65740 , n65741 );
buf ( n65743 , n65742 );
buf ( n65744 , n65743 );
not ( n65745 , n31437 );
buf ( n65746 , RI15b52ae8_686);
and ( n65747 , n65745 , n65746 );
not ( n65748 , n45766 );
and ( n65749 , n65748 , n45745 );
xor ( n65750 , n45886 , n45893 );
and ( n65751 , n65750 , n45766 );
or ( n65752 , n65749 , n65751 );
and ( n65753 , n65752 , n31437 );
or ( n65754 , n65747 , n65753 );
and ( n65755 , n65754 , n31468 );
not ( n65756 , n44817 );
and ( n65757 , n65756 , n65746 );
and ( n65758 , n45026 , n44817 );
or ( n65759 , n65757 , n65758 );
and ( n65760 , n65759 , n31521 );
and ( n65761 , n65746 , n42158 );
or ( n65762 , n65755 , n65760 , n65761 );
and ( n65763 , n65762 , n31557 );
and ( n65764 , n65746 , n40154 );
or ( n65765 , C0 , n65763 , n65764 );
buf ( n65766 , n65765 );
buf ( n65767 , n65766 );
and ( n65768 , n31740 , n50275 );
buf ( n65769 , n31740 );
and ( n65770 , n65769 , n32421 );
buf ( n65771 , n31740 );
and ( n65772 , n65771 , n32419 );
buf ( n65773 , n31740 );
and ( n65774 , n65773 , n32417 );
buf ( n65775 , n31740 );
and ( n65776 , n65775 , n32415 );
not ( n65777 , n47331 );
and ( n65778 , n65777 , n31740 );
and ( n65779 , n32035 , n47331 );
or ( n65780 , n65778 , n65779 );
and ( n65781 , n65780 , n32413 );
not ( n65782 , n50067 );
and ( n65783 , n65782 , n31740 );
and ( n65784 , n32035 , n50067 );
or ( n65785 , n65783 , n65784 );
and ( n65786 , n65785 , n32411 );
not ( n65787 , n31728 );
and ( n65788 , n65787 , n31740 );
xor ( n65789 , n32035 , n32068 );
and ( n65790 , n65789 , n31728 );
or ( n65791 , n65788 , n65790 );
and ( n65792 , n65791 , n32253 );
not ( n65793 , n32283 );
and ( n65794 , n65793 , n31740 );
not ( n65795 , n31823 );
xor ( n65796 , n31740 , n32068 );
and ( n65797 , n65795 , n65796 );
xor ( n65798 , n32368 , n32369 );
and ( n65799 , n65798 , n31823 );
or ( n65800 , n65797 , n65799 );
and ( n65801 , n65800 , n32283 );
or ( n65802 , n65794 , n65801 );
and ( n65803 , n65802 , n32398 );
and ( n65804 , n32368 , n50334 );
or ( n65805 , n65768 , n65770 , n65772 , n65774 , n65776 , n65781 , n65786 , n65792 , n65803 , n65804 );
and ( n65806 , n65805 , n32456 );
and ( n65807 , n35213 , n32489 );
and ( n65808 , n31740 , n50345 );
or ( n65809 , C0 , n65806 , n65807 , n65808 );
buf ( n65810 , n65809 );
buf ( n65811 , n65810 );
buf ( n65812 , n31655 );
buf ( n65813 , n30987 );
buf ( n65814 , n30987 );
not ( n65815 , n36587 );
and ( n65816 , n65815 , n36362 );
xor ( n65817 , n50179 , n50208 );
and ( n65818 , n65817 , n36587 );
or ( n65819 , n65816 , n65818 );
and ( n65820 , n65819 , n36596 );
not ( n65821 , n37485 );
and ( n65822 , n65821 , n37264 );
xor ( n65823 , n50229 , n50258 );
and ( n65824 , n65823 , n37485 );
or ( n65825 , n65822 , n65824 );
and ( n65826 , n65825 , n37494 );
and ( n65827 , n41855 , n37506 );
or ( n65828 , n65820 , n65826 , n65827 );
buf ( n65829 , n65828 );
buf ( n65830 , n65829 );
buf ( n65831 , n31655 );
and ( n65832 , n50407 , n50438 );
xor ( n65833 , n55565 , n65832 );
and ( n65834 , n65833 , n50275 );
not ( n65835 , n50278 );
and ( n65836 , n65835 , n55565 );
and ( n65837 , n65833 , n50278 );
or ( n65838 , n65836 , n65837 );
and ( n65839 , n65838 , n32421 );
not ( n65840 , n50002 );
and ( n65841 , n65840 , n55565 );
and ( n65842 , n65833 , n50002 );
or ( n65843 , n65841 , n65842 );
and ( n65844 , n65843 , n32419 );
not ( n65845 , n50289 );
and ( n65846 , n65845 , n55565 );
and ( n65847 , n65833 , n50289 );
or ( n65848 , n65846 , n65847 );
and ( n65849 , n65848 , n32417 );
not ( n65850 , n50008 );
and ( n65851 , n65850 , n55565 );
and ( n65852 , n65833 , n50008 );
or ( n65853 , n65851 , n65852 );
and ( n65854 , n65853 , n32415 );
not ( n65855 , n47331 );
and ( n65856 , n65855 , n55565 );
and ( n65857 , n50407 , n50416 );
xor ( n65858 , n55565 , n65857 );
and ( n65859 , n65858 , n47331 );
or ( n65860 , n65856 , n65859 );
and ( n65861 , n65860 , n32413 );
not ( n65862 , n50067 );
and ( n65863 , n65862 , n55565 );
and ( n65864 , n65858 , n50067 );
or ( n65865 , n65863 , n65864 );
and ( n65866 , n65865 , n32411 );
not ( n65867 , n31728 );
and ( n65868 , n65867 , n55565 );
and ( n65869 , n50417 , n50426 );
xor ( n65870 , n65858 , n65869 );
and ( n65871 , n65870 , n31728 );
or ( n65872 , n65868 , n65871 );
and ( n65873 , n65872 , n32253 );
not ( n65874 , n32283 );
and ( n65875 , n65874 , n55565 );
not ( n65876 , n31823 );
and ( n65877 , n50439 , n50448 );
xor ( n65878 , n65833 , n65877 );
and ( n65879 , n65876 , n65878 );
and ( n65880 , n50407 , n50455 );
xor ( n65881 , n55565 , n65880 );
or ( n65882 , n50456 , n50465 );
xnor ( n65883 , n65881 , n65882 );
and ( n65884 , n65883 , n31823 );
or ( n65885 , n65879 , n65884 );
and ( n65886 , n65885 , n32283 );
or ( n65887 , n65875 , n65886 );
and ( n65888 , n65887 , n32398 );
and ( n65889 , n65881 , n50334 );
or ( n65890 , n65834 , n65839 , n65844 , n65849 , n65854 , n65861 , n65866 , n65873 , n65888 , n65889 );
and ( n65891 , n65890 , n32456 );
and ( n65892 , n37512 , n32489 );
and ( n65893 , n55565 , n50345 );
or ( n65894 , C0 , n65891 , n65892 , n65893 );
buf ( n65895 , n65894 );
buf ( n65896 , n65895 );
buf ( n65897 , n31655 );
buf ( n65898 , n30987 );
not ( n65899 , n43755 );
and ( n65900 , n65899 , n43309 );
xor ( n65901 , n43761 , n43767 );
and ( n65902 , n65901 , n43755 );
or ( n65903 , n65900 , n65902 );
and ( n65904 , n65903 , n43774 );
not ( n65905 , n44663 );
and ( n65906 , n65905 , n44221 );
xor ( n65907 , n44669 , n44675 );
and ( n65908 , n65907 , n44663 );
or ( n65909 , n65906 , n65908 );
and ( n65910 , n65909 , n44682 );
buf ( n65911 , RI15b451e0_223);
and ( n65912 , n65911 , n44695 );
or ( n65913 , n65904 , n65910 , n65912 );
buf ( n65914 , n65913 );
buf ( n65915 , n65914 );
buf ( n65916 , n30987 );
buf ( n65917 , n31655 );
not ( n65918 , n36587 );
and ( n65919 , n65918 , n35700 );
xor ( n65920 , n36591 , n36091 );
and ( n65921 , n65920 , n36587 );
or ( n65922 , n65919 , n65921 );
and ( n65923 , n65922 , n36596 );
not ( n65924 , n37485 );
and ( n65925 , n65924 , n36615 );
xor ( n65926 , n37489 , n36993 );
and ( n65927 , n65926 , n37485 );
or ( n65928 , n65925 , n65927 );
and ( n65929 , n65928 , n37494 );
and ( n65930 , n41840 , n37506 );
or ( n65931 , n65923 , n65929 , n65930 );
buf ( n65932 , n65931 );
buf ( n65933 , n65932 );
not ( n65934 , n38443 );
and ( n65935 , n65934 , n37963 );
xor ( n65936 , n53484 , n53485 );
and ( n65937 , n65936 , n38443 );
or ( n65938 , n65935 , n65937 );
and ( n65939 , n65938 , n38450 );
not ( n65940 , n39339 );
and ( n65941 , n65940 , n38863 );
xor ( n65942 , n53540 , n53541 );
and ( n65943 , n65942 , n39339 );
or ( n65944 , n65941 , n65943 );
and ( n65945 , n65944 , n39346 );
and ( n65946 , n40200 , n39359 );
or ( n65947 , n65939 , n65945 , n65946 );
buf ( n65948 , n65947 );
buf ( n65949 , n65948 );
buf ( n65950 , n30987 );
buf ( n65951 , n31655 );
and ( n65952 , n41284 , n32500 );
not ( n65953 , n35211 );
and ( n65954 , n65953 , n37573 );
buf ( n65955 , n65954 );
and ( n65956 , n65955 , n32421 );
not ( n65957 , n35245 );
and ( n65958 , n65957 , n37573 );
buf ( n65959 , n65958 );
and ( n65960 , n65959 , n32419 );
not ( n65961 , n35278 );
and ( n65962 , n65961 , n37573 );
not ( n65963 , n35295 );
and ( n65964 , n65963 , n47284 );
xor ( n65965 , n37573 , n49529 );
and ( n65966 , n65965 , n35295 );
or ( n65967 , n65964 , n65966 );
and ( n65968 , n65967 , n35278 );
or ( n65969 , n65962 , n65968 );
and ( n65970 , n65969 , n32417 );
not ( n65971 , n35331 );
and ( n65972 , n65971 , n37573 );
not ( n65973 , n35294 );
not ( n65974 , n45995 );
and ( n65975 , n65974 , n47284 );
xor ( n65976 , n49602 , n49615 );
and ( n65977 , n65976 , n45995 );
or ( n65978 , n65975 , n65977 );
and ( n65979 , n65973 , n65978 );
and ( n65980 , n65965 , n35294 );
or ( n65981 , n65979 , n65980 );
and ( n65982 , n65981 , n35331 );
or ( n65983 , n65972 , n65982 );
and ( n65984 , n65983 , n32415 );
and ( n65985 , n37573 , n35354 );
or ( n65986 , n65956 , n65960 , n65970 , n65984 , n65985 );
and ( n65987 , n65986 , n32456 );
not ( n65988 , n32475 );
not ( n65989 , n46060 );
and ( n65990 , n65989 , n41315 );
xor ( n65991 , n49693 , n49709 );
and ( n65992 , n65991 , n46060 );
or ( n65993 , n65990 , n65992 );
and ( n65994 , n65988 , n65993 );
and ( n65995 , n37573 , n32475 );
or ( n65996 , n65994 , n65995 );
and ( n65997 , n65996 , n32486 );
buf ( n65998 , n32489 );
and ( n65999 , n37573 , n35367 );
or ( n66000 , C0 , n65952 , n65987 , n65997 , n65998 , n65999 );
buf ( n66001 , n66000 );
buf ( n66002 , n66001 );
buf ( n66003 , n30987 );
not ( n66004 , n48765 );
and ( n66005 , n66004 , n33212 );
and ( n66006 , n49022 , n48765 );
or ( n66007 , n66005 , n66006 );
and ( n66008 , n66007 , n33180 );
not ( n66009 , n49054 );
and ( n66010 , n66009 , n33212 );
and ( n66011 , n49264 , n49054 );
or ( n66012 , n66010 , n66011 );
and ( n66013 , n66012 , n33178 );
and ( n66014 , n33212 , n49774 );
or ( n66015 , n66008 , n66013 , n66014 );
and ( n66016 , n66015 , n33208 );
and ( n66017 , n33275 , n33375 );
not ( n66018 , n32968 );
and ( n66019 , n66018 , n33275 );
and ( n66020 , n33216 , n59702 );
and ( n66021 , n33215 , n66020 );
and ( n66022 , n33214 , n66021 );
and ( n66023 , n33213 , n66022 );
xor ( n66024 , n33212 , n66023 );
and ( n66025 , n66024 , n32968 );
or ( n66026 , n66019 , n66025 );
and ( n66027 , n66026 , n33370 );
and ( n66028 , n32975 , n35056 );
and ( n66029 , n33212 , n49794 );
or ( n66030 , C0 , n66016 , n66017 , n66027 , n66028 , n66029 );
buf ( n66031 , n66030 );
buf ( n66032 , n66031 );
buf ( n66033 , n30987 );
buf ( n66034 , n31655 );
not ( n66035 , n35542 );
and ( n66036 , n66035 , n41861 );
and ( n66037 , n52964 , n35542 );
or ( n66038 , n66036 , n66037 );
buf ( n66039 , n66038 );
buf ( n66040 , n66039 );
buf ( n66041 , n31655 );
buf ( n66042 , RI15b52548_674);
and ( n66043 , n66042 , n31645 );
not ( n66044 , n45274 );
and ( n66045 , n66044 , n54960 );
buf ( n66046 , n66045 );
and ( n66047 , n66046 , n31373 );
not ( n66048 , n45280 );
and ( n66049 , n66048 , n54960 );
not ( n66050 , n45766 );
and ( n66051 , n66050 , n45541 );
xor ( n66052 , n45777 , n45779 );
and ( n66053 , n66052 , n45766 );
or ( n66054 , n66051 , n66053 );
and ( n66055 , n66054 , n45280 );
or ( n66056 , n66049 , n66055 );
and ( n66057 , n66056 , n31468 );
and ( n66058 , n54960 , n45802 );
or ( n66059 , n66047 , n66057 , n66058 );
and ( n66060 , n66059 , n31557 );
and ( n66061 , n54960 , n45808 );
or ( n66062 , C0 , n66043 , n66060 , n66061 );
buf ( n66063 , n66062 );
buf ( n66064 , n66063 );
not ( n66065 , n40163 );
and ( n66066 , n66065 , n31869 );
not ( n66067 , n54629 );
and ( n66068 , n66067 , n31869 );
and ( n66069 , n32218 , n54629 );
or ( n66070 , n66068 , n66069 );
and ( n66071 , n66070 , n40163 );
or ( n66072 , n66066 , n66071 );
and ( n66073 , n66072 , n32498 );
not ( n66074 , n54637 );
not ( n66075 , n54629 );
and ( n66076 , n66075 , n31869 );
and ( n66077 , n42255 , n54629 );
or ( n66078 , n66076 , n66077 );
and ( n66079 , n66074 , n66078 );
and ( n66080 , n42255 , n54637 );
or ( n66081 , n66079 , n66080 );
and ( n66082 , n66081 , n32473 );
not ( n66083 , n32475 );
not ( n66084 , n54637 );
not ( n66085 , n54629 );
and ( n66086 , n66085 , n31869 );
and ( n66087 , n42255 , n54629 );
or ( n66088 , n66086 , n66087 );
and ( n66089 , n66084 , n66088 );
and ( n66090 , n42255 , n54637 );
or ( n66091 , n66089 , n66090 );
and ( n66092 , n66083 , n66091 );
not ( n66093 , n54657 );
not ( n66094 , n54659 );
and ( n66095 , n66094 , n66091 );
and ( n66096 , n42283 , n54659 );
or ( n66097 , n66095 , n66096 );
and ( n66098 , n66093 , n66097 );
and ( n66099 , n42291 , n54657 );
or ( n66100 , n66098 , n66099 );
and ( n66101 , n66100 , n32475 );
or ( n66102 , n66092 , n66101 );
and ( n66103 , n66102 , n32486 );
and ( n66104 , n31869 , n41278 );
or ( n66105 , C0 , n66073 , n66082 , n66103 , n66104 );
buf ( n66106 , n66105 );
buf ( n66107 , n66106 );
buf ( n66108 , n30987 );
buf ( n66109 , n31655 );
buf ( n66110 , n31655 );
not ( n66111 , n34150 );
and ( n66112 , n66111 , n32637 );
not ( n66113 , n56413 );
and ( n66114 , n66113 , n32637 );
and ( n66115 , n32655 , n56413 );
or ( n66116 , n66114 , n66115 );
and ( n66117 , n66116 , n34150 );
or ( n66118 , n66112 , n66117 );
and ( n66119 , n66118 , n33381 );
not ( n66120 , n56421 );
not ( n66121 , n56413 );
and ( n66122 , n66121 , n32637 );
and ( n66123 , n56044 , n56413 );
or ( n66124 , n66122 , n66123 );
and ( n66125 , n66120 , n66124 );
and ( n66126 , n56044 , n56421 );
or ( n66127 , n66125 , n66126 );
and ( n66128 , n66127 , n33375 );
not ( n66129 , n32968 );
not ( n66130 , n56421 );
not ( n66131 , n56413 );
and ( n66132 , n66131 , n32637 );
and ( n66133 , n56044 , n56413 );
or ( n66134 , n66132 , n66133 );
and ( n66135 , n66130 , n66134 );
and ( n66136 , n56044 , n56421 );
or ( n66137 , n66135 , n66136 );
and ( n66138 , n66129 , n66137 );
not ( n66139 , n56441 );
not ( n66140 , n56443 );
and ( n66141 , n66140 , n66137 );
and ( n66142 , n56068 , n56443 );
or ( n66143 , n66141 , n66142 );
and ( n66144 , n66139 , n66143 );
and ( n66145 , n56076 , n56441 );
or ( n66146 , n66144 , n66145 );
and ( n66147 , n66146 , n32968 );
or ( n66148 , n66138 , n66147 );
and ( n66149 , n66148 , n33370 );
and ( n66150 , n32637 , n35062 );
or ( n66151 , C0 , n66119 , n66128 , n66149 , n66150 );
buf ( n66152 , n66151 );
buf ( n66153 , n66152 );
not ( n66154 , n34150 );
and ( n66155 , n66154 , n32530 );
buf ( n66156 , n66155 );
and ( n66157 , n66156 , n33381 );
not ( n66158 , n56687 );
not ( n66159 , n56464 );
and ( n66160 , n66159 , n32530 );
buf ( n66161 , n66160 );
and ( n66162 , n66158 , n66161 );
buf ( n66163 , n66162 );
and ( n66164 , n66163 , n33379 );
and ( n66165 , n32530 , n56699 );
or ( n66166 , C0 , n66157 , n66164 , C0 , C0 , n66165 );
buf ( n66167 , n66166 );
buf ( n66168 , n66167 );
buf ( n66169 , n31655 );
buf ( n66170 , n30987 );
buf ( n66171 , n30987 );
not ( n66172 , n50828 );
not ( n66173 , n50834 );
and ( n66174 , n66173 , n40639 );
and ( n66175 , n64906 , n50834 );
or ( n66176 , n66174 , n66175 );
and ( n66177 , n66172 , n66176 );
buf ( n66178 , RI15b60030_1141);
and ( n66179 , n66178 , n50828 );
or ( n66180 , n66177 , n66179 );
buf ( n66181 , n66180 );
buf ( n66182 , n66181 );
buf ( n66183 , n31655 );
buf ( n66184 , n30987 );
buf ( n66185 , n30987 );
buf ( n66186 , n31655 );
xor ( n66187 , n33093 , n58387 );
and ( n66188 , n66187 , n33201 );
not ( n66189 , n41576 );
and ( n66190 , n66189 , n33093 );
and ( n66191 , n64891 , n41576 );
or ( n66192 , n66190 , n66191 );
and ( n66193 , n66192 , n33189 );
and ( n66194 , n33093 , n41592 );
or ( n66195 , n66188 , n66193 , n66194 );
and ( n66196 , n66195 , n33208 );
and ( n66197 , n33093 , n39805 );
or ( n66198 , C0 , n66196 , n66197 );
buf ( n66199 , n66198 );
buf ( n66200 , n66199 );
buf ( n66201 , n31655 );
buf ( n66202 , n30987 );
and ( n66203 , n33222 , n32528 );
not ( n66204 , n32598 );
and ( n66205 , n66204 , n32985 );
buf ( n66206 , n66205 );
and ( n66207 , n66206 , n32890 );
not ( n66208 , n32919 );
and ( n66209 , n66208 , n32985 );
buf ( n66210 , n66209 );
and ( n66211 , n66210 , n32924 );
not ( n66212 , n32953 );
and ( n66213 , n66212 , n32985 );
not ( n66214 , n32971 );
and ( n66215 , n66214 , n33095 );
xor ( n66216 , n32985 , n33020 );
and ( n66217 , n66216 , n32971 );
or ( n66218 , n66215 , n66217 );
and ( n66219 , n66218 , n32953 );
or ( n66220 , n66213 , n66219 );
and ( n66221 , n66220 , n33038 );
not ( n66222 , n33067 );
and ( n66223 , n66222 , n32985 );
not ( n66224 , n32970 );
not ( n66225 , n33071 );
and ( n66226 , n66225 , n33095 );
xor ( n66227 , n33096 , n33152 );
and ( n66228 , n66227 , n33071 );
or ( n66229 , n66226 , n66228 );
and ( n66230 , n66224 , n66229 );
and ( n66231 , n66216 , n32970 );
or ( n66232 , n66230 , n66231 );
and ( n66233 , n66232 , n33067 );
or ( n66234 , n66223 , n66233 );
and ( n66235 , n66234 , n33172 );
and ( n66236 , n32985 , n33204 );
or ( n66237 , n66207 , n66211 , n66221 , n66235 , n66236 );
and ( n66238 , n66237 , n33208 );
not ( n66239 , n32968 );
not ( n66240 , n33270 );
and ( n66241 , n66240 , n33295 );
xor ( n66242 , n33296 , n33352 );
and ( n66243 , n66242 , n33270 );
or ( n66244 , n66241 , n66243 );
and ( n66245 , n66239 , n66244 );
and ( n66246 , n32985 , n32968 );
or ( n66247 , n66245 , n66246 );
and ( n66248 , n66247 , n33370 );
buf ( n66249 , n35056 );
and ( n66250 , n32985 , n33382 );
or ( n66251 , C0 , n66203 , n66238 , n66248 , n66249 , n66250 );
buf ( n66252 , n66251 );
buf ( n66253 , n66252 );
buf ( n66254 , n30987 );
buf ( n66255 , n31655 );
not ( n66256 , n31728 );
and ( n66257 , n66256 , n46028 );
and ( n66258 , n61912 , n31728 );
or ( n66259 , n66257 , n66258 );
and ( n66260 , n66259 , n32253 );
not ( n66261 , n32283 );
and ( n66262 , n66261 , n46028 );
and ( n66263 , n61923 , n32283 );
or ( n66264 , n66262 , n66263 );
and ( n66265 , n66264 , n32398 );
and ( n66266 , n46028 , n32436 );
or ( n66267 , n66260 , n66265 , n66266 );
and ( n66268 , n66267 , n32456 );
and ( n66269 , n49673 , n32473 );
not ( n66270 , n32475 );
and ( n66271 , n66270 , n49673 );
xor ( n66272 , n46028 , n47758 );
and ( n66273 , n66272 , n32475 );
or ( n66274 , n66271 , n66273 );
and ( n66275 , n66274 , n32486 );
and ( n66276 , n37553 , n32489 );
and ( n66277 , n46028 , n32501 );
or ( n66278 , C0 , n66268 , n66269 , n66275 , n66276 , n66277 );
buf ( n66279 , n66278 );
buf ( n66280 , n66279 );
buf ( n66281 , n31655 );
buf ( n66282 , n31655 );
buf ( n66283 , n30987 );
xor ( n66284 , n47285 , n47297 );
and ( n66285 , n66284 , n32433 );
not ( n66286 , n47331 );
and ( n66287 , n66286 , n47285 );
and ( n66288 , n32036 , n47357 );
and ( n66289 , n32038 , n47359 );
and ( n66290 , n32040 , n47361 );
and ( n66291 , n32042 , n47363 );
and ( n66292 , n32044 , n47365 );
and ( n66293 , n32046 , n47367 );
and ( n66294 , n32048 , n47369 );
and ( n66295 , n32050 , n47371 );
and ( n66296 , n32052 , n47373 );
and ( n66297 , n32054 , n47375 );
and ( n66298 , n32056 , n47377 );
and ( n66299 , n32058 , n47379 );
and ( n66300 , n32060 , n47381 );
and ( n66301 , n32062 , n47383 );
and ( n66302 , n32064 , n47385 );
and ( n66303 , n32066 , n47387 );
or ( n66304 , n66288 , n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , n66301 , n66302 , n66303 );
and ( n66305 , n66304 , n47331 );
or ( n66306 , n66287 , n66305 );
and ( n66307 , n66306 , n32413 );
and ( n66308 , n47285 , n47402 );
or ( n66309 , n66285 , n66307 , n66308 );
and ( n66310 , n66309 , n32456 );
and ( n66311 , n47285 , n47409 );
or ( n66312 , C0 , n66310 , n66311 );
buf ( n66313 , n66312 );
buf ( n66314 , n66313 );
not ( n66315 , n35542 );
and ( n66316 , n66315 , n41855 );
buf ( n66317 , RI15b457f8_236);
and ( n66318 , n66317 , n35542 );
or ( n66319 , n66316 , n66318 );
buf ( n66320 , n66319 );
buf ( n66321 , n66320 );
not ( n66322 , n46356 );
and ( n66323 , n66322 , n31126 );
not ( n66324 , n49427 );
and ( n66325 , n66324 , n31126 );
and ( n66326 , n31138 , n49427 );
or ( n66327 , n66325 , n66326 );
and ( n66328 , n66327 , n46356 );
or ( n66329 , n66323 , n66328 );
and ( n66330 , n66329 , n31649 );
not ( n66331 , n49435 );
not ( n66332 , n49427 );
and ( n66333 , n66332 , n31126 );
and ( n66334 , n56920 , n49427 );
or ( n66335 , n66333 , n66334 );
and ( n66336 , n66331 , n66335 );
and ( n66337 , n56920 , n49435 );
or ( n66338 , n66336 , n66337 );
and ( n66339 , n66338 , n31643 );
not ( n66340 , n31452 );
not ( n66341 , n49435 );
not ( n66342 , n49427 );
and ( n66343 , n66342 , n31126 );
and ( n66344 , n56920 , n49427 );
or ( n66345 , n66343 , n66344 );
and ( n66346 , n66341 , n66345 );
and ( n66347 , n56920 , n49435 );
or ( n66348 , n66346 , n66347 );
and ( n66349 , n66340 , n66348 );
not ( n66350 , n49460 );
not ( n66351 , n49462 );
and ( n66352 , n66351 , n66348 );
and ( n66353 , n56946 , n49462 );
or ( n66354 , n66352 , n66353 );
and ( n66355 , n66350 , n66354 );
and ( n66356 , n56954 , n49460 );
or ( n66357 , n66355 , n66356 );
and ( n66358 , n66357 , n31452 );
or ( n66359 , n66349 , n66358 );
and ( n66360 , n66359 , n31638 );
and ( n66361 , n31126 , n47277 );
or ( n66362 , C0 , n66330 , n66339 , n66360 , n66361 );
buf ( n66363 , n66362 );
buf ( n66364 , n66363 );
not ( n66365 , n34150 );
and ( n66366 , n66365 , n32634 );
not ( n66367 , n56836 );
and ( n66368 , n66367 , n32634 );
and ( n66369 , n32655 , n56836 );
or ( n66370 , n66368 , n66369 );
and ( n66371 , n66370 , n34150 );
or ( n66372 , n66366 , n66371 );
and ( n66373 , n66372 , n33381 );
not ( n66374 , n56844 );
not ( n66375 , n56836 );
and ( n66376 , n66375 , n32634 );
and ( n66377 , n56044 , n56836 );
or ( n66378 , n66376 , n66377 );
and ( n66379 , n66374 , n66378 );
and ( n66380 , n56044 , n56844 );
or ( n66381 , n66379 , n66380 );
and ( n66382 , n66381 , n33375 );
not ( n66383 , n32968 );
not ( n66384 , n56844 );
not ( n66385 , n56836 );
and ( n66386 , n66385 , n32634 );
and ( n66387 , n56044 , n56836 );
or ( n66388 , n66386 , n66387 );
and ( n66389 , n66384 , n66388 );
and ( n66390 , n56044 , n56844 );
or ( n66391 , n66389 , n66390 );
and ( n66392 , n66383 , n66391 );
not ( n66393 , n56864 );
not ( n66394 , n56866 );
and ( n66395 , n66394 , n66391 );
and ( n66396 , n56068 , n56866 );
or ( n66397 , n66395 , n66396 );
and ( n66398 , n66393 , n66397 );
and ( n66399 , n56076 , n56864 );
or ( n66400 , n66398 , n66399 );
and ( n66401 , n66400 , n32968 );
or ( n66402 , n66392 , n66401 );
and ( n66403 , n66402 , n33370 );
and ( n66404 , n32634 , n35062 );
or ( n66405 , C0 , n66373 , n66382 , n66403 , n66404 );
buf ( n66406 , n66405 );
buf ( n66407 , n66406 );
buf ( n66408 , n31655 );
buf ( n66409 , n31655 );
not ( n66410 , n35542 );
and ( n66411 , n66410 , n41842 );
and ( n66412 , n65911 , n35542 );
or ( n66413 , n66411 , n66412 );
buf ( n66414 , n66413 );
buf ( n66415 , n66414 );
buf ( n66416 , n30987 );
buf ( n66417 , n30987 );
buf ( n66418 , n30987 );
buf ( n66419 , n31655 );
buf ( n66420 , n31655 );
buf ( n66421 , n30987 );
buf ( n66422 , n42734 );
buf ( n66423 , n66422 );
and ( n66424 , n66423 , n42771 );
buf ( n66425 , n42734 );
buf ( n66426 , n42810 );
or ( n66427 , C0 , n66425 , C0 , C0 , n66426 );
and ( n66428 , n66427 , n42806 );
buf ( n66429 , n42734 );
nor ( n66430 , n42721 , n42728 , n42733 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n66431 , n66430 );
buf ( n66432 , n42810 );
or ( n66433 , C0 , n66429 , C0 , n66431 , n66432 );
and ( n66434 , n66433 , n42842 );
or ( n66435 , C0 , n66424 , n66428 , n66434 );
buf ( n66436 , n66435 );
buf ( n66437 , n66436 );
and ( n66438 , n31774 , n40163 );
buf ( n66439 , n66438 );
and ( n66440 , n66439 , n32498 );
and ( n66441 , n55718 , n32496 );
and ( n66442 , n47355 , n50275 );
not ( n66443 , n50278 );
and ( n66444 , n66443 , n31662 );
and ( n66445 , n47355 , n50278 );
or ( n66446 , n66444 , n66445 );
and ( n66447 , n66446 , n32421 );
not ( n66448 , n50002 );
and ( n66449 , n66448 , n31662 );
and ( n66450 , n47351 , n50002 );
or ( n66451 , n66449 , n66450 );
and ( n66452 , n66451 , n32419 );
not ( n66453 , n50289 );
and ( n66454 , n66453 , n31662 );
and ( n66455 , n47355 , n50289 );
or ( n66456 , n66454 , n66455 );
and ( n66457 , n66456 , n32417 );
not ( n66458 , n50008 );
and ( n66459 , n66458 , n31662 );
and ( n66460 , n47355 , n50008 );
or ( n66461 , n66459 , n66460 );
and ( n66462 , n66461 , n32415 );
not ( n66463 , n47331 );
and ( n66464 , n66463 , n31662 );
or ( n66465 , n31666 , n64621 );
xor ( n66466 , n31662 , n66465 );
not ( n66467 , n66466 );
buf ( n66468 , n66467 );
buf ( n66469 , n66468 );
not ( n66470 , n66469 );
and ( n66471 , n66470 , n47331 );
or ( n66472 , n66464 , n66471 );
and ( n66473 , n66472 , n32413 );
not ( n66474 , n50067 );
and ( n66475 , n66474 , n31662 );
and ( n66476 , n66470 , n50067 );
or ( n66477 , n66475 , n66476 );
and ( n66478 , n66477 , n32411 );
and ( n66479 , n31662 , n63978 );
and ( n66480 , n31774 , n50334 );
or ( n66481 , n66442 , n66447 , n66452 , n66457 , n66462 , n66473 , n66478 , n66479 , n66480 );
and ( n66482 , n66481 , n32456 );
and ( n66483 , n31662 , n63983 );
or ( n66484 , C0 , n66440 , n66441 , n66482 , n66483 );
buf ( n66485 , n66484 );
buf ( n66486 , n66485 );
buf ( n66487 , n31655 );
not ( n66488 , n36587 );
and ( n66489 , n66488 , n36294 );
xor ( n66490 , n50183 , n50204 );
and ( n66491 , n66490 , n36587 );
or ( n66492 , n66489 , n66491 );
and ( n66493 , n66492 , n36596 );
not ( n66494 , n37485 );
and ( n66495 , n66494 , n37196 );
xor ( n66496 , n50233 , n50254 );
and ( n66497 , n66496 , n37485 );
or ( n66498 , n66495 , n66497 );
and ( n66499 , n66498 , n37494 );
and ( n66500 , n41851 , n37506 );
or ( n66501 , n66493 , n66499 , n66500 );
buf ( n66502 , n66501 );
buf ( n66503 , n66502 );
buf ( n66504 , n30987 );
not ( n66505 , n36587 );
and ( n66506 , n66505 , n36158 );
xor ( n66507 , n50191 , n50196 );
and ( n66508 , n66507 , n36587 );
or ( n66509 , n66506 , n66508 );
and ( n66510 , n66509 , n36596 );
not ( n66511 , n37485 );
and ( n66512 , n66511 , n37060 );
xor ( n66513 , n50241 , n50246 );
and ( n66514 , n66513 , n37485 );
or ( n66515 , n66512 , n66514 );
and ( n66516 , n66515 , n37494 );
and ( n66517 , n41843 , n37506 );
or ( n66518 , n66510 , n66516 , n66517 );
buf ( n66519 , n66518 );
buf ( n66520 , n66519 );
buf ( n66521 , n30987 );
buf ( n66522 , RI15b60990_1161);
and ( n66523 , n66522 , n48531 );
and ( n66524 , n50824 , n39359 );
or ( n66525 , n66523 , n66524 );
buf ( n66526 , n66525 );
buf ( n66527 , n66526 );
buf ( n66528 , n31655 );
buf ( n66529 , n31655 );
buf ( n66530 , n31655 );
buf ( n66531 , n30987 );
not ( n66532 , n33419 );
and ( n66533 , n66532 , n31571 );
xor ( n66534 , n33465 , n33700 );
and ( n66535 , n66534 , n33419 );
or ( n66536 , n66533 , n66535 );
and ( n66537 , n66536 , n31529 );
not ( n66538 , n33734 );
and ( n66539 , n66538 , n31571 );
not ( n66540 , n33533 );
xor ( n66541 , n33758 , n33818 );
and ( n66542 , n66540 , n66541 );
xnor ( n66543 , n33843 , n33920 );
and ( n66544 , n66543 , n33533 );
or ( n66545 , n66542 , n66544 );
and ( n66546 , n66545 , n33734 );
or ( n66547 , n66539 , n66546 );
and ( n66548 , n66547 , n31527 );
and ( n66549 , n31571 , n33942 );
or ( n66550 , n66537 , n66548 , n66549 );
and ( n66551 , n66550 , n31557 );
and ( n66552 , n35497 , n31643 );
not ( n66553 , n31452 );
and ( n66554 , n66553 , n35497 );
xor ( n66555 , n31571 , n33966 );
and ( n66556 , n66555 , n31452 );
or ( n66557 , n66554 , n66556 );
and ( n66558 , n66557 , n31638 );
and ( n66559 , n35396 , n33973 );
and ( n66560 , n31571 , n33978 );
or ( n66561 , C0 , n66551 , n66552 , n66558 , n66559 , n66560 );
buf ( n66562 , n66561 );
buf ( n66563 , n66562 );
and ( n66564 , n31573 , n31007 );
not ( n66565 , n31077 );
and ( n66566 , n66565 , n35398 );
buf ( n66567 , n66566 );
and ( n66568 , n66567 , n31373 );
not ( n66569 , n31402 );
and ( n66570 , n66569 , n35398 );
buf ( n66571 , n66570 );
and ( n66572 , n66571 , n31408 );
not ( n66573 , n31437 );
and ( n66574 , n66573 , n35398 );
not ( n66575 , n31455 );
and ( n66576 , n66575 , n35447 );
xor ( n66577 , n35398 , n35399 );
and ( n66578 , n66577 , n31455 );
or ( n66579 , n66576 , n66578 );
and ( n66580 , n66579 , n31437 );
or ( n66581 , n66574 , n66580 );
and ( n66582 , n66581 , n31468 );
not ( n66583 , n31497 );
and ( n66584 , n66583 , n35398 );
not ( n66585 , n31454 );
not ( n66586 , n31501 );
and ( n66587 , n66586 , n35447 );
xor ( n66588 , n35448 , n35449 );
and ( n66589 , n66588 , n31501 );
or ( n66590 , n66587 , n66589 );
and ( n66591 , n66585 , n66590 );
and ( n66592 , n66577 , n31454 );
or ( n66593 , n66591 , n66592 );
and ( n66594 , n66593 , n31497 );
or ( n66595 , n66584 , n66594 );
and ( n66596 , n66595 , n31521 );
and ( n66597 , n35398 , n31553 );
or ( n66598 , n66568 , n66572 , n66582 , n66596 , n66597 );
and ( n66599 , n66598 , n31557 );
not ( n66600 , n31452 );
not ( n66601 , n31619 );
and ( n66602 , n66601 , n35501 );
xor ( n66603 , n35502 , n35503 );
and ( n66604 , n66603 , n31619 );
or ( n66605 , n66602 , n66604 );
and ( n66606 , n66600 , n66605 );
and ( n66607 , n35398 , n31452 );
or ( n66608 , n66606 , n66607 );
and ( n66609 , n66608 , n31638 );
buf ( n66610 , n33973 );
and ( n66611 , n35398 , n31650 );
or ( n66612 , C0 , n66564 , n66599 , n66609 , n66610 , n66611 );
buf ( n66613 , n66612 );
buf ( n66614 , n66613 );
buf ( n66615 , n30987 );
buf ( n66616 , n31655 );
not ( n66617 , n46356 );
and ( n66618 , n66617 , n31226 );
not ( n66619 , n64746 );
and ( n66620 , n66619 , n31226 );
and ( n66621 , n31238 , n64746 );
or ( n66622 , n66620 , n66621 );
and ( n66623 , n66622 , n46356 );
or ( n66624 , n66618 , n66623 );
and ( n66625 , n66624 , n31649 );
not ( n66626 , n64754 );
not ( n66627 , n64746 );
and ( n66628 , n66627 , n31226 );
and ( n66629 , n49901 , n64746 );
or ( n66630 , n66628 , n66629 );
and ( n66631 , n66626 , n66630 );
and ( n66632 , n49901 , n64754 );
or ( n66633 , n66631 , n66632 );
and ( n66634 , n66633 , n31643 );
not ( n66635 , n31452 );
not ( n66636 , n64754 );
not ( n66637 , n64746 );
and ( n66638 , n66637 , n31226 );
and ( n66639 , n49901 , n64746 );
or ( n66640 , n66638 , n66639 );
and ( n66641 , n66636 , n66640 );
and ( n66642 , n49901 , n64754 );
or ( n66643 , n66641 , n66642 );
and ( n66644 , n66635 , n66643 );
not ( n66645 , n64774 );
not ( n66646 , n64776 );
and ( n66647 , n66646 , n66643 );
and ( n66648 , n49925 , n64776 );
or ( n66649 , n66647 , n66648 );
and ( n66650 , n66645 , n66649 );
and ( n66651 , n49933 , n64774 );
or ( n66652 , n66650 , n66651 );
and ( n66653 , n66652 , n31452 );
or ( n66654 , n66644 , n66653 );
and ( n66655 , n66654 , n31638 );
and ( n66656 , n31226 , n47277 );
or ( n66657 , C0 , n66625 , n66634 , n66655 , n66656 );
buf ( n66658 , n66657 );
buf ( n66659 , n66658 );
buf ( n66660 , n31655 );
xor ( n66661 , n50965 , n64714 );
and ( n66662 , n66661 , n32431 );
not ( n66663 , n50002 );
and ( n66664 , n66663 , n50965 );
and ( n66665 , n40620 , n50002 );
or ( n66666 , n66664 , n66665 );
and ( n66667 , n66666 , n32419 );
not ( n66668 , n50008 );
and ( n66669 , n66668 , n50965 );
not ( n66670 , n51594 );
and ( n66671 , n66670 , n51482 );
xor ( n66672 , n51598 , n51608 );
and ( n66673 , n66672 , n51594 );
or ( n66674 , n66671 , n66673 );
and ( n66675 , n66674 , n50008 );
or ( n66676 , n66669 , n66675 );
and ( n66677 , n66676 , n32415 );
not ( n66678 , n50067 );
and ( n66679 , n66678 , n50965 );
and ( n66680 , n31861 , n60510 );
and ( n66681 , n31863 , n60512 );
and ( n66682 , n31865 , n60514 );
and ( n66683 , n31867 , n60516 );
and ( n66684 , n31869 , n60518 );
and ( n66685 , n31871 , n60520 );
and ( n66686 , n31873 , n60522 );
and ( n66687 , n31875 , n60524 );
and ( n66688 , n31877 , n60526 );
and ( n66689 , n31879 , n60528 );
and ( n66690 , n31881 , n60530 );
and ( n66691 , n31883 , n60532 );
and ( n66692 , n31885 , n60534 );
and ( n66693 , n31887 , n60536 );
and ( n66694 , n31889 , n60538 );
and ( n66695 , n31891 , n60540 );
or ( n66696 , n66680 , n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , n66695 );
and ( n66697 , n66696 , n50067 );
or ( n66698 , n66679 , n66697 );
and ( n66699 , n66698 , n32411 );
and ( n66700 , n50965 , n50098 );
or ( n66701 , n66662 , n66667 , n66677 , n66699 , n66700 );
and ( n66702 , n66701 , n32456 );
and ( n66703 , n50965 , n47409 );
or ( n66704 , C0 , n66702 , n66703 );
buf ( n66705 , n66704 );
buf ( n66706 , n66705 );
buf ( n66707 , n30987 );
buf ( n66708 , n31655 );
not ( n66709 , n50828 );
not ( n66710 , n50834 );
and ( n66711 , n66710 , n40455 );
buf ( n66712 , RI15b53ad8_720);
and ( n66713 , n66712 , n50834 );
or ( n66714 , n66711 , n66713 );
and ( n66715 , n66709 , n66714 );
buf ( n66716 , RI15b5ff40_1139);
and ( n66717 , n66716 , n50828 );
or ( n66718 , n66715 , n66717 );
buf ( n66719 , n66718 );
buf ( n66720 , n66719 );
buf ( n66721 , n30987 );
buf ( n66722 , n30987 );
xor ( n66723 , n33089 , n58389 );
and ( n66724 , n66723 , n33201 );
not ( n66725 , n41576 );
and ( n66726 , n66725 , n33089 );
and ( n66727 , n32824 , n55215 );
and ( n66728 , n32826 , n55217 );
and ( n66729 , n32828 , n55219 );
and ( n66730 , n32830 , n55221 );
and ( n66731 , n32832 , n55223 );
and ( n66732 , n32834 , n55225 );
and ( n66733 , n32836 , n55227 );
and ( n66734 , n32838 , n55229 );
and ( n66735 , n32840 , n55231 );
and ( n66736 , n32842 , n55233 );
and ( n66737 , n32844 , n55235 );
and ( n66738 , n32846 , n55237 );
and ( n66739 , n32848 , n55239 );
and ( n66740 , n32850 , n55241 );
and ( n66741 , n32852 , n55243 );
and ( n66742 , n32854 , n55245 );
or ( n66743 , n66727 , n66728 , n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , n66741 , n66742 );
and ( n66744 , n66743 , n41576 );
or ( n66745 , n66726 , n66744 );
and ( n66746 , n66745 , n33189 );
and ( n66747 , n33089 , n41592 );
or ( n66748 , n66724 , n66746 , n66747 );
and ( n66749 , n66748 , n33208 );
and ( n66750 , n33089 , n39805 );
or ( n66751 , C0 , n66749 , n66750 );
buf ( n66752 , n66751 );
buf ( n66753 , n66752 );
buf ( n66754 , n31655 );
buf ( n66755 , n31655 );
not ( n66756 , n43755 );
and ( n66757 , n66756 , n43428 );
xor ( n66758 , n50499 , n50506 );
and ( n66759 , n66758 , n43755 );
or ( n66760 , n66757 , n66759 );
and ( n66761 , n66760 , n43774 );
not ( n66762 , n44663 );
and ( n66763 , n66762 , n44340 );
xor ( n66764 , n50517 , n50524 );
and ( n66765 , n66764 , n44663 );
or ( n66766 , n66763 , n66765 );
and ( n66767 , n66766 , n44682 );
buf ( n66768 , RI15b45528_230);
and ( n66769 , n66768 , n44695 );
or ( n66770 , n66761 , n66767 , n66769 );
buf ( n66771 , n66770 );
buf ( n66772 , n66771 );
buf ( n66773 , n30987 );
buf ( n66774 , n30987 );
buf ( n66775 , n31655 );
buf ( n66776 , n31655 );
buf ( n66777 , n30987 );
not ( n66778 , n48765 );
and ( n66779 , n66778 , n33240 );
xor ( n66780 , n48942 , n48959 );
xor ( n66781 , n66780 , n48979 );
and ( n66782 , n66781 , n48765 );
or ( n66783 , n66779 , n66782 );
and ( n66784 , n66783 , n33180 );
not ( n66785 , n49054 );
and ( n66786 , n66785 , n33240 );
not ( n66787 , n48845 );
xor ( n66788 , n49091 , n48959 );
xor ( n66789 , n66788 , n49093 );
and ( n66790 , n66787 , n66789 );
xor ( n66791 , n49212 , n49214 );
xor ( n66792 , n66791 , n49219 );
and ( n66793 , n66792 , n48845 );
or ( n66794 , n66790 , n66793 );
and ( n66795 , n66794 , n49054 );
or ( n66796 , n66786 , n66795 );
and ( n66797 , n66796 , n33178 );
and ( n66798 , n33240 , n49774 );
or ( n66799 , n66784 , n66797 , n66798 );
and ( n66800 , n66799 , n33208 );
and ( n66801 , n33331 , n33375 );
not ( n66802 , n32968 );
and ( n66803 , n66802 , n33331 );
and ( n66804 , n33240 , n32968 );
or ( n66805 , n66803 , n66804 );
and ( n66806 , n66805 , n33370 );
and ( n66807 , n33003 , n35056 );
and ( n66808 , n33240 , n49794 );
or ( n66809 , C0 , n66800 , n66801 , n66806 , n66807 , n66808 );
buf ( n66810 , n66809 );
buf ( n66811 , n66810 );
buf ( n66812 , n30987 );
not ( n66813 , n50828 );
not ( n66814 , n50834 );
and ( n66815 , n66814 , n40321 );
and ( n66816 , n56336 , n50834 );
or ( n66817 , n66815 , n66816 );
and ( n66818 , n66813 , n66817 );
buf ( n66819 , RI15b5fa18_1128);
and ( n66820 , n66819 , n50828 );
or ( n66821 , n66818 , n66820 );
buf ( n66822 , n66821 );
buf ( n66823 , n66822 );
buf ( n66824 , n31655 );
buf ( n66825 , n31655 );
xor ( n66826 , n49595 , n60308 );
and ( n66827 , n66826 , n32433 );
not ( n66828 , n47331 );
and ( n66829 , n66828 , n49595 );
and ( n66830 , n63386 , n47331 );
or ( n66831 , n66829 , n66830 );
and ( n66832 , n66831 , n32413 );
and ( n66833 , n49595 , n47402 );
or ( n66834 , n66827 , n66832 , n66833 );
and ( n66835 , n66834 , n32456 );
and ( n66836 , n49595 , n47409 );
or ( n66837 , C0 , n66835 , n66836 );
buf ( n66838 , n66837 );
buf ( n66839 , n66838 );
buf ( n66840 , n30987 );
buf ( n66841 , n50814 );
not ( n66842 , n46356 );
and ( n66843 , n66842 , n31232 );
not ( n66844 , n47423 );
and ( n66845 , n66844 , n31232 );
and ( n66846 , n31238 , n47423 );
or ( n66847 , n66845 , n66846 );
and ( n66848 , n66847 , n46356 );
or ( n66849 , n66843 , n66848 );
and ( n66850 , n66849 , n31649 );
not ( n66851 , n47431 );
not ( n66852 , n47423 );
and ( n66853 , n66852 , n31232 );
and ( n66854 , n49901 , n47423 );
or ( n66855 , n66853 , n66854 );
and ( n66856 , n66851 , n66855 );
and ( n66857 , n49901 , n47431 );
or ( n66858 , n66856 , n66857 );
and ( n66859 , n66858 , n31643 );
not ( n66860 , n31452 );
not ( n66861 , n47431 );
not ( n66862 , n47423 );
and ( n66863 , n66862 , n31232 );
and ( n66864 , n49901 , n47423 );
or ( n66865 , n66863 , n66864 );
and ( n66866 , n66861 , n66865 );
and ( n66867 , n49901 , n47431 );
or ( n66868 , n66866 , n66867 );
and ( n66869 , n66860 , n66868 );
not ( n66870 , n47466 );
not ( n66871 , n47468 );
and ( n66872 , n66871 , n66868 );
and ( n66873 , n49925 , n47468 );
or ( n66874 , n66872 , n66873 );
and ( n66875 , n66870 , n66874 );
and ( n66876 , n49933 , n47466 );
or ( n66877 , n66875 , n66876 );
and ( n66878 , n66877 , n31452 );
or ( n66879 , n66869 , n66878 );
and ( n66880 , n66879 , n31638 );
and ( n66881 , n31232 , n47277 );
or ( n66882 , C0 , n66850 , n66859 , n66880 , n66881 );
buf ( n66883 , n66882 );
buf ( n66884 , n66883 );
buf ( n66885 , n31655 );
not ( n66886 , n50828 );
not ( n66887 , n50834 );
and ( n66888 , n66887 , n40232 );
buf ( n66889 , RI15b53358_704);
and ( n66890 , n66889 , n50834 );
or ( n66891 , n66888 , n66890 );
and ( n66892 , n66886 , n66891 );
buf ( n66893 , RI15b5f7c0_1123);
and ( n66894 , n66893 , n50828 );
or ( n66895 , n66892 , n66894 );
buf ( n66896 , n66895 );
buf ( n66897 , n66896 );
buf ( n66898 , n30987 );
buf ( n66899 , n31655 );
not ( n66900 , n48765 );
and ( n66901 , n66900 , n33235 );
xor ( n66902 , n48847 , n48864 );
xor ( n66903 , n66902 , n48994 );
and ( n66904 , n66903 , n48765 );
or ( n66905 , n66901 , n66904 );
and ( n66906 , n66905 , n33180 );
not ( n66907 , n49054 );
and ( n66908 , n66907 , n33235 );
not ( n66909 , n48845 );
xor ( n66910 , n49081 , n48864 );
xor ( n66911 , n66910 , n49108 );
and ( n66912 , n66909 , n66911 );
xor ( n66913 , n49192 , n49194 );
xor ( n66914 , n66913 , n49234 );
and ( n66915 , n66914 , n48845 );
or ( n66916 , n66912 , n66915 );
and ( n66917 , n66916 , n49054 );
or ( n66918 , n66908 , n66917 );
and ( n66919 , n66918 , n33178 );
and ( n66920 , n33235 , n49774 );
or ( n66921 , n66906 , n66919 , n66920 );
and ( n66922 , n66921 , n33208 );
and ( n66923 , n33321 , n33375 );
not ( n66924 , n32968 );
and ( n66925 , n66924 , n33321 );
xor ( n66926 , n33235 , n49783 );
and ( n66927 , n66926 , n32968 );
or ( n66928 , n66925 , n66927 );
and ( n66929 , n66928 , n33370 );
and ( n66930 , n32998 , n35056 );
and ( n66931 , n33235 , n49794 );
or ( n66932 , C0 , n66922 , n66923 , n66929 , n66930 , n66931 );
buf ( n66933 , n66932 );
buf ( n66934 , n66933 );
buf ( n66935 , n31655 );
buf ( n66936 , n30987 );
buf ( n66937 , n31655 );
buf ( n66938 , n30987 );
not ( n66939 , n32953 );
buf ( n66940 , RI15b462c0_259);
and ( n66941 , n66939 , n66940 );
not ( n66942 , n54581 );
and ( n66943 , n66942 , n54424 );
xor ( n66944 , n64017 , n64024 );
and ( n66945 , n66944 , n54581 );
or ( n66946 , n66943 , n66945 );
and ( n66947 , n66946 , n32953 );
or ( n66948 , n66941 , n66947 );
and ( n66949 , n66948 , n33038 );
not ( n66950 , n48660 );
and ( n66951 , n66950 , n66940 );
and ( n66952 , n55184 , n48660 );
or ( n66953 , n66951 , n66952 );
and ( n66954 , n66953 , n33172 );
and ( n66955 , n66940 , n39795 );
or ( n66956 , n66949 , n66954 , n66955 );
and ( n66957 , n66956 , n33208 );
and ( n66958 , n66940 , n39805 );
or ( n66959 , C0 , n66957 , n66958 );
buf ( n66960 , n66959 );
buf ( n66961 , n66960 );
buf ( n66962 , n30987 );
buf ( n66963 , n31655 );
buf ( n66964 , n30987 );
buf ( n66965 , n31655 );
buf ( n66966 , n31655 );
buf ( n66967 , n30987 );
and ( n66968 , n31570 , n31007 );
not ( n66969 , n31077 );
and ( n66970 , n66969 , n33972 );
buf ( n66971 , n66970 );
and ( n66972 , n66971 , n31373 );
not ( n66973 , n31402 );
and ( n66974 , n66973 , n33972 );
buf ( n66975 , n66974 );
and ( n66976 , n66975 , n31408 );
not ( n66977 , n31437 );
and ( n66978 , n66977 , n33972 );
not ( n66979 , n31455 );
and ( n66980 , n66979 , n35441 );
xor ( n66981 , n33972 , n35402 );
and ( n66982 , n66981 , n31455 );
or ( n66983 , n66980 , n66982 );
and ( n66984 , n66983 , n31437 );
or ( n66985 , n66978 , n66984 );
and ( n66986 , n66985 , n31468 );
not ( n66987 , n31497 );
and ( n66988 , n66987 , n33972 );
not ( n66989 , n31454 );
not ( n66990 , n31501 );
and ( n66991 , n66990 , n35441 );
xor ( n66992 , n35442 , n35452 );
and ( n66993 , n66992 , n31501 );
or ( n66994 , n66991 , n66993 );
and ( n66995 , n66989 , n66994 );
and ( n66996 , n66981 , n31454 );
or ( n66997 , n66995 , n66996 );
and ( n66998 , n66997 , n31497 );
or ( n66999 , n66988 , n66998 );
and ( n67000 , n66999 , n31521 );
and ( n67001 , n33972 , n31553 );
or ( n67002 , n66972 , n66976 , n66986 , n67000 , n67001 );
and ( n67003 , n67002 , n31557 );
not ( n67004 , n31452 );
not ( n67005 , n31619 );
and ( n67006 , n67005 , n33946 );
xor ( n67007 , n35496 , n35506 );
and ( n67008 , n67007 , n31619 );
or ( n67009 , n67006 , n67008 );
and ( n67010 , n67004 , n67009 );
and ( n67011 , n33972 , n31452 );
or ( n67012 , n67010 , n67011 );
and ( n67013 , n67012 , n31638 );
and ( n67014 , n33972 , n31650 );
or ( n67015 , C0 , n66968 , n67003 , n67013 , C0 , n67014 );
buf ( n67016 , n67015 );
buf ( n67017 , n67016 );
not ( n67018 , n33419 );
and ( n67019 , n67018 , n31574 );
and ( n67020 , n63269 , n33419 );
or ( n67021 , n67019 , n67020 );
and ( n67022 , n67021 , n31529 );
not ( n67023 , n33734 );
and ( n67024 , n67023 , n31574 );
and ( n67025 , n63280 , n33734 );
or ( n67026 , n67024 , n67025 );
and ( n67027 , n67026 , n31527 );
and ( n67028 , n31574 , n33942 );
or ( n67029 , n67022 , n67027 , n67028 );
and ( n67030 , n67029 , n31557 );
and ( n67031 , n34092 , n31643 );
not ( n67032 , n31452 );
and ( n67033 , n67032 , n34092 );
xor ( n67034 , n31574 , n33963 );
and ( n67035 , n67034 , n31452 );
or ( n67036 , n67033 , n67035 );
and ( n67037 , n67036 , n31638 );
and ( n67038 , n33986 , n33973 );
and ( n67039 , n31574 , n33978 );
or ( n67040 , C0 , n67030 , n67031 , n67037 , n67038 , n67039 );
buf ( n67041 , n67040 );
buf ( n67042 , n67041 );
buf ( n67043 , n31655 );
buf ( n67044 , n30987 );
not ( n67045 , n34150 );
and ( n67046 , n67045 , n32681 );
not ( n67047 , n56093 );
and ( n67048 , n67047 , n32681 );
and ( n67049 , n32689 , n56093 );
or ( n67050 , n67048 , n67049 );
and ( n67051 , n67050 , n34150 );
or ( n67052 , n67046 , n67051 );
and ( n67053 , n67052 , n33381 );
not ( n67054 , n56101 );
not ( n67055 , n56093 );
and ( n67056 , n67055 , n32681 );
and ( n67057 , n50682 , n56093 );
or ( n67058 , n67056 , n67057 );
and ( n67059 , n67054 , n67058 );
and ( n67060 , n50682 , n56101 );
or ( n67061 , n67059 , n67060 );
and ( n67062 , n67061 , n33375 );
not ( n67063 , n32968 );
not ( n67064 , n56101 );
not ( n67065 , n56093 );
and ( n67066 , n67065 , n32681 );
and ( n67067 , n50682 , n56093 );
or ( n67068 , n67066 , n67067 );
and ( n67069 , n67064 , n67068 );
and ( n67070 , n50682 , n56101 );
or ( n67071 , n67069 , n67070 );
and ( n67072 , n67063 , n67071 );
not ( n67073 , n56121 );
not ( n67074 , n56123 );
and ( n67075 , n67074 , n67071 );
and ( n67076 , n50706 , n56123 );
or ( n67077 , n67075 , n67076 );
and ( n67078 , n67073 , n67077 );
and ( n67079 , n50714 , n56121 );
or ( n67080 , n67078 , n67079 );
and ( n67081 , n67080 , n32968 );
or ( n67082 , n67072 , n67081 );
and ( n67083 , n67082 , n33370 );
and ( n67084 , n32681 , n35062 );
or ( n67085 , C0 , n67053 , n67062 , n67083 , n67084 );
buf ( n67086 , n67085 );
buf ( n67087 , n67086 );
not ( n67088 , n34150 );
and ( n67089 , n67088 , n32852 );
not ( n67090 , n56140 );
and ( n67091 , n67090 , n32852 );
and ( n67092 , n32856 , n56140 );
or ( n67093 , n67091 , n67092 );
and ( n67094 , n67093 , n34150 );
or ( n67095 , n67089 , n67094 );
and ( n67096 , n67095 , n33381 );
not ( n67097 , n56148 );
not ( n67098 , n56140 );
and ( n67099 , n67098 , n32852 );
and ( n67100 , n48160 , n56140 );
or ( n67101 , n67099 , n67100 );
and ( n67102 , n67097 , n67101 );
and ( n67103 , n48160 , n56148 );
or ( n67104 , n67102 , n67103 );
and ( n67105 , n67104 , n33375 );
not ( n67106 , n32968 );
not ( n67107 , n56148 );
not ( n67108 , n56140 );
and ( n67109 , n67108 , n32852 );
and ( n67110 , n48160 , n56140 );
or ( n67111 , n67109 , n67110 );
and ( n67112 , n67107 , n67111 );
and ( n67113 , n48160 , n56148 );
or ( n67114 , n67112 , n67113 );
and ( n67115 , n67106 , n67114 );
not ( n67116 , n56168 );
not ( n67117 , n56170 );
and ( n67118 , n67117 , n67114 );
and ( n67119 , n48186 , n56170 );
or ( n67120 , n67118 , n67119 );
and ( n67121 , n67116 , n67120 );
and ( n67122 , n48196 , n56168 );
or ( n67123 , n67121 , n67122 );
and ( n67124 , n67123 , n32968 );
or ( n67125 , n67115 , n67124 );
and ( n67126 , n67125 , n33370 );
and ( n67127 , n32852 , n35062 );
or ( n67128 , C0 , n67096 , n67105 , n67126 , n67127 );
buf ( n67129 , n67128 );
buf ( n67130 , n67129 );
buf ( n67131 , n30987 );
buf ( n67132 , n31655 );
not ( n67133 , n40163 );
and ( n67134 , n67133 , n32036 );
not ( n67135 , n56988 );
and ( n67136 , n67135 , n32036 );
and ( n67137 , n32130 , n56988 );
or ( n67138 , n67136 , n67137 );
and ( n67139 , n67138 , n40163 );
or ( n67140 , n67134 , n67139 );
and ( n67141 , n67140 , n32498 );
not ( n67142 , n56996 );
not ( n67143 , n56988 );
and ( n67144 , n67143 , n32036 );
and ( n67145 , n45833 , n56988 );
or ( n67146 , n67144 , n67145 );
and ( n67147 , n67142 , n67146 );
and ( n67148 , n45833 , n56996 );
or ( n67149 , n67147 , n67148 );
and ( n67150 , n67149 , n32473 );
not ( n67151 , n32475 );
not ( n67152 , n56996 );
not ( n67153 , n56988 );
and ( n67154 , n67153 , n32036 );
and ( n67155 , n45833 , n56988 );
or ( n67156 , n67154 , n67155 );
and ( n67157 , n67152 , n67156 );
and ( n67158 , n45833 , n56996 );
or ( n67159 , n67157 , n67158 );
and ( n67160 , n67151 , n67159 );
not ( n67161 , n57016 );
not ( n67162 , n57018 );
and ( n67163 , n67162 , n67159 );
and ( n67164 , n45857 , n57018 );
or ( n67165 , n67163 , n67164 );
and ( n67166 , n67161 , n67165 );
and ( n67167 , n45865 , n57016 );
or ( n67168 , n67166 , n67167 );
and ( n67169 , n67168 , n32475 );
or ( n67170 , n67160 , n67169 );
and ( n67171 , n67170 , n32486 );
and ( n67172 , n32036 , n41278 );
or ( n67173 , C0 , n67141 , n67150 , n67171 , n67172 );
buf ( n67174 , n67173 );
buf ( n67175 , n67174 );
buf ( n67176 , n30987 );
buf ( n67177 , n31655 );
not ( n67178 , n31437 );
and ( n67179 , n67178 , n65187 );
and ( n67180 , n65196 , n31437 );
or ( n67181 , n67179 , n67180 );
and ( n67182 , n67181 , n31468 );
not ( n67183 , n41837 );
and ( n67184 , n67183 , n65187 );
not ( n67185 , n42124 );
and ( n67186 , n67185 , n41976 );
xor ( n67187 , n42129 , n42141 );
and ( n67188 , n67187 , n42124 );
or ( n67189 , n67186 , n67188 );
and ( n67190 , n67189 , n41837 );
or ( n67191 , n67184 , n67190 );
and ( n67192 , n67191 , n31521 );
and ( n67193 , n65187 , n42158 );
or ( n67194 , n67182 , n67192 , n67193 );
and ( n67195 , n67194 , n31557 );
and ( n67196 , n65187 , n40154 );
or ( n67197 , C0 , n67195 , n67196 );
buf ( n67198 , n67197 );
buf ( n67199 , n67198 );
buf ( n67200 , n30987 );
xor ( n67201 , n41678 , n44781 );
and ( n67202 , n67201 , n31548 );
not ( n67203 , n44807 );
and ( n67204 , n67203 , n41678 );
and ( n67205 , n41966 , n44807 );
or ( n67206 , n67204 , n67205 );
and ( n67207 , n67206 , n31408 );
not ( n67208 , n44817 );
and ( n67209 , n67208 , n41678 );
not ( n67210 , n41835 );
and ( n67211 , n67210 , n65187 );
and ( n67212 , n67189 , n41835 );
or ( n67213 , n67211 , n67212 );
and ( n67214 , n67213 , n44817 );
or ( n67215 , n67209 , n67214 );
and ( n67216 , n67215 , n31521 );
not ( n67217 , n45059 );
and ( n67218 , n67217 , n41678 );
and ( n67219 , n33552 , n45059 );
or ( n67220 , n67218 , n67219 );
and ( n67221 , n67220 , n31536 );
and ( n67222 , n41678 , n45148 );
or ( n67223 , n67202 , n67207 , n67216 , n67221 , n67222 );
and ( n67224 , n67223 , n31557 );
and ( n67225 , n41678 , n40154 );
or ( n67226 , C0 , n67224 , n67225 );
buf ( n67227 , n67226 );
buf ( n67228 , n67227 );
buf ( n67229 , n31655 );
not ( n67230 , n40163 );
and ( n67231 , n67230 , n31982 );
not ( n67232 , n50540 );
and ( n67233 , n67232 , n31982 );
and ( n67234 , n32165 , n50540 );
or ( n67235 , n67233 , n67234 );
and ( n67236 , n67235 , n40163 );
or ( n67237 , n67231 , n67236 );
and ( n67238 , n67237 , n32498 );
not ( n67239 , n50548 );
not ( n67240 , n50540 );
and ( n67241 , n67240 , n31982 );
and ( n67242 , n59005 , n50540 );
or ( n67243 , n67241 , n67242 );
and ( n67244 , n67239 , n67243 );
and ( n67245 , n59005 , n50548 );
or ( n67246 , n67244 , n67245 );
and ( n67247 , n67246 , n32473 );
not ( n67248 , n32475 );
not ( n67249 , n50548 );
not ( n67250 , n50540 );
and ( n67251 , n67250 , n31982 );
and ( n67252 , n59005 , n50540 );
or ( n67253 , n67251 , n67252 );
and ( n67254 , n67249 , n67253 );
and ( n67255 , n59005 , n50548 );
or ( n67256 , n67254 , n67255 );
and ( n67257 , n67248 , n67256 );
not ( n67258 , n50568 );
not ( n67259 , n50570 );
and ( n67260 , n67259 , n67256 );
and ( n67261 , n59029 , n50570 );
or ( n67262 , n67260 , n67261 );
and ( n67263 , n67258 , n67262 );
and ( n67264 , n59037 , n50568 );
or ( n67265 , n67263 , n67264 );
and ( n67266 , n67265 , n32475 );
or ( n67267 , n67257 , n67266 );
and ( n67268 , n67267 , n32486 );
and ( n67269 , n31982 , n41278 );
or ( n67270 , C0 , n67238 , n67247 , n67268 , n67269 );
buf ( n67271 , n67270 );
buf ( n67272 , n67271 );
buf ( n67273 , n30987 );
buf ( n67274 , n31655 );
buf ( n67275 , n53756 );
buf ( n67276 , n53758 );
nor ( n67277 , n53743 , n53750 , n53755 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n67278 , n67277 );
or ( n67279 , n67275 , n67276 , n67278 , C0 );
and ( n67280 , n67279 , n53793 );
buf ( n67281 , n53756 );
buf ( n67282 , n53758 );
buf ( n67283 , n67277 );
or ( n67284 , C0 , n67281 , n67282 , n67283 , C0 );
and ( n67285 , n67284 , n53828 );
buf ( n67286 , n53756 );
buf ( n67287 , n53758 );
buf ( n67288 , n67277 );
or ( n67289 , C0 , n67286 , n67287 , n67288 , C0 );
and ( n67290 , n67289 , n53864 );
or ( n67291 , C0 , n67280 , n67285 , n67290 );
buf ( n67292 , n67291 );
buf ( n67293 , n67292 );
buf ( n67294 , n30987 );
buf ( n67295 , n30987 );
not ( n67296 , n40163 );
and ( n67297 , n67296 , n31978 );
not ( n67298 , n52903 );
and ( n67299 , n67298 , n31978 );
and ( n67300 , n32165 , n52903 );
or ( n67301 , n67299 , n67300 );
and ( n67302 , n67301 , n40163 );
or ( n67303 , n67297 , n67302 );
and ( n67304 , n67303 , n32498 );
not ( n67305 , n52911 );
not ( n67306 , n52903 );
and ( n67307 , n67306 , n31978 );
and ( n67308 , n59005 , n52903 );
or ( n67309 , n67307 , n67308 );
and ( n67310 , n67305 , n67309 );
and ( n67311 , n59005 , n52911 );
or ( n67312 , n67310 , n67311 );
and ( n67313 , n67312 , n32473 );
not ( n67314 , n32475 );
not ( n67315 , n52911 );
not ( n67316 , n52903 );
and ( n67317 , n67316 , n31978 );
and ( n67318 , n59005 , n52903 );
or ( n67319 , n67317 , n67318 );
and ( n67320 , n67315 , n67319 );
and ( n67321 , n59005 , n52911 );
or ( n67322 , n67320 , n67321 );
and ( n67323 , n67314 , n67322 );
not ( n67324 , n52931 );
not ( n67325 , n52933 );
and ( n67326 , n67325 , n67322 );
and ( n67327 , n59029 , n52933 );
or ( n67328 , n67326 , n67327 );
and ( n67329 , n67324 , n67328 );
and ( n67330 , n59037 , n52931 );
or ( n67331 , n67329 , n67330 );
and ( n67332 , n67331 , n32475 );
or ( n67333 , n67323 , n67332 );
and ( n67334 , n67333 , n32486 );
and ( n67335 , n31978 , n41278 );
or ( n67336 , C0 , n67304 , n67313 , n67334 , n67335 );
buf ( n67337 , n67336 );
buf ( n67338 , n67337 );
buf ( n67339 , n31655 );
buf ( n67340 , n30987 );
not ( n67341 , n43755 );
and ( n67342 , n67341 , n43377 );
xor ( n67343 , n50502 , n50503 );
and ( n67344 , n67343 , n43755 );
or ( n67345 , n67342 , n67344 );
and ( n67346 , n67345 , n43774 );
not ( n67347 , n44663 );
and ( n67348 , n67347 , n44289 );
xor ( n67349 , n50520 , n50521 );
and ( n67350 , n67349 , n44663 );
or ( n67351 , n67348 , n67350 );
and ( n67352 , n67351 , n44682 );
buf ( n67353 , RI15b453c0_227);
and ( n67354 , n67353 , n44695 );
or ( n67355 , n67346 , n67352 , n67354 );
buf ( n67356 , n67355 );
buf ( n67357 , n67356 );
buf ( n67358 , n30987 );
buf ( n67359 , n31655 );
and ( n67360 , n50959 , n65295 );
xor ( n67361 , n50957 , n67360 );
and ( n67362 , n67361 , n32431 );
not ( n67363 , n50002 );
and ( n67364 , n67363 , n50957 );
and ( n67365 , n40592 , n50002 );
or ( n67366 , n67364 , n67365 );
and ( n67367 , n67366 , n32419 );
not ( n67368 , n50008 );
and ( n67369 , n67368 , n50957 );
not ( n67370 , n51594 );
and ( n67371 , n67370 , n51530 );
xor ( n67372 , n59228 , n59233 );
and ( n67373 , n67372 , n51594 );
or ( n67374 , n67371 , n67373 );
and ( n67375 , n67374 , n50008 );
or ( n67376 , n67369 , n67375 );
and ( n67377 , n67376 , n32415 );
not ( n67378 , n50067 );
and ( n67379 , n67378 , n50957 );
and ( n67380 , n60467 , n65310 );
xor ( n67381 , n60450 , n67380 );
and ( n67382 , n67381 , n50067 );
or ( n67383 , n67379 , n67382 );
and ( n67384 , n67383 , n32411 );
and ( n67385 , n50957 , n50098 );
or ( n67386 , n67362 , n67367 , n67377 , n67384 , n67385 );
and ( n67387 , n67386 , n32456 );
and ( n67388 , n50957 , n47409 );
or ( n67389 , C0 , n67387 , n67388 );
buf ( n67390 , n67389 );
buf ( n67391 , n67390 );
buf ( n67392 , n31655 );
not ( n67393 , n46356 );
and ( n67394 , n67393 , n31362 );
not ( n67395 , n56904 );
and ( n67396 , n67395 , n31362 );
and ( n67397 , n31372 , n56904 );
or ( n67398 , n67396 , n67397 );
and ( n67399 , n67398 , n46356 );
or ( n67400 , n67394 , n67399 );
and ( n67401 , n67400 , n31649 );
not ( n67402 , n56912 );
not ( n67403 , n56904 );
and ( n67404 , n67403 , n31362 );
and ( n67405 , n47849 , n56904 );
or ( n67406 , n67404 , n67405 );
and ( n67407 , n67402 , n67406 );
and ( n67408 , n47849 , n56912 );
or ( n67409 , n67407 , n67408 );
and ( n67410 , n67409 , n31643 );
not ( n67411 , n31452 );
not ( n67412 , n56912 );
not ( n67413 , n56904 );
and ( n67414 , n67413 , n31362 );
and ( n67415 , n47849 , n56904 );
or ( n67416 , n67414 , n67415 );
and ( n67417 , n67412 , n67416 );
and ( n67418 , n47849 , n56912 );
or ( n67419 , n67417 , n67418 );
and ( n67420 , n67411 , n67419 );
not ( n67421 , n56937 );
not ( n67422 , n56939 );
and ( n67423 , n67422 , n67419 );
and ( n67424 , n47877 , n56939 );
or ( n67425 , n67423 , n67424 );
and ( n67426 , n67421 , n67425 );
and ( n67427 , n47887 , n56937 );
or ( n67428 , n67426 , n67427 );
and ( n67429 , n67428 , n31452 );
or ( n67430 , n67420 , n67429 );
and ( n67431 , n67430 , n31638 );
and ( n67432 , n31362 , n47277 );
or ( n67433 , C0 , n67401 , n67410 , n67431 , n67432 );
buf ( n67434 , n67433 );
buf ( n67435 , n67434 );
buf ( n67436 , n31655 );
buf ( n67437 , n65459 );
buf ( n67438 , n30987 );
buf ( n67439 , n31655 );
not ( n67440 , n43755 );
and ( n67441 , n67440 , n43547 );
xor ( n67442 , n52310 , n52319 );
and ( n67443 , n67442 , n43755 );
or ( n67444 , n67441 , n67443 );
and ( n67445 , n67444 , n43774 );
not ( n67446 , n44663 );
and ( n67447 , n67446 , n44459 );
xor ( n67448 , n52348 , n52357 );
and ( n67449 , n67448 , n44663 );
or ( n67450 , n67447 , n67449 );
and ( n67451 , n67450 , n44682 );
buf ( n67452 , RI15b45870_237);
and ( n67453 , n67452 , n44695 );
or ( n67454 , n67445 , n67451 , n67453 );
buf ( n67455 , n67454 );
buf ( n67456 , n67455 );
buf ( n67457 , n30987 );
buf ( n67458 , n30987 );
buf ( n67459 , n31655 );
buf ( n67460 , n31655 );
buf ( n67461 , n31655 );
not ( n67462 , n34150 );
and ( n67463 , n67462 , n32665 );
not ( n67464 , n59105 );
and ( n67465 , n67464 , n32665 );
and ( n67466 , n32689 , n59105 );
or ( n67467 , n67465 , n67466 );
and ( n67468 , n67467 , n34150 );
or ( n67469 , n67463 , n67468 );
and ( n67470 , n67469 , n33381 );
not ( n67471 , n59113 );
not ( n67472 , n59105 );
and ( n67473 , n67472 , n32665 );
and ( n67474 , n50682 , n59105 );
or ( n67475 , n67473 , n67474 );
and ( n67476 , n67471 , n67475 );
and ( n67477 , n50682 , n59113 );
or ( n67478 , n67476 , n67477 );
and ( n67479 , n67478 , n33375 );
not ( n67480 , n32968 );
not ( n67481 , n59113 );
not ( n67482 , n59105 );
and ( n67483 , n67482 , n32665 );
and ( n67484 , n50682 , n59105 );
or ( n67485 , n67483 , n67484 );
and ( n67486 , n67481 , n67485 );
and ( n67487 , n50682 , n59113 );
or ( n67488 , n67486 , n67487 );
and ( n67489 , n67480 , n67488 );
not ( n67490 , n59133 );
not ( n67491 , n59135 );
and ( n67492 , n67491 , n67488 );
and ( n67493 , n50706 , n59135 );
or ( n67494 , n67492 , n67493 );
and ( n67495 , n67490 , n67494 );
and ( n67496 , n50714 , n59133 );
or ( n67497 , n67495 , n67496 );
and ( n67498 , n67497 , n32968 );
or ( n67499 , n67489 , n67498 );
and ( n67500 , n67499 , n33370 );
and ( n67501 , n32665 , n35062 );
or ( n67502 , C0 , n67470 , n67479 , n67500 , n67501 );
buf ( n67503 , n67502 );
buf ( n67504 , n67503 );
buf ( n67505 , n30987 );
buf ( n67506 , n30987 );
buf ( n67507 , n31655 );
buf ( n67508 , n30987 );
not ( n67509 , n32953 );
buf ( n67510 , RI15b46518_264);
and ( n67511 , n67509 , n67510 );
not ( n67512 , n54581 );
and ( n67513 , n67512 , n54509 );
xor ( n67514 , n54509 , n54340 );
and ( n67515 , n65079 , n65080 );
xor ( n67516 , n67514 , n67515 );
and ( n67517 , n67516 , n54581 );
or ( n67518 , n67513 , n67517 );
and ( n67519 , n67518 , n32953 );
or ( n67520 , n67511 , n67519 );
and ( n67521 , n67520 , n33038 );
not ( n67522 , n48660 );
and ( n67523 , n67522 , n67510 );
not ( n67524 , n55168 );
and ( n67525 , n67524 , n55116 );
xor ( n67526 , n55116 , n34193 );
and ( n67527 , n65091 , n65092 );
xor ( n67528 , n67526 , n67527 );
and ( n67529 , n67528 , n55168 );
or ( n67530 , n67525 , n67529 );
and ( n67531 , n67530 , n48660 );
or ( n67532 , n67523 , n67531 );
and ( n67533 , n67532 , n33172 );
and ( n67534 , n67510 , n39795 );
or ( n67535 , n67521 , n67533 , n67534 );
and ( n67536 , n67535 , n33208 );
and ( n67537 , n67510 , n39805 );
or ( n67538 , C0 , n67536 , n67537 );
buf ( n67539 , n67538 );
buf ( n67540 , n67539 );
buf ( n67541 , n30987 );
buf ( n67542 , n31655 );
buf ( n67543 , n30987 );
buf ( n67544 , n30987 );
buf ( n67545 , n31655 );
buf ( n67546 , RI15b47058_288);
buf ( n67547 , n67546 );
not ( n67548 , n34150 );
and ( n67549 , n67548 , n32873 );
not ( n67550 , n57038 );
and ( n67551 , n67550 , n32873 );
and ( n67552 , n32889 , n57038 );
or ( n67553 , n67551 , n67552 );
and ( n67554 , n67553 , n34150 );
or ( n67555 , n67549 , n67554 );
and ( n67556 , n67555 , n33381 );
not ( n67557 , n57046 );
not ( n67558 , n57038 );
and ( n67559 , n67558 , n32873 );
and ( n67560 , n52819 , n57038 );
or ( n67561 , n67559 , n67560 );
and ( n67562 , n67557 , n67561 );
and ( n67563 , n52819 , n57046 );
or ( n67564 , n67562 , n67563 );
and ( n67565 , n67564 , n33375 );
not ( n67566 , n32968 );
not ( n67567 , n57046 );
not ( n67568 , n57038 );
and ( n67569 , n67568 , n32873 );
and ( n67570 , n52819 , n57038 );
or ( n67571 , n67569 , n67570 );
and ( n67572 , n67567 , n67571 );
and ( n67573 , n52819 , n57046 );
or ( n67574 , n67572 , n67573 );
and ( n67575 , n67566 , n67574 );
not ( n67576 , n57066 );
not ( n67577 , n57068 );
and ( n67578 , n67577 , n67574 );
and ( n67579 , n52845 , n57068 );
or ( n67580 , n67578 , n67579 );
and ( n67581 , n67576 , n67580 );
and ( n67582 , n52855 , n57066 );
or ( n67583 , n67581 , n67582 );
and ( n67584 , n67583 , n32968 );
or ( n67585 , n67575 , n67584 );
and ( n67586 , n67585 , n33370 );
and ( n67587 , n32873 , n35062 );
or ( n67588 , C0 , n67556 , n67565 , n67586 , n67587 );
buf ( n67589 , n67588 );
buf ( n67590 , n67589 );
buf ( n67591 , n31655 );
buf ( n67592 , n31655 );
buf ( n67593 , n35213 );
not ( n67594 , n67593 );
buf ( n67595 , n67594 );
not ( n67596 , n67595 );
not ( n67597 , n37512 );
and ( n67598 , n67597 , n37514 );
not ( n67599 , n37514 );
not ( n67600 , n35213 );
xor ( n67601 , n67599 , n67600 );
and ( n67602 , n67601 , n37512 );
or ( n67603 , n67598 , n67602 );
not ( n67604 , n67603 );
buf ( n67605 , n67604 );
buf ( n67606 , n67605 );
not ( n67607 , n67606 );
or ( n67608 , n67596 , n67607 );
buf ( n67609 , n67608 );
buf ( n67610 , n67609 );
and ( n67611 , n67610 , n37512 );
not ( n67612 , n67611 );
and ( n67613 , n67612 , n67596 );
xor ( n67614 , n67596 , n37512 );
xor ( n67615 , n67614 , n37512 );
and ( n67616 , n67615 , n67611 );
or ( n67617 , n67613 , n67616 );
not ( n67618 , n67617 );
not ( n67619 , n67611 );
and ( n67620 , n67619 , n67607 );
xor ( n67621 , n67607 , n37512 );
and ( n67622 , n67614 , n37512 );
xor ( n67623 , n67621 , n67622 );
and ( n67624 , n67623 , n67611 );
or ( n67625 , n67620 , n67624 );
not ( n67626 , n67625 );
and ( n67627 , n67621 , n67622 );
buf ( n67628 , n67627 );
and ( n67629 , n67628 , n67611 );
buf ( n67630 , n67629 );
nor ( n67631 , n67618 , n67626 , n67630 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n67632 , n67631 );
buf ( n67633 , n67632 );
not ( n67634 , n32475 );
buf ( n67635 , RI15b60b70_1165);
buf ( n67636 , n67635 );
buf ( n67637 , n67635 );
buf ( n67638 , n67635 );
buf ( n67639 , n67635 );
buf ( n67640 , n67635 );
buf ( n67641 , n67635 );
buf ( n67642 , n67635 );
buf ( n67643 , n67635 );
buf ( n67644 , n67635 );
buf ( n67645 , n67635 );
buf ( n67646 , n67635 );
buf ( n67647 , n67635 );
buf ( n67648 , n67635 );
buf ( n67649 , n67635 );
buf ( n67650 , n67635 );
buf ( n67651 , n67635 );
buf ( n67652 , n67635 );
buf ( n67653 , n67635 );
buf ( n67654 , n67635 );
buf ( n67655 , n67635 );
buf ( n67656 , n67635 );
buf ( n67657 , n67635 );
buf ( n67658 , n67635 );
buf ( n67659 , n67635 );
buf ( n67660 , n67635 );
buf ( n67661 , n67635 );
buf ( n67662 , n67635 );
buf ( n67663 , n67635 );
buf ( n67664 , n67635 );
nor ( n67665 , n58110 , n67634 , n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , n67661 , n67662 , n67663 , n67664 );
and ( n67666 , n67633 , n67665 );
buf ( n67667 , n67631 );
nor ( n67668 , n67617 , n67625 , n67630 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n67669 , n67668 );
or ( n67670 , C0 , n67667 , C0 , C0 , n67669 );
not ( n67671 , n58110 );
buf ( n67672 , n67635 );
buf ( n67673 , n67635 );
buf ( n67674 , n67635 );
buf ( n67675 , n67635 );
buf ( n67676 , n67635 );
buf ( n67677 , n67635 );
buf ( n67678 , n67635 );
buf ( n67679 , n67635 );
buf ( n67680 , n67635 );
buf ( n67681 , n67635 );
buf ( n67682 , n67635 );
buf ( n67683 , n67635 );
buf ( n67684 , n67635 );
buf ( n67685 , n67635 );
buf ( n67686 , n67635 );
buf ( n67687 , n67635 );
buf ( n67688 , n67635 );
buf ( n67689 , n67635 );
buf ( n67690 , n67635 );
buf ( n67691 , n67635 );
buf ( n67692 , n67635 );
buf ( n67693 , n67635 );
buf ( n67694 , n67635 );
buf ( n67695 , n67635 );
buf ( n67696 , n67635 );
buf ( n67697 , n67635 );
buf ( n67698 , n67635 );
buf ( n67699 , n67635 );
buf ( n67700 , n67635 );
nor ( n67701 , n67671 , n32475 , n67635 , n67672 , n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , n67699 , n67700 );
and ( n67702 , n67670 , n67701 );
buf ( n67703 , n67631 );
nor ( n67704 , n67618 , n67625 , n67630 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n67705 , n67704 );
buf ( n67706 , n67668 );
or ( n67707 , C0 , n67703 , C0 , n67705 , n67706 );
buf ( n67708 , n67635 );
buf ( n67709 , n67635 );
buf ( n67710 , n67635 );
buf ( n67711 , n67635 );
buf ( n67712 , n67635 );
buf ( n67713 , n67635 );
buf ( n67714 , n67635 );
buf ( n67715 , n67635 );
buf ( n67716 , n67635 );
buf ( n67717 , n67635 );
buf ( n67718 , n67635 );
buf ( n67719 , n67635 );
buf ( n67720 , n67635 );
buf ( n67721 , n67635 );
buf ( n67722 , n67635 );
buf ( n67723 , n67635 );
buf ( n67724 , n67635 );
buf ( n67725 , n67635 );
buf ( n67726 , n67635 );
buf ( n67727 , n67635 );
buf ( n67728 , n67635 );
buf ( n67729 , n67635 );
buf ( n67730 , n67635 );
buf ( n67731 , n67635 );
buf ( n67732 , n67635 );
buf ( n67733 , n67635 );
buf ( n67734 , n67635 );
buf ( n67735 , n67635 );
buf ( n67736 , n67635 );
nor ( n67737 , n58110 , n32475 , n67635 , n67708 , n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , n67735 , n67736 );
and ( n67738 , n67707 , n67737 );
or ( n67739 , C0 , n67666 , n67702 , n67738 );
buf ( n67740 , n67739 );
buf ( n67741 , n67740 );
not ( n67742 , n46356 );
and ( n67743 , n67742 , n31354 );
not ( n67744 , n48214 );
and ( n67745 , n67744 , n31354 );
and ( n67746 , n31372 , n48214 );
or ( n67747 , n67745 , n67746 );
and ( n67748 , n67747 , n46356 );
or ( n67749 , n67743 , n67748 );
and ( n67750 , n67749 , n31649 );
not ( n67751 , n48223 );
not ( n67752 , n48214 );
and ( n67753 , n67752 , n31354 );
and ( n67754 , n47849 , n48214 );
or ( n67755 , n67753 , n67754 );
and ( n67756 , n67751 , n67755 );
and ( n67757 , n47849 , n48223 );
or ( n67758 , n67756 , n67757 );
and ( n67759 , n67758 , n31643 );
not ( n67760 , n31452 );
not ( n67761 , n48223 );
not ( n67762 , n48214 );
and ( n67763 , n67762 , n31354 );
and ( n67764 , n47849 , n48214 );
or ( n67765 , n67763 , n67764 );
and ( n67766 , n67761 , n67765 );
and ( n67767 , n47849 , n48223 );
or ( n67768 , n67766 , n67767 );
and ( n67769 , n67760 , n67768 );
not ( n67770 , n48244 );
not ( n67771 , n48247 );
and ( n67772 , n67771 , n67768 );
and ( n67773 , n47877 , n48247 );
or ( n67774 , n67772 , n67773 );
and ( n67775 , n67770 , n67774 );
and ( n67776 , n47887 , n48244 );
or ( n67777 , n67775 , n67776 );
and ( n67778 , n67777 , n31452 );
or ( n67779 , n67769 , n67778 );
and ( n67780 , n67779 , n31638 );
and ( n67781 , n31354 , n47277 );
or ( n67782 , C0 , n67750 , n67759 , n67780 , n67781 );
buf ( n67783 , n67782 );
buf ( n67784 , n67783 );
buf ( n67785 , n30987 );
buf ( n67786 , n31655 );
buf ( n67787 , n30987 );
buf ( n67788 , n31655 );
not ( n67789 , n38443 );
and ( n67790 , n67789 , n38354 );
xor ( n67791 , n53461 , n53508 );
and ( n67792 , n67791 , n38443 );
or ( n67793 , n67790 , n67792 );
and ( n67794 , n67793 , n38450 );
not ( n67795 , n39339 );
and ( n67796 , n67795 , n39254 );
xor ( n67797 , n53517 , n53564 );
and ( n67798 , n67797 , n39339 );
or ( n67799 , n67796 , n67798 );
and ( n67800 , n67799 , n39346 );
and ( n67801 , n40223 , n39359 );
or ( n67802 , n67794 , n67800 , n67801 );
buf ( n67803 , n67802 );
buf ( n67804 , n67803 );
and ( n67805 , n42405 , n48455 );
not ( n67806 , n48457 );
and ( n67807 , n67806 , n42378 );
and ( n67808 , n42405 , n48457 );
or ( n67809 , n67807 , n67808 );
and ( n67810 , n67809 , n31373 );
not ( n67811 , n44807 );
and ( n67812 , n67811 , n42378 );
and ( n67813 , n42405 , n44807 );
or ( n67814 , n67812 , n67813 );
and ( n67815 , n67814 , n31408 );
not ( n67816 , n48468 );
and ( n67817 , n67816 , n42378 );
and ( n67818 , n42405 , n48468 );
or ( n67819 , n67817 , n67818 );
and ( n67820 , n67819 , n31468 );
not ( n67821 , n44817 );
and ( n67822 , n67821 , n42378 );
and ( n67823 , n42405 , n44817 );
or ( n67824 , n67822 , n67823 );
and ( n67825 , n67824 , n31521 );
not ( n67826 , n39979 );
and ( n67827 , n67826 , n42378 );
and ( n67828 , n42386 , n39979 );
or ( n67829 , n67827 , n67828 );
and ( n67830 , n67829 , n31538 );
not ( n67831 , n45059 );
and ( n67832 , n67831 , n42378 );
and ( n67833 , n42386 , n45059 );
or ( n67834 , n67832 , n67833 );
and ( n67835 , n67834 , n31536 );
not ( n67836 , n33419 );
and ( n67837 , n67836 , n42378 );
xor ( n67838 , n42386 , n42389 );
and ( n67839 , n67838 , n33419 );
or ( n67840 , n67837 , n67839 );
and ( n67841 , n67840 , n31529 );
not ( n67842 , n33734 );
and ( n67843 , n67842 , n42378 );
not ( n67844 , n33533 );
xor ( n67845 , n42405 , n42408 );
and ( n67846 , n67844 , n67845 );
xnor ( n67847 , n42419 , n42422 );
and ( n67848 , n67847 , n33533 );
or ( n67849 , n67846 , n67848 );
and ( n67850 , n67849 , n33734 );
or ( n67851 , n67843 , n67850 );
and ( n67852 , n67851 , n31527 );
and ( n67853 , n42419 , n48513 );
or ( n67854 , n67805 , n67810 , n67815 , n67820 , n67825 , n67830 , n67835 , n67841 , n67852 , n67853 );
and ( n67855 , n67854 , n31557 );
and ( n67856 , n35394 , n33973 );
and ( n67857 , n42378 , n48524 );
or ( n67858 , C0 , n67855 , n67856 , n67857 );
buf ( n67859 , n67858 );
buf ( n67860 , n67859 );
not ( n67861 , n40163 );
and ( n67862 , n67861 , n31910 );
not ( n67863 , n52120 );
and ( n67864 , n67863 , n31910 );
and ( n67865 , n32200 , n52120 );
or ( n67866 , n67864 , n67865 );
and ( n67867 , n67866 , n40163 );
or ( n67868 , n67862 , n67867 );
and ( n67869 , n67868 , n32498 );
not ( n67870 , n52128 );
not ( n67871 , n52120 );
and ( n67872 , n67871 , n31910 );
and ( n67873 , n53243 , n52120 );
or ( n67874 , n67872 , n67873 );
and ( n67875 , n67870 , n67874 );
and ( n67876 , n53243 , n52128 );
or ( n67877 , n67875 , n67876 );
and ( n67878 , n67877 , n32473 );
not ( n67879 , n32475 );
not ( n67880 , n52128 );
not ( n67881 , n52120 );
and ( n67882 , n67881 , n31910 );
and ( n67883 , n53243 , n52120 );
or ( n67884 , n67882 , n67883 );
and ( n67885 , n67880 , n67884 );
and ( n67886 , n53243 , n52128 );
or ( n67887 , n67885 , n67886 );
and ( n67888 , n67879 , n67887 );
not ( n67889 , n52148 );
not ( n67890 , n52150 );
and ( n67891 , n67890 , n67887 );
and ( n67892 , n53269 , n52150 );
or ( n67893 , n67891 , n67892 );
and ( n67894 , n67889 , n67893 );
and ( n67895 , n53277 , n52148 );
or ( n67896 , n67894 , n67895 );
and ( n67897 , n67896 , n32475 );
or ( n67898 , n67888 , n67897 );
and ( n67899 , n67898 , n32486 );
and ( n67900 , n31910 , n41278 );
or ( n67901 , C0 , n67869 , n67878 , n67899 , n67900 );
buf ( n67902 , n67901 );
buf ( n67903 , n67902 );
buf ( n67904 , n31655 );
or ( n67905 , n37496 , n37494 );
or ( n67906 , n67905 , n37503 );
or ( n67907 , n67906 , n36596 );
or ( n67908 , n67907 , n37505 );
and ( n67909 , n53763 , n67908 );
buf ( n67910 , n67909 );
buf ( n67911 , n67910 );
buf ( n67912 , n30987 );
buf ( n67913 , n30987 );
buf ( n67914 , n31655 );
and ( n67915 , n33482 , n46356 );
buf ( n67916 , n67915 );
and ( n67917 , n67916 , n31649 );
and ( n67918 , n52594 , n31647 );
and ( n67919 , n63762 , n31557 );
and ( n67920 , n31026 , n61220 );
or ( n67921 , C0 , n67917 , n67918 , n67919 , n67920 );
buf ( n67922 , n67921 );
buf ( n67923 , n67922 );
not ( n67924 , n38443 );
and ( n67925 , n67924 , n38201 );
xor ( n67926 , n53470 , n53499 );
and ( n67927 , n67926 , n38443 );
or ( n67928 , n67925 , n67927 );
and ( n67929 , n67928 , n38450 );
not ( n67930 , n39339 );
and ( n67931 , n67930 , n39101 );
xor ( n67932 , n53526 , n53555 );
and ( n67933 , n67932 , n39339 );
or ( n67934 , n67931 , n67933 );
and ( n67935 , n67934 , n39346 );
and ( n67936 , n40214 , n39359 );
or ( n67937 , n67929 , n67935 , n67936 );
buf ( n67938 , n67937 );
buf ( n67939 , n67938 );
buf ( n67940 , n30987 );
not ( n67941 , n34150 );
and ( n67942 , n67941 , n32663 );
not ( n67943 , n59574 );
and ( n67944 , n67943 , n32663 );
and ( n67945 , n32689 , n59574 );
or ( n67946 , n67944 , n67945 );
and ( n67947 , n67946 , n34150 );
or ( n67948 , n67942 , n67947 );
and ( n67949 , n67948 , n33381 );
not ( n67950 , n59582 );
not ( n67951 , n59574 );
and ( n67952 , n67951 , n32663 );
and ( n67953 , n50682 , n59574 );
or ( n67954 , n67952 , n67953 );
and ( n67955 , n67950 , n67954 );
and ( n67956 , n50682 , n59582 );
or ( n67957 , n67955 , n67956 );
and ( n67958 , n67957 , n33375 );
not ( n67959 , n32968 );
not ( n67960 , n59582 );
not ( n67961 , n59574 );
and ( n67962 , n67961 , n32663 );
and ( n67963 , n50682 , n59574 );
or ( n67964 , n67962 , n67963 );
and ( n67965 , n67960 , n67964 );
and ( n67966 , n50682 , n59582 );
or ( n67967 , n67965 , n67966 );
and ( n67968 , n67959 , n67967 );
not ( n67969 , n59602 );
not ( n67970 , n59604 );
and ( n67971 , n67970 , n67967 );
and ( n67972 , n50706 , n59604 );
or ( n67973 , n67971 , n67972 );
and ( n67974 , n67969 , n67973 );
and ( n67975 , n50714 , n59602 );
or ( n67976 , n67974 , n67975 );
and ( n67977 , n67976 , n32968 );
or ( n67978 , n67968 , n67977 );
and ( n67979 , n67978 , n33370 );
and ( n67980 , n32663 , n35062 );
or ( n67981 , C0 , n67949 , n67958 , n67979 , n67980 );
buf ( n67982 , n67981 );
buf ( n67983 , n67982 );
buf ( n67984 , n31655 );
buf ( n67985 , n30987 );
buf ( n67986 , n30987 );
buf ( n67987 , n31655 );
buf ( n67988 , n30987 );
buf ( n67989 , n30987 );
buf ( n67990 , n31655 );
not ( n67991 , n34150 );
and ( n67992 , n67991 , n32702 );
not ( n67993 , n57872 );
and ( n67994 , n67993 , n32702 );
and ( n67995 , n32722 , n57872 );
or ( n67996 , n67994 , n67995 );
and ( n67997 , n67996 , n34150 );
or ( n67998 , n67992 , n67997 );
and ( n67999 , n67998 , n33381 );
not ( n68000 , n57880 );
not ( n68001 , n57872 );
and ( n68002 , n68001 , n32702 );
and ( n68003 , n42565 , n57872 );
or ( n68004 , n68002 , n68003 );
and ( n68005 , n68000 , n68004 );
and ( n68006 , n42565 , n57880 );
or ( n68007 , n68005 , n68006 );
and ( n68008 , n68007 , n33375 );
not ( n68009 , n32968 );
not ( n68010 , n57880 );
not ( n68011 , n57872 );
and ( n68012 , n68011 , n32702 );
and ( n68013 , n42565 , n57872 );
or ( n68014 , n68012 , n68013 );
and ( n68015 , n68010 , n68014 );
and ( n68016 , n42565 , n57880 );
or ( n68017 , n68015 , n68016 );
and ( n68018 , n68009 , n68017 );
not ( n68019 , n57900 );
not ( n68020 , n57902 );
and ( n68021 , n68020 , n68017 );
and ( n68022 , n42589 , n57902 );
or ( n68023 , n68021 , n68022 );
and ( n68024 , n68019 , n68023 );
and ( n68025 , n42597 , n57900 );
or ( n68026 , n68024 , n68025 );
and ( n68027 , n68026 , n32968 );
or ( n68028 , n68018 , n68027 );
and ( n68029 , n68028 , n33370 );
and ( n68030 , n32702 , n35062 );
or ( n68031 , C0 , n67999 , n68008 , n68029 , n68030 );
buf ( n68032 , n68031 );
buf ( n68033 , n68032 );
buf ( n68034 , n31655 );
buf ( n68035 , n31655 );
buf ( n68036 , n30987 );
not ( n68037 , n46356 );
and ( n68038 , n68037 , n31230 );
not ( n68039 , n49427 );
and ( n68040 , n68039 , n31230 );
and ( n68041 , n31238 , n49427 );
or ( n68042 , n68040 , n68041 );
and ( n68043 , n68042 , n46356 );
or ( n68044 , n68038 , n68043 );
and ( n68045 , n68044 , n31649 );
not ( n68046 , n49435 );
not ( n68047 , n49427 );
and ( n68048 , n68047 , n31230 );
and ( n68049 , n49901 , n49427 );
or ( n68050 , n68048 , n68049 );
and ( n68051 , n68046 , n68050 );
and ( n68052 , n49901 , n49435 );
or ( n68053 , n68051 , n68052 );
and ( n68054 , n68053 , n31643 );
not ( n68055 , n31452 );
not ( n68056 , n49435 );
not ( n68057 , n49427 );
and ( n68058 , n68057 , n31230 );
and ( n68059 , n49901 , n49427 );
or ( n68060 , n68058 , n68059 );
and ( n68061 , n68056 , n68060 );
and ( n68062 , n49901 , n49435 );
or ( n68063 , n68061 , n68062 );
and ( n68064 , n68055 , n68063 );
not ( n68065 , n49460 );
not ( n68066 , n49462 );
and ( n68067 , n68066 , n68063 );
and ( n68068 , n49925 , n49462 );
or ( n68069 , n68067 , n68068 );
and ( n68070 , n68065 , n68069 );
and ( n68071 , n49933 , n49460 );
or ( n68072 , n68070 , n68071 );
and ( n68073 , n68072 , n31452 );
or ( n68074 , n68064 , n68073 );
and ( n68075 , n68074 , n31638 );
and ( n68076 , n31230 , n47277 );
or ( n68077 , C0 , n68045 , n68054 , n68075 , n68076 );
buf ( n68078 , n68077 );
buf ( n68079 , n68078 );
not ( n68080 , n35542 );
and ( n68081 , n68080 , n41867 );
and ( n68082 , n52373 , n35542 );
or ( n68083 , n68081 , n68082 );
buf ( n68084 , n68083 );
buf ( n68085 , n68084 );
xor ( n68086 , n47288 , n47294 );
and ( n68087 , n68086 , n32433 );
not ( n68088 , n47331 );
and ( n68089 , n68088 , n47288 );
buf ( n68090 , n31891 );
and ( n68091 , n68090 , n47331 );
or ( n68092 , n68089 , n68091 );
and ( n68093 , n68092 , n32413 );
and ( n68094 , n47288 , n47402 );
or ( n68095 , n68087 , n68093 , n68094 );
and ( n68096 , n68095 , n32456 );
and ( n68097 , n47288 , n47409 );
or ( n68098 , C0 , n68096 , n68097 );
buf ( n68099 , n68098 );
buf ( n68100 , n68099 );
buf ( n68101 , n31655 );
buf ( n68102 , n31655 );
buf ( n68103 , n30987 );
not ( n68104 , n46356 );
and ( n68105 , n68104 , n31364 );
not ( n68106 , n49427 );
and ( n68107 , n68106 , n31364 );
and ( n68108 , n31372 , n49427 );
or ( n68109 , n68107 , n68108 );
and ( n68110 , n68109 , n46356 );
or ( n68111 , n68105 , n68110 );
and ( n68112 , n68111 , n31649 );
not ( n68113 , n49435 );
not ( n68114 , n49427 );
and ( n68115 , n68114 , n31364 );
and ( n68116 , n47849 , n49427 );
or ( n68117 , n68115 , n68116 );
and ( n68118 , n68113 , n68117 );
and ( n68119 , n47849 , n49435 );
or ( n68120 , n68118 , n68119 );
and ( n68121 , n68120 , n31643 );
not ( n68122 , n31452 );
not ( n68123 , n49435 );
not ( n68124 , n49427 );
and ( n68125 , n68124 , n31364 );
and ( n68126 , n47849 , n49427 );
or ( n68127 , n68125 , n68126 );
and ( n68128 , n68123 , n68127 );
and ( n68129 , n47849 , n49435 );
or ( n68130 , n68128 , n68129 );
and ( n68131 , n68122 , n68130 );
not ( n68132 , n49460 );
not ( n68133 , n49462 );
and ( n68134 , n68133 , n68130 );
and ( n68135 , n47877 , n49462 );
or ( n68136 , n68134 , n68135 );
and ( n68137 , n68132 , n68136 );
and ( n68138 , n47887 , n49460 );
or ( n68139 , n68137 , n68138 );
and ( n68140 , n68139 , n31452 );
or ( n68141 , n68131 , n68140 );
and ( n68142 , n68141 , n31638 );
and ( n68143 , n31364 , n47277 );
or ( n68144 , C0 , n68112 , n68121 , n68142 , n68143 );
buf ( n68145 , n68144 );
buf ( n68146 , n68145 );
buf ( n68147 , n40213 );
buf ( n68148 , n31655 );
xor ( n68149 , n45999 , n35297 );
and ( n68150 , n68149 , n32433 );
not ( n68151 , n47331 );
and ( n68152 , n68151 , n45999 );
buf ( n68153 , n32031 );
and ( n68154 , n68153 , n47331 );
or ( n68155 , n68152 , n68154 );
and ( n68156 , n68155 , n32413 );
and ( n68157 , n45999 , n47402 );
or ( n68158 , n68150 , n68156 , n68157 );
and ( n68159 , n68158 , n32456 );
and ( n68160 , n45999 , n47409 );
or ( n68161 , C0 , n68159 , n68160 );
buf ( n68162 , n68161 );
buf ( n68163 , n68162 );
not ( n68164 , n43755 );
and ( n68165 , n68164 , n43666 );
xor ( n68166 , n52303 , n52326 );
and ( n68167 , n68166 , n43755 );
or ( n68168 , n68165 , n68167 );
and ( n68169 , n68168 , n43774 );
not ( n68170 , n44663 );
and ( n68171 , n68170 , n44578 );
xor ( n68172 , n52341 , n52364 );
and ( n68173 , n68172 , n44663 );
or ( n68174 , n68171 , n68173 );
and ( n68175 , n68174 , n44682 );
buf ( n68176 , RI15b45bb8_244);
and ( n68177 , n68176 , n44695 );
or ( n68178 , n68169 , n68175 , n68177 );
buf ( n68179 , n68178 );
buf ( n68180 , n68179 );
buf ( n68181 , n30987 );
buf ( n68182 , n31655 );
buf ( n68183 , n31655 );
buf ( n68184 , n30987 );
xor ( n68185 , n33123 , n52217 );
and ( n68186 , n68185 , n33201 );
not ( n68187 , n41576 );
and ( n68188 , n68187 , n33123 );
buf ( n68189 , n32821 );
and ( n68190 , n68189 , n41576 );
or ( n68191 , n68188 , n68190 );
and ( n68192 , n68191 , n33189 );
and ( n68193 , n33123 , n41592 );
or ( n68194 , n68186 , n68192 , n68193 );
and ( n68195 , n68194 , n33208 );
and ( n68196 , n33123 , n39805 );
or ( n68197 , C0 , n68195 , n68196 );
buf ( n68198 , n68197 );
buf ( n68199 , n68198 );
buf ( n68200 , n30987 );
buf ( n68201 , n31655 );
not ( n68202 , n41532 );
and ( n68203 , n68202 , n34195 );
buf ( n68204 , RI15b533d0_705);
and ( n68205 , n68204 , n41532 );
or ( n68206 , n68203 , n68205 );
buf ( n68207 , n68206 );
buf ( n68208 , n68207 );
buf ( n68209 , n31655 );
buf ( n68210 , n30987 );
buf ( n68211 , n30987 );
not ( n68212 , n36587 );
and ( n68213 , n68212 , n36379 );
xor ( n68214 , n50178 , n50209 );
and ( n68215 , n68214 , n36587 );
or ( n68216 , n68213 , n68215 );
and ( n68217 , n68216 , n36596 );
not ( n68218 , n37485 );
and ( n68219 , n68218 , n37281 );
xor ( n68220 , n50228 , n50259 );
and ( n68221 , n68220 , n37485 );
or ( n68222 , n68219 , n68221 );
and ( n68223 , n68222 , n37494 );
and ( n68224 , n41856 , n37506 );
or ( n68225 , n68217 , n68223 , n68224 );
buf ( n68226 , n68225 );
buf ( n68227 , n68226 );
buf ( n68228 , n31655 );
and ( n68229 , n50439 , n50275 );
not ( n68230 , n50278 );
and ( n68231 , n68230 , n50407 );
and ( n68232 , n50439 , n50278 );
or ( n68233 , n68231 , n68232 );
and ( n68234 , n68233 , n32421 );
not ( n68235 , n50002 );
and ( n68236 , n68235 , n50407 );
and ( n68237 , n50439 , n50002 );
or ( n68238 , n68236 , n68237 );
and ( n68239 , n68238 , n32419 );
not ( n68240 , n50289 );
and ( n68241 , n68240 , n50407 );
and ( n68242 , n50439 , n50289 );
or ( n68243 , n68241 , n68242 );
and ( n68244 , n68243 , n32417 );
not ( n68245 , n50008 );
and ( n68246 , n68245 , n50407 );
and ( n68247 , n50439 , n50008 );
or ( n68248 , n68246 , n68247 );
and ( n68249 , n68248 , n32415 );
not ( n68250 , n47331 );
and ( n68251 , n68250 , n50407 );
and ( n68252 , n50417 , n47331 );
or ( n68253 , n68251 , n68252 );
and ( n68254 , n68253 , n32413 );
not ( n68255 , n50067 );
and ( n68256 , n68255 , n50407 );
and ( n68257 , n50417 , n50067 );
or ( n68258 , n68256 , n68257 );
and ( n68259 , n68258 , n32411 );
not ( n68260 , n31728 );
and ( n68261 , n68260 , n50407 );
and ( n68262 , n50427 , n31728 );
or ( n68263 , n68261 , n68262 );
and ( n68264 , n68263 , n32253 );
not ( n68265 , n32283 );
and ( n68266 , n68265 , n50407 );
and ( n68267 , n50468 , n32283 );
or ( n68268 , n68266 , n68267 );
and ( n68269 , n68268 , n32398 );
and ( n68270 , n50456 , n50334 );
or ( n68271 , n68229 , n68234 , n68239 , n68244 , n68249 , n68254 , n68259 , n68264 , n68269 , n68270 );
and ( n68272 , n68271 , n32456 );
and ( n68273 , n37531 , n32489 );
and ( n68274 , n50407 , n50345 );
or ( n68275 , C0 , n68272 , n68273 , n68274 );
buf ( n68276 , n68275 );
buf ( n68277 , n68276 );
buf ( n68278 , n30987 );
buf ( n68279 , n31655 );
buf ( n68280 , n31655 );
buf ( n68281 , RI15b47e68_318);
and ( n68282 , n32966 , n68281 );
not ( n68283 , n48265 );
and ( n68284 , n68282 , n68283 );
not ( n68285 , n68284 );
and ( n68286 , n32967 , n48265 );
not ( n68287 , n68286 );
and ( n68288 , n32967 , n68283 );
and ( n68289 , n68288 , n68281 );
not ( n68290 , n68289 );
not ( n68291 , n68281 );
and ( n68292 , n68288 , n68291 );
not ( n68293 , n68292 );
and ( n68294 , n68290 , n68293 );
buf ( n68295 , n68294 );
and ( n68296 , n68287 , n68295 );
buf ( n68297 , n68286 );
or ( n68298 , n68296 , n68297 );
and ( n68299 , n68285 , n68298 );
buf ( n68300 , n68284 );
or ( n68301 , n68299 , n68300 );
and ( n68302 , n68301 , n44694 );
buf ( n68303 , n43774 );
and ( n68304 , n68281 , n68283 );
not ( n68305 , n68304 );
and ( n68306 , n68291 , n68283 );
not ( n68307 , n68306 );
and ( n68308 , n68305 , n68307 );
buf ( n68309 , n68308 );
and ( n68310 , n68309 , n44692 );
not ( n68311 , n48294 );
and ( n68312 , n68311 , n68283 );
and ( n68313 , n68312 , n68281 );
not ( n68314 , n68313 );
or ( n68315 , n48265 , n68291 );
and ( n68316 , n68311 , n68315 );
not ( n68317 , n68316 );
not ( n68318 , n48294 );
and ( n68319 , n68317 , n68318 );
buf ( n68320 , n68316 );
or ( n68321 , n68319 , n68320 );
and ( n68322 , n68314 , n68321 );
buf ( n68323 , n68313 );
or ( n68324 , n68322 , n68323 );
and ( n68325 , n68324 , n44690 );
not ( n68326 , n68289 );
and ( n68327 , n32966 , n48294 );
not ( n68328 , n68327 );
or ( n68329 , n68281 , n48265 );
and ( n68330 , n32966 , n68311 );
and ( n68331 , n68329 , n68330 );
not ( n68332 , n68331 );
and ( n68333 , n68304 , n32966 );
and ( n68334 , n68333 , n68311 );
not ( n68335 , n68334 );
and ( n68336 , n68306 , n32967 );
not ( n68337 , n68336 );
and ( n68338 , n48265 , n32966 );
and ( n68339 , n68337 , n68338 );
buf ( n68340 , n68339 );
and ( n68341 , n68335 , n68340 );
buf ( n68342 , n68334 );
or ( n68343 , n68341 , n68342 );
and ( n68344 , n68332 , n68343 );
buf ( n68345 , n68331 );
or ( n68346 , n68344 , n68345 );
and ( n68347 , n68328 , n68346 );
and ( n68348 , n32959 , n68327 );
or ( n68349 , n68347 , n68348 );
and ( n68350 , n68326 , n68349 );
buf ( n68351 , n68350 );
and ( n68352 , n68351 , n44688 );
not ( n68353 , n68281 );
and ( n68354 , n68353 , n48265 );
buf ( n68355 , n68354 );
and ( n68356 , n68355 , n44685 );
or ( n68357 , n68302 , n68303 , n68310 , n68325 , n68352 , C0 , n68356 , C0 );
buf ( n68358 , n68357 );
buf ( n68359 , n68358 );
buf ( n68360 , n30987 );
not ( n68361 , n40163 );
and ( n68362 , n68361 , n31891 );
not ( n68363 , n40166 );
and ( n68364 , n68363 , n31891 );
and ( n68365 , n32218 , n40166 );
or ( n68366 , n68364 , n68365 );
and ( n68367 , n68366 , n40163 );
or ( n68368 , n68362 , n68367 );
and ( n68369 , n68368 , n32498 );
not ( n68370 , n40195 );
not ( n68371 , n40166 );
and ( n68372 , n68371 , n31891 );
and ( n68373 , n42255 , n40166 );
or ( n68374 , n68372 , n68373 );
and ( n68375 , n68370 , n68374 );
and ( n68376 , n42255 , n40195 );
or ( n68377 , n68375 , n68376 );
and ( n68378 , n68377 , n32473 );
not ( n68379 , n32475 );
not ( n68380 , n40195 );
not ( n68381 , n40166 );
and ( n68382 , n68381 , n31891 );
and ( n68383 , n42255 , n40166 );
or ( n68384 , n68382 , n68383 );
and ( n68385 , n68380 , n68384 );
and ( n68386 , n42255 , n40195 );
or ( n68387 , n68385 , n68386 );
and ( n68388 , n68379 , n68387 );
not ( n68389 , n40446 );
not ( n68390 , n40448 );
and ( n68391 , n68390 , n68387 );
and ( n68392 , n42283 , n40448 );
or ( n68393 , n68391 , n68392 );
and ( n68394 , n68389 , n68393 );
and ( n68395 , n42291 , n40446 );
or ( n68396 , n68394 , n68395 );
and ( n68397 , n68396 , n32475 );
or ( n68398 , n68388 , n68397 );
and ( n68399 , n68398 , n32486 );
and ( n68400 , n31891 , n41278 );
or ( n68401 , C0 , n68369 , n68378 , n68399 , n68400 );
buf ( n68402 , n68401 );
buf ( n68403 , n68402 );
xor ( n68404 , n35429 , n62854 );
and ( n68405 , n68404 , n31550 );
not ( n68406 , n39979 );
and ( n68407 , n68406 , n35429 );
and ( n68408 , n45129 , n59502 );
xor ( n68409 , n45112 , n68408 );
and ( n68410 , n68409 , n39979 );
or ( n68411 , n68407 , n68410 );
and ( n68412 , n68411 , n31538 );
and ( n68413 , n35429 , n40143 );
or ( n68414 , n68405 , n68412 , n68413 );
and ( n68415 , n68414 , n31557 );
and ( n68416 , n35429 , n40154 );
or ( n68417 , C0 , n68415 , n68416 );
buf ( n68418 , n68417 );
buf ( n68419 , n68418 );
buf ( n68420 , n30987 );
buf ( n68421 , n40218 );
buf ( n68422 , n31655 );
buf ( n68423 , n30987 );
buf ( n68424 , n31655 );
buf ( n68425 , n30987 );
not ( n68426 , n46356 );
and ( n68427 , n68426 , n31013 );
and ( n68428 , n46392 , n46356 );
or ( n68429 , n68427 , n68428 );
and ( n68430 , n68429 , n31649 );
not ( n68431 , n52614 );
not ( n68432 , n44702 );
and ( n68433 , n68432 , n31013 );
buf ( n68434 , n68433 );
and ( n68435 , n68431 , n68434 );
buf ( n68436 , n68435 );
and ( n68437 , n68436 , n31647 );
and ( n68438 , n46544 , n31643 );
not ( n68439 , n31452 );
and ( n68440 , n68439 , n46544 );
and ( n68441 , n46539 , n62675 );
xor ( n68442 , n46549 , n68441 );
not ( n68443 , n68442 );
buf ( n68444 , n68443 );
not ( n68445 , n68444 );
and ( n68446 , n68445 , n31452 );
or ( n68447 , n68440 , n68446 );
and ( n68448 , n68447 , n31638 );
and ( n68449 , n31013 , n52626 );
or ( n68450 , C0 , n68430 , n68437 , n68438 , n68448 , n68449 );
buf ( n68451 , n68450 );
buf ( n68452 , n68451 );
buf ( n68453 , n30987 );
buf ( n68454 , n31655 );
not ( n68455 , n31728 );
and ( n68456 , n68455 , n32463 );
xor ( n68457 , n31965 , n31998 );
xor ( n68458 , n68457 , n32072 );
and ( n68459 , n68458 , n31728 );
or ( n68460 , n68456 , n68459 );
and ( n68461 , n68460 , n32253 );
not ( n68462 , n32283 );
and ( n68463 , n68462 , n32463 );
not ( n68464 , n31823 );
xor ( n68465 , n32304 , n31998 );
xor ( n68466 , n68465 , n32311 );
and ( n68467 , n68464 , n68466 );
xor ( n68468 , n32360 , n32362 );
xor ( n68469 , n68468 , n32374 );
and ( n68470 , n68469 , n31823 );
or ( n68471 , n68467 , n68470 );
and ( n68472 , n68471 , n32283 );
or ( n68473 , n68463 , n68472 );
and ( n68474 , n68473 , n32398 );
and ( n68475 , n32463 , n32436 );
or ( n68476 , n68461 , n68474 , n68475 );
and ( n68477 , n68476 , n32456 );
and ( n68478 , n46062 , n32473 );
not ( n68479 , n32475 );
and ( n68480 , n68479 , n46062 );
not ( n68481 , n32463 );
and ( n68482 , n68481 , n32475 );
or ( n68483 , n68480 , n68482 );
and ( n68484 , n68483 , n32486 );
and ( n68485 , n37585 , n32489 );
and ( n68486 , n32463 , n32501 );
or ( n68487 , C0 , n68477 , n68478 , n68484 , n68485 , n68486 );
buf ( n68488 , n68487 );
buf ( n68489 , n68488 );
not ( n68490 , n46356 );
and ( n68491 , n68490 , n31286 );
not ( n68492 , n52734 );
and ( n68493 , n68492 , n31286 );
and ( n68494 , n31306 , n52734 );
or ( n68495 , n68493 , n68494 );
and ( n68496 , n68495 , n46356 );
or ( n68497 , n68491 , n68496 );
and ( n68498 , n68497 , n31649 );
not ( n68499 , n52742 );
not ( n68500 , n52734 );
and ( n68501 , n68500 , n31286 );
and ( n68502 , n58061 , n52734 );
or ( n68503 , n68501 , n68502 );
and ( n68504 , n68499 , n68503 );
and ( n68505 , n58061 , n52742 );
or ( n68506 , n68504 , n68505 );
and ( n68507 , n68506 , n31643 );
not ( n68508 , n31452 );
not ( n68509 , n52742 );
not ( n68510 , n52734 );
and ( n68511 , n68510 , n31286 );
and ( n68512 , n58061 , n52734 );
or ( n68513 , n68511 , n68512 );
and ( n68514 , n68509 , n68513 );
and ( n68515 , n58061 , n52742 );
or ( n68516 , n68514 , n68515 );
and ( n68517 , n68508 , n68516 );
not ( n68518 , n52762 );
not ( n68519 , n52764 );
and ( n68520 , n68519 , n68516 );
and ( n68521 , n58085 , n52764 );
or ( n68522 , n68520 , n68521 );
and ( n68523 , n68518 , n68522 );
and ( n68524 , n58093 , n52762 );
or ( n68525 , n68523 , n68524 );
and ( n68526 , n68525 , n31452 );
or ( n68527 , n68517 , n68526 );
and ( n68528 , n68527 , n31638 );
and ( n68529 , n31286 , n47277 );
or ( n68530 , C0 , n68498 , n68507 , n68528 , n68529 );
buf ( n68531 , n68530 );
buf ( n68532 , n68531 );
buf ( n68533 , n30987 );
or ( n68534 , n32496 , n32498 );
or ( n68535 , n68534 , n32500 );
and ( n68536 , n48263 , n68535 );
not ( n68537 , n35292 );
and ( n68538 , n48263 , n68537 );
and ( n68539 , n68538 , n32494 );
not ( n68540 , n35211 );
and ( n68541 , n68540 , n48263 );
not ( n68542 , n35288 );
buf ( n68543 , n68542 );
and ( n68544 , n35291 , n35288 );
or ( n68545 , n68543 , n68544 );
and ( n68546 , n68545 , n35211 );
or ( n68547 , n68541 , n68546 );
and ( n68548 , n68547 , n32421 );
not ( n68549 , n35245 );
and ( n68550 , n68549 , n48263 );
and ( n68551 , n35291 , n35245 );
or ( n68552 , n68550 , n68551 );
and ( n68553 , n68552 , n32419 );
not ( n68554 , n35278 );
and ( n68555 , n68554 , n48263 );
not ( n68556 , n50277 );
buf ( n68557 , n68556 );
and ( n68558 , n35293 , n50277 );
or ( n68559 , n68557 , n68558 );
and ( n68560 , n68559 , n35278 );
or ( n68561 , n68555 , n68560 );
and ( n68562 , n68561 , n32417 );
not ( n68563 , n35331 );
and ( n68564 , n68563 , n48263 );
not ( n68565 , n35292 );
buf ( n68566 , n68565 );
buf ( n68567 , n68566 );
and ( n68568 , n68567 , n35331 );
or ( n68569 , n68564 , n68568 );
and ( n68570 , n68569 , n32415 );
and ( n68571 , n48263 , n35354 );
or ( n68572 , n68548 , n68553 , n68562 , n68570 , n68571 );
and ( n68573 , n68572 , n32456 );
or ( n68574 , n32489 , n32491 );
or ( n68575 , n68574 , n32492 );
buf ( n68576 , n68575 );
or ( n68577 , C0 , n68536 , n68539 , n68573 , C0 , n68576 );
buf ( n68578 , n68577 );
buf ( n68579 , n68578 );
buf ( n68580 , n31655 );
buf ( n68581 , n31655 );
buf ( n68582 , n30987 );
buf ( n68583 , n31655 );
and ( n68584 , n48805 , n34150 );
buf ( n68585 , n68584 );
and ( n68586 , n68585 , n33381 );
and ( n68587 , n56609 , n33379 );
and ( n68588 , n57670 , n33208 );
and ( n68589 , n32539 , n61311 );
or ( n68590 , C0 , n68586 , n68587 , n68588 , n68589 );
buf ( n68591 , n68590 );
buf ( n68592 , n68591 );
buf ( n68593 , n31655 );
buf ( n68594 , n30987 );
buf ( n68595 , n31655 );
buf ( n68596 , n30987 );
not ( n68597 , n40163 );
and ( n68598 , n68597 , n32054 );
not ( n68599 , n49298 );
and ( n68600 , n68599 , n32054 );
and ( n68601 , n32130 , n49298 );
or ( n68602 , n68600 , n68601 );
and ( n68603 , n68602 , n40163 );
or ( n68604 , n68598 , n68603 );
and ( n68605 , n68604 , n32498 );
not ( n68606 , n49306 );
not ( n68607 , n49298 );
and ( n68608 , n68607 , n32054 );
and ( n68609 , n45833 , n49298 );
or ( n68610 , n68608 , n68609 );
and ( n68611 , n68606 , n68610 );
and ( n68612 , n45833 , n49306 );
or ( n68613 , n68611 , n68612 );
and ( n68614 , n68613 , n32473 );
not ( n68615 , n32475 );
not ( n68616 , n49306 );
not ( n68617 , n49298 );
and ( n68618 , n68617 , n32054 );
and ( n68619 , n45833 , n49298 );
or ( n68620 , n68618 , n68619 );
and ( n68621 , n68616 , n68620 );
and ( n68622 , n45833 , n49306 );
or ( n68623 , n68621 , n68622 );
and ( n68624 , n68615 , n68623 );
not ( n68625 , n49331 );
not ( n68626 , n49333 );
and ( n68627 , n68626 , n68623 );
and ( n68628 , n45857 , n49333 );
or ( n68629 , n68627 , n68628 );
and ( n68630 , n68625 , n68629 );
and ( n68631 , n45865 , n49331 );
or ( n68632 , n68630 , n68631 );
and ( n68633 , n68632 , n32475 );
or ( n68634 , n68624 , n68633 );
and ( n68635 , n68634 , n32486 );
and ( n68636 , n32054 , n41278 );
or ( n68637 , C0 , n68605 , n68614 , n68635 , n68636 );
buf ( n68638 , n68637 );
buf ( n68639 , n68638 );
xor ( n68640 , n44776 , n44791 );
and ( n68641 , n68640 , n31548 );
not ( n68642 , n44807 );
and ( n68643 , n68642 , n44776 );
and ( n68644 , n46561 , n44807 );
or ( n68645 , n68643 , n68644 );
and ( n68646 , n68645 , n31408 );
not ( n68647 , n44817 );
and ( n68648 , n68647 , n44776 );
and ( n68649 , n65510 , n44817 );
or ( n68650 , n68648 , n68649 );
and ( n68651 , n68650 , n31521 );
not ( n68652 , n45059 );
and ( n68653 , n68652 , n44776 );
and ( n68654 , n31086 , n40095 );
and ( n68655 , n31090 , n40097 );
and ( n68656 , n31094 , n40099 );
and ( n68657 , n31098 , n40101 );
and ( n68658 , n31101 , n40103 );
and ( n68659 , n31105 , n40105 );
and ( n68660 , n31108 , n40107 );
and ( n68661 , n31111 , n40109 );
and ( n68662 , n31114 , n40111 );
and ( n68663 , n31117 , n40113 );
and ( n68664 , n31120 , n40115 );
and ( n68665 , n31123 , n40117 );
and ( n68666 , n31126 , n40119 );
and ( n68667 , n31129 , n40121 );
and ( n68668 , n31132 , n40123 );
and ( n68669 , n31135 , n40125 );
or ( n68670 , n68654 , n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , n68661 , n68662 , n68663 , n68664 , n68665 , n68666 , n68667 , n68668 , n68669 );
and ( n68671 , n68670 , n45059 );
or ( n68672 , n68653 , n68671 );
and ( n68673 , n68672 , n31536 );
and ( n68674 , n44776 , n45148 );
or ( n68675 , n68641 , n68646 , n68651 , n68673 , n68674 );
and ( n68676 , n68675 , n31557 );
and ( n68677 , n44776 , n40154 );
or ( n68678 , C0 , n68676 , n68677 );
buf ( n68679 , n68678 );
buf ( n68680 , n68679 );
buf ( n68681 , n30987 );
and ( n68682 , n51807 , n31645 );
not ( n68683 , n45274 );
and ( n68684 , n68683 , n60249 );
not ( n68685 , n41809 );
and ( n68686 , n68685 , n41753 );
xor ( n68687 , n62435 , n62436 );
and ( n68688 , n68687 , n41809 );
or ( n68689 , n68686 , n68688 );
and ( n68690 , n68689 , n45274 );
or ( n68691 , n68684 , n68690 );
and ( n68692 , n68691 , n31373 );
not ( n68693 , n45280 );
and ( n68694 , n68693 , n60249 );
and ( n68695 , n68689 , n45280 );
or ( n68696 , n68694 , n68695 );
and ( n68697 , n68696 , n31468 );
and ( n68698 , n60249 , n45802 );
or ( n68699 , n68692 , n68697 , n68698 );
and ( n68700 , n68699 , n31557 );
and ( n68701 , n60249 , n45808 );
or ( n68702 , C0 , n68682 , n68700 , n68701 );
buf ( n68703 , n68702 );
buf ( n68704 , n68703 );
buf ( n68705 , n30987 );
buf ( n68706 , n31655 );
not ( n68707 , n40163 );
and ( n68708 , n68707 , n31937 );
not ( n68709 , n53227 );
and ( n68710 , n68709 , n31937 );
and ( n68711 , n32183 , n53227 );
or ( n68712 , n68710 , n68711 );
and ( n68713 , n68712 , n40163 );
or ( n68714 , n68708 , n68713 );
and ( n68715 , n68714 , n32498 );
not ( n68716 , n53235 );
not ( n68717 , n53227 );
and ( n68718 , n68717 , n31937 );
and ( n68719 , n45178 , n53227 );
or ( n68720 , n68718 , n68719 );
and ( n68721 , n68716 , n68720 );
and ( n68722 , n45178 , n53235 );
or ( n68723 , n68721 , n68722 );
and ( n68724 , n68723 , n32473 );
not ( n68725 , n32475 );
not ( n68726 , n53235 );
not ( n68727 , n53227 );
and ( n68728 , n68727 , n31937 );
and ( n68729 , n45178 , n53227 );
or ( n68730 , n68728 , n68729 );
and ( n68731 , n68726 , n68730 );
and ( n68732 , n45178 , n53235 );
or ( n68733 , n68731 , n68732 );
and ( n68734 , n68725 , n68733 );
not ( n68735 , n53260 );
not ( n68736 , n53262 );
and ( n68737 , n68736 , n68733 );
and ( n68738 , n45206 , n53262 );
or ( n68739 , n68737 , n68738 );
and ( n68740 , n68735 , n68739 );
and ( n68741 , n45214 , n53260 );
or ( n68742 , n68740 , n68741 );
and ( n68743 , n68742 , n32475 );
or ( n68744 , n68734 , n68743 );
and ( n68745 , n68744 , n32486 );
and ( n68746 , n31937 , n41278 );
or ( n68747 , C0 , n68715 , n68724 , n68745 , n68746 );
buf ( n68748 , n68747 );
buf ( n68749 , n68748 );
buf ( n68750 , n31655 );
buf ( n68751 , n30987 );
buf ( n68752 , n31655 );
buf ( n68753 , n30987 );
not ( n68754 , n32598 );
and ( n68755 , n58206 , n68754 );
and ( n68756 , n68755 , n32890 );
not ( n68757 , n32919 );
and ( n68758 , n58206 , n68757 );
and ( n68759 , n68758 , n32924 );
not ( n68760 , n32953 );
and ( n68761 , n68760 , n58206 );
buf ( n68762 , n32953 );
or ( n68763 , n68761 , n68762 );
and ( n68764 , n68763 , n33038 );
not ( n68765 , n33067 );
and ( n68766 , n68765 , n58206 );
buf ( n68767 , n33067 );
or ( n68768 , n68766 , n68767 );
and ( n68769 , n68768 , n33172 );
and ( n68770 , n58206 , n33204 );
or ( n68771 , n68756 , n68759 , n68764 , n68769 , n68770 );
and ( n68772 , n68771 , n33208 );
and ( n68773 , n58206 , n58908 );
buf ( n68774 , n58910 );
or ( n68775 , C0 , n68772 , n68773 , n68774 );
buf ( n68776 , n68775 );
buf ( n68777 , n68776 );
and ( n68778 , n32459 , n32500 );
not ( n68779 , n35211 );
and ( n68780 , n68779 , n37577 );
buf ( n68781 , n68780 );
and ( n68782 , n68781 , n32421 );
not ( n68783 , n35245 );
and ( n68784 , n68783 , n37577 );
buf ( n68785 , n68784 );
and ( n68786 , n68785 , n32419 );
not ( n68787 , n35278 );
and ( n68788 , n68787 , n37577 );
not ( n68789 , n35295 );
and ( n68790 , n68789 , n47287 );
xor ( n68791 , n37577 , n49526 );
and ( n68792 , n68791 , n35295 );
or ( n68793 , n68790 , n68792 );
and ( n68794 , n68793 , n35278 );
or ( n68795 , n68788 , n68794 );
and ( n68796 , n68795 , n32417 );
not ( n68797 , n35331 );
and ( n68798 , n68797 , n37577 );
not ( n68799 , n35294 );
not ( n68800 , n45995 );
and ( n68801 , n68800 , n47287 );
xor ( n68802 , n49605 , n49612 );
and ( n68803 , n68802 , n45995 );
or ( n68804 , n68801 , n68803 );
and ( n68805 , n68799 , n68804 );
and ( n68806 , n68791 , n35294 );
or ( n68807 , n68805 , n68806 );
and ( n68808 , n68807 , n35331 );
or ( n68809 , n68798 , n68808 );
and ( n68810 , n68809 , n32415 );
and ( n68811 , n37577 , n35354 );
or ( n68812 , n68782 , n68786 , n68796 , n68810 , n68811 );
and ( n68813 , n68812 , n32456 );
not ( n68814 , n32475 );
not ( n68815 , n46060 );
and ( n68816 , n68815 , n44750 );
xor ( n68817 , n49696 , n49706 );
and ( n68818 , n68817 , n46060 );
or ( n68819 , n68816 , n68818 );
and ( n68820 , n68814 , n68819 );
and ( n68821 , n37577 , n32475 );
or ( n68822 , n68820 , n68821 );
and ( n68823 , n68822 , n32486 );
buf ( n68824 , n32489 );
and ( n68825 , n37577 , n35367 );
or ( n68826 , C0 , n68778 , n68813 , n68823 , n68824 , n68825 );
buf ( n68827 , n68826 );
buf ( n68828 , n68827 );
buf ( n68829 , n30987 );
buf ( n68830 , n31655 );
not ( n68831 , n35542 );
and ( n68832 , n68831 , n41849 );
and ( n68833 , n66768 , n35542 );
or ( n68834 , n68832 , n68833 );
buf ( n68835 , n68834 );
buf ( n68836 , n68835 );
buf ( n68837 , n31655 );
and ( n68838 , n33333 , n32528 );
not ( n68839 , n32598 );
and ( n68840 , n68839 , n42695 );
and ( n68841 , n48790 , n32598 );
or ( n68842 , n68840 , n68841 );
and ( n68843 , n68842 , n32890 );
not ( n68844 , n32919 );
and ( n68845 , n68844 , n42695 );
and ( n68846 , n48790 , n32919 );
or ( n68847 , n68845 , n68846 );
and ( n68848 , n68847 , n32924 );
not ( n68849 , n32953 );
and ( n68850 , n68849 , n42695 );
not ( n68851 , n32971 );
and ( n68852 , n68851 , n33133 );
and ( n68853 , n42695 , n32971 );
or ( n68854 , n68852 , n68853 );
and ( n68855 , n68854 , n32953 );
or ( n68856 , n68850 , n68855 );
and ( n68857 , n68856 , n33038 );
not ( n68858 , n33067 );
and ( n68859 , n68858 , n42695 );
not ( n68860 , n32970 );
buf ( n68861 , n33133 );
and ( n68862 , n68860 , n68861 );
and ( n68863 , n42695 , n32970 );
or ( n68864 , n68862 , n68863 );
and ( n68865 , n68864 , n33067 );
or ( n68866 , n68859 , n68865 );
and ( n68867 , n68866 , n33172 );
and ( n68868 , n42695 , n33204 );
or ( n68869 , n68843 , n68848 , n68857 , n68867 , n68868 );
and ( n68870 , n68869 , n33208 );
not ( n68871 , n32968 );
buf ( n68872 , n33333 );
and ( n68873 , n68871 , n68872 );
and ( n68874 , n42695 , n32968 );
or ( n68875 , n68873 , n68874 );
and ( n68876 , n68875 , n33370 );
and ( n68877 , n42695 , n33382 );
or ( n68878 , C0 , n68838 , n68870 , n68876 , C0 , n68877 );
buf ( n68879 , n68878 );
buf ( n68880 , n68879 );
buf ( n68881 , n30987 );
buf ( n68882 , n31655 );
not ( n68883 , n46356 );
and ( n68884 , n68883 , n31260 );
not ( n68885 , n64746 );
and ( n68886 , n68885 , n31260 );
and ( n68887 , n31272 , n64746 );
or ( n68888 , n68886 , n68887 );
and ( n68889 , n68888 , n46356 );
or ( n68890 , n68884 , n68889 );
and ( n68891 , n68890 , n31649 );
not ( n68892 , n64754 );
not ( n68893 , n64746 );
and ( n68894 , n68893 , n31260 );
and ( n68895 , n49443 , n64746 );
or ( n68896 , n68894 , n68895 );
and ( n68897 , n68892 , n68896 );
and ( n68898 , n49443 , n64754 );
or ( n68899 , n68897 , n68898 );
and ( n68900 , n68899 , n31643 );
not ( n68901 , n31452 );
not ( n68902 , n64754 );
not ( n68903 , n64746 );
and ( n68904 , n68903 , n31260 );
and ( n68905 , n49443 , n64746 );
or ( n68906 , n68904 , n68905 );
and ( n68907 , n68902 , n68906 );
and ( n68908 , n49443 , n64754 );
or ( n68909 , n68907 , n68908 );
and ( n68910 , n68901 , n68909 );
not ( n68911 , n64774 );
not ( n68912 , n64776 );
and ( n68913 , n68912 , n68909 );
and ( n68914 , n49469 , n64776 );
or ( n68915 , n68913 , n68914 );
and ( n68916 , n68911 , n68915 );
and ( n68917 , n49477 , n64774 );
or ( n68918 , n68916 , n68917 );
and ( n68919 , n68918 , n31452 );
or ( n68920 , n68910 , n68919 );
and ( n68921 , n68920 , n31638 );
and ( n68922 , n31260 , n47277 );
or ( n68923 , C0 , n68891 , n68900 , n68921 , n68922 );
buf ( n68924 , n68923 );
buf ( n68925 , n68924 );
buf ( n68926 , n31655 );
xor ( n68927 , n50967 , n64713 );
and ( n68928 , n68927 , n32431 );
not ( n68929 , n50002 );
and ( n68930 , n68929 , n50967 );
and ( n68931 , n40627 , n50002 );
or ( n68932 , n68930 , n68931 );
and ( n68933 , n68932 , n32419 );
not ( n68934 , n50008 );
and ( n68935 , n68934 , n50967 );
not ( n68936 , n51594 );
and ( n68937 , n68936 , n51470 );
xor ( n68938 , n51599 , n51607 );
and ( n68939 , n68938 , n51594 );
or ( n68940 , n68937 , n68939 );
and ( n68941 , n68940 , n50008 );
or ( n68942 , n68935 , n68941 );
and ( n68943 , n68942 , n32415 );
not ( n68944 , n50067 );
and ( n68945 , n68944 , n50967 );
and ( n68946 , n31896 , n60510 );
and ( n68947 , n31898 , n60512 );
and ( n68948 , n31900 , n60514 );
and ( n68949 , n31902 , n60516 );
and ( n68950 , n31904 , n60518 );
and ( n68951 , n31906 , n60520 );
and ( n68952 , n31908 , n60522 );
and ( n68953 , n31910 , n60524 );
and ( n68954 , n31912 , n60526 );
and ( n68955 , n31914 , n60528 );
and ( n68956 , n31916 , n60530 );
and ( n68957 , n31918 , n60532 );
and ( n68958 , n31920 , n60534 );
and ( n68959 , n31922 , n60536 );
and ( n68960 , n31924 , n60538 );
and ( n68961 , n31926 , n60540 );
or ( n68962 , n68946 , n68947 , n68948 , n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , n68961 );
and ( n68963 , n68962 , n50067 );
or ( n68964 , n68945 , n68963 );
and ( n68965 , n68964 , n32411 );
and ( n68966 , n50967 , n50098 );
or ( n68967 , n68928 , n68933 , n68943 , n68965 , n68966 );
and ( n68968 , n68967 , n32456 );
and ( n68969 , n50967 , n47409 );
or ( n68970 , C0 , n68968 , n68969 );
buf ( n68971 , n68970 );
buf ( n68972 , n68971 );
buf ( n68973 , n30987 );
buf ( n68974 , n31655 );
buf ( n68975 , n30987 );
xor ( n68976 , n44773 , n44794 );
and ( n68977 , n68976 , n31548 );
not ( n68978 , n44807 );
and ( n68979 , n68978 , n44773 );
and ( n68980 , n46662 , n44807 );
or ( n68981 , n68979 , n68980 );
and ( n68982 , n68981 , n31408 );
not ( n68983 , n44817 );
and ( n68984 , n68983 , n44773 );
not ( n68985 , n44994 );
and ( n68986 , n68985 , n44858 );
xor ( n68987 , n45007 , n45013 );
and ( n68988 , n68987 , n44994 );
or ( n68989 , n68986 , n68988 );
and ( n68990 , n68989 , n44817 );
or ( n68991 , n68984 , n68990 );
and ( n68992 , n68991 , n31521 );
not ( n68993 , n45059 );
and ( n68994 , n68993 , n44773 );
and ( n68995 , n31206 , n40095 );
and ( n68996 , n31208 , n40097 );
and ( n68997 , n31210 , n40099 );
and ( n68998 , n31212 , n40101 );
and ( n68999 , n31214 , n40103 );
and ( n69000 , n31216 , n40105 );
and ( n69001 , n31218 , n40107 );
and ( n69002 , n31220 , n40109 );
and ( n69003 , n31222 , n40111 );
and ( n69004 , n31224 , n40113 );
and ( n69005 , n31226 , n40115 );
and ( n69006 , n31228 , n40117 );
and ( n69007 , n31230 , n40119 );
and ( n69008 , n31232 , n40121 );
and ( n69009 , n31234 , n40123 );
and ( n69010 , n31236 , n40125 );
or ( n69011 , n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , n69010 );
and ( n69012 , n69011 , n45059 );
or ( n69013 , n68994 , n69012 );
and ( n69014 , n69013 , n31536 );
and ( n69015 , n44773 , n45148 );
or ( n69016 , n68977 , n68982 , n68992 , n69014 , n69015 );
and ( n69017 , n69016 , n31557 );
and ( n69018 , n44773 , n40154 );
or ( n69019 , C0 , n69017 , n69018 );
buf ( n69020 , n69019 );
buf ( n69021 , n69020 );
not ( n69022 , n40163 );
and ( n69023 , n69022 , n31881 );
not ( n69024 , n55888 );
and ( n69025 , n69024 , n31881 );
and ( n69026 , n32218 , n55888 );
or ( n69027 , n69025 , n69026 );
and ( n69028 , n69027 , n40163 );
or ( n69029 , n69023 , n69028 );
and ( n69030 , n69029 , n32498 );
not ( n69031 , n55896 );
not ( n69032 , n55888 );
and ( n69033 , n69032 , n31881 );
and ( n69034 , n42255 , n55888 );
or ( n69035 , n69033 , n69034 );
and ( n69036 , n69031 , n69035 );
and ( n69037 , n42255 , n55896 );
or ( n69038 , n69036 , n69037 );
and ( n69039 , n69038 , n32473 );
not ( n69040 , n32475 );
not ( n69041 , n55896 );
not ( n69042 , n55888 );
and ( n69043 , n69042 , n31881 );
and ( n69044 , n42255 , n55888 );
or ( n69045 , n69043 , n69044 );
and ( n69046 , n69041 , n69045 );
and ( n69047 , n42255 , n55896 );
or ( n69048 , n69046 , n69047 );
and ( n69049 , n69040 , n69048 );
not ( n69050 , n55916 );
not ( n69051 , n55918 );
and ( n69052 , n69051 , n69048 );
and ( n69053 , n42283 , n55918 );
or ( n69054 , n69052 , n69053 );
and ( n69055 , n69050 , n69054 );
and ( n69056 , n42291 , n55916 );
or ( n69057 , n69055 , n69056 );
and ( n69058 , n69057 , n32475 );
or ( n69059 , n69049 , n69058 );
and ( n69060 , n69059 , n32486 );
and ( n69061 , n31881 , n41278 );
or ( n69062 , C0 , n69030 , n69039 , n69060 , n69061 );
buf ( n69063 , n69062 );
buf ( n69064 , n69063 );
buf ( n69065 , n30987 );
xor ( n69066 , n34052 , n39931 );
and ( n69067 , n69066 , n31550 );
not ( n69068 , n39979 );
and ( n69069 , n69068 , n34052 );
and ( n69070 , n31140 , n42330 );
and ( n69071 , n31142 , n42332 );
and ( n69072 , n31144 , n42334 );
and ( n69073 , n31146 , n42336 );
and ( n69074 , n31148 , n42338 );
and ( n69075 , n31150 , n42340 );
and ( n69076 , n31152 , n42342 );
and ( n69077 , n31154 , n42344 );
and ( n69078 , n31156 , n42346 );
and ( n69079 , n31158 , n42348 );
and ( n69080 , n31160 , n42350 );
and ( n69081 , n31162 , n42352 );
and ( n69082 , n31164 , n42354 );
and ( n69083 , n31166 , n42356 );
and ( n69084 , n31168 , n42358 );
and ( n69085 , n31170 , n42360 );
or ( n69086 , n69070 , n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , n69085 );
and ( n69087 , n69086 , n39979 );
or ( n69088 , n69069 , n69087 );
and ( n69089 , n69088 , n31538 );
and ( n69090 , n34052 , n40143 );
or ( n69091 , n69067 , n69089 , n69090 );
and ( n69092 , n69091 , n31557 );
and ( n69093 , n34052 , n40154 );
or ( n69094 , C0 , n69092 , n69093 );
buf ( n69095 , n69094 );
buf ( n69096 , n69095 );
not ( n69097 , n40163 );
and ( n69098 , n69097 , n31814 );
not ( n69099 , n42238 );
and ( n69100 , n69099 , n31814 );
and ( n69101 , n32252 , n42238 );
or ( n69102 , n69100 , n69101 );
and ( n69103 , n69102 , n40163 );
or ( n69104 , n69098 , n69103 );
and ( n69105 , n69104 , n32498 );
not ( n69106 , n42247 );
not ( n69107 , n42238 );
and ( n69108 , n69107 , n31814 );
and ( n69109 , n40393 , n42238 );
or ( n69110 , n69108 , n69109 );
and ( n69111 , n69106 , n69110 );
and ( n69112 , n40393 , n42247 );
or ( n69113 , n69111 , n69112 );
and ( n69114 , n69113 , n32473 );
not ( n69115 , n32475 );
not ( n69116 , n42247 );
not ( n69117 , n42238 );
and ( n69118 , n69117 , n31814 );
and ( n69119 , n40393 , n42238 );
or ( n69120 , n69118 , n69119 );
and ( n69121 , n69116 , n69120 );
and ( n69122 , n40393 , n42247 );
or ( n69123 , n69121 , n69122 );
and ( n69124 , n69115 , n69123 );
not ( n69125 , n42273 );
not ( n69126 , n42276 );
and ( n69127 , n69126 , n69123 );
and ( n69128 , n40972 , n42276 );
or ( n69129 , n69127 , n69128 );
and ( n69130 , n69125 , n69129 );
and ( n69131 , n41267 , n42273 );
or ( n69132 , n69130 , n69131 );
and ( n69133 , n69132 , n32475 );
or ( n69134 , n69124 , n69133 );
and ( n69135 , n69134 , n32486 );
and ( n69136 , n31814 , n41278 );
or ( n69137 , C0 , n69105 , n69114 , n69135 , n69136 );
buf ( n69138 , n69137 );
buf ( n69139 , n69138 );
buf ( n69140 , n30987 );
buf ( n69141 , n31655 );
buf ( n69142 , n30987 );
buf ( n69143 , n30987 );
buf ( n69144 , n31655 );
buf ( n69145 , n31655 );
buf ( n69146 , n30987 );
buf ( n69147 , RI15b47fd0_321);
not ( n69148 , n69147 );
and ( n69149 , n69148 , n58207 );
buf ( n69150 , n44686 );
or ( n69151 , n44685 , n44688 );
or ( n69152 , n69151 , n44690 );
or ( n69153 , n69152 , n44692 );
or ( n69154 , n69153 , n44694 );
and ( n69155 , n54728 , n69154 );
or ( n69156 , n69149 , n69150 , n69155 );
buf ( n69157 , n69156 );
buf ( n69158 , n69157 );
and ( n69159 , n55561 , n32496 );
not ( n69160 , n50278 );
and ( n69161 , n69160 , n31658 );
buf ( n69162 , n69161 );
and ( n69163 , n69162 , n32421 );
not ( n69164 , n50002 );
and ( n69165 , n69164 , n31658 );
and ( n69166 , n31662 , n47350 );
xor ( n69167 , n31658 , n69166 );
and ( n69168 , n69167 , n50002 );
or ( n69169 , n69165 , n69168 );
and ( n69170 , n69169 , n32419 );
not ( n69171 , n50289 );
and ( n69172 , n69171 , n31658 );
buf ( n69173 , n69172 );
and ( n69174 , n69173 , n32417 );
not ( n69175 , n50008 );
and ( n69176 , n69175 , n31658 );
buf ( n69177 , n69176 );
and ( n69178 , n69177 , n32415 );
not ( n69179 , n47331 );
and ( n69180 , n69179 , n31658 );
buf ( n69181 , n69180 );
and ( n69182 , n69181 , n32413 );
not ( n69183 , n50067 );
and ( n69184 , n69183 , n31658 );
buf ( n69185 , n69184 );
and ( n69186 , n69185 , n32411 );
and ( n69187 , n31658 , n63978 );
or ( n69188 , C0 , n69163 , n69170 , n69174 , n69178 , n69182 , n69186 , n69187 , C0 );
and ( n69189 , n69188 , n32456 );
and ( n69190 , n31658 , n63983 );
or ( n69191 , C0 , C0 , n69159 , n69189 , n69190 );
buf ( n69192 , n69191 );
buf ( n69193 , n69192 );
buf ( n69194 , n31655 );
not ( n69195 , n36587 );
and ( n69196 , n69195 , n36277 );
xor ( n69197 , n50184 , n50203 );
and ( n69198 , n69197 , n36587 );
or ( n69199 , n69196 , n69198 );
and ( n69200 , n69199 , n36596 );
not ( n69201 , n37485 );
and ( n69202 , n69201 , n37179 );
xor ( n69203 , n50234 , n50253 );
and ( n69204 , n69203 , n37485 );
or ( n69205 , n69202 , n69204 );
and ( n69206 , n69205 , n37494 );
and ( n69207 , n41850 , n37506 );
or ( n69208 , n69200 , n69206 , n69207 );
buf ( n69209 , n69208 );
buf ( n69210 , n69209 );
buf ( n69211 , n30987 );
buf ( n69212 , n30987 );
not ( n69213 , n34150 );
and ( n69214 , n69213 , n32881 );
not ( n69215 , n56093 );
and ( n69216 , n69215 , n32881 );
and ( n69217 , n32889 , n56093 );
or ( n69218 , n69216 , n69217 );
and ( n69219 , n69218 , n34150 );
or ( n69220 , n69214 , n69219 );
and ( n69221 , n69220 , n33381 );
not ( n69222 , n56101 );
not ( n69223 , n56093 );
and ( n69224 , n69223 , n32881 );
and ( n69225 , n52819 , n56093 );
or ( n69226 , n69224 , n69225 );
and ( n69227 , n69222 , n69226 );
and ( n69228 , n52819 , n56101 );
or ( n69229 , n69227 , n69228 );
and ( n69230 , n69229 , n33375 );
not ( n69231 , n32968 );
not ( n69232 , n56101 );
not ( n69233 , n56093 );
and ( n69234 , n69233 , n32881 );
and ( n69235 , n52819 , n56093 );
or ( n69236 , n69234 , n69235 );
and ( n69237 , n69232 , n69236 );
and ( n69238 , n52819 , n56101 );
or ( n69239 , n69237 , n69238 );
and ( n69240 , n69231 , n69239 );
not ( n69241 , n56121 );
not ( n69242 , n56123 );
and ( n69243 , n69242 , n69239 );
and ( n69244 , n52845 , n56123 );
or ( n69245 , n69243 , n69244 );
and ( n69246 , n69241 , n69245 );
and ( n69247 , n52855 , n56121 );
or ( n69248 , n69246 , n69247 );
and ( n69249 , n69248 , n32968 );
or ( n69250 , n69240 , n69249 );
and ( n69251 , n69250 , n33370 );
and ( n69252 , n32881 , n35062 );
or ( n69253 , C0 , n69221 , n69230 , n69251 , n69252 );
buf ( n69254 , n69253 );
buf ( n69255 , n69254 );
not ( n69256 , n34150 );
and ( n69257 , n69256 , n32649 );
not ( n69258 , n56140 );
and ( n69259 , n69258 , n32649 );
and ( n69260 , n32655 , n56140 );
or ( n69261 , n69259 , n69260 );
and ( n69262 , n69261 , n34150 );
or ( n69263 , n69257 , n69262 );
and ( n69264 , n69263 , n33381 );
not ( n69265 , n56148 );
not ( n69266 , n56140 );
and ( n69267 , n69266 , n32649 );
and ( n69268 , n56044 , n56140 );
or ( n69269 , n69267 , n69268 );
and ( n69270 , n69265 , n69269 );
and ( n69271 , n56044 , n56148 );
or ( n69272 , n69270 , n69271 );
and ( n69273 , n69272 , n33375 );
not ( n69274 , n32968 );
not ( n69275 , n56148 );
not ( n69276 , n56140 );
and ( n69277 , n69276 , n32649 );
and ( n69278 , n56044 , n56140 );
or ( n69279 , n69277 , n69278 );
and ( n69280 , n69275 , n69279 );
and ( n69281 , n56044 , n56148 );
or ( n69282 , n69280 , n69281 );
and ( n69283 , n69274 , n69282 );
not ( n69284 , n56168 );
not ( n69285 , n56170 );
and ( n69286 , n69285 , n69282 );
and ( n69287 , n56068 , n56170 );
or ( n69288 , n69286 , n69287 );
and ( n69289 , n69284 , n69288 );
and ( n69290 , n56076 , n56168 );
or ( n69291 , n69289 , n69290 );
and ( n69292 , n69291 , n32968 );
or ( n69293 , n69283 , n69292 );
and ( n69294 , n69293 , n33370 );
and ( n69295 , n32649 , n35062 );
or ( n69296 , C0 , n69264 , n69273 , n69294 , n69295 );
buf ( n69297 , n69296 );
buf ( n69298 , n69297 );
buf ( n69299 , n30987 );
buf ( n69300 , n31655 );
buf ( n69301 , n31655 );
not ( n69302 , n35278 );
and ( n69303 , n69302 , n60901 );
and ( n69304 , n60910 , n35278 );
or ( n69305 , n69303 , n69304 );
and ( n69306 , n69305 , n32417 );
not ( n69307 , n47912 );
and ( n69308 , n69307 , n60901 );
not ( n69309 , n48101 );
and ( n69310 , n69309 , n48061 );
xor ( n69311 , n50018 , n50027 );
and ( n69312 , n69311 , n48101 );
or ( n69313 , n69310 , n69312 );
and ( n69314 , n69313 , n47912 );
or ( n69315 , n69308 , n69314 );
and ( n69316 , n69315 , n32415 );
and ( n69317 , n60901 , n48133 );
or ( n69318 , n69306 , n69316 , n69317 );
and ( n69319 , n69318 , n32456 );
and ( n69320 , n60901 , n47409 );
or ( n69321 , C0 , n69319 , n69320 );
buf ( n69322 , n69321 );
buf ( n69323 , n69322 );
buf ( n69324 , n31655 );
buf ( n69325 , n30987 );
buf ( n69326 , n31655 );
not ( n69327 , n46356 );
and ( n69328 , n69327 , n31175 );
not ( n69329 , n47831 );
and ( n69330 , n69329 , n31175 );
and ( n69331 , n31205 , n47831 );
or ( n69332 , n69330 , n69331 );
and ( n69333 , n69332 , n46356 );
or ( n69334 , n69328 , n69333 );
and ( n69335 , n69334 , n31649 );
not ( n69336 , n47839 );
not ( n69337 , n47831 );
and ( n69338 , n69337 , n31175 );
and ( n69339 , n50125 , n47831 );
or ( n69340 , n69338 , n69339 );
and ( n69341 , n69336 , n69340 );
and ( n69342 , n50125 , n47839 );
or ( n69343 , n69341 , n69342 );
and ( n69344 , n69343 , n31643 );
not ( n69345 , n31452 );
not ( n69346 , n47839 );
not ( n69347 , n47831 );
and ( n69348 , n69347 , n31175 );
and ( n69349 , n50125 , n47831 );
or ( n69350 , n69348 , n69349 );
and ( n69351 , n69346 , n69350 );
and ( n69352 , n50125 , n47839 );
or ( n69353 , n69351 , n69352 );
and ( n69354 , n69345 , n69353 );
not ( n69355 , n47866 );
not ( n69356 , n47868 );
and ( n69357 , n69356 , n69353 );
and ( n69358 , n50151 , n47868 );
or ( n69359 , n69357 , n69358 );
and ( n69360 , n69355 , n69359 );
and ( n69361 , n50159 , n47866 );
or ( n69362 , n69360 , n69361 );
and ( n69363 , n69362 , n31452 );
or ( n69364 , n69354 , n69363 );
and ( n69365 , n69364 , n31638 );
and ( n69366 , n31175 , n47277 );
or ( n69367 , C0 , n69335 , n69344 , n69365 , n69366 );
buf ( n69368 , n69367 );
buf ( n69369 , n69368 );
buf ( n69370 , n31655 );
not ( n69371 , n43755 );
and ( n69372 , n69371 , n43513 );
xor ( n69373 , n52312 , n52317 );
and ( n69374 , n69373 , n43755 );
or ( n69375 , n69372 , n69374 );
and ( n69376 , n69375 , n43774 );
not ( n69377 , n44663 );
and ( n69378 , n69377 , n44425 );
xor ( n69379 , n52350 , n52355 );
and ( n69380 , n69379 , n44663 );
or ( n69381 , n69378 , n69380 );
and ( n69382 , n69381 , n44682 );
and ( n69383 , n56827 , n44695 );
or ( n69384 , n69376 , n69382 , n69383 );
buf ( n69385 , n69384 );
buf ( n69386 , n69385 );
buf ( n69387 , n30987 );
buf ( n69388 , n30987 );
buf ( n69389 , n31655 );
buf ( n69390 , n31655 );
buf ( n69391 , RI15b5f568_1118);
and ( n69392 , n69391 , n32494 );
not ( n69393 , n46083 );
and ( n69394 , n69393 , n60253 );
not ( n69395 , n46290 );
and ( n69396 , n69395 , n46234 );
xor ( n69397 , n46295 , n46317 );
and ( n69398 , n69397 , n46290 );
or ( n69399 , n69396 , n69398 );
and ( n69400 , n69399 , n46083 );
or ( n69401 , n69394 , n69400 );
and ( n69402 , n69401 , n32421 );
not ( n69403 , n46326 );
and ( n69404 , n69403 , n60253 );
and ( n69405 , n69399 , n46326 );
or ( n69406 , n69404 , n69405 );
and ( n69407 , n69406 , n32417 );
and ( n69408 , n60253 , n46340 );
or ( n69409 , n69402 , n69407 , n69408 );
and ( n69410 , n69409 , n32456 );
and ( n69411 , n60253 , n46349 );
or ( n69412 , C0 , n69392 , n69410 , n69411 );
buf ( n69413 , n69412 );
buf ( n69414 , n69413 );
buf ( n69415 , n31655 );
buf ( n69416 , n30987 );
not ( n69417 , n46356 );
and ( n69418 , n69417 , n31212 );
not ( n69419 , n46362 );
and ( n69420 , n69419 , n31212 );
and ( n69421 , n31238 , n46362 );
or ( n69422 , n69420 , n69421 );
and ( n69423 , n69422 , n46356 );
or ( n69424 , n69418 , n69423 );
and ( n69425 , n69424 , n31649 );
not ( n69426 , n46393 );
not ( n69427 , n46362 );
and ( n69428 , n69427 , n31212 );
and ( n69429 , n49901 , n46362 );
or ( n69430 , n69428 , n69429 );
and ( n69431 , n69426 , n69430 );
and ( n69432 , n49901 , n46393 );
or ( n69433 , n69431 , n69432 );
and ( n69434 , n69433 , n31643 );
not ( n69435 , n31452 );
not ( n69436 , n46393 );
not ( n69437 , n46362 );
and ( n69438 , n69437 , n31212 );
and ( n69439 , n49901 , n46362 );
or ( n69440 , n69438 , n69439 );
and ( n69441 , n69436 , n69440 );
and ( n69442 , n49901 , n46393 );
or ( n69443 , n69441 , n69442 );
and ( n69444 , n69435 , n69443 );
not ( n69445 , n46550 );
not ( n69446 , n46554 );
and ( n69447 , n69446 , n69443 );
and ( n69448 , n49925 , n46554 );
or ( n69449 , n69447 , n69448 );
and ( n69450 , n69445 , n69449 );
and ( n69451 , n49933 , n46550 );
or ( n69452 , n69450 , n69451 );
and ( n69453 , n69452 , n31452 );
or ( n69454 , n69444 , n69453 );
and ( n69455 , n69454 , n31638 );
and ( n69456 , n31212 , n47277 );
or ( n69457 , C0 , n69425 , n69434 , n69455 , n69456 );
buf ( n69458 , n69457 );
buf ( n69459 , n69458 );
buf ( n69460 , n30987 );
buf ( n69461 , n31655 );
buf ( n69462 , RI15b480c0_323);
and ( n69463 , n69462 , n58207 );
and ( n69464 , n54735 , n44695 );
or ( n69465 , n69463 , n69464 );
buf ( n69466 , n69465 );
buf ( n69467 , n69466 );
buf ( n69468 , n31655 );
buf ( n69469 , n30987 );
buf ( n69470 , n30987 );
buf ( n69471 , n31655 );
buf ( n69472 , n31655 );
buf ( n69473 , n30987 );
buf ( n69474 , n40208 );
not ( n69475 , n34150 );
and ( n69476 , n69475 , n32673 );
not ( n69477 , n57038 );
and ( n69478 , n69477 , n32673 );
and ( n69479 , n32689 , n57038 );
or ( n69480 , n69478 , n69479 );
and ( n69481 , n69480 , n34150 );
or ( n69482 , n69476 , n69481 );
and ( n69483 , n69482 , n33381 );
not ( n69484 , n57046 );
not ( n69485 , n57038 );
and ( n69486 , n69485 , n32673 );
and ( n69487 , n50682 , n57038 );
or ( n69488 , n69486 , n69487 );
and ( n69489 , n69484 , n69488 );
and ( n69490 , n50682 , n57046 );
or ( n69491 , n69489 , n69490 );
and ( n69492 , n69491 , n33375 );
not ( n69493 , n32968 );
not ( n69494 , n57046 );
not ( n69495 , n57038 );
and ( n69496 , n69495 , n32673 );
and ( n69497 , n50682 , n57038 );
or ( n69498 , n69496 , n69497 );
and ( n69499 , n69494 , n69498 );
and ( n69500 , n50682 , n57046 );
or ( n69501 , n69499 , n69500 );
and ( n69502 , n69493 , n69501 );
not ( n69503 , n57066 );
not ( n69504 , n57068 );
and ( n69505 , n69504 , n69501 );
and ( n69506 , n50706 , n57068 );
or ( n69507 , n69505 , n69506 );
and ( n69508 , n69503 , n69507 );
and ( n69509 , n50714 , n57066 );
or ( n69510 , n69508 , n69509 );
and ( n69511 , n69510 , n32968 );
or ( n69512 , n69502 , n69511 );
and ( n69513 , n69512 , n33370 );
and ( n69514 , n32673 , n35062 );
or ( n69515 , C0 , n69483 , n69492 , n69513 , n69514 );
buf ( n69516 , n69515 );
buf ( n69517 , n69516 );
buf ( n69518 , n30987 );
buf ( n69519 , n31655 );
buf ( n69520 , n31655 );
buf ( n69521 , n30987 );
not ( n69522 , n43755 );
and ( n69523 , n69522 , n43717 );
xor ( n69524 , n52300 , n52329 );
and ( n69525 , n69524 , n43755 );
or ( n69526 , n69523 , n69525 );
and ( n69527 , n69526 , n43774 );
not ( n69528 , n44663 );
and ( n69529 , n69528 , n44629 );
xor ( n69530 , n52338 , n52367 );
and ( n69531 , n69530 , n44663 );
or ( n69532 , n69529 , n69531 );
and ( n69533 , n69532 , n44682 );
and ( n69534 , n58705 , n44695 );
or ( n69535 , n69527 , n69533 , n69534 );
buf ( n69536 , n69535 );
buf ( n69537 , n69536 );
not ( n69538 , n43755 );
and ( n69539 , n69538 , n43581 );
xor ( n69540 , n52308 , n52321 );
and ( n69541 , n69540 , n43755 );
or ( n69542 , n69539 , n69541 );
and ( n69543 , n69542 , n43774 );
not ( n69544 , n44663 );
and ( n69545 , n69544 , n44493 );
xor ( n69546 , n52346 , n52359 );
and ( n69547 , n69546 , n44663 );
or ( n69548 , n69545 , n69547 );
and ( n69549 , n69548 , n44682 );
buf ( n69550 , RI15b45960_239);
and ( n69551 , n69550 , n44695 );
or ( n69552 , n69543 , n69549 , n69551 );
buf ( n69553 , n69552 );
buf ( n69554 , n69553 );
buf ( n69555 , n31655 );
buf ( n69556 , n30987 );
buf ( n69557 , n30987 );
buf ( n69558 , n31655 );
buf ( n69559 , n31655 );
buf ( n69560 , n30987 );
and ( n69561 , n32302 , n50275 );
not ( n69562 , n50278 );
and ( n69563 , n69562 , n31737 );
and ( n69564 , n32302 , n50278 );
or ( n69565 , n69563 , n69564 );
and ( n69566 , n69565 , n32421 );
not ( n69567 , n50002 );
and ( n69568 , n69567 , n31737 );
and ( n69569 , n32302 , n50002 );
or ( n69570 , n69568 , n69569 );
and ( n69571 , n69570 , n32419 );
not ( n69572 , n50289 );
and ( n69573 , n69572 , n31737 );
and ( n69574 , n32302 , n50289 );
or ( n69575 , n69573 , n69574 );
and ( n69576 , n69575 , n32417 );
not ( n69577 , n50008 );
and ( n69578 , n69577 , n31737 );
and ( n69579 , n32302 , n50008 );
or ( n69580 , n69578 , n69579 );
and ( n69581 , n69580 , n32415 );
not ( n69582 , n47331 );
and ( n69583 , n69582 , n31737 );
and ( n69584 , n31930 , n47331 );
or ( n69585 , n69583 , n69584 );
and ( n69586 , n69585 , n32413 );
not ( n69587 , n50067 );
and ( n69588 , n69587 , n31737 );
and ( n69589 , n31930 , n50067 );
or ( n69590 , n69588 , n69589 );
and ( n69591 , n69590 , n32411 );
not ( n69592 , n31728 );
and ( n69593 , n69592 , n31737 );
and ( n69594 , n62692 , n31728 );
or ( n69595 , n69593 , n69594 );
and ( n69596 , n69595 , n32253 );
not ( n69597 , n32283 );
and ( n69598 , n69597 , n31737 );
and ( n69599 , n62705 , n32283 );
or ( n69600 , n69598 , n69599 );
and ( n69601 , n69600 , n32398 );
and ( n69602 , n32356 , n50334 );
or ( n69603 , n69561 , n69566 , n69571 , n69576 , n69581 , n69586 , n69591 , n69596 , n69601 , n69602 );
and ( n69604 , n69603 , n32456 );
and ( n69605 , n37583 , n32489 );
and ( n69606 , n31737 , n50345 );
or ( n69607 , C0 , n69604 , n69605 , n69606 );
buf ( n69608 , n69607 );
buf ( n69609 , n69608 );
not ( n69610 , n31437 );
buf ( n69611 , RI15b52980_683);
and ( n69612 , n69610 , n69611 );
not ( n69613 , n45766 );
and ( n69614 , n69613 , n45694 );
xor ( n69615 , n45889 , n45890 );
and ( n69616 , n69615 , n45766 );
or ( n69617 , n69614 , n69616 );
and ( n69618 , n69617 , n31437 );
or ( n69619 , n69612 , n69618 );
and ( n69620 , n69619 , n31468 );
not ( n69621 , n44817 );
and ( n69622 , n69621 , n69611 );
not ( n69623 , n44994 );
and ( n69624 , n69623 , n44942 );
xor ( n69625 , n45000 , n45020 );
and ( n69626 , n69625 , n44994 );
or ( n69627 , n69624 , n69626 );
and ( n69628 , n69627 , n44817 );
or ( n69629 , n69622 , n69628 );
and ( n69630 , n69629 , n31521 );
and ( n69631 , n69611 , n42158 );
or ( n69632 , n69620 , n69630 , n69631 );
and ( n69633 , n69632 , n31557 );
and ( n69634 , n69611 , n40154 );
or ( n69635 , C0 , n69633 , n69634 );
buf ( n69636 , n69635 );
buf ( n69637 , n69636 );
buf ( n69638 , n30987 );
not ( n69639 , n34150 );
and ( n69640 , n69639 , n32607 );
not ( n69641 , n50731 );
and ( n69642 , n69641 , n32607 );
and ( n69643 , n32655 , n50731 );
or ( n69644 , n69642 , n69643 );
and ( n69645 , n69644 , n34150 );
or ( n69646 , n69640 , n69645 );
and ( n69647 , n69646 , n33381 );
not ( n69648 , n50739 );
not ( n69649 , n50731 );
and ( n69650 , n69649 , n32607 );
and ( n69651 , n56044 , n50731 );
or ( n69652 , n69650 , n69651 );
and ( n69653 , n69648 , n69652 );
and ( n69654 , n56044 , n50739 );
or ( n69655 , n69653 , n69654 );
and ( n69656 , n69655 , n33375 );
not ( n69657 , n32968 );
not ( n69658 , n50739 );
not ( n69659 , n50731 );
and ( n69660 , n69659 , n32607 );
and ( n69661 , n56044 , n50731 );
or ( n69662 , n69660 , n69661 );
and ( n69663 , n69658 , n69662 );
and ( n69664 , n56044 , n50739 );
or ( n69665 , n69663 , n69664 );
and ( n69666 , n69657 , n69665 );
not ( n69667 , n50759 );
not ( n69668 , n50761 );
and ( n69669 , n69668 , n69665 );
and ( n69670 , n56068 , n50761 );
or ( n69671 , n69669 , n69670 );
and ( n69672 , n69667 , n69671 );
and ( n69673 , n56076 , n50759 );
or ( n69674 , n69672 , n69673 );
and ( n69675 , n69674 , n32968 );
or ( n69676 , n69666 , n69675 );
and ( n69677 , n69676 , n33370 );
and ( n69678 , n32607 , n35062 );
or ( n69679 , C0 , n69647 , n69656 , n69677 , n69678 );
buf ( n69680 , n69679 );
buf ( n69681 , n69680 );
buf ( n69682 , n30987 );
buf ( n69683 , n31655 );
buf ( n69684 , n31655 );
not ( n69685 , n50828 );
not ( n69686 , n50834 );
and ( n69687 , n69686 , n40625 );
buf ( n69688 , RI15b53cb8_724);
and ( n69689 , n69688 , n50834 );
or ( n69690 , n69687 , n69689 );
and ( n69691 , n69685 , n69690 );
buf ( n69692 , RI15b60120_1143);
and ( n69693 , n69692 , n50828 );
or ( n69694 , n69691 , n69693 );
buf ( n69695 , n69694 );
buf ( n69696 , n69695 );
buf ( n69697 , n31655 );
buf ( n69698 , n30987 );
buf ( n69699 , n30987 );
buf ( n69700 , n31655 );
xor ( n69701 , n33097 , n58385 );
and ( n69702 , n69701 , n33201 );
not ( n69703 , n41576 );
and ( n69704 , n69703 , n33097 );
and ( n69705 , n32690 , n55215 );
and ( n69706 , n32692 , n55217 );
and ( n69707 , n32694 , n55219 );
and ( n69708 , n32696 , n55221 );
and ( n69709 , n32698 , n55223 );
and ( n69710 , n32700 , n55225 );
and ( n69711 , n32702 , n55227 );
and ( n69712 , n32704 , n55229 );
and ( n69713 , n32706 , n55231 );
and ( n69714 , n32708 , n55233 );
and ( n69715 , n32710 , n55235 );
and ( n69716 , n32712 , n55237 );
and ( n69717 , n32714 , n55239 );
and ( n69718 , n32716 , n55241 );
and ( n69719 , n32718 , n55243 );
and ( n69720 , n32720 , n55245 );
or ( n69721 , n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n69719 , n69720 );
and ( n69722 , n69721 , n41576 );
or ( n69723 , n69704 , n69722 );
and ( n69724 , n69723 , n33189 );
and ( n69725 , n33097 , n41592 );
or ( n69726 , n69702 , n69724 , n69725 );
and ( n69727 , n69726 , n33208 );
and ( n69728 , n33097 , n39805 );
or ( n69729 , C0 , n69727 , n69728 );
buf ( n69730 , n69729 );
buf ( n69731 , n69730 );
not ( n69732 , n35278 );
buf ( n69733 , RI15b5f4f0_1117);
and ( n69734 , n69732 , n69733 );
not ( n69735 , n46290 );
and ( n69736 , n69735 , n46221 );
xor ( n69737 , n46296 , n46316 );
and ( n69738 , n69737 , n46290 );
or ( n69739 , n69736 , n69738 );
and ( n69740 , n69739 , n35278 );
or ( n69741 , n69734 , n69740 );
and ( n69742 , n69741 , n32417 );
not ( n69743 , n47912 );
and ( n69744 , n69743 , n69733 );
not ( n69745 , n48101 );
and ( n69746 , n69745 , n48037 );
xor ( n69747 , n50020 , n50025 );
and ( n69748 , n69747 , n48101 );
or ( n69749 , n69746 , n69748 );
and ( n69750 , n69749 , n47912 );
or ( n69751 , n69744 , n69750 );
and ( n69752 , n69751 , n32415 );
and ( n69753 , n69733 , n48133 );
or ( n69754 , n69742 , n69752 , n69753 );
and ( n69755 , n69754 , n32456 );
and ( n69756 , n69733 , n47409 );
or ( n69757 , C0 , n69755 , n69756 );
buf ( n69758 , n69757 );
buf ( n69759 , n69758 );
buf ( n69760 , n30987 );
not ( n69761 , n46356 );
and ( n69762 , n69761 , n31242 );
not ( n69763 , n47831 );
and ( n69764 , n69763 , n31242 );
and ( n69765 , n31272 , n47831 );
or ( n69766 , n69764 , n69765 );
and ( n69767 , n69766 , n46356 );
or ( n69768 , n69762 , n69767 );
and ( n69769 , n69768 , n31649 );
not ( n69770 , n47839 );
not ( n69771 , n47831 );
and ( n69772 , n69771 , n31242 );
and ( n69773 , n49443 , n47831 );
or ( n69774 , n69772 , n69773 );
and ( n69775 , n69770 , n69774 );
and ( n69776 , n49443 , n47839 );
or ( n69777 , n69775 , n69776 );
and ( n69778 , n69777 , n31643 );
not ( n69779 , n31452 );
not ( n69780 , n47839 );
not ( n69781 , n47831 );
and ( n69782 , n69781 , n31242 );
and ( n69783 , n49443 , n47831 );
or ( n69784 , n69782 , n69783 );
and ( n69785 , n69780 , n69784 );
and ( n69786 , n49443 , n47839 );
or ( n69787 , n69785 , n69786 );
and ( n69788 , n69779 , n69787 );
not ( n69789 , n47866 );
not ( n69790 , n47868 );
and ( n69791 , n69790 , n69787 );
and ( n69792 , n49469 , n47868 );
or ( n69793 , n69791 , n69792 );
and ( n69794 , n69789 , n69793 );
and ( n69795 , n49477 , n47866 );
or ( n69796 , n69794 , n69795 );
and ( n69797 , n69796 , n31452 );
or ( n69798 , n69788 , n69797 );
and ( n69799 , n69798 , n31638 );
and ( n69800 , n31242 , n47277 );
or ( n69801 , C0 , n69769 , n69778 , n69799 , n69800 );
buf ( n69802 , n69801 );
buf ( n69803 , n69802 );
buf ( n69804 , n31655 );
buf ( n69805 , n31655 );
buf ( n69806 , n30987 );
not ( n69807 , n32953 );
buf ( n69808 , RI15b46248_258);
and ( n69809 , n69807 , n69808 );
not ( n69810 , n54581 );
and ( n69811 , n69810 , n54407 );
xor ( n69812 , n64018 , n64023 );
and ( n69813 , n69812 , n54581 );
or ( n69814 , n69811 , n69813 );
and ( n69815 , n69814 , n32953 );
or ( n69816 , n69809 , n69815 );
and ( n69817 , n69816 , n33038 );
not ( n69818 , n48660 );
and ( n69819 , n69818 , n69808 );
and ( n69820 , n64869 , n48660 );
or ( n69821 , n69819 , n69820 );
and ( n69822 , n69821 , n33172 );
and ( n69823 , n69808 , n39795 );
or ( n69824 , n69817 , n69822 , n69823 );
and ( n69825 , n69824 , n33208 );
and ( n69826 , n69808 , n39805 );
or ( n69827 , C0 , n69825 , n69826 );
buf ( n69828 , n69827 );
buf ( n69829 , n69828 );
buf ( n69830 , n30987 );
buf ( n69831 , n31655 );
and ( n69832 , n31582 , n31007 );
not ( n69833 , n31077 );
and ( n69834 , n69833 , n34006 );
buf ( n69835 , n69834 );
and ( n69836 , n69835 , n31373 );
not ( n69837 , n31402 );
and ( n69838 , n69837 , n34006 );
buf ( n69839 , n69838 );
and ( n69840 , n69839 , n31408 );
not ( n69841 , n31437 );
and ( n69842 , n69841 , n34006 );
not ( n69843 , n31455 );
and ( n69844 , n69843 , n34052 );
xor ( n69845 , n34006 , n34017 );
and ( n69846 , n69845 , n31455 );
or ( n69847 , n69844 , n69846 );
and ( n69848 , n69847 , n31437 );
or ( n69849 , n69842 , n69848 );
and ( n69850 , n69849 , n31468 );
not ( n69851 , n31497 );
and ( n69852 , n69851 , n34006 );
not ( n69853 , n31454 );
not ( n69854 , n31501 );
and ( n69855 , n69854 , n34052 );
xor ( n69856 , n34053 , n34069 );
and ( n69857 , n69856 , n31501 );
or ( n69858 , n69855 , n69857 );
and ( n69859 , n69853 , n69858 );
and ( n69860 , n69845 , n31454 );
or ( n69861 , n69859 , n69860 );
and ( n69862 , n69861 , n31497 );
or ( n69863 , n69852 , n69862 );
and ( n69864 , n69863 , n31521 );
and ( n69865 , n34006 , n31553 );
or ( n69866 , n69836 , n69840 , n69850 , n69864 , n69865 );
and ( n69867 , n69866 , n31557 );
not ( n69868 , n31452 );
not ( n69869 , n31619 );
and ( n69870 , n69869 , n34109 );
xor ( n69871 , n34110 , n34126 );
and ( n69872 , n69871 , n31619 );
or ( n69873 , n69870 , n69872 );
and ( n69874 , n69868 , n69873 );
and ( n69875 , n34006 , n31452 );
or ( n69876 , n69874 , n69875 );
and ( n69877 , n69876 , n31638 );
buf ( n69878 , n33973 );
and ( n69879 , n34006 , n31650 );
or ( n69880 , C0 , n69832 , n69867 , n69877 , n69878 , n69879 );
buf ( n69881 , n69880 );
buf ( n69882 , n69881 );
buf ( n69883 , n31655 );
buf ( n69884 , n31655 );
not ( n69885 , n33419 );
and ( n69886 , n69885 , n31562 );
and ( n69887 , n57507 , n33419 );
or ( n69888 , n69886 , n69887 );
and ( n69889 , n69888 , n31529 );
not ( n69890 , n33734 );
and ( n69891 , n69890 , n31562 );
and ( n69892 , n57532 , n33734 );
or ( n69893 , n69891 , n69892 );
and ( n69894 , n69893 , n31527 );
and ( n69895 , n31562 , n33942 );
or ( n69896 , n69889 , n69894 , n69895 );
and ( n69897 , n69896 , n31557 );
and ( n69898 , n35480 , n31643 );
not ( n69899 , n31452 );
and ( n69900 , n69899 , n35480 );
xor ( n69901 , n31562 , n59438 );
and ( n69902 , n69901 , n31452 );
or ( n69903 , n69900 , n69902 );
and ( n69904 , n69903 , n31638 );
and ( n69905 , n35388 , n33973 );
and ( n69906 , n31562 , n33978 );
or ( n69907 , C0 , n69897 , n69898 , n69904 , n69905 , n69906 );
buf ( n69908 , n69907 );
buf ( n69909 , n69908 );
buf ( n69910 , n30987 );
buf ( n69911 , n30987 );
buf ( n69912 , n31655 );
not ( n69913 , n38443 );
and ( n69914 , n69913 , n38439 );
xor ( n69915 , n38439 , n37947 );
xor ( n69916 , n38422 , n37947 );
xor ( n69917 , n38405 , n37947 );
xor ( n69918 , n38388 , n37947 );
and ( n69919 , n53460 , n53509 );
and ( n69920 , n69918 , n69919 );
and ( n69921 , n69917 , n69920 );
and ( n69922 , n69916 , n69921 );
xor ( n69923 , n69915 , n69922 );
and ( n69924 , n69923 , n38443 );
or ( n69925 , n69914 , n69924 );
and ( n69926 , n69925 , n38450 );
not ( n69927 , n39339 );
and ( n69928 , n69927 , n39335 );
xor ( n69929 , n39335 , n38847 );
xor ( n69930 , n39322 , n38847 );
xor ( n69931 , n39305 , n38847 );
xor ( n69932 , n39288 , n38847 );
and ( n69933 , n53516 , n53565 );
and ( n69934 , n69932 , n69933 );
and ( n69935 , n69931 , n69934 );
and ( n69936 , n69930 , n69935 );
xor ( n69937 , n69929 , n69936 );
and ( n69938 , n69937 , n39339 );
or ( n69939 , n69928 , n69938 );
and ( n69940 , n69939 , n39346 );
and ( n69941 , n40199 , n39359 );
or ( n69942 , n69926 , n69940 , n69941 );
buf ( n69943 , n69942 );
buf ( n69944 , n69943 );
buf ( n69945 , n30987 );
and ( n69946 , n33760 , n48455 );
not ( n69947 , n48457 );
and ( n69948 , n69947 , n33425 );
and ( n69949 , n33760 , n48457 );
or ( n69950 , n69948 , n69949 );
and ( n69951 , n69950 , n31373 );
not ( n69952 , n44807 );
and ( n69953 , n69952 , n33425 );
and ( n69954 , n33760 , n44807 );
or ( n69955 , n69953 , n69954 );
and ( n69956 , n69955 , n31408 );
not ( n69957 , n48468 );
and ( n69958 , n69957 , n33425 );
and ( n69959 , n33760 , n48468 );
or ( n69960 , n69958 , n69959 );
and ( n69961 , n69960 , n31468 );
not ( n69962 , n44817 );
and ( n69963 , n69962 , n33425 );
and ( n69964 , n33760 , n44817 );
or ( n69965 , n69963 , n69964 );
and ( n69966 , n69965 , n31521 );
not ( n69967 , n39979 );
and ( n69968 , n69967 , n33425 );
and ( n69969 , n33467 , n39979 );
or ( n69970 , n69968 , n69969 );
and ( n69971 , n69970 , n31538 );
not ( n69972 , n45059 );
and ( n69973 , n69972 , n33425 );
and ( n69974 , n33467 , n45059 );
or ( n69975 , n69973 , n69974 );
and ( n69976 , n69975 , n31536 );
not ( n69977 , n33419 );
and ( n69978 , n69977 , n33425 );
xor ( n69979 , n33467 , n33698 );
and ( n69980 , n69979 , n33419 );
or ( n69981 , n69978 , n69980 );
and ( n69982 , n69981 , n31529 );
not ( n69983 , n33734 );
and ( n69984 , n69983 , n33425 );
not ( n69985 , n33533 );
xor ( n69986 , n33760 , n33816 );
and ( n69987 , n69985 , n69986 );
xnor ( n69988 , n33845 , n33918 );
and ( n69989 , n69988 , n33533 );
or ( n69990 , n69987 , n69989 );
and ( n69991 , n69990 , n33734 );
or ( n69992 , n69984 , n69991 );
and ( n69993 , n69992 , n31527 );
and ( n69994 , n33845 , n48513 );
or ( n69995 , n69946 , n69951 , n69956 , n69961 , n69966 , n69971 , n69976 , n69982 , n69993 , n69994 );
and ( n69996 , n69995 , n31557 );
and ( n69997 , n35398 , n33973 );
and ( n69998 , n33425 , n48524 );
or ( n69999 , C0 , n69996 , n69997 , n69998 );
buf ( n70000 , n69999 );
buf ( n70001 , n70000 );
not ( n70002 , n41532 );
and ( n70003 , n70002 , n34419 );
and ( n70004 , n61591 , n41532 );
or ( n70005 , n70003 , n70004 );
buf ( n70006 , n70005 );
buf ( n70007 , n70006 );
xor ( n70008 , n39480 , n54972 );
and ( n70009 , n70008 , n33199 );
not ( n70010 , n48648 );
and ( n70011 , n70010 , n39480 );
and ( n70012 , n34377 , n48648 );
or ( n70013 , n70011 , n70012 );
and ( n70014 , n70013 , n32924 );
not ( n70015 , n48660 );
and ( n70016 , n70015 , n39480 );
not ( n70017 , n39584 );
and ( n70018 , n70017 , n51913 );
and ( n70019 , n51929 , n39584 );
or ( n70020 , n70018 , n70019 );
and ( n70021 , n70020 , n48660 );
or ( n70022 , n70016 , n70021 );
and ( n70023 , n70022 , n33172 );
not ( n70024 , n48730 );
and ( n70025 , n70024 , n39480 );
and ( n70026 , n61574 , n48730 );
or ( n70027 , n70025 , n70026 );
and ( n70028 , n70027 , n33187 );
and ( n70029 , n39480 , n54713 );
or ( n70030 , n70009 , n70014 , n70023 , n70028 , n70029 );
and ( n70031 , n70030 , n33208 );
and ( n70032 , n39480 , n39805 );
or ( n70033 , C0 , n70031 , n70032 );
buf ( n70034 , n70033 );
buf ( n70035 , n70034 );
buf ( n70036 , n30987 );
buf ( n70037 , n31655 );
buf ( n70038 , n31655 );
buf ( n70039 , n30987 );
and ( n70040 , n50957 , n67360 );
xor ( n70041 , n50955 , n70040 );
and ( n70042 , n70041 , n32431 );
not ( n70043 , n50002 );
and ( n70044 , n70043 , n50955 );
and ( n70045 , n40585 , n50002 );
or ( n70046 , n70044 , n70045 );
and ( n70047 , n70046 , n32419 );
not ( n70048 , n50008 );
and ( n70049 , n70048 , n50955 );
not ( n70050 , n51594 );
and ( n70051 , n70050 , n51542 );
xor ( n70052 , n59227 , n59234 );
and ( n70053 , n70052 , n51594 );
or ( n70054 , n70051 , n70053 );
and ( n70055 , n70054 , n50008 );
or ( n70056 , n70049 , n70055 );
and ( n70057 , n70056 , n32415 );
not ( n70058 , n50067 );
and ( n70059 , n70058 , n50955 );
and ( n70060 , n60450 , n67380 );
xor ( n70061 , n60433 , n70060 );
and ( n70062 , n70061 , n50067 );
or ( n70063 , n70059 , n70062 );
and ( n70064 , n70063 , n32411 );
and ( n70065 , n50955 , n50098 );
or ( n70066 , n70042 , n70047 , n70057 , n70064 , n70065 );
and ( n70067 , n70066 , n32456 );
and ( n70068 , n50955 , n47409 );
or ( n70069 , C0 , n70067 , n70068 );
buf ( n70070 , n70069 );
buf ( n70071 , n70070 );
buf ( n70072 , n31655 );
not ( n70073 , n46356 );
and ( n70074 , n70073 , n31329 );
not ( n70075 , n56904 );
and ( n70076 , n70075 , n31329 );
and ( n70077 , n31339 , n56904 );
or ( n70078 , n70076 , n70077 );
and ( n70079 , n70078 , n46356 );
or ( n70080 , n70074 , n70079 );
and ( n70081 , n70080 , n31649 );
not ( n70082 , n56912 );
not ( n70083 , n56904 );
and ( n70084 , n70083 , n31329 );
and ( n70085 , n47449 , n56904 );
or ( n70086 , n70084 , n70085 );
and ( n70087 , n70082 , n70086 );
and ( n70088 , n47449 , n56912 );
or ( n70089 , n70087 , n70088 );
and ( n70090 , n70089 , n31643 );
not ( n70091 , n31452 );
not ( n70092 , n56912 );
not ( n70093 , n56904 );
and ( n70094 , n70093 , n31329 );
and ( n70095 , n47449 , n56904 );
or ( n70096 , n70094 , n70095 );
and ( n70097 , n70092 , n70096 );
and ( n70098 , n47449 , n56912 );
or ( n70099 , n70097 , n70098 );
and ( n70100 , n70091 , n70099 );
not ( n70101 , n56937 );
not ( n70102 , n56939 );
and ( n70103 , n70102 , n70099 );
and ( n70104 , n47485 , n56939 );
or ( n70105 , n70103 , n70104 );
and ( n70106 , n70101 , n70105 );
and ( n70107 , n47503 , n56937 );
or ( n70108 , n70106 , n70107 );
and ( n70109 , n70108 , n31452 );
or ( n70110 , n70100 , n70109 );
and ( n70111 , n70110 , n31638 );
and ( n70112 , n31329 , n47277 );
or ( n70113 , C0 , n70081 , n70090 , n70111 , n70112 );
buf ( n70114 , n70113 );
buf ( n70115 , n70114 );
buf ( n70116 , n31655 );
buf ( n70117 , n61693 );
buf ( n70118 , n30987 );
xor ( n70119 , n39558 , n54978 );
and ( n70120 , n70119 , n33199 );
not ( n70121 , n48648 );
and ( n70122 , n70121 , n39558 );
and ( n70123 , n34365 , n48648 );
or ( n70124 , n70122 , n70123 );
and ( n70125 , n70124 , n32924 );
not ( n70126 , n48660 );
and ( n70127 , n70126 , n39558 );
not ( n70128 , n39584 );
buf ( n70129 , RI15b46e78_284);
and ( n70130 , n70128 , n70129 );
not ( n70131 , n39775 );
and ( n70132 , n70131 , n39771 );
xor ( n70133 , n39771 , n34193 );
and ( n70134 , n42650 , n42675 );
xor ( n70135 , n70133 , n70134 );
and ( n70136 , n70135 , n39775 );
or ( n70137 , n70132 , n70136 );
and ( n70138 , n70137 , n39584 );
or ( n70139 , n70130 , n70138 );
and ( n70140 , n70139 , n48660 );
or ( n70141 , n70127 , n70140 );
and ( n70142 , n70141 , n33172 );
not ( n70143 , n48730 );
and ( n70144 , n70143 , n39558 );
and ( n70145 , n56383 , n48730 );
or ( n70146 , n70144 , n70145 );
and ( n70147 , n70146 , n33187 );
and ( n70148 , n39558 , n54713 );
or ( n70149 , n70120 , n70125 , n70142 , n70147 , n70148 );
and ( n70150 , n70149 , n33208 );
and ( n70151 , n39558 , n39805 );
or ( n70152 , C0 , n70150 , n70151 );
buf ( n70153 , n70152 );
buf ( n70154 , n70153 );
buf ( n70155 , n30987 );
not ( n70156 , n41532 );
and ( n70157 , n70156 , n34431 );
and ( n70158 , n56397 , n41532 );
or ( n70159 , n70157 , n70158 );
buf ( n70160 , n70159 );
buf ( n70161 , n70160 );
buf ( n70162 , n31655 );
buf ( n70163 , n31655 );
buf ( n70164 , n30987 );
buf ( n70165 , n31655 );
buf ( n70166 , n31655 );
buf ( n70167 , n30987 );
not ( n70168 , n34150 );
and ( n70169 , n70168 , n32622 );
not ( n70170 , n58762 );
and ( n70171 , n70170 , n32622 );
and ( n70172 , n32655 , n58762 );
or ( n70173 , n70171 , n70172 );
and ( n70174 , n70173 , n34150 );
or ( n70175 , n70169 , n70174 );
and ( n70176 , n70175 , n33381 );
not ( n70177 , n58770 );
not ( n70178 , n58762 );
and ( n70179 , n70178 , n32622 );
and ( n70180 , n56044 , n58762 );
or ( n70181 , n70179 , n70180 );
and ( n70182 , n70177 , n70181 );
and ( n70183 , n56044 , n58770 );
or ( n70184 , n70182 , n70183 );
and ( n70185 , n70184 , n33375 );
not ( n70186 , n32968 );
not ( n70187 , n58770 );
not ( n70188 , n58762 );
and ( n70189 , n70188 , n32622 );
and ( n70190 , n56044 , n58762 );
or ( n70191 , n70189 , n70190 );
and ( n70192 , n70187 , n70191 );
and ( n70193 , n56044 , n58770 );
or ( n70194 , n70192 , n70193 );
and ( n70195 , n70186 , n70194 );
not ( n70196 , n58790 );
not ( n70197 , n58792 );
and ( n70198 , n70197 , n70194 );
and ( n70199 , n56068 , n58792 );
or ( n70200 , n70198 , n70199 );
and ( n70201 , n70196 , n70200 );
and ( n70202 , n56076 , n58790 );
or ( n70203 , n70201 , n70202 );
and ( n70204 , n70203 , n32968 );
or ( n70205 , n70195 , n70204 );
and ( n70206 , n70205 , n33370 );
and ( n70207 , n32622 , n35062 );
or ( n70208 , C0 , n70176 , n70185 , n70206 , n70207 );
buf ( n70209 , n70208 );
buf ( n70210 , n70209 );
buf ( n70211 , n30987 );
not ( n70212 , n48765 );
and ( n70213 , n70212 , n33220 );
and ( n70214 , n62911 , n48765 );
or ( n70215 , n70213 , n70214 );
and ( n70216 , n70215 , n33180 );
not ( n70217 , n49054 );
and ( n70218 , n70217 , n33220 );
and ( n70219 , n62922 , n49054 );
or ( n70220 , n70218 , n70219 );
and ( n70221 , n70220 , n33178 );
and ( n70222 , n33220 , n49774 );
or ( n70223 , n70216 , n70221 , n70222 );
and ( n70224 , n70223 , n33208 );
and ( n70225 , n33291 , n33375 );
not ( n70226 , n32968 );
and ( n70227 , n70226 , n33291 );
xor ( n70228 , n33220 , n59698 );
and ( n70229 , n70228 , n32968 );
or ( n70230 , n70227 , n70229 );
and ( n70231 , n70230 , n33370 );
and ( n70232 , n32983 , n35056 );
and ( n70233 , n33220 , n49794 );
or ( n70234 , C0 , n70224 , n70225 , n70231 , n70232 , n70233 );
buf ( n70235 , n70234 );
buf ( n70236 , n70235 );
buf ( n70237 , n31655 );
buf ( n70238 , n30987 );
and ( n70239 , n46030 , n32500 );
not ( n70240 , n35211 );
and ( n70241 , n70240 , n37557 );
buf ( n70242 , n70241 );
and ( n70243 , n70242 , n32421 );
not ( n70244 , n35245 );
and ( n70245 , n70244 , n37557 );
buf ( n70246 , n70245 );
and ( n70247 , n70246 , n32419 );
not ( n70248 , n35278 );
and ( n70249 , n70248 , n37557 );
not ( n70250 , n35295 );
and ( n70251 , n70250 , n49587 );
xor ( n70252 , n37557 , n49537 );
and ( n70253 , n70252 , n35295 );
or ( n70254 , n70251 , n70253 );
and ( n70255 , n70254 , n35278 );
or ( n70256 , n70249 , n70255 );
and ( n70257 , n70256 , n32417 );
not ( n70258 , n35331 );
and ( n70259 , n70258 , n37557 );
not ( n70260 , n35294 );
not ( n70261 , n45995 );
and ( n70262 , n70261 , n49587 );
xor ( n70263 , n49588 , n49623 );
and ( n70264 , n70263 , n45995 );
or ( n70265 , n70262 , n70264 );
and ( n70266 , n70260 , n70265 );
and ( n70267 , n70252 , n35294 );
or ( n70268 , n70266 , n70267 );
and ( n70269 , n70268 , n35331 );
or ( n70270 , n70259 , n70269 );
and ( n70271 , n70270 , n32415 );
and ( n70272 , n37557 , n35354 );
or ( n70273 , n70243 , n70247 , n70257 , n70271 , n70272 );
and ( n70274 , n70273 , n32456 );
not ( n70275 , n32475 );
not ( n70276 , n46060 );
and ( n70277 , n70276 , n49677 );
xor ( n70278 , n49678 , n49717 );
and ( n70279 , n70278 , n46060 );
or ( n70280 , n70277 , n70279 );
and ( n70281 , n70275 , n70280 );
and ( n70282 , n37557 , n32475 );
or ( n70283 , n70281 , n70282 );
and ( n70284 , n70283 , n32486 );
buf ( n70285 , n32489 );
and ( n70286 , n37557 , n35367 );
or ( n70287 , C0 , n70239 , n70274 , n70284 , n70285 , n70286 );
buf ( n70288 , n70287 );
buf ( n70289 , n70288 );
buf ( n70290 , n40223 );
buf ( n70291 , n30987 );
buf ( n70292 , n31655 );
buf ( n70293 , n30987 );
and ( n70294 , n33226 , n32528 );
not ( n70295 , n32598 );
and ( n70296 , n70295 , n32989 );
buf ( n70297 , n70296 );
and ( n70298 , n70297 , n32890 );
not ( n70299 , n32919 );
and ( n70300 , n70299 , n32989 );
buf ( n70301 , n70300 );
and ( n70302 , n70301 , n32924 );
not ( n70303 , n32953 );
and ( n70304 , n70303 , n32989 );
not ( n70305 , n32971 );
and ( n70306 , n70305 , n33103 );
xor ( n70307 , n32989 , n33016 );
and ( n70308 , n70307 , n32971 );
or ( n70309 , n70306 , n70308 );
and ( n70310 , n70309 , n32953 );
or ( n70311 , n70304 , n70310 );
and ( n70312 , n70311 , n33038 );
not ( n70313 , n33067 );
and ( n70314 , n70313 , n32989 );
not ( n70315 , n32970 );
not ( n70316 , n33071 );
and ( n70317 , n70316 , n33103 );
xor ( n70318 , n33104 , n33148 );
and ( n70319 , n70318 , n33071 );
or ( n70320 , n70317 , n70319 );
and ( n70321 , n70315 , n70320 );
and ( n70322 , n70307 , n32970 );
or ( n70323 , n70321 , n70322 );
and ( n70324 , n70323 , n33067 );
or ( n70325 , n70314 , n70324 );
and ( n70326 , n70325 , n33172 );
and ( n70327 , n32989 , n33204 );
or ( n70328 , n70298 , n70302 , n70312 , n70326 , n70327 );
and ( n70329 , n70328 , n33208 );
not ( n70330 , n32968 );
not ( n70331 , n33270 );
and ( n70332 , n70331 , n33303 );
xor ( n70333 , n33304 , n33348 );
and ( n70334 , n70333 , n33270 );
or ( n70335 , n70332 , n70334 );
and ( n70336 , n70330 , n70335 );
and ( n70337 , n32989 , n32968 );
or ( n70338 , n70336 , n70337 );
and ( n70339 , n70338 , n33370 );
buf ( n70340 , n35056 );
and ( n70341 , n32989 , n33382 );
or ( n70342 , C0 , n70294 , n70329 , n70339 , n70340 , n70341 );
buf ( n70343 , n70342 );
buf ( n70344 , n70343 );
not ( n70345 , n31728 );
and ( n70346 , n70345 , n46024 );
and ( n70347 , n63455 , n31728 );
or ( n70348 , n70346 , n70347 );
and ( n70349 , n70348 , n32253 );
not ( n70350 , n32283 );
and ( n70351 , n70350 , n46024 );
and ( n70352 , n63466 , n32283 );
or ( n70353 , n70351 , n70352 );
and ( n70354 , n70353 , n32398 );
and ( n70355 , n46024 , n32436 );
or ( n70356 , n70349 , n70354 , n70355 );
and ( n70357 , n70356 , n32456 );
and ( n70358 , n49665 , n32473 );
not ( n70359 , n32475 );
and ( n70360 , n70359 , n49665 );
xor ( n70361 , n46024 , n47762 );
and ( n70362 , n70361 , n32475 );
or ( n70363 , n70360 , n70362 );
and ( n70364 , n70363 , n32486 );
and ( n70365 , n37545 , n32489 );
and ( n70366 , n46024 , n32501 );
or ( n70367 , C0 , n70357 , n70358 , n70364 , n70365 , n70366 );
buf ( n70368 , n70367 );
buf ( n70369 , n70368 );
buf ( n70370 , n30987 );
buf ( n70371 , n31655 );
buf ( n70372 , n31655 );
not ( n70373 , n34150 );
and ( n70374 , n70373 , n32723 );
not ( n70375 , n56708 );
and ( n70376 , n70375 , n32723 );
and ( n70377 , n32755 , n56708 );
or ( n70378 , n70376 , n70377 );
and ( n70379 , n70378 , n34150 );
or ( n70380 , n70374 , n70379 );
and ( n70381 , n70380 , n33381 );
not ( n70382 , n56716 );
not ( n70383 , n56708 );
and ( n70384 , n70383 , n32723 );
and ( n70385 , n35083 , n56708 );
or ( n70386 , n70384 , n70385 );
and ( n70387 , n70382 , n70386 );
and ( n70388 , n35083 , n56716 );
or ( n70389 , n70387 , n70388 );
and ( n70390 , n70389 , n33375 );
not ( n70391 , n32968 );
not ( n70392 , n56716 );
not ( n70393 , n56708 );
and ( n70394 , n70393 , n32723 );
and ( n70395 , n35083 , n56708 );
or ( n70396 , n70394 , n70395 );
and ( n70397 , n70392 , n70396 );
and ( n70398 , n35083 , n56716 );
or ( n70399 , n70397 , n70398 );
and ( n70400 , n70391 , n70399 );
not ( n70401 , n56736 );
not ( n70402 , n56738 );
and ( n70403 , n70402 , n70399 );
and ( n70404 , n35107 , n56738 );
or ( n70405 , n70403 , n70404 );
and ( n70406 , n70401 , n70405 );
and ( n70407 , n35115 , n56736 );
or ( n70408 , n70406 , n70407 );
and ( n70409 , n70408 , n32968 );
or ( n70410 , n70400 , n70409 );
and ( n70411 , n70410 , n33370 );
and ( n70412 , n32723 , n35062 );
or ( n70413 , C0 , n70381 , n70390 , n70411 , n70412 );
buf ( n70414 , n70413 );
buf ( n70415 , n70414 );
buf ( n70416 , n30987 );
buf ( n70417 , n31655 );
buf ( n70418 , n31655 );
buf ( n70419 , n30987 );
buf ( n70420 , n30987 );
or ( n70421 , n31647 , n31649 );
or ( n70422 , n70421 , n31007 );
and ( n70423 , n54792 , n70422 );
not ( n70424 , n31451 );
and ( n70425 , n54792 , n70424 );
and ( n70426 , n70425 , n31645 );
not ( n70427 , n31077 );
and ( n70428 , n70427 , n54792 );
not ( n70429 , n31447 );
buf ( n70430 , n70429 );
and ( n70431 , n31450 , n31447 );
or ( n70432 , n70430 , n70431 );
and ( n70433 , n70432 , n31077 );
or ( n70434 , n70428 , n70433 );
and ( n70435 , n70434 , n31373 );
not ( n70436 , n31402 );
and ( n70437 , n70436 , n54792 );
and ( n70438 , n31450 , n31402 );
or ( n70439 , n70437 , n70438 );
and ( n70440 , n70439 , n31408 );
not ( n70441 , n31437 );
and ( n70442 , n70441 , n54792 );
not ( n70443 , n44703 );
buf ( n70444 , n70443 );
and ( n70445 , n31453 , n44703 );
or ( n70446 , n70444 , n70445 );
and ( n70447 , n70446 , n31437 );
or ( n70448 , n70442 , n70447 );
and ( n70449 , n70448 , n31468 );
not ( n70450 , n31497 );
and ( n70451 , n70450 , n54792 );
not ( n70452 , n31451 );
buf ( n70453 , n70452 );
buf ( n70454 , n70453 );
and ( n70455 , n70454 , n31497 );
or ( n70456 , n70451 , n70455 );
and ( n70457 , n70456 , n31521 );
and ( n70458 , n54792 , n31553 );
or ( n70459 , n70435 , n70440 , n70449 , n70457 , n70458 );
and ( n70460 , n70459 , n31557 );
or ( n70461 , n52896 , n31641 );
buf ( n70462 , n70461 );
or ( n70463 , C0 , n70423 , n70426 , n70460 , C0 , n70462 );
buf ( n70464 , n70463 );
buf ( n70465 , n70464 );
not ( n70466 , n40163 );
and ( n70467 , n70466 , n31838 );
not ( n70468 , n52903 );
and ( n70469 , n70468 , n31838 );
and ( n70470 , n32235 , n52903 );
or ( n70471 , n70469 , n70470 );
and ( n70472 , n70471 , n40163 );
or ( n70473 , n70467 , n70472 );
and ( n70474 , n70473 , n32498 );
not ( n70475 , n52911 );
not ( n70476 , n52903 );
and ( n70477 , n70476 , n31838 );
and ( n70478 , n42188 , n52903 );
or ( n70479 , n70477 , n70478 );
and ( n70480 , n70475 , n70479 );
and ( n70481 , n42188 , n52911 );
or ( n70482 , n70480 , n70481 );
and ( n70483 , n70482 , n32473 );
not ( n70484 , n32475 );
not ( n70485 , n52911 );
not ( n70486 , n52903 );
and ( n70487 , n70486 , n31838 );
and ( n70488 , n42188 , n52903 );
or ( n70489 , n70487 , n70488 );
and ( n70490 , n70485 , n70489 );
and ( n70491 , n42188 , n52911 );
or ( n70492 , n70490 , n70491 );
and ( n70493 , n70484 , n70492 );
not ( n70494 , n52931 );
not ( n70495 , n52933 );
and ( n70496 , n70495 , n70492 );
and ( n70497 , n42216 , n52933 );
or ( n70498 , n70496 , n70497 );
and ( n70499 , n70494 , n70498 );
and ( n70500 , n42224 , n52931 );
or ( n70501 , n70499 , n70500 );
and ( n70502 , n70501 , n32475 );
or ( n70503 , n70493 , n70502 );
and ( n70504 , n70503 , n32486 );
and ( n70505 , n31838 , n41278 );
or ( n70506 , C0 , n70474 , n70483 , n70504 , n70505 );
buf ( n70507 , n70506 );
buf ( n70508 , n70507 );
buf ( n70509 , n30987 );
buf ( n70510 , n31655 );
buf ( n70511 , n31655 );
buf ( n70512 , n30987 );
buf ( n70513 , n30987 );
buf ( n70514 , n31655 );
and ( n70515 , n49076 , n48639 );
not ( n70516 , n48642 );
and ( n70517 , n70516 , n48601 );
and ( n70518 , n49076 , n48642 );
or ( n70519 , n70517 , n70518 );
and ( n70520 , n70519 , n32890 );
not ( n70521 , n48648 );
and ( n70522 , n70521 , n48601 );
and ( n70523 , n49076 , n48648 );
or ( n70524 , n70522 , n70523 );
and ( n70525 , n70524 , n32924 );
not ( n70526 , n48654 );
and ( n70527 , n70526 , n48601 );
and ( n70528 , n49076 , n48654 );
or ( n70529 , n70527 , n70528 );
and ( n70530 , n70529 , n33038 );
not ( n70531 , n48660 );
and ( n70532 , n70531 , n48601 );
and ( n70533 , n49076 , n48660 );
or ( n70534 , n70532 , n70533 );
and ( n70535 , n70534 , n33172 );
not ( n70536 , n41576 );
and ( n70537 , n70536 , n48601 );
and ( n70538 , n48786 , n41576 );
or ( n70539 , n70537 , n70538 );
and ( n70540 , n70539 , n33189 );
not ( n70541 , n48730 );
and ( n70542 , n70541 , n48601 );
and ( n70543 , n48786 , n48730 );
or ( n70544 , n70542 , n70543 );
and ( n70545 , n70544 , n33187 );
not ( n70546 , n48765 );
and ( n70547 , n70546 , n48601 );
xor ( n70548 , n48786 , n49002 );
and ( n70549 , n70548 , n48765 );
or ( n70550 , n70547 , n70549 );
and ( n70551 , n70550 , n33180 );
not ( n70552 , n49054 );
and ( n70553 , n70552 , n48601 );
not ( n70554 , n48845 );
xor ( n70555 , n49076 , n49116 );
and ( n70556 , n70554 , n70555 );
xnor ( n70557 , n49185 , n49242 );
and ( n70558 , n70557 , n48845 );
or ( n70559 , n70556 , n70558 );
and ( n70560 , n70559 , n49054 );
or ( n70561 , n70553 , n70560 );
and ( n70562 , n70561 , n33178 );
and ( n70563 , n49185 , n49275 );
or ( n70564 , n70515 , n70520 , n70525 , n70530 , n70535 , n70540 , n70545 , n70551 , n70562 , n70563 );
and ( n70565 , n70564 , n33208 );
and ( n70566 , n32994 , n35056 );
and ( n70567 , n48601 , n49286 );
or ( n70568 , C0 , n70565 , n70566 , n70567 );
buf ( n70569 , n70568 );
buf ( n70570 , n70569 );
buf ( n70571 , n30987 );
buf ( n70572 , n30987 );
and ( n70573 , n31563 , n31007 );
not ( n70574 , n31077 );
and ( n70575 , n70574 , n35389 );
buf ( n70576 , n70575 );
and ( n70577 , n70576 , n31373 );
not ( n70578 , n31402 );
and ( n70579 , n70578 , n35389 );
buf ( n70580 , n70579 );
and ( n70581 , n70580 , n31408 );
not ( n70582 , n31437 );
and ( n70583 , n70582 , n35389 );
not ( n70584 , n31455 );
and ( n70585 , n70584 , n35427 );
xor ( n70586 , n35389 , n35409 );
and ( n70587 , n70586 , n31455 );
or ( n70588 , n70585 , n70587 );
and ( n70589 , n70588 , n31437 );
or ( n70590 , n70583 , n70589 );
and ( n70591 , n70590 , n31468 );
not ( n70592 , n31497 );
and ( n70593 , n70592 , n35389 );
not ( n70594 , n31454 );
not ( n70595 , n31501 );
and ( n70596 , n70595 , n35427 );
xor ( n70597 , n35428 , n35459 );
and ( n70598 , n70597 , n31501 );
or ( n70599 , n70596 , n70598 );
and ( n70600 , n70594 , n70599 );
and ( n70601 , n70586 , n31454 );
or ( n70602 , n70600 , n70601 );
and ( n70603 , n70602 , n31497 );
or ( n70604 , n70593 , n70603 );
and ( n70605 , n70604 , n31521 );
and ( n70606 , n35389 , n31553 );
or ( n70607 , n70577 , n70581 , n70591 , n70605 , n70606 );
and ( n70608 , n70607 , n31557 );
not ( n70609 , n31452 );
not ( n70610 , n31619 );
and ( n70611 , n70610 , n35482 );
xor ( n70612 , n35483 , n35513 );
and ( n70613 , n70612 , n31619 );
or ( n70614 , n70611 , n70613 );
and ( n70615 , n70609 , n70614 );
and ( n70616 , n35389 , n31452 );
or ( n70617 , n70615 , n70616 );
and ( n70618 , n70617 , n31638 );
and ( n70619 , n35389 , n31650 );
or ( n70620 , C0 , n70573 , n70608 , n70618 , C0 , n70619 );
buf ( n70621 , n70620 );
buf ( n70622 , n70621 );
buf ( n70623 , n31655 );
buf ( n70624 , n31655 );
not ( n70625 , n33419 );
and ( n70626 , n70625 , n31581 );
xor ( n70627 , n33475 , n33690 );
and ( n70628 , n70627 , n33419 );
or ( n70629 , n70626 , n70628 );
and ( n70630 , n70629 , n31529 );
not ( n70631 , n33734 );
and ( n70632 , n70631 , n31581 );
not ( n70633 , n33533 );
xor ( n70634 , n33768 , n33808 );
and ( n70635 , n70633 , n70634 );
xnor ( n70636 , n33853 , n33910 );
and ( n70637 , n70636 , n33533 );
or ( n70638 , n70635 , n70637 );
and ( n70639 , n70638 , n33734 );
or ( n70640 , n70632 , n70639 );
and ( n70641 , n70640 , n31527 );
and ( n70642 , n31581 , n33942 );
or ( n70643 , n70630 , n70641 , n70642 );
and ( n70644 , n70643 , n31557 );
and ( n70645 , n34107 , n31643 );
not ( n70646 , n31452 );
and ( n70647 , n70646 , n34107 );
xor ( n70648 , n31581 , n33956 );
and ( n70649 , n70648 , n31452 );
or ( n70650 , n70647 , n70649 );
and ( n70651 , n70650 , n31638 );
and ( n70652 , n34005 , n33973 );
and ( n70653 , n31581 , n33978 );
or ( n70654 , C0 , n70644 , n70645 , n70651 , n70652 , n70653 );
buf ( n70655 , n70654 );
buf ( n70656 , n70655 );
buf ( n70657 , n31655 );
buf ( n70658 , n30987 );
not ( n70659 , n32953 );
buf ( n70660 , RI15b46590_265);
and ( n70661 , n70659 , n70660 );
not ( n70662 , n54581 );
and ( n70663 , n70662 , n54526 );
xor ( n70664 , n54526 , n54340 );
and ( n70665 , n67514 , n67515 );
xor ( n70666 , n70664 , n70665 );
and ( n70667 , n70666 , n54581 );
or ( n70668 , n70663 , n70667 );
and ( n70669 , n70668 , n32953 );
or ( n70670 , n70661 , n70669 );
and ( n70671 , n70670 , n33038 );
not ( n70672 , n48660 );
and ( n70673 , n70672 , n70660 );
not ( n70674 , n55168 );
and ( n70675 , n70674 , n55128 );
xor ( n70676 , n55128 , n34193 );
and ( n70677 , n67526 , n67527 );
xor ( n70678 , n70676 , n70677 );
and ( n70679 , n70678 , n55168 );
or ( n70680 , n70675 , n70679 );
and ( n70681 , n70680 , n48660 );
or ( n70682 , n70673 , n70681 );
and ( n70683 , n70682 , n33172 );
and ( n70684 , n70660 , n39795 );
or ( n70685 , n70671 , n70683 , n70684 );
and ( n70686 , n70685 , n33208 );
and ( n70687 , n70660 , n39805 );
or ( n70688 , C0 , n70686 , n70687 );
buf ( n70689 , n70688 );
buf ( n70690 , n70689 );
buf ( n70691 , n30987 );
buf ( n70692 , n31655 );
not ( n70693 , n31451 );
and ( n70694 , n70693 , n30994 );
buf ( n70695 , n31451 );
or ( n70696 , n70694 , n70695 );
and ( n70697 , n70696 , n31645 );
not ( n70698 , n63845 );
not ( n70699 , n63847 );
and ( n70700 , n70699 , n30994 );
buf ( n70701 , n63847 );
or ( n70702 , n70700 , n70701 );
and ( n70703 , n70702 , n31468 );
and ( n70704 , n30994 , n63859 );
or ( n70705 , n70703 , n70704 );
and ( n70706 , n70698 , n70705 );
buf ( n70707 , n63845 );
or ( n70708 , n70706 , n70707 );
and ( n70709 , n70708 , n31557 );
buf ( n70710 , n31643 );
not ( n70711 , n59060 );
and ( n70712 , n70711 , n31641 );
and ( n70713 , n31452 , n31638 );
or ( n70714 , C0 , C0 , C0 , n70697 , n70709 , n70710 , n70712 , n70713 , C0 , C0 );
buf ( n70715 , n70714 );
buf ( n70716 , n70715 );
buf ( n70717 , n31655 );
buf ( n70718 , n30987 );
not ( n70719 , n38443 );
and ( n70720 , n70719 , n38065 );
xor ( n70721 , n53478 , n53491 );
and ( n70722 , n70721 , n38443 );
or ( n70723 , n70720 , n70722 );
and ( n70724 , n70723 , n38450 );
not ( n70725 , n39339 );
and ( n70726 , n70725 , n38965 );
xor ( n70727 , n53534 , n53547 );
and ( n70728 , n70727 , n39339 );
or ( n70729 , n70726 , n70728 );
and ( n70730 , n70729 , n39346 );
and ( n70731 , n40206 , n39359 );
or ( n70732 , n70724 , n70730 , n70731 );
buf ( n70733 , n70732 );
buf ( n70734 , n70733 );
buf ( n70735 , n31655 );
not ( n70736 , n50828 );
not ( n70737 , n50834 );
and ( n70738 , n70737 , n40470 );
and ( n70739 , n62428 , n50834 );
or ( n70740 , n70738 , n70739 );
and ( n70741 , n70736 , n70740 );
buf ( n70742 , RI15b5fe50_1137);
and ( n70743 , n70742 , n50828 );
or ( n70744 , n70741 , n70743 );
buf ( n70745 , n70744 );
buf ( n70746 , n70745 );
buf ( n70747 , n30987 );
buf ( n70748 , n30987 );
xor ( n70749 , n33085 , n58391 );
and ( n70750 , n70749 , n33201 );
not ( n70751 , n41576 );
and ( n70752 , n70751 , n33085 );
xor ( n70753 , n58557 , n58592 );
and ( n70754 , n70753 , n41576 );
or ( n70755 , n70752 , n70754 );
and ( n70756 , n70755 , n33189 );
and ( n70757 , n33085 , n41592 );
or ( n70758 , n70750 , n70756 , n70757 );
and ( n70759 , n70758 , n33208 );
and ( n70760 , n33085 , n39805 );
or ( n70761 , C0 , n70759 , n70760 );
buf ( n70762 , n70761 );
buf ( n70763 , n70762 );
buf ( n70764 , n31655 );
buf ( n70765 , n31655 );
buf ( n70766 , n30987 );
not ( n70767 , n31437 );
and ( n70768 , n70767 , n50596 );
not ( n70769 , n41809 );
and ( n70770 , n70769 , n41623 );
xor ( n70771 , n41819 , n41821 );
and ( n70772 , n70771 , n41809 );
or ( n70773 , n70770 , n70772 );
and ( n70774 , n70773 , n31437 );
or ( n70775 , n70768 , n70774 );
and ( n70776 , n70775 , n31468 );
not ( n70777 , n41837 );
and ( n70778 , n70777 , n50596 );
and ( n70779 , n50602 , n41837 );
or ( n70780 , n70778 , n70779 );
and ( n70781 , n70780 , n31521 );
and ( n70782 , n50596 , n42158 );
or ( n70783 , n70776 , n70781 , n70782 );
and ( n70784 , n70783 , n31557 );
and ( n70785 , n50596 , n40154 );
or ( n70786 , C0 , n70784 , n70785 );
buf ( n70787 , n70786 );
buf ( n70788 , n70787 );
not ( n70789 , n40163 );
and ( n70790 , n70789 , n31861 );
not ( n70791 , n56988 );
and ( n70792 , n70791 , n31861 );
and ( n70793 , n32218 , n56988 );
or ( n70794 , n70792 , n70793 );
and ( n70795 , n70794 , n40163 );
or ( n70796 , n70790 , n70795 );
and ( n70797 , n70796 , n32498 );
not ( n70798 , n56996 );
not ( n70799 , n56988 );
and ( n70800 , n70799 , n31861 );
and ( n70801 , n42255 , n56988 );
or ( n70802 , n70800 , n70801 );
and ( n70803 , n70798 , n70802 );
and ( n70804 , n42255 , n56996 );
or ( n70805 , n70803 , n70804 );
and ( n70806 , n70805 , n32473 );
not ( n70807 , n32475 );
not ( n70808 , n56996 );
not ( n70809 , n56988 );
and ( n70810 , n70809 , n31861 );
and ( n70811 , n42255 , n56988 );
or ( n70812 , n70810 , n70811 );
and ( n70813 , n70808 , n70812 );
and ( n70814 , n42255 , n56996 );
or ( n70815 , n70813 , n70814 );
and ( n70816 , n70807 , n70815 );
not ( n70817 , n57016 );
not ( n70818 , n57018 );
and ( n70819 , n70818 , n70815 );
and ( n70820 , n42283 , n57018 );
or ( n70821 , n70819 , n70820 );
and ( n70822 , n70817 , n70821 );
and ( n70823 , n42291 , n57016 );
or ( n70824 , n70822 , n70823 );
and ( n70825 , n70824 , n32475 );
or ( n70826 , n70816 , n70825 );
and ( n70827 , n70826 , n32486 );
and ( n70828 , n31861 , n41278 );
or ( n70829 , C0 , n70797 , n70806 , n70827 , n70828 );
buf ( n70830 , n70829 );
buf ( n70831 , n70830 );
buf ( n70832 , n30987 );
buf ( n70833 , n30987 );
buf ( n70834 , n31655 );
buf ( n70835 , n31655 );
and ( n70836 , n65075 , n33377 );
not ( n70837 , n48545 );
buf ( n70838 , RI15b47aa8_310);
and ( n70839 , n70837 , n70838 );
buf ( n70840 , n70839 );
and ( n70841 , n70840 , n32890 );
not ( n70842 , n48557 );
and ( n70843 , n70842 , n70838 );
and ( n70844 , n65083 , n48557 );
or ( n70845 , n70843 , n70844 );
and ( n70846 , n70845 , n33038 );
and ( n70847 , n70838 , n48571 );
or ( n70848 , n70841 , n70846 , n70847 );
and ( n70849 , n70848 , n33208 );
and ( n70850 , n70838 , n48577 );
or ( n70851 , C0 , n70836 , n70849 , n70850 );
buf ( n70852 , n70851 );
buf ( n70853 , n70852 );
buf ( n70854 , n31655 );
buf ( n70855 , n30987 );
buf ( n70856 , n30987 );
and ( n70857 , n49068 , n48639 );
not ( n70858 , n48642 );
and ( n70859 , n70858 , n48593 );
and ( n70860 , n49068 , n48642 );
or ( n70861 , n70859 , n70860 );
and ( n70862 , n70861 , n32890 );
not ( n70863 , n48648 );
and ( n70864 , n70863 , n48593 );
and ( n70865 , n49068 , n48648 );
or ( n70866 , n70864 , n70865 );
and ( n70867 , n70866 , n32924 );
not ( n70868 , n48654 );
and ( n70869 , n70868 , n48593 );
and ( n70870 , n49068 , n48654 );
or ( n70871 , n70869 , n70870 );
and ( n70872 , n70871 , n33038 );
not ( n70873 , n48660 );
and ( n70874 , n70873 , n48593 );
and ( n70875 , n49068 , n48660 );
or ( n70876 , n70874 , n70875 );
and ( n70877 , n70876 , n33172 );
not ( n70878 , n41576 );
and ( n70879 , n70878 , n48593 );
and ( n70880 , n48778 , n41576 );
or ( n70881 , n70879 , n70880 );
and ( n70882 , n70881 , n33189 );
not ( n70883 , n48730 );
and ( n70884 , n70883 , n48593 );
and ( n70885 , n48778 , n48730 );
or ( n70886 , n70884 , n70885 );
and ( n70887 , n70886 , n33187 );
not ( n70888 , n48765 );
and ( n70889 , n70888 , n48593 );
xor ( n70890 , n48778 , n49010 );
and ( n70891 , n70890 , n48765 );
or ( n70892 , n70889 , n70891 );
and ( n70893 , n70892 , n33180 );
not ( n70894 , n49054 );
and ( n70895 , n70894 , n48593 );
not ( n70896 , n48845 );
xor ( n70897 , n49068 , n49124 );
and ( n70898 , n70896 , n70897 );
xnor ( n70899 , n49177 , n49250 );
and ( n70900 , n70899 , n48845 );
or ( n70901 , n70898 , n70900 );
and ( n70902 , n70901 , n49054 );
or ( n70903 , n70895 , n70902 );
and ( n70904 , n70903 , n33178 );
and ( n70905 , n49177 , n49275 );
or ( n70906 , n70857 , n70862 , n70867 , n70872 , n70877 , n70882 , n70887 , n70893 , n70904 , n70905 );
and ( n70907 , n70906 , n33208 );
and ( n70908 , n32986 , n35056 );
and ( n70909 , n48593 , n49286 );
or ( n70910 , C0 , n70907 , n70908 , n70909 );
buf ( n70911 , n70910 );
buf ( n70912 , n70911 );
buf ( n70913 , n31655 );
buf ( n70914 , n30987 );
not ( n70915 , n40163 );
and ( n70916 , n70915 , n32011 );
not ( n70917 , n45227 );
and ( n70918 , n70917 , n32011 );
and ( n70919 , n32147 , n45227 );
or ( n70920 , n70918 , n70919 );
and ( n70921 , n70920 , n40163 );
or ( n70922 , n70916 , n70921 );
and ( n70923 , n70922 , n32498 );
not ( n70924 , n45235 );
not ( n70925 , n45227 );
and ( n70926 , n70925 , n32011 );
and ( n70927 , n49314 , n45227 );
or ( n70928 , n70926 , n70927 );
and ( n70929 , n70924 , n70928 );
and ( n70930 , n49314 , n45235 );
or ( n70931 , n70929 , n70930 );
and ( n70932 , n70931 , n32473 );
not ( n70933 , n32475 );
not ( n70934 , n45235 );
not ( n70935 , n45227 );
and ( n70936 , n70935 , n32011 );
and ( n70937 , n49314 , n45227 );
or ( n70938 , n70936 , n70937 );
and ( n70939 , n70934 , n70938 );
and ( n70940 , n49314 , n45235 );
or ( n70941 , n70939 , n70940 );
and ( n70942 , n70933 , n70941 );
not ( n70943 , n45255 );
not ( n70944 , n45257 );
and ( n70945 , n70944 , n70941 );
and ( n70946 , n49340 , n45257 );
or ( n70947 , n70945 , n70946 );
and ( n70948 , n70943 , n70947 );
and ( n70949 , n49348 , n45255 );
or ( n70950 , n70948 , n70949 );
and ( n70951 , n70950 , n32475 );
or ( n70952 , n70942 , n70951 );
and ( n70953 , n70952 , n32486 );
and ( n70954 , n32011 , n41278 );
or ( n70955 , C0 , n70923 , n70932 , n70953 , n70954 );
buf ( n70956 , n70955 );
buf ( n70957 , n70956 );
and ( n70958 , n65746 , n31645 );
not ( n70959 , n45274 );
and ( n70960 , n70959 , n61591 );
buf ( n70961 , n70960 );
and ( n70962 , n70961 , n31373 );
not ( n70963 , n45280 );
and ( n70964 , n70963 , n61591 );
and ( n70965 , n65752 , n45280 );
or ( n70966 , n70964 , n70965 );
and ( n70967 , n70966 , n31468 );
and ( n70968 , n61591 , n45802 );
or ( n70969 , n70962 , n70967 , n70968 );
and ( n70970 , n70969 , n31557 );
and ( n70971 , n61591 , n45808 );
or ( n70972 , C0 , n70958 , n70970 , n70971 );
buf ( n70973 , n70972 );
buf ( n70974 , n70973 );
buf ( n70975 , n30987 );
buf ( n70976 , n31655 );
buf ( n70977 , n30987 );
buf ( n70978 , n30987 );
buf ( n70979 , n31655 );
and ( n70980 , n67510 , n33377 );
not ( n70981 , n48545 );
buf ( n70982 , RI15b47b20_311);
and ( n70983 , n70981 , n70982 );
buf ( n70984 , n70983 );
and ( n70985 , n70984 , n32890 );
not ( n70986 , n48557 );
and ( n70987 , n70986 , n70982 );
and ( n70988 , n67518 , n48557 );
or ( n70989 , n70987 , n70988 );
and ( n70990 , n70989 , n33038 );
and ( n70991 , n70982 , n48571 );
or ( n70992 , n70985 , n70990 , n70991 );
and ( n70993 , n70992 , n33208 );
and ( n70994 , n70982 , n48577 );
or ( n70995 , C0 , n70980 , n70993 , n70994 );
buf ( n70996 , n70995 );
buf ( n70997 , n70996 );
buf ( n70998 , n31655 );
xor ( n70999 , n49583 , n60314 );
and ( n71000 , n70999 , n32433 );
not ( n71001 , n47331 );
and ( n71002 , n71001 , n49583 );
and ( n71003 , n31931 , n60510 );
and ( n71004 , n31933 , n60512 );
and ( n71005 , n31935 , n60514 );
and ( n71006 , n31937 , n60516 );
and ( n71007 , n31939 , n60518 );
and ( n71008 , n31941 , n60520 );
and ( n71009 , n31943 , n60522 );
and ( n71010 , n31945 , n60524 );
and ( n71011 , n31947 , n60526 );
and ( n71012 , n31949 , n60528 );
and ( n71013 , n31951 , n60530 );
and ( n71014 , n31953 , n60532 );
and ( n71015 , n31955 , n60534 );
and ( n71016 , n31957 , n60536 );
and ( n71017 , n31959 , n60538 );
and ( n71018 , n31961 , n60540 );
or ( n71019 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 );
and ( n71020 , n71019 , n47331 );
or ( n71021 , n71002 , n71020 );
and ( n71022 , n71021 , n32413 );
and ( n71023 , n49583 , n47402 );
or ( n71024 , n71000 , n71022 , n71023 );
and ( n71025 , n71024 , n32456 );
and ( n71026 , n49583 , n47409 );
or ( n71027 , C0 , n71025 , n71026 );
buf ( n71028 , n71027 );
buf ( n71029 , n71028 );
buf ( n71030 , n31655 );
buf ( n71031 , n30987 );
buf ( n71032 , n30987 );
buf ( n71033 , n31655 );
not ( n71034 , n46356 );
and ( n71035 , n71034 , n31302 );
not ( n71036 , n61975 );
and ( n71037 , n71036 , n31302 );
and ( n71038 , n31306 , n61975 );
or ( n71039 , n71037 , n71038 );
and ( n71040 , n71039 , n46356 );
or ( n71041 , n71035 , n71040 );
and ( n71042 , n71041 , n31649 );
not ( n71043 , n61983 );
not ( n71044 , n61975 );
and ( n71045 , n71044 , n31302 );
and ( n71046 , n58061 , n61975 );
or ( n71047 , n71045 , n71046 );
and ( n71048 , n71043 , n71047 );
and ( n71049 , n58061 , n61983 );
or ( n71050 , n71048 , n71049 );
and ( n71051 , n71050 , n31643 );
not ( n71052 , n31452 );
not ( n71053 , n61983 );
not ( n71054 , n61975 );
and ( n71055 , n71054 , n31302 );
and ( n71056 , n58061 , n61975 );
or ( n71057 , n71055 , n71056 );
and ( n71058 , n71053 , n71057 );
and ( n71059 , n58061 , n61983 );
or ( n71060 , n71058 , n71059 );
and ( n71061 , n71052 , n71060 );
not ( n71062 , n62003 );
not ( n71063 , n62005 );
and ( n71064 , n71063 , n71060 );
and ( n71065 , n58085 , n62005 );
or ( n71066 , n71064 , n71065 );
and ( n71067 , n71062 , n71066 );
and ( n71068 , n58093 , n62003 );
or ( n71069 , n71067 , n71068 );
and ( n71070 , n71069 , n31452 );
or ( n71071 , n71061 , n71070 );
and ( n71072 , n71071 , n31638 );
and ( n71073 , n31302 , n47277 );
or ( n71074 , C0 , n71042 , n71051 , n71072 , n71073 );
buf ( n71075 , n71074 );
buf ( n71076 , n71075 );
not ( n71077 , n34150 );
and ( n71078 , n71077 , n32694 );
not ( n71079 , n60126 );
and ( n71080 , n71079 , n32694 );
and ( n71081 , n32722 , n60126 );
or ( n71082 , n71080 , n71081 );
and ( n71083 , n71082 , n34150 );
or ( n71084 , n71078 , n71083 );
and ( n71085 , n71084 , n33381 );
not ( n71086 , n60134 );
not ( n71087 , n60126 );
and ( n71088 , n71087 , n32694 );
and ( n71089 , n42565 , n60126 );
or ( n71090 , n71088 , n71089 );
and ( n71091 , n71086 , n71090 );
and ( n71092 , n42565 , n60134 );
or ( n71093 , n71091 , n71092 );
and ( n71094 , n71093 , n33375 );
not ( n71095 , n32968 );
not ( n71096 , n60134 );
not ( n71097 , n60126 );
and ( n71098 , n71097 , n32694 );
and ( n71099 , n42565 , n60126 );
or ( n71100 , n71098 , n71099 );
and ( n71101 , n71096 , n71100 );
and ( n71102 , n42565 , n60134 );
or ( n71103 , n71101 , n71102 );
and ( n71104 , n71095 , n71103 );
not ( n71105 , n60154 );
not ( n71106 , n60156 );
and ( n71107 , n71106 , n71103 );
and ( n71108 , n42589 , n60156 );
or ( n71109 , n71107 , n71108 );
and ( n71110 , n71105 , n71109 );
and ( n71111 , n42597 , n60154 );
or ( n71112 , n71110 , n71111 );
and ( n71113 , n71112 , n32968 );
or ( n71114 , n71104 , n71113 );
and ( n71115 , n71114 , n33370 );
and ( n71116 , n32694 , n35062 );
or ( n71117 , C0 , n71085 , n71094 , n71115 , n71116 );
buf ( n71118 , n71117 );
buf ( n71119 , n71118 );
buf ( n71120 , n30987 );
buf ( n71121 , n31655 );
buf ( n71122 , n31655 );
buf ( n71123 , n30987 );
buf ( n71124 , n31655 );
buf ( n71125 , n30987 );
and ( n71126 , n33217 , n32528 );
not ( n71127 , n32598 );
and ( n71128 , n71127 , n32980 );
buf ( n71129 , n71128 );
and ( n71130 , n71129 , n32890 );
not ( n71131 , n32919 );
and ( n71132 , n71131 , n32980 );
buf ( n71133 , n71132 );
and ( n71134 , n71133 , n32924 );
not ( n71135 , n32953 );
and ( n71136 , n71135 , n32980 );
not ( n71137 , n32971 );
and ( n71138 , n71137 , n33085 );
xor ( n71139 , n32980 , n33025 );
and ( n71140 , n71139 , n32971 );
or ( n71141 , n71138 , n71140 );
and ( n71142 , n71141 , n32953 );
or ( n71143 , n71136 , n71142 );
and ( n71144 , n71143 , n33038 );
not ( n71145 , n33067 );
and ( n71146 , n71145 , n32980 );
not ( n71147 , n32970 );
not ( n71148 , n33071 );
and ( n71149 , n71148 , n33085 );
xor ( n71150 , n33086 , n33157 );
and ( n71151 , n71150 , n33071 );
or ( n71152 , n71149 , n71151 );
and ( n71153 , n71147 , n71152 );
and ( n71154 , n71139 , n32970 );
or ( n71155 , n71153 , n71154 );
and ( n71156 , n71155 , n33067 );
or ( n71157 , n71146 , n71156 );
and ( n71158 , n71157 , n33172 );
and ( n71159 , n32980 , n33204 );
or ( n71160 , n71130 , n71134 , n71144 , n71158 , n71159 );
and ( n71161 , n71160 , n33208 );
not ( n71162 , n32968 );
not ( n71163 , n33270 );
and ( n71164 , n71163 , n33285 );
xor ( n71165 , n33286 , n33357 );
and ( n71166 , n71165 , n33270 );
or ( n71167 , n71164 , n71166 );
and ( n71168 , n71162 , n71167 );
and ( n71169 , n32980 , n32968 );
or ( n71170 , n71168 , n71169 );
and ( n71171 , n71170 , n33370 );
and ( n71172 , n32980 , n33382 );
or ( n71173 , C0 , n71126 , n71161 , n71171 , C0 , n71172 );
buf ( n71174 , n71173 );
buf ( n71175 , n71174 );
buf ( n71176 , n30987 );
buf ( n71177 , n31655 );
not ( n71178 , n31728 );
and ( n71179 , n71178 , n46033 );
xor ( n71180 , n47610 , n47619 );
and ( n71181 , n71180 , n31728 );
or ( n71182 , n71179 , n71181 );
and ( n71183 , n71182 , n32253 );
not ( n71184 , n32283 );
and ( n71185 , n71184 , n46033 );
not ( n71186 , n31823 );
xor ( n71187 , n47665 , n47674 );
and ( n71188 , n71186 , n71187 );
xnor ( n71189 , n47715 , n47724 );
and ( n71190 , n71189 , n31823 );
or ( n71191 , n71188 , n71190 );
and ( n71192 , n71191 , n32283 );
or ( n71193 , n71185 , n71192 );
and ( n71194 , n71193 , n32398 );
and ( n71195 , n46033 , n32436 );
or ( n71196 , n71183 , n71194 , n71195 );
and ( n71197 , n71196 , n32456 );
and ( n71198 , n49683 , n32473 );
not ( n71199 , n32475 );
and ( n71200 , n71199 , n49683 );
xor ( n71201 , n46033 , n47753 );
and ( n71202 , n71201 , n32475 );
or ( n71203 , n71200 , n71202 );
and ( n71204 , n71203 , n32486 );
and ( n71205 , n37563 , n32489 );
and ( n71206 , n46033 , n32501 );
or ( n71207 , C0 , n71197 , n71198 , n71204 , n71205 , n71206 );
buf ( n71208 , n71207 );
buf ( n71209 , n71208 );
not ( n71210 , n46356 );
and ( n71211 , n71210 , n31340 );
not ( n71212 , n63024 );
and ( n71213 , n71212 , n31340 );
and ( n71214 , n31372 , n63024 );
or ( n71215 , n71213 , n71214 );
and ( n71216 , n71215 , n46356 );
or ( n71217 , n71211 , n71216 );
and ( n71218 , n71217 , n31649 );
not ( n71219 , n63032 );
not ( n71220 , n63024 );
and ( n71221 , n71220 , n31340 );
and ( n71222 , n47849 , n63024 );
or ( n71223 , n71221 , n71222 );
and ( n71224 , n71219 , n71223 );
and ( n71225 , n47849 , n63032 );
or ( n71226 , n71224 , n71225 );
and ( n71227 , n71226 , n31643 );
not ( n71228 , n31452 );
not ( n71229 , n63032 );
not ( n71230 , n63024 );
and ( n71231 , n71230 , n31340 );
and ( n71232 , n47849 , n63024 );
or ( n71233 , n71231 , n71232 );
and ( n71234 , n71229 , n71233 );
and ( n71235 , n47849 , n63032 );
or ( n71236 , n71234 , n71235 );
and ( n71237 , n71228 , n71236 );
not ( n71238 , n63052 );
not ( n71239 , n63054 );
and ( n71240 , n71239 , n71236 );
and ( n71241 , n47877 , n63054 );
or ( n71242 , n71240 , n71241 );
and ( n71243 , n71238 , n71242 );
and ( n71244 , n47887 , n63052 );
or ( n71245 , n71243 , n71244 );
and ( n71246 , n71245 , n31452 );
or ( n71247 , n71237 , n71246 );
and ( n71248 , n71247 , n31638 );
and ( n71249 , n31340 , n47277 );
or ( n71250 , C0 , n71218 , n71227 , n71248 , n71249 );
buf ( n71251 , n71250 );
buf ( n71252 , n71251 );
not ( n71253 , n35278 );
buf ( n71254 , RI15b5efc8_1106);
and ( n71255 , n71253 , n71254 );
not ( n71256 , n51396 );
and ( n71257 , n71256 , n51392 );
xor ( n71258 , n51392 , n51155 );
and ( n71259 , n59210 , n59213 );
xor ( n71260 , n71258 , n71259 );
and ( n71261 , n71260 , n51396 );
or ( n71262 , n71257 , n71261 );
and ( n71263 , n71262 , n35278 );
or ( n71264 , n71255 , n71263 );
and ( n71265 , n71264 , n32417 );
not ( n71266 , n50008 );
and ( n71267 , n71266 , n71254 );
not ( n71268 , n51594 );
and ( n71269 , n71268 , n51590 );
xor ( n71270 , n51590 , n40244 );
and ( n71271 , n59224 , n59237 );
xor ( n71272 , n71270 , n71271 );
and ( n71273 , n71272 , n51594 );
or ( n71274 , n71269 , n71273 );
and ( n71275 , n71274 , n50008 );
or ( n71276 , n71267 , n71275 );
and ( n71277 , n71276 , n32415 );
and ( n71278 , n71254 , n48133 );
or ( n71279 , n71265 , n71277 , n71278 );
and ( n71280 , n71279 , n32456 );
and ( n71281 , n71254 , n47409 );
or ( n71282 , C0 , n71280 , n71281 );
buf ( n71283 , n71282 );
buf ( n71284 , n71283 );
buf ( n71285 , n31655 );
buf ( n71286 , n30987 );
buf ( n71287 , n30987 );
not ( n71288 , n31728 );
and ( n71289 , n71288 , n46021 );
xor ( n71290 , n50421 , n50422 );
and ( n71291 , n71290 , n31728 );
or ( n71292 , n71289 , n71291 );
and ( n71293 , n71292 , n32253 );
not ( n71294 , n32283 );
and ( n71295 , n71294 , n46021 );
not ( n71296 , n31823 );
xor ( n71297 , n50443 , n50444 );
and ( n71298 , n71296 , n71297 );
xnor ( n71299 , n50460 , n50461 );
and ( n71300 , n71299 , n31823 );
or ( n71301 , n71298 , n71300 );
and ( n71302 , n71301 , n32283 );
or ( n71303 , n71295 , n71302 );
and ( n71304 , n71303 , n32398 );
and ( n71305 , n46021 , n32436 );
or ( n71306 , n71293 , n71304 , n71305 );
and ( n71307 , n71306 , n32456 );
and ( n71308 , n49660 , n32473 );
not ( n71309 , n32475 );
and ( n71310 , n71309 , n49660 );
xor ( n71311 , n46021 , n50478 );
and ( n71312 , n71311 , n32475 );
or ( n71313 , n71310 , n71312 );
and ( n71314 , n71313 , n32486 );
and ( n71315 , n37539 , n32489 );
and ( n71316 , n46021 , n32501 );
or ( n71317 , C0 , n71307 , n71308 , n71314 , n71315 , n71316 );
buf ( n71318 , n71317 );
buf ( n71319 , n71318 );
and ( n71320 , n33229 , n32528 );
not ( n71321 , n32598 );
and ( n71322 , n71321 , n32992 );
buf ( n71323 , n71322 );
and ( n71324 , n71323 , n32890 );
not ( n71325 , n32919 );
and ( n71326 , n71325 , n32992 );
buf ( n71327 , n71326 );
and ( n71328 , n71327 , n32924 );
not ( n71329 , n32953 );
and ( n71330 , n71329 , n32992 );
not ( n71331 , n32971 );
and ( n71332 , n71331 , n33109 );
xor ( n71333 , n32992 , n33013 );
and ( n71334 , n71333 , n32971 );
or ( n71335 , n71332 , n71334 );
and ( n71336 , n71335 , n32953 );
or ( n71337 , n71330 , n71336 );
and ( n71338 , n71337 , n33038 );
not ( n71339 , n33067 );
and ( n71340 , n71339 , n32992 );
not ( n71341 , n32970 );
not ( n71342 , n33071 );
and ( n71343 , n71342 , n33109 );
xor ( n71344 , n33110 , n33145 );
and ( n71345 , n71344 , n33071 );
or ( n71346 , n71343 , n71345 );
and ( n71347 , n71341 , n71346 );
and ( n71348 , n71333 , n32970 );
or ( n71349 , n71347 , n71348 );
and ( n71350 , n71349 , n33067 );
or ( n71351 , n71340 , n71350 );
and ( n71352 , n71351 , n33172 );
and ( n71353 , n32992 , n33204 );
or ( n71354 , n71324 , n71328 , n71338 , n71352 , n71353 );
and ( n71355 , n71354 , n33208 );
not ( n71356 , n32968 );
not ( n71357 , n33270 );
and ( n71358 , n71357 , n33309 );
xor ( n71359 , n33310 , n33345 );
and ( n71360 , n71359 , n33270 );
or ( n71361 , n71358 , n71360 );
and ( n71362 , n71356 , n71361 );
and ( n71363 , n32992 , n32968 );
or ( n71364 , n71362 , n71363 );
and ( n71365 , n71364 , n33370 );
buf ( n71366 , n35056 );
and ( n71367 , n32992 , n33382 );
or ( n71368 , C0 , n71320 , n71355 , n71365 , n71366 , n71367 );
buf ( n71369 , n71368 );
buf ( n71370 , n71369 );
buf ( n71371 , n30987 );
buf ( n71372 , n31655 );
buf ( n71373 , n31655 );
buf ( n71374 , n30987 );
buf ( n71375 , n30987 );
buf ( n71376 , n31655 );
and ( n71377 , n31565 , n31007 );
not ( n71378 , n31077 );
and ( n71379 , n71378 , n35391 );
buf ( n71380 , n71379 );
and ( n71381 , n71380 , n31373 );
not ( n71382 , n31402 );
and ( n71383 , n71382 , n35391 );
buf ( n71384 , n71383 );
and ( n71385 , n71384 , n31408 );
not ( n71386 , n31437 );
and ( n71387 , n71386 , n35391 );
not ( n71388 , n31455 );
and ( n71389 , n71388 , n35431 );
xor ( n71390 , n35391 , n35407 );
and ( n71391 , n71390 , n31455 );
or ( n71392 , n71389 , n71391 );
and ( n71393 , n71392 , n31437 );
or ( n71394 , n71387 , n71393 );
and ( n71395 , n71394 , n31468 );
not ( n71396 , n31497 );
and ( n71397 , n71396 , n35391 );
not ( n71398 , n31454 );
not ( n71399 , n31501 );
and ( n71400 , n71399 , n35431 );
xor ( n71401 , n35432 , n35457 );
and ( n71402 , n71401 , n31501 );
or ( n71403 , n71400 , n71402 );
and ( n71404 , n71398 , n71403 );
and ( n71405 , n71390 , n31454 );
or ( n71406 , n71404 , n71405 );
and ( n71407 , n71406 , n31497 );
or ( n71408 , n71397 , n71407 );
and ( n71409 , n71408 , n31521 );
and ( n71410 , n35391 , n31553 );
or ( n71411 , n71381 , n71385 , n71395 , n71409 , n71410 );
and ( n71412 , n71411 , n31557 );
not ( n71413 , n31452 );
not ( n71414 , n31619 );
and ( n71415 , n71414 , n35486 );
xor ( n71416 , n35487 , n35511 );
and ( n71417 , n71416 , n31619 );
or ( n71418 , n71415 , n71417 );
and ( n71419 , n71413 , n71418 );
and ( n71420 , n35391 , n31452 );
or ( n71421 , n71419 , n71420 );
and ( n71422 , n71421 , n31638 );
and ( n71423 , n35391 , n31650 );
or ( n71424 , C0 , n71377 , n71412 , n71422 , C0 , n71423 );
buf ( n71425 , n71424 );
buf ( n71426 , n71425 );
not ( n71427 , n33419 );
and ( n71428 , n71427 , n31579 );
xor ( n71429 , n33473 , n33692 );
and ( n71430 , n71429 , n33419 );
or ( n71431 , n71428 , n71430 );
and ( n71432 , n71431 , n31529 );
not ( n71433 , n33734 );
and ( n71434 , n71433 , n31579 );
not ( n71435 , n33533 );
xor ( n71436 , n33766 , n33810 );
and ( n71437 , n71435 , n71436 );
xnor ( n71438 , n33851 , n33912 );
and ( n71439 , n71438 , n33533 );
or ( n71440 , n71437 , n71439 );
and ( n71441 , n71440 , n33734 );
or ( n71442 , n71434 , n71441 );
and ( n71443 , n71442 , n31527 );
and ( n71444 , n31579 , n33942 );
or ( n71445 , n71432 , n71443 , n71444 );
and ( n71446 , n71445 , n31557 );
and ( n71447 , n34103 , n31643 );
not ( n71448 , n31452 );
and ( n71449 , n71448 , n34103 );
xor ( n71450 , n31579 , n33958 );
and ( n71451 , n71450 , n31452 );
or ( n71452 , n71449 , n71451 );
and ( n71453 , n71452 , n31638 );
and ( n71454 , n34003 , n33973 );
and ( n71455 , n31579 , n33978 );
or ( n71456 , C0 , n71446 , n71447 , n71453 , n71454 , n71455 );
buf ( n71457 , n71456 );
buf ( n71458 , n71457 );
buf ( n71459 , n31655 );
buf ( n71460 , n31655 );
buf ( n71461 , n30987 );
not ( n71462 , n32953 );
and ( n71463 , n71462 , n54688 );
not ( n71464 , n39572 );
and ( n71465 , n71464 , n39412 );
xor ( n71466 , n42625 , n42628 );
and ( n71467 , n71466 , n39572 );
or ( n71468 , n71465 , n71467 );
and ( n71469 , n71468 , n32953 );
or ( n71470 , n71463 , n71469 );
and ( n71471 , n71470 , n33038 );
not ( n71472 , n39586 );
and ( n71473 , n71472 , n54688 );
and ( n71474 , n54694 , n39586 );
or ( n71475 , n71473 , n71474 );
and ( n71476 , n71475 , n33172 );
and ( n71477 , n54688 , n39795 );
or ( n71478 , n71471 , n71476 , n71477 );
and ( n71479 , n71478 , n33208 );
and ( n71480 , n54688 , n39805 );
or ( n71481 , C0 , n71479 , n71480 );
buf ( n71482 , n71481 );
buf ( n71483 , n71482 );
buf ( n71484 , n30987 );
buf ( n71485 , n31655 );
buf ( n71486 , n30987 );
not ( n71487 , n36587 );
and ( n71488 , n71487 , n36396 );
xor ( n71489 , n50177 , n50210 );
and ( n71490 , n71489 , n36587 );
or ( n71491 , n71488 , n71490 );
and ( n71492 , n71491 , n36596 );
not ( n71493 , n37485 );
and ( n71494 , n71493 , n37298 );
xor ( n71495 , n50227 , n50260 );
and ( n71496 , n71495 , n37485 );
or ( n71497 , n71494 , n71496 );
and ( n71498 , n71497 , n37494 );
and ( n71499 , n41857 , n37506 );
or ( n71500 , n71492 , n71498 , n71499 );
buf ( n71501 , n71500 );
buf ( n71502 , n71501 );
buf ( n71503 , n31655 );
and ( n71504 , n50440 , n50275 );
not ( n71505 , n50278 );
and ( n71506 , n71505 , n50408 );
and ( n71507 , n50440 , n50278 );
or ( n71508 , n71506 , n71507 );
and ( n71509 , n71508 , n32421 );
not ( n71510 , n50002 );
and ( n71511 , n71510 , n50408 );
and ( n71512 , n50440 , n50002 );
or ( n71513 , n71511 , n71512 );
and ( n71514 , n71513 , n32419 );
not ( n71515 , n50289 );
and ( n71516 , n71515 , n50408 );
and ( n71517 , n50440 , n50289 );
or ( n71518 , n71516 , n71517 );
and ( n71519 , n71518 , n32417 );
not ( n71520 , n50008 );
and ( n71521 , n71520 , n50408 );
and ( n71522 , n50440 , n50008 );
or ( n71523 , n71521 , n71522 );
and ( n71524 , n71523 , n32415 );
not ( n71525 , n47331 );
and ( n71526 , n71525 , n50408 );
and ( n71527 , n50418 , n47331 );
or ( n71528 , n71526 , n71527 );
and ( n71529 , n71528 , n32413 );
not ( n71530 , n50067 );
and ( n71531 , n71530 , n50408 );
and ( n71532 , n50418 , n50067 );
or ( n71533 , n71531 , n71532 );
and ( n71534 , n71533 , n32411 );
not ( n71535 , n31728 );
and ( n71536 , n71535 , n50408 );
xor ( n71537 , n50418 , n50425 );
and ( n71538 , n71537 , n31728 );
or ( n71539 , n71536 , n71538 );
and ( n71540 , n71539 , n32253 );
not ( n71541 , n32283 );
and ( n71542 , n71541 , n50408 );
not ( n71543 , n31823 );
xor ( n71544 , n50440 , n50447 );
and ( n71545 , n71543 , n71544 );
xnor ( n71546 , n50457 , n50464 );
and ( n71547 , n71546 , n31823 );
or ( n71548 , n71545 , n71547 );
and ( n71549 , n71548 , n32283 );
or ( n71550 , n71542 , n71549 );
and ( n71551 , n71550 , n32398 );
and ( n71552 , n50457 , n50334 );
or ( n71553 , n71504 , n71509 , n71514 , n71519 , n71524 , n71529 , n71534 , n71540 , n71551 , n71552 );
and ( n71554 , n71553 , n32456 );
and ( n71555 , n37533 , n32489 );
and ( n71556 , n50408 , n50345 );
or ( n71557 , C0 , n71554 , n71555 , n71556 );
buf ( n71558 , n71557 );
buf ( n71559 , n71558 );
buf ( n71560 , n30987 );
buf ( n71561 , n31655 );
buf ( n71562 , n31655 );
buf ( n71563 , n30987 );
xor ( n71564 , n33107 , n56360 );
and ( n71565 , n71564 , n33201 );
not ( n71566 , n41576 );
and ( n71567 , n71566 , n33107 );
and ( n71568 , n32791 , n52252 );
and ( n71569 , n32793 , n52254 );
and ( n71570 , n32795 , n52256 );
and ( n71571 , n32797 , n52258 );
and ( n71572 , n32799 , n52260 );
and ( n71573 , n32801 , n52262 );
and ( n71574 , n32803 , n52264 );
and ( n71575 , n32805 , n52266 );
and ( n71576 , n32807 , n52268 );
and ( n71577 , n32809 , n52270 );
and ( n71578 , n32811 , n52272 );
and ( n71579 , n32813 , n52274 );
and ( n71580 , n32815 , n52276 );
and ( n71581 , n32817 , n52278 );
and ( n71582 , n32819 , n52280 );
and ( n71583 , n32821 , n52282 );
or ( n71584 , n71568 , n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , n71581 , n71582 , n71583 );
and ( n71585 , n71584 , n41576 );
or ( n71586 , n71567 , n71585 );
and ( n71587 , n71586 , n33189 );
and ( n71588 , n33107 , n41592 );
or ( n71589 , n71565 , n71587 , n71588 );
and ( n71590 , n71589 , n33208 );
and ( n71591 , n33107 , n39805 );
or ( n71592 , C0 , n71590 , n71591 );
buf ( n71593 , n71592 );
buf ( n71594 , n71593 );
not ( n71595 , n50828 );
not ( n71596 , n50834 );
and ( n71597 , n71596 , n40590 );
and ( n71598 , n45276 , n50834 );
or ( n71599 , n71597 , n71598 );
and ( n71600 , n71595 , n71599 );
buf ( n71601 , RI15b60378_1148);
and ( n71602 , n71601 , n50828 );
or ( n71603 , n71600 , n71602 );
buf ( n71604 , n71603 );
buf ( n71605 , n71604 );
buf ( n71606 , n30987 );
buf ( n71607 , n30987 );
buf ( n71608 , n31655 );
and ( n71609 , n64057 , n33377 );
not ( n71610 , n48545 );
and ( n71611 , n71610 , n64792 );
buf ( n71612 , n71611 );
and ( n71613 , n71612 , n32890 );
not ( n71614 , n48557 );
and ( n71615 , n71614 , n64792 );
and ( n71616 , n64065 , n48557 );
or ( n71617 , n71615 , n71616 );
and ( n71618 , n71617 , n33038 );
and ( n71619 , n64792 , n48571 );
or ( n71620 , n71613 , n71618 , n71619 );
and ( n71621 , n71620 , n33208 );
and ( n71622 , n64792 , n48577 );
or ( n71623 , C0 , n71609 , n71621 , n71622 );
buf ( n71624 , n71623 );
buf ( n71625 , n71624 );
buf ( n71626 , n31655 );
buf ( n71627 , n30987 );
buf ( n71628 , n31655 );
xor ( n71629 , n49565 , n60323 );
and ( n71630 , n71629 , n32433 );
not ( n71631 , n47331 );
and ( n71632 , n71631 , n49565 );
xor ( n71633 , n60399 , n60547 );
and ( n71634 , n71633 , n47331 );
or ( n71635 , n71632 , n71634 );
and ( n71636 , n71635 , n32413 );
and ( n71637 , n49565 , n47402 );
or ( n71638 , n71630 , n71636 , n71637 );
and ( n71639 , n71638 , n32456 );
and ( n71640 , n49565 , n47409 );
or ( n71641 , C0 , n71639 , n71640 );
buf ( n71642 , n71641 );
buf ( n71643 , n71642 );
buf ( n71644 , n31655 );
buf ( n71645 , n30987 );
not ( n71646 , n46356 );
and ( n71647 , n71646 , n31270 );
not ( n71648 , n60564 );
and ( n71649 , n71648 , n31270 );
and ( n71650 , n31272 , n60564 );
or ( n71651 , n71649 , n71650 );
and ( n71652 , n71651 , n46356 );
or ( n71653 , n71647 , n71652 );
and ( n71654 , n71653 , n31649 );
not ( n71655 , n60572 );
not ( n71656 , n60564 );
and ( n71657 , n71656 , n31270 );
and ( n71658 , n49443 , n60564 );
or ( n71659 , n71657 , n71658 );
and ( n71660 , n71655 , n71659 );
and ( n71661 , n49443 , n60572 );
or ( n71662 , n71660 , n71661 );
and ( n71663 , n71662 , n31643 );
not ( n71664 , n31452 );
not ( n71665 , n60572 );
not ( n71666 , n60564 );
and ( n71667 , n71666 , n31270 );
and ( n71668 , n49443 , n60564 );
or ( n71669 , n71667 , n71668 );
and ( n71670 , n71665 , n71669 );
and ( n71671 , n49443 , n60572 );
or ( n71672 , n71670 , n71671 );
and ( n71673 , n71664 , n71672 );
not ( n71674 , n60592 );
not ( n71675 , n60594 );
and ( n71676 , n71675 , n71672 );
and ( n71677 , n49469 , n60594 );
or ( n71678 , n71676 , n71677 );
and ( n71679 , n71674 , n71678 );
and ( n71680 , n49477 , n60592 );
or ( n71681 , n71679 , n71680 );
and ( n71682 , n71681 , n31452 );
or ( n71683 , n71673 , n71682 );
and ( n71684 , n71683 , n31638 );
and ( n71685 , n31270 , n47277 );
or ( n71686 , C0 , n71654 , n71663 , n71684 , n71685 );
buf ( n71687 , n71686 );
buf ( n71688 , n71687 );
not ( n71689 , n46356 );
and ( n71690 , n71689 , n31294 );
not ( n71691 , n64746 );
and ( n71692 , n71691 , n31294 );
and ( n71693 , n31306 , n64746 );
or ( n71694 , n71692 , n71693 );
and ( n71695 , n71694 , n46356 );
or ( n71696 , n71690 , n71695 );
and ( n71697 , n71696 , n31649 );
not ( n71698 , n64754 );
not ( n71699 , n64746 );
and ( n71700 , n71699 , n31294 );
and ( n71701 , n58061 , n64746 );
or ( n71702 , n71700 , n71701 );
and ( n71703 , n71698 , n71702 );
and ( n71704 , n58061 , n64754 );
or ( n71705 , n71703 , n71704 );
and ( n71706 , n71705 , n31643 );
not ( n71707 , n31452 );
not ( n71708 , n64754 );
not ( n71709 , n64746 );
and ( n71710 , n71709 , n31294 );
and ( n71711 , n58061 , n64746 );
or ( n71712 , n71710 , n71711 );
and ( n71713 , n71708 , n71712 );
and ( n71714 , n58061 , n64754 );
or ( n71715 , n71713 , n71714 );
and ( n71716 , n71707 , n71715 );
not ( n71717 , n64774 );
not ( n71718 , n64776 );
and ( n71719 , n71718 , n71715 );
and ( n71720 , n58085 , n64776 );
or ( n71721 , n71719 , n71720 );
and ( n71722 , n71717 , n71721 );
and ( n71723 , n58093 , n64774 );
or ( n71724 , n71722 , n71723 );
and ( n71725 , n71724 , n31452 );
or ( n71726 , n71716 , n71725 );
and ( n71727 , n71726 , n31638 );
and ( n71728 , n31294 , n47277 );
or ( n71729 , C0 , n71697 , n71706 , n71727 , n71728 );
buf ( n71730 , n71729 );
buf ( n71731 , n71730 );
buf ( n71732 , n31655 );
xor ( n71733 , n50969 , n64712 );
and ( n71734 , n71733 , n32431 );
not ( n71735 , n50002 );
and ( n71736 , n71735 , n50969 );
and ( n71737 , n40634 , n50002 );
or ( n71738 , n71736 , n71737 );
and ( n71739 , n71738 , n32419 );
not ( n71740 , n50008 );
and ( n71741 , n71740 , n50969 );
not ( n71742 , n51594 );
and ( n71743 , n71742 , n51458 );
xor ( n71744 , n51600 , n51606 );
and ( n71745 , n71744 , n51594 );
or ( n71746 , n71743 , n71745 );
and ( n71747 , n71746 , n50008 );
or ( n71748 , n71741 , n71747 );
and ( n71749 , n71748 , n32415 );
not ( n71750 , n50067 );
and ( n71751 , n71750 , n50969 );
and ( n71752 , n71019 , n50067 );
or ( n71753 , n71751 , n71752 );
and ( n71754 , n71753 , n32411 );
and ( n71755 , n50969 , n50098 );
or ( n71756 , n71734 , n71739 , n71749 , n71754 , n71755 );
and ( n71757 , n71756 , n32456 );
and ( n71758 , n50969 , n47409 );
or ( n71759 , C0 , n71757 , n71758 );
buf ( n71760 , n71759 );
buf ( n71761 , n71760 );
buf ( n71762 , n30987 );
buf ( n71763 , n31655 );
buf ( n71764 , n30987 );
buf ( n71765 , n30987 );
xor ( n71766 , n44766 , n44801 );
and ( n71767 , n71766 , n31548 );
not ( n71768 , n44807 );
and ( n71769 , n71768 , n44766 );
and ( n71770 , n46627 , n44807 );
or ( n71771 , n71769 , n71770 );
and ( n71772 , n71771 , n31408 );
not ( n71773 , n44817 );
and ( n71774 , n71773 , n44766 );
and ( n71775 , n69627 , n44817 );
or ( n71776 , n71774 , n71775 );
and ( n71777 , n71776 , n31521 );
not ( n71778 , n45059 );
and ( n71779 , n71778 , n44766 );
xor ( n71780 , n45129 , n45132 );
and ( n71781 , n71780 , n45059 );
or ( n71782 , n71779 , n71781 );
and ( n71783 , n71782 , n31536 );
and ( n71784 , n44766 , n45148 );
or ( n71785 , n71767 , n71772 , n71777 , n71783 , n71784 );
and ( n71786 , n71785 , n31557 );
and ( n71787 , n44766 , n40154 );
or ( n71788 , C0 , n71786 , n71787 );
buf ( n71789 , n71788 );
buf ( n71790 , n71789 );
buf ( n71791 , n31655 );
not ( n71792 , n40163 );
and ( n71793 , n71792 , n31848 );
not ( n71794 , n45161 );
and ( n71795 , n71794 , n31848 );
and ( n71796 , n32235 , n45161 );
or ( n71797 , n71795 , n71796 );
and ( n71798 , n71797 , n40163 );
or ( n71799 , n71793 , n71798 );
and ( n71800 , n71799 , n32498 );
not ( n71801 , n45170 );
not ( n71802 , n45161 );
and ( n71803 , n71802 , n31848 );
and ( n71804 , n42188 , n45161 );
or ( n71805 , n71803 , n71804 );
and ( n71806 , n71801 , n71805 );
and ( n71807 , n42188 , n45170 );
or ( n71808 , n71806 , n71807 );
and ( n71809 , n71808 , n32473 );
not ( n71810 , n32475 );
not ( n71811 , n45170 );
not ( n71812 , n45161 );
and ( n71813 , n71812 , n31848 );
and ( n71814 , n42188 , n45161 );
or ( n71815 , n71813 , n71814 );
and ( n71816 , n71811 , n71815 );
and ( n71817 , n42188 , n45170 );
or ( n71818 , n71816 , n71817 );
and ( n71819 , n71810 , n71818 );
not ( n71820 , n45196 );
not ( n71821 , n45199 );
and ( n71822 , n71821 , n71818 );
and ( n71823 , n42216 , n45199 );
or ( n71824 , n71822 , n71823 );
and ( n71825 , n71820 , n71824 );
and ( n71826 , n42224 , n45196 );
or ( n71827 , n71825 , n71826 );
and ( n71828 , n71827 , n32475 );
or ( n71829 , n71819 , n71828 );
and ( n71830 , n71829 , n32486 );
and ( n71831 , n31848 , n41278 );
or ( n71832 , C0 , n71800 , n71809 , n71830 , n71831 );
buf ( n71833 , n71832 );
buf ( n71834 , n71833 );
and ( n71835 , n33777 , n48455 );
not ( n71836 , n48457 );
and ( n71837 , n71836 , n33439 );
and ( n71838 , n33777 , n48457 );
or ( n71839 , n71837 , n71838 );
and ( n71840 , n71839 , n31373 );
not ( n71841 , n44807 );
and ( n71842 , n71841 , n33439 );
and ( n71843 , n33777 , n44807 );
or ( n71844 , n71842 , n71843 );
and ( n71845 , n71844 , n31408 );
not ( n71846 , n48468 );
and ( n71847 , n71846 , n33439 );
and ( n71848 , n33777 , n48468 );
or ( n71849 , n71847 , n71848 );
and ( n71850 , n71849 , n31468 );
not ( n71851 , n44817 );
and ( n71852 , n71851 , n33439 );
and ( n71853 , n33777 , n44817 );
or ( n71854 , n71852 , n71853 );
and ( n71855 , n71854 , n31521 );
not ( n71856 , n39979 );
and ( n71857 , n71856 , n33439 );
and ( n71858 , n33573 , n39979 );
or ( n71859 , n71857 , n71858 );
and ( n71860 , n71859 , n31538 );
not ( n71861 , n45059 );
and ( n71862 , n71861 , n33439 );
and ( n71863 , n33573 , n45059 );
or ( n71864 , n71862 , n71863 );
and ( n71865 , n71864 , n31536 );
not ( n71866 , n33419 );
and ( n71867 , n71866 , n33439 );
xor ( n71868 , n33573 , n33590 );
xor ( n71869 , n71868 , n33676 );
and ( n71870 , n71869 , n33419 );
or ( n71871 , n71867 , n71870 );
and ( n71872 , n71871 , n31529 );
not ( n71873 , n33734 );
and ( n71874 , n71873 , n33439 );
not ( n71875 , n33533 );
xor ( n71876 , n33777 , n33590 );
xor ( n71877 , n71876 , n33794 );
and ( n71878 , n71875 , n71877 );
xor ( n71879 , n33868 , n33870 );
xor ( n71880 , n71879 , n33896 );
and ( n71881 , n71880 , n33533 );
or ( n71882 , n71878 , n71881 );
and ( n71883 , n71882 , n33734 );
or ( n71884 , n71874 , n71883 );
and ( n71885 , n71884 , n31527 );
and ( n71886 , n33868 , n48513 );
or ( n71887 , n71835 , n71840 , n71845 , n71850 , n71855 , n71860 , n71865 , n71872 , n71885 , n71886 );
and ( n71888 , n71887 , n31557 );
and ( n71889 , n34011 , n33973 );
and ( n71890 , n33439 , n48524 );
or ( n71891 , C0 , n71888 , n71889 , n71890 );
buf ( n71892 , n71891 );
buf ( n71893 , n71892 );
not ( n71894 , n35278 );
buf ( n71895 , RI15b5ed70_1101);
and ( n71896 , n71894 , n71895 );
not ( n71897 , n51396 );
and ( n71898 , n71897 , n51307 );
xor ( n71899 , n53329 , n53334 );
and ( n71900 , n71899 , n51396 );
or ( n71901 , n71898 , n71900 );
and ( n71902 , n71901 , n35278 );
or ( n71903 , n71896 , n71902 );
and ( n71904 , n71903 , n32417 );
not ( n71905 , n50008 );
and ( n71906 , n71905 , n71895 );
and ( n71907 , n67374 , n50008 );
or ( n71908 , n71906 , n71907 );
and ( n71909 , n71908 , n32415 );
and ( n71910 , n71895 , n48133 );
or ( n71911 , n71904 , n71909 , n71910 );
and ( n71912 , n71911 , n32456 );
and ( n71913 , n71895 , n47409 );
or ( n71914 , C0 , n71912 , n71913 );
buf ( n71915 , n71914 );
buf ( n71916 , n71915 );
buf ( n71917 , n30987 );
buf ( n71918 , n31655 );
buf ( n71919 , n30987 );
buf ( n71920 , n31655 );
buf ( n71921 , n40203 );
buf ( n71922 , n31655 );
and ( n71923 , n46035 , n32500 );
not ( n71924 , n35211 );
and ( n71925 , n71924 , n37567 );
buf ( n71926 , n71925 );
and ( n71927 , n71926 , n32421 );
not ( n71928 , n35245 );
and ( n71929 , n71928 , n37567 );
buf ( n71930 , n71929 );
and ( n71931 , n71930 , n32419 );
not ( n71932 , n35278 );
and ( n71933 , n71932 , n37567 );
not ( n71934 , n35295 );
and ( n71935 , n71934 , n49597 );
xor ( n71936 , n37567 , n49532 );
and ( n71937 , n71936 , n35295 );
or ( n71938 , n71935 , n71937 );
and ( n71939 , n71938 , n35278 );
or ( n71940 , n71933 , n71939 );
and ( n71941 , n71940 , n32417 );
not ( n71942 , n35331 );
and ( n71943 , n71942 , n37567 );
not ( n71944 , n35294 );
not ( n71945 , n45995 );
and ( n71946 , n71945 , n49597 );
xor ( n71947 , n49598 , n49618 );
and ( n71948 , n71947 , n45995 );
or ( n71949 , n71946 , n71948 );
and ( n71950 , n71944 , n71949 );
and ( n71951 , n71936 , n35294 );
or ( n71952 , n71950 , n71951 );
and ( n71953 , n71952 , n35331 );
or ( n71954 , n71943 , n71953 );
and ( n71955 , n71954 , n32415 );
and ( n71956 , n37567 , n35354 );
or ( n71957 , n71927 , n71931 , n71941 , n71955 , n71956 );
and ( n71958 , n71957 , n32456 );
not ( n71959 , n32475 );
not ( n71960 , n46060 );
and ( n71961 , n71960 , n49687 );
xor ( n71962 , n49688 , n49712 );
and ( n71963 , n71962 , n46060 );
or ( n71964 , n71961 , n71963 );
and ( n71965 , n71959 , n71964 );
and ( n71966 , n37567 , n32475 );
or ( n71967 , n71965 , n71966 );
and ( n71968 , n71967 , n32486 );
buf ( n71969 , n32489 );
and ( n71970 , n37567 , n35367 );
or ( n71971 , C0 , n71923 , n71958 , n71968 , n71969 , n71970 );
buf ( n71972 , n71971 );
buf ( n71973 , n71972 );
buf ( n71974 , n30987 );
not ( n71975 , n48765 );
and ( n71976 , n71975 , n33215 );
xor ( n71977 , n48770 , n49018 );
and ( n71978 , n71977 , n48765 );
or ( n71979 , n71976 , n71978 );
and ( n71980 , n71979 , n33180 );
not ( n71981 , n49054 );
and ( n71982 , n71981 , n33215 );
not ( n71983 , n48845 );
xor ( n71984 , n49060 , n49132 );
and ( n71985 , n71983 , n71984 );
xnor ( n71986 , n49169 , n49258 );
and ( n71987 , n71986 , n48845 );
or ( n71988 , n71985 , n71987 );
and ( n71989 , n71988 , n49054 );
or ( n71990 , n71982 , n71989 );
and ( n71991 , n71990 , n33178 );
and ( n71992 , n33215 , n49774 );
or ( n71993 , n71980 , n71991 , n71992 );
and ( n71994 , n71993 , n33208 );
and ( n71995 , n33281 , n33375 );
not ( n71996 , n32968 );
and ( n71997 , n71996 , n33281 );
xor ( n71998 , n33215 , n66020 );
and ( n71999 , n71998 , n32968 );
or ( n72000 , n71997 , n71999 );
and ( n72001 , n72000 , n33370 );
and ( n72002 , n32978 , n35056 );
and ( n72003 , n33215 , n49794 );
or ( n72004 , C0 , n71994 , n71995 , n72001 , n72002 , n72003 );
buf ( n72005 , n72004 );
buf ( n72006 , n72005 );
buf ( n72007 , n30987 );
buf ( n72008 , n30987 );
buf ( n72009 , n31655 );
and ( n72010 , n70660 , n33377 );
not ( n72011 , n48545 );
and ( n72012 , n72011 , n41510 );
buf ( n72013 , n72012 );
and ( n72014 , n72013 , n32890 );
not ( n72015 , n48557 );
and ( n72016 , n72015 , n41510 );
and ( n72017 , n70668 , n48557 );
or ( n72018 , n72016 , n72017 );
and ( n72019 , n72018 , n33038 );
and ( n72020 , n41510 , n48571 );
or ( n72021 , n72014 , n72019 , n72020 );
and ( n72022 , n72021 , n33208 );
and ( n72023 , n41510 , n48577 );
or ( n72024 , C0 , n72010 , n72022 , n72023 );
buf ( n72025 , n72024 );
buf ( n72026 , n72025 );
buf ( n72027 , n31655 );
buf ( n72028 , n31655 );
buf ( n72029 , n30987 );
buf ( n72030 , n31655 );
not ( n72031 , n46356 );
and ( n72032 , n72031 , n31090 );
not ( n72033 , n47831 );
and ( n72034 , n72033 , n31090 );
and ( n72035 , n31138 , n47831 );
or ( n72036 , n72034 , n72035 );
and ( n72037 , n72036 , n46356 );
or ( n72038 , n72032 , n72037 );
and ( n72039 , n72038 , n31649 );
not ( n72040 , n47839 );
not ( n72041 , n47831 );
and ( n72042 , n72041 , n31090 );
and ( n72043 , n56920 , n47831 );
or ( n72044 , n72042 , n72043 );
and ( n72045 , n72040 , n72044 );
and ( n72046 , n56920 , n47839 );
or ( n72047 , n72045 , n72046 );
and ( n72048 , n72047 , n31643 );
not ( n72049 , n31452 );
not ( n72050 , n47839 );
not ( n72051 , n47831 );
and ( n72052 , n72051 , n31090 );
and ( n72053 , n56920 , n47831 );
or ( n72054 , n72052 , n72053 );
and ( n72055 , n72050 , n72054 );
and ( n72056 , n56920 , n47839 );
or ( n72057 , n72055 , n72056 );
and ( n72058 , n72049 , n72057 );
not ( n72059 , n47866 );
not ( n72060 , n47868 );
and ( n72061 , n72060 , n72057 );
and ( n72062 , n56946 , n47868 );
or ( n72063 , n72061 , n72062 );
and ( n72064 , n72059 , n72063 );
and ( n72065 , n56954 , n47866 );
or ( n72066 , n72064 , n72065 );
and ( n72067 , n72066 , n31452 );
or ( n72068 , n72058 , n72067 );
and ( n72069 , n72068 , n31638 );
and ( n72070 , n31090 , n47277 );
or ( n72071 , C0 , n72039 , n72048 , n72069 , n72070 );
buf ( n72072 , n72071 );
buf ( n72073 , n72072 );
not ( n72074 , n35278 );
and ( n72075 , n72074 , n50012 );
not ( n72076 , n46290 );
and ( n72077 , n72076 , n46273 );
xor ( n72078 , n46273 , n46092 );
and ( n72079 , n46293 , n46319 );
xor ( n72080 , n72078 , n72079 );
and ( n72081 , n72080 , n46290 );
or ( n72082 , n72077 , n72081 );
and ( n72083 , n72082 , n35278 );
or ( n72084 , n72075 , n72083 );
and ( n72085 , n72084 , n32417 );
not ( n72086 , n47912 );
and ( n72087 , n72086 , n50012 );
and ( n72088 , n50032 , n47912 );
or ( n72089 , n72087 , n72088 );
and ( n72090 , n72089 , n32415 );
and ( n72091 , n50012 , n48133 );
or ( n72092 , n72085 , n72090 , n72091 );
and ( n72093 , n72092 , n32456 );
and ( n72094 , n50012 , n47409 );
or ( n72095 , C0 , n72093 , n72094 );
buf ( n72096 , n72095 );
buf ( n72097 , n72096 );
buf ( n72098 , n31655 );
buf ( n72099 , n31655 );
buf ( n72100 , n30987 );
not ( n72101 , n32953 );
buf ( n72102 , RI15b46c20_279);
and ( n72103 , n72101 , n72102 );
not ( n72104 , n39572 );
and ( n72105 , n72104 , n39503 );
xor ( n72106 , n42618 , n42635 );
and ( n72107 , n72106 , n39572 );
or ( n72108 , n72105 , n72107 );
and ( n72109 , n72108 , n32953 );
or ( n72110 , n72103 , n72109 );
and ( n72111 , n72110 , n33038 );
not ( n72112 , n39586 );
and ( n72113 , n72112 , n72102 );
not ( n72114 , n39775 );
and ( n72115 , n72114 , n39711 );
xor ( n72116 , n42654 , n42671 );
and ( n72117 , n72116 , n39775 );
or ( n72118 , n72115 , n72117 );
and ( n72119 , n72118 , n39586 );
or ( n72120 , n72113 , n72119 );
and ( n72121 , n72120 , n33172 );
and ( n72122 , n72102 , n39795 );
or ( n72123 , n72111 , n72121 , n72122 );
and ( n72124 , n72123 , n33208 );
and ( n72125 , n72102 , n39805 );
or ( n72126 , C0 , n72124 , n72125 );
buf ( n72127 , n72126 );
buf ( n72128 , n72127 );
buf ( n72129 , n30987 );
buf ( n72130 , n31655 );
not ( n72131 , n40163 );
and ( n72132 , n72131 , n32017 );
not ( n72133 , n50540 );
and ( n72134 , n72133 , n32017 );
and ( n72135 , n32147 , n50540 );
or ( n72136 , n72134 , n72135 );
and ( n72137 , n72136 , n40163 );
or ( n72138 , n72132 , n72137 );
and ( n72139 , n72138 , n32498 );
not ( n72140 , n50548 );
not ( n72141 , n50540 );
and ( n72142 , n72141 , n32017 );
and ( n72143 , n49314 , n50540 );
or ( n72144 , n72142 , n72143 );
and ( n72145 , n72140 , n72144 );
and ( n72146 , n49314 , n50548 );
or ( n72147 , n72145 , n72146 );
and ( n72148 , n72147 , n32473 );
not ( n72149 , n32475 );
not ( n72150 , n50548 );
not ( n72151 , n50540 );
and ( n72152 , n72151 , n32017 );
and ( n72153 , n49314 , n50540 );
or ( n72154 , n72152 , n72153 );
and ( n72155 , n72150 , n72154 );
and ( n72156 , n49314 , n50548 );
or ( n72157 , n72155 , n72156 );
and ( n72158 , n72149 , n72157 );
not ( n72159 , n50568 );
not ( n72160 , n50570 );
and ( n72161 , n72160 , n72157 );
and ( n72162 , n49340 , n50570 );
or ( n72163 , n72161 , n72162 );
and ( n72164 , n72159 , n72163 );
and ( n72165 , n49348 , n50568 );
or ( n72166 , n72164 , n72165 );
and ( n72167 , n72166 , n32475 );
or ( n72168 , n72158 , n72167 );
and ( n72169 , n72168 , n32486 );
and ( n72170 , n32017 , n41278 );
or ( n72171 , C0 , n72139 , n72148 , n72169 , n72170 );
buf ( n72172 , n72171 );
buf ( n72173 , n72172 );
buf ( n72174 , n30987 );
buf ( n72175 , n30987 );
xor ( n72176 , n41691 , n44782 );
and ( n72177 , n72176 , n31548 );
not ( n72178 , n44807 );
and ( n72179 , n72178 , n41691 );
and ( n72180 , n41982 , n44807 );
or ( n72181 , n72179 , n72180 );
and ( n72182 , n72181 , n31408 );
not ( n72183 , n44817 );
and ( n72184 , n72183 , n41691 );
not ( n72185 , n41835 );
and ( n72186 , n72185 , n58809 );
and ( n72187 , n58825 , n41835 );
or ( n72188 , n72186 , n72187 );
and ( n72189 , n72188 , n44817 );
or ( n72190 , n72184 , n72189 );
and ( n72191 , n72190 , n31521 );
not ( n72192 , n45059 );
and ( n72193 , n72192 , n41691 );
and ( n72194 , n33533 , n45059 );
or ( n72195 , n72193 , n72194 );
and ( n72196 , n72195 , n31536 );
and ( n72197 , n41691 , n45148 );
or ( n72198 , n72177 , n72182 , n72191 , n72196 , n72197 );
and ( n72199 , n72198 , n31557 );
and ( n72200 , n41691 , n40154 );
or ( n72201 , C0 , n72199 , n72200 );
buf ( n72202 , n72201 );
buf ( n72203 , n72202 );
not ( n72204 , n35211 );
buf ( n72205 , n72204 );
buf ( n72206 , RI15b5d510_1049);
not ( n72207 , n50277 );
and ( n72208 , n72206 , n72207 );
and ( n72209 , n72208 , n35211 );
or ( n72210 , n72205 , n72209 );
and ( n72211 , n72210 , n32421 );
not ( n72212 , n35245 );
buf ( n72213 , n72212 );
not ( n72214 , n35292 );
and ( n72215 , n72206 , n72214 );
and ( n72216 , n72215 , n35245 );
or ( n72217 , n72213 , n72216 );
and ( n72218 , n72217 , n32419 );
not ( n72219 , n35278 );
buf ( n72220 , n72219 );
and ( n72221 , n72208 , n35278 );
or ( n72222 , n72220 , n72221 );
and ( n72223 , n72222 , n32417 );
not ( n72224 , n35331 );
buf ( n72225 , n72224 );
and ( n72226 , n72215 , n35331 );
or ( n72227 , n72225 , n72226 );
and ( n72228 , n72227 , n32415 );
not ( n72229 , n47331 );
and ( n72230 , n72229 , n32413 );
not ( n72231 , n50067 );
and ( n72232 , n72231 , n32411 );
not ( n72233 , n31728 );
and ( n72234 , n72233 , n32253 );
not ( n72235 , n32283 );
and ( n72236 , n72235 , n32398 );
or ( n72237 , n72211 , n72218 , n72223 , n72228 , n72230 , n72232 , n72234 , n72236 , C0 );
and ( n72238 , n72237 , n32456 );
and ( n72239 , n72206 , n47409 );
or ( n72240 , C0 , n72238 , n72239 );
buf ( n72241 , n72240 );
buf ( n72242 , n72241 );
buf ( n72243 , n31655 );
not ( n72244 , n36587 );
and ( n72245 , n72244 , n36260 );
xor ( n72246 , n50185 , n50202 );
and ( n72247 , n72246 , n36587 );
or ( n72248 , n72245 , n72247 );
and ( n72249 , n72248 , n36596 );
not ( n72250 , n37485 );
and ( n72251 , n72250 , n37162 );
xor ( n72252 , n50235 , n50252 );
and ( n72253 , n72252 , n37485 );
or ( n72254 , n72251 , n72253 );
and ( n72255 , n72254 , n37494 );
and ( n72256 , n41849 , n37506 );
or ( n72257 , n72249 , n72255 , n72256 );
buf ( n72258 , n72257 );
buf ( n72259 , n72258 );
buf ( n72260 , n30987 );
not ( n72261 , n46356 );
and ( n72262 , n72261 , n31150 );
not ( n72263 , n53353 );
and ( n72264 , n72263 , n31150 );
and ( n72265 , n31172 , n53353 );
or ( n72266 , n72264 , n72265 );
and ( n72267 , n72266 , n46356 );
or ( n72268 , n72262 , n72267 );
and ( n72269 , n72268 , n31649 );
not ( n72270 , n53361 );
not ( n72271 , n53353 );
and ( n72272 , n72271 , n31150 );
and ( n72273 , n46495 , n53353 );
or ( n72274 , n72272 , n72273 );
and ( n72275 , n72270 , n72274 );
and ( n72276 , n46495 , n53361 );
or ( n72277 , n72275 , n72276 );
and ( n72278 , n72277 , n31643 );
not ( n72279 , n31452 );
not ( n72280 , n53361 );
not ( n72281 , n53353 );
and ( n72282 , n72281 , n31150 );
and ( n72283 , n46495 , n53353 );
or ( n72284 , n72282 , n72283 );
and ( n72285 , n72280 , n72284 );
and ( n72286 , n46495 , n53361 );
or ( n72287 , n72285 , n72286 );
and ( n72288 , n72279 , n72287 );
not ( n72289 , n53381 );
not ( n72290 , n53383 );
and ( n72291 , n72290 , n72287 );
and ( n72292 , n46984 , n53383 );
or ( n72293 , n72291 , n72292 );
and ( n72294 , n72289 , n72293 );
and ( n72295 , n47267 , n53381 );
or ( n72296 , n72294 , n72295 );
and ( n72297 , n72296 , n31452 );
or ( n72298 , n72288 , n72297 );
and ( n72299 , n72298 , n31638 );
and ( n72300 , n31150 , n47277 );
or ( n72301 , C0 , n72269 , n72278 , n72299 , n72300 );
buf ( n72302 , n72301 );
buf ( n72303 , n72302 );
buf ( n72304 , n30987 );
buf ( n72305 , n31655 );
and ( n72306 , n59206 , n32494 );
not ( n72307 , n46083 );
and ( n72308 , n72307 , n61595 );
buf ( n72309 , n72308 );
and ( n72310 , n72309 , n32421 );
not ( n72311 , n46326 );
and ( n72312 , n72311 , n61595 );
and ( n72313 , n59216 , n46326 );
or ( n72314 , n72312 , n72313 );
and ( n72315 , n72314 , n32417 );
and ( n72316 , n61595 , n46340 );
or ( n72317 , n72310 , n72315 , n72316 );
and ( n72318 , n72317 , n32456 );
and ( n72319 , n61595 , n46349 );
or ( n72320 , C0 , n72306 , n72318 , n72319 );
buf ( n72321 , n72320 );
buf ( n72322 , n72321 );
buf ( n72323 , n31655 );
buf ( n72324 , n30987 );
buf ( n72325 , n31655 );
buf ( n72326 , n31655 );
buf ( n72327 , n30987 );
and ( n72328 , n49091 , n48639 );
not ( n72329 , n48642 );
and ( n72330 , n72329 , n48610 );
and ( n72331 , n49091 , n48642 );
or ( n72332 , n72330 , n72331 );
and ( n72333 , n72332 , n32890 );
not ( n72334 , n48648 );
and ( n72335 , n72334 , n48610 );
and ( n72336 , n49091 , n48648 );
or ( n72337 , n72335 , n72336 );
and ( n72338 , n72337 , n32924 );
not ( n72339 , n48654 );
and ( n72340 , n72339 , n48610 );
and ( n72341 , n49091 , n48654 );
or ( n72342 , n72340 , n72341 );
and ( n72343 , n72342 , n33038 );
not ( n72344 , n48660 );
and ( n72345 , n72344 , n48610 );
and ( n72346 , n49091 , n48660 );
or ( n72347 , n72345 , n72346 );
and ( n72348 , n72347 , n33172 );
not ( n72349 , n41576 );
and ( n72350 , n72349 , n48610 );
and ( n72351 , n48942 , n41576 );
or ( n72352 , n72350 , n72351 );
and ( n72353 , n72352 , n33189 );
not ( n72354 , n48730 );
and ( n72355 , n72354 , n48610 );
and ( n72356 , n48942 , n48730 );
or ( n72357 , n72355 , n72356 );
and ( n72358 , n72357 , n33187 );
not ( n72359 , n48765 );
and ( n72360 , n72359 , n48610 );
and ( n72361 , n66781 , n48765 );
or ( n72362 , n72360 , n72361 );
and ( n72363 , n72362 , n33180 );
not ( n72364 , n49054 );
and ( n72365 , n72364 , n48610 );
and ( n72366 , n66794 , n49054 );
or ( n72367 , n72365 , n72366 );
and ( n72368 , n72367 , n33178 );
and ( n72369 , n49212 , n49275 );
or ( n72370 , n72328 , n72333 , n72338 , n72343 , n72348 , n72353 , n72358 , n72363 , n72368 , n72369 );
and ( n72371 , n72370 , n33208 );
and ( n72372 , n33003 , n35056 );
and ( n72373 , n48610 , n49286 );
or ( n72374 , C0 , n72371 , n72372 , n72373 );
buf ( n72375 , n72374 );
buf ( n72376 , n72375 );
not ( n72377 , n34150 );
and ( n72378 , n72377 , n32714 );
not ( n72379 , n56093 );
and ( n72380 , n72379 , n32714 );
and ( n72381 , n32722 , n56093 );
or ( n72382 , n72380 , n72381 );
and ( n72383 , n72382 , n34150 );
or ( n72384 , n72378 , n72383 );
and ( n72385 , n72384 , n33381 );
not ( n72386 , n56101 );
not ( n72387 , n56093 );
and ( n72388 , n72387 , n32714 );
and ( n72389 , n42565 , n56093 );
or ( n72390 , n72388 , n72389 );
and ( n72391 , n72386 , n72390 );
and ( n72392 , n42565 , n56101 );
or ( n72393 , n72391 , n72392 );
and ( n72394 , n72393 , n33375 );
not ( n72395 , n32968 );
not ( n72396 , n56101 );
not ( n72397 , n56093 );
and ( n72398 , n72397 , n32714 );
and ( n72399 , n42565 , n56093 );
or ( n72400 , n72398 , n72399 );
and ( n72401 , n72396 , n72400 );
and ( n72402 , n42565 , n56101 );
or ( n72403 , n72401 , n72402 );
and ( n72404 , n72395 , n72403 );
not ( n72405 , n56121 );
not ( n72406 , n56123 );
and ( n72407 , n72406 , n72403 );
and ( n72408 , n42589 , n56123 );
or ( n72409 , n72407 , n72408 );
and ( n72410 , n72405 , n72409 );
and ( n72411 , n42597 , n56121 );
or ( n72412 , n72410 , n72411 );
and ( n72413 , n72412 , n32968 );
or ( n72414 , n72404 , n72413 );
and ( n72415 , n72414 , n33370 );
and ( n72416 , n32714 , n35062 );
or ( n72417 , C0 , n72385 , n72394 , n72415 , n72416 );
buf ( n72418 , n72417 );
buf ( n72419 , n72418 );
not ( n72420 , n34150 );
and ( n72421 , n72420 , n32819 );
not ( n72422 , n56140 );
and ( n72423 , n72422 , n32819 );
and ( n72424 , n32823 , n56140 );
or ( n72425 , n72423 , n72424 );
and ( n72426 , n72425 , n34150 );
or ( n72427 , n72421 , n72426 );
and ( n72428 , n72427 , n33381 );
not ( n72429 , n56148 );
not ( n72430 , n56140 );
and ( n72431 , n72430 , n32819 );
and ( n72432 , n41464 , n56140 );
or ( n72433 , n72431 , n72432 );
and ( n72434 , n72429 , n72433 );
and ( n72435 , n41464 , n56148 );
or ( n72436 , n72434 , n72435 );
and ( n72437 , n72436 , n33375 );
not ( n72438 , n32968 );
not ( n72439 , n56148 );
not ( n72440 , n56140 );
and ( n72441 , n72440 , n32819 );
and ( n72442 , n41464 , n56140 );
or ( n72443 , n72441 , n72442 );
and ( n72444 , n72439 , n72443 );
and ( n72445 , n41464 , n56148 );
or ( n72446 , n72444 , n72445 );
and ( n72447 , n72438 , n72446 );
not ( n72448 , n56168 );
not ( n72449 , n56170 );
and ( n72450 , n72449 , n72446 );
and ( n72451 , n41490 , n56170 );
or ( n72452 , n72450 , n72451 );
and ( n72453 , n72448 , n72452 );
and ( n72454 , n41500 , n56168 );
or ( n72455 , n72453 , n72454 );
and ( n72456 , n72455 , n32968 );
or ( n72457 , n72447 , n72456 );
and ( n72458 , n72457 , n33370 );
and ( n72459 , n32819 , n35062 );
or ( n72460 , C0 , n72428 , n72437 , n72458 , n72459 );
buf ( n72461 , n72460 );
buf ( n72462 , n72461 );
buf ( n72463 , n30987 );
buf ( n72464 , n31655 );
buf ( n72465 , n31655 );
buf ( n72466 , n30987 );
buf ( n72467 , n31655 );
buf ( n72468 , n30987 );
not ( n72469 , n32953 );
and ( n72470 , n72469 , n61336 );
not ( n72471 , n39572 );
and ( n72472 , n72471 , n39464 );
xor ( n72473 , n42621 , n42632 );
and ( n72474 , n72473 , n39572 );
or ( n72475 , n72472 , n72474 );
and ( n72476 , n72475 , n32953 );
or ( n72477 , n72470 , n72476 );
and ( n72478 , n72477 , n33038 );
not ( n72479 , n39586 );
and ( n72480 , n72479 , n61336 );
and ( n72481 , n61342 , n39586 );
or ( n72482 , n72480 , n72481 );
and ( n72483 , n72482 , n33172 );
and ( n72484 , n61336 , n39795 );
or ( n72485 , n72478 , n72483 , n72484 );
and ( n72486 , n72485 , n33208 );
and ( n72487 , n61336 , n39805 );
or ( n72488 , C0 , n72486 , n72487 );
buf ( n72489 , n72488 );
buf ( n72490 , n72489 );
buf ( n72491 , n30987 );
buf ( n72492 , n31655 );
buf ( n72493 , n30987 );
buf ( n72494 , n31655 );
xor ( n72495 , n44768 , n44799 );
and ( n72496 , n72495 , n31548 );
not ( n72497 , n44807 );
and ( n72498 , n72497 , n44768 );
and ( n72499 , n46637 , n44807 );
or ( n72500 , n72498 , n72499 );
and ( n72501 , n72500 , n31408 );
not ( n72502 , n44817 );
and ( n72503 , n72502 , n44768 );
and ( n72504 , n60757 , n44817 );
or ( n72505 , n72503 , n72504 );
and ( n72506 , n72505 , n31521 );
not ( n72507 , n45059 );
and ( n72508 , n72507 , n44768 );
xor ( n72509 , n40052 , n45130 );
and ( n72510 , n72509 , n45059 );
or ( n72511 , n72508 , n72510 );
and ( n72512 , n72511 , n31536 );
and ( n72513 , n44768 , n45148 );
or ( n72514 , n72496 , n72501 , n72506 , n72512 , n72513 );
and ( n72515 , n72514 , n31557 );
and ( n72516 , n44768 , n40154 );
or ( n72517 , C0 , n72515 , n72516 );
buf ( n72518 , n72517 );
buf ( n72519 , n72518 );
not ( n72520 , n40163 );
and ( n72521 , n72520 , n32056 );
not ( n72522 , n55888 );
and ( n72523 , n72522 , n32056 );
and ( n72524 , n32130 , n55888 );
or ( n72525 , n72523 , n72524 );
and ( n72526 , n72525 , n40163 );
or ( n72527 , n72521 , n72526 );
and ( n72528 , n72527 , n32498 );
not ( n72529 , n55896 );
not ( n72530 , n55888 );
and ( n72531 , n72530 , n32056 );
and ( n72532 , n45833 , n55888 );
or ( n72533 , n72531 , n72532 );
and ( n72534 , n72529 , n72533 );
and ( n72535 , n45833 , n55896 );
or ( n72536 , n72534 , n72535 );
and ( n72537 , n72536 , n32473 );
not ( n72538 , n32475 );
not ( n72539 , n55896 );
not ( n72540 , n55888 );
and ( n72541 , n72540 , n32056 );
and ( n72542 , n45833 , n55888 );
or ( n72543 , n72541 , n72542 );
and ( n72544 , n72539 , n72543 );
and ( n72545 , n45833 , n55896 );
or ( n72546 , n72544 , n72545 );
and ( n72547 , n72538 , n72546 );
not ( n72548 , n55916 );
not ( n72549 , n55918 );
and ( n72550 , n72549 , n72546 );
and ( n72551 , n45857 , n55918 );
or ( n72552 , n72550 , n72551 );
and ( n72553 , n72548 , n72552 );
and ( n72554 , n45865 , n55916 );
or ( n72555 , n72553 , n72554 );
and ( n72556 , n72555 , n32475 );
or ( n72557 , n72547 , n72556 );
and ( n72558 , n72557 , n32486 );
and ( n72559 , n32056 , n41278 );
or ( n72560 , C0 , n72528 , n72537 , n72558 , n72559 );
buf ( n72561 , n72560 );
buf ( n72562 , n72561 );
buf ( n72563 , n30987 );
not ( n72564 , n52719 );
not ( n72565 , n72564 );
or ( n72566 , n37499 , n37501 );
and ( n72567 , n72565 , n72566 );
buf ( n72568 , n37497 );
and ( n72569 , n31452 , n67908 );
or ( n72570 , n72567 , n72568 , n72569 );
buf ( n72571 , n72570 );
buf ( n72572 , n72571 );
buf ( n72573 , n30987 );
buf ( n72574 , n30987 );
not ( n72575 , n40163 );
and ( n72576 , n72575 , n31875 );
not ( n72577 , n52120 );
and ( n72578 , n72577 , n31875 );
and ( n72579 , n32218 , n52120 );
or ( n72580 , n72578 , n72579 );
and ( n72581 , n72580 , n40163 );
or ( n72582 , n72576 , n72581 );
and ( n72583 , n72582 , n32498 );
not ( n72584 , n52128 );
not ( n72585 , n52120 );
and ( n72586 , n72585 , n31875 );
and ( n72587 , n42255 , n52120 );
or ( n72588 , n72586 , n72587 );
and ( n72589 , n72584 , n72588 );
and ( n72590 , n42255 , n52128 );
or ( n72591 , n72589 , n72590 );
and ( n72592 , n72591 , n32473 );
not ( n72593 , n32475 );
not ( n72594 , n52128 );
not ( n72595 , n52120 );
and ( n72596 , n72595 , n31875 );
and ( n72597 , n42255 , n52120 );
or ( n72598 , n72596 , n72597 );
and ( n72599 , n72594 , n72598 );
and ( n72600 , n42255 , n52128 );
or ( n72601 , n72599 , n72600 );
and ( n72602 , n72593 , n72601 );
not ( n72603 , n52148 );
not ( n72604 , n52150 );
and ( n72605 , n72604 , n72601 );
and ( n72606 , n42283 , n52150 );
or ( n72607 , n72605 , n72606 );
and ( n72608 , n72603 , n72607 );
and ( n72609 , n42291 , n52148 );
or ( n72610 , n72608 , n72609 );
and ( n72611 , n72610 , n32475 );
or ( n72612 , n72602 , n72611 );
and ( n72613 , n72612 , n32486 );
and ( n72614 , n31875 , n41278 );
or ( n72615 , C0 , n72583 , n72592 , n72613 , n72614 );
buf ( n72616 , n72615 );
buf ( n72617 , n72616 );
buf ( n72618 , n31655 );
buf ( n72619 , n31655 );
and ( n72620 , n48799 , n34150 );
buf ( n72621 , n72620 );
and ( n72622 , n72621 , n33381 );
and ( n72623 , n56683 , n33379 );
and ( n72624 , n57711 , n33208 );
and ( n72625 , n32543 , n61311 );
or ( n72626 , C0 , n72622 , n72623 , n72624 , n72625 );
buf ( n72627 , n72626 );
buf ( n72628 , n72627 );
buf ( n72629 , n31655 );
buf ( n72630 , n30987 );
buf ( n72631 , n30987 );
buf ( n72632 , n30987 );
xor ( n72633 , n49599 , n60306 );
and ( n72634 , n72633 , n32433 );
not ( n72635 , n47331 );
and ( n72636 , n72635 , n49599 );
and ( n72637 , n31931 , n47357 );
and ( n72638 , n31933 , n47359 );
and ( n72639 , n31935 , n47361 );
and ( n72640 , n31937 , n47363 );
and ( n72641 , n31939 , n47365 );
and ( n72642 , n31941 , n47367 );
and ( n72643 , n31943 , n47369 );
and ( n72644 , n31945 , n47371 );
and ( n72645 , n31947 , n47373 );
and ( n72646 , n31949 , n47375 );
and ( n72647 , n31951 , n47377 );
and ( n72648 , n31953 , n47379 );
and ( n72649 , n31955 , n47381 );
and ( n72650 , n31957 , n47383 );
and ( n72651 , n31959 , n47385 );
and ( n72652 , n31961 , n47387 );
or ( n72653 , n72637 , n72638 , n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , n72651 , n72652 );
and ( n72654 , n72653 , n47331 );
or ( n72655 , n72636 , n72654 );
and ( n72656 , n72655 , n32413 );
and ( n72657 , n49599 , n47402 );
or ( n72658 , n72634 , n72656 , n72657 );
and ( n72659 , n72658 , n32456 );
and ( n72660 , n49599 , n47409 );
or ( n72661 , C0 , n72659 , n72660 );
buf ( n72662 , n72661 );
buf ( n72663 , n72662 );
not ( n72664 , n35542 );
and ( n72665 , n72664 , n41843 );
buf ( n72666 , RI15b45258_224);
and ( n72667 , n72666 , n35542 );
or ( n72668 , n72665 , n72667 );
buf ( n72669 , n72668 );
buf ( n72670 , n72669 );
not ( n72671 , n46356 );
and ( n72672 , n72671 , n31300 );
not ( n72673 , n47423 );
and ( n72674 , n72673 , n31300 );
and ( n72675 , n31306 , n47423 );
or ( n72676 , n72674 , n72675 );
and ( n72677 , n72676 , n46356 );
or ( n72678 , n72672 , n72677 );
and ( n72679 , n72678 , n31649 );
not ( n72680 , n47431 );
not ( n72681 , n47423 );
and ( n72682 , n72681 , n31300 );
and ( n72683 , n58061 , n47423 );
or ( n72684 , n72682 , n72683 );
and ( n72685 , n72680 , n72684 );
and ( n72686 , n58061 , n47431 );
or ( n72687 , n72685 , n72686 );
and ( n72688 , n72687 , n31643 );
not ( n72689 , n31452 );
not ( n72690 , n47431 );
not ( n72691 , n47423 );
and ( n72692 , n72691 , n31300 );
and ( n72693 , n58061 , n47423 );
or ( n72694 , n72692 , n72693 );
and ( n72695 , n72690 , n72694 );
and ( n72696 , n58061 , n47431 );
or ( n72697 , n72695 , n72696 );
and ( n72698 , n72689 , n72697 );
not ( n72699 , n47466 );
not ( n72700 , n47468 );
and ( n72701 , n72700 , n72697 );
and ( n72702 , n58085 , n47468 );
or ( n72703 , n72701 , n72702 );
and ( n72704 , n72699 , n72703 );
and ( n72705 , n58093 , n47466 );
or ( n72706 , n72704 , n72705 );
and ( n72707 , n72706 , n31452 );
or ( n72708 , n72698 , n72707 );
and ( n72709 , n72708 , n31638 );
and ( n72710 , n31300 , n47277 );
or ( n72711 , C0 , n72679 , n72688 , n72709 , n72710 );
buf ( n72712 , n72711 );
buf ( n72713 , n72712 );
buf ( n72714 , n31655 );
buf ( n72715 , n31655 );
and ( n72716 , n39367 , n33377 );
not ( n72717 , n48545 );
buf ( n72718 , RI15b46f68_286);
and ( n72719 , n72717 , n72718 );
and ( n72720 , n39580 , n48545 );
or ( n72721 , n72719 , n72720 );
and ( n72722 , n72721 , n32890 );
not ( n72723 , n48557 );
and ( n72724 , n72723 , n72718 );
and ( n72725 , n39580 , n48557 );
or ( n72726 , n72724 , n72725 );
and ( n72727 , n72726 , n33038 );
and ( n72728 , n72718 , n48571 );
or ( n72729 , n72722 , n72727 , n72728 );
and ( n72730 , n72729 , n33208 );
and ( n72731 , n72718 , n48577 );
or ( n72732 , C0 , n72716 , n72730 , n72731 );
buf ( n72733 , n72732 );
buf ( n72734 , n72733 );
buf ( n72735 , n31655 );
buf ( n72736 , n31655 );
buf ( n72737 , n30987 );
buf ( n72738 , n30987 );
buf ( n72739 , n30987 );
buf ( n72740 , n31655 );
buf ( n72741 , n40199 );
not ( n72742 , n34150 );
and ( n72743 , n72742 , n32840 );
not ( n72744 , n57038 );
and ( n72745 , n72744 , n32840 );
and ( n72746 , n32856 , n57038 );
or ( n72747 , n72745 , n72746 );
and ( n72748 , n72747 , n34150 );
or ( n72749 , n72743 , n72748 );
and ( n72750 , n72749 , n33381 );
not ( n72751 , n57046 );
not ( n72752 , n57038 );
and ( n72753 , n72752 , n32840 );
and ( n72754 , n48160 , n57038 );
or ( n72755 , n72753 , n72754 );
and ( n72756 , n72751 , n72755 );
and ( n72757 , n48160 , n57046 );
or ( n72758 , n72756 , n72757 );
and ( n72759 , n72758 , n33375 );
not ( n72760 , n32968 );
not ( n72761 , n57046 );
not ( n72762 , n57038 );
and ( n72763 , n72762 , n32840 );
and ( n72764 , n48160 , n57038 );
or ( n72765 , n72763 , n72764 );
and ( n72766 , n72761 , n72765 );
and ( n72767 , n48160 , n57046 );
or ( n72768 , n72766 , n72767 );
and ( n72769 , n72760 , n72768 );
not ( n72770 , n57066 );
not ( n72771 , n57068 );
and ( n72772 , n72771 , n72768 );
and ( n72773 , n48186 , n57068 );
or ( n72774 , n72772 , n72773 );
and ( n72775 , n72770 , n72774 );
and ( n72776 , n48196 , n57066 );
or ( n72777 , n72775 , n72776 );
and ( n72778 , n72777 , n32968 );
or ( n72779 , n72769 , n72778 );
and ( n72780 , n72779 , n33370 );
and ( n72781 , n32840 , n35062 );
or ( n72782 , C0 , n72750 , n72759 , n72780 , n72781 );
buf ( n72783 , n72782 );
buf ( n72784 , n72783 );
buf ( n72785 , n31655 );
buf ( n72786 , n30987 );
buf ( n72787 , n30987 );
and ( n72788 , n31561 , n31007 );
not ( n72789 , n31077 );
and ( n72790 , n72789 , n35387 );
buf ( n72791 , n72790 );
and ( n72792 , n72791 , n31373 );
not ( n72793 , n31402 );
and ( n72794 , n72793 , n35387 );
buf ( n72795 , n72794 );
and ( n72796 , n72795 , n31408 );
not ( n72797 , n31437 );
and ( n72798 , n72797 , n35387 );
not ( n72799 , n31455 );
and ( n72800 , n72799 , n35423 );
xor ( n72801 , n35387 , n35411 );
and ( n72802 , n72801 , n31455 );
or ( n72803 , n72800 , n72802 );
and ( n72804 , n72803 , n31437 );
or ( n72805 , n72798 , n72804 );
and ( n72806 , n72805 , n31468 );
not ( n72807 , n31497 );
and ( n72808 , n72807 , n35387 );
not ( n72809 , n31454 );
not ( n72810 , n31501 );
and ( n72811 , n72810 , n35423 );
xor ( n72812 , n35424 , n35461 );
and ( n72813 , n72812 , n31501 );
or ( n72814 , n72811 , n72813 );
and ( n72815 , n72809 , n72814 );
and ( n72816 , n72801 , n31454 );
or ( n72817 , n72815 , n72816 );
and ( n72818 , n72817 , n31497 );
or ( n72819 , n72808 , n72818 );
and ( n72820 , n72819 , n31521 );
and ( n72821 , n35387 , n31553 );
or ( n72822 , n72792 , n72796 , n72806 , n72820 , n72821 );
and ( n72823 , n72822 , n31557 );
not ( n72824 , n31452 );
not ( n72825 , n31619 );
and ( n72826 , n72825 , n35478 );
xor ( n72827 , n35479 , n35515 );
and ( n72828 , n72827 , n31619 );
or ( n72829 , n72826 , n72828 );
and ( n72830 , n72824 , n72829 );
and ( n72831 , n35387 , n31452 );
or ( n72832 , n72830 , n72831 );
and ( n72833 , n72832 , n31638 );
and ( n72834 , n35387 , n31650 );
or ( n72835 , C0 , n72788 , n72823 , n72833 , C0 , n72834 );
buf ( n72836 , n72835 );
buf ( n72837 , n72836 );
buf ( n72838 , n54726 );
buf ( n72839 , n31655 );
not ( n72840 , n33419 );
and ( n72841 , n72840 , n31583 );
xor ( n72842 , n33477 , n33688 );
and ( n72843 , n72842 , n33419 );
or ( n72844 , n72841 , n72843 );
and ( n72845 , n72844 , n31529 );
not ( n72846 , n33734 );
and ( n72847 , n72846 , n31583 );
not ( n72848 , n33533 );
xor ( n72849 , n33770 , n33806 );
and ( n72850 , n72848 , n72849 );
xnor ( n72851 , n33855 , n33908 );
and ( n72852 , n72851 , n33533 );
or ( n72853 , n72850 , n72852 );
and ( n72854 , n72853 , n33734 );
or ( n72855 , n72847 , n72854 );
and ( n72856 , n72855 , n31527 );
and ( n72857 , n31583 , n33942 );
or ( n72858 , n72845 , n72856 , n72857 );
and ( n72859 , n72858 , n31557 );
and ( n72860 , n34111 , n31643 );
not ( n72861 , n31452 );
and ( n72862 , n72861 , n34111 );
xor ( n72863 , n31583 , n33954 );
and ( n72864 , n72863 , n31452 );
or ( n72865 , n72862 , n72864 );
and ( n72866 , n72865 , n31638 );
and ( n72867 , n34007 , n33973 );
and ( n72868 , n31583 , n33978 );
or ( n72869 , C0 , n72859 , n72860 , n72866 , n72867 , n72868 );
buf ( n72870 , n72869 );
buf ( n72871 , n72870 );
buf ( n72872 , n30987 );
buf ( n72873 , n31655 );
buf ( n72874 , n30987 );
not ( n72875 , n32953 );
buf ( n72876 , RI15b461d0_257);
and ( n72877 , n72875 , n72876 );
not ( n72878 , n54581 );
and ( n72879 , n72878 , n54390 );
xor ( n72880 , n64019 , n64022 );
and ( n72881 , n72880 , n54581 );
or ( n72882 , n72879 , n72881 );
and ( n72883 , n72882 , n32953 );
or ( n72884 , n72877 , n72883 );
and ( n72885 , n72884 , n33038 );
not ( n72886 , n48660 );
and ( n72887 , n72886 , n72876 );
not ( n72888 , n55168 );
and ( n72889 , n72888 , n55032 );
xor ( n72890 , n55173 , n55179 );
and ( n72891 , n72890 , n55168 );
or ( n72892 , n72889 , n72891 );
and ( n72893 , n72892 , n48660 );
or ( n72894 , n72887 , n72893 );
and ( n72895 , n72894 , n33172 );
and ( n72896 , n72876 , n39795 );
or ( n72897 , n72885 , n72895 , n72896 );
and ( n72898 , n72897 , n33208 );
and ( n72899 , n72876 , n39805 );
or ( n72900 , C0 , n72898 , n72899 );
buf ( n72901 , n72900 );
buf ( n72902 , n72901 );
buf ( n72903 , n30987 );
buf ( n72904 , n31655 );
buf ( n72905 , n30987 );
buf ( n72906 , n30987 );
buf ( n72907 , n31655 );
and ( n72908 , n64011 , n33377 );
not ( n72909 , n48545 );
and ( n72910 , n72909 , n41384 );
buf ( n72911 , n72910 );
and ( n72912 , n72911 , n32890 );
not ( n72913 , n48557 );
and ( n72914 , n72913 , n41384 );
and ( n72915 , n64029 , n48557 );
or ( n72916 , n72914 , n72915 );
and ( n72917 , n72916 , n33038 );
and ( n72918 , n41384 , n48571 );
or ( n72919 , n72912 , n72917 , n72918 );
and ( n72920 , n72919 , n33208 );
and ( n72921 , n41384 , n48577 );
or ( n72922 , C0 , n72908 , n72920 , n72921 );
buf ( n72923 , n72922 );
buf ( n72924 , n72923 );
buf ( n72925 , n31655 );
not ( n72926 , n46356 );
and ( n72927 , n72926 , n31296 );
not ( n72928 , n56904 );
and ( n72929 , n72928 , n31296 );
and ( n72930 , n31306 , n56904 );
or ( n72931 , n72929 , n72930 );
and ( n72932 , n72931 , n46356 );
or ( n72933 , n72927 , n72932 );
and ( n72934 , n72933 , n31649 );
not ( n72935 , n56912 );
not ( n72936 , n56904 );
and ( n72937 , n72936 , n31296 );
and ( n72938 , n58061 , n56904 );
or ( n72939 , n72937 , n72938 );
and ( n72940 , n72935 , n72939 );
and ( n72941 , n58061 , n56912 );
or ( n72942 , n72940 , n72941 );
and ( n72943 , n72942 , n31643 );
not ( n72944 , n31452 );
not ( n72945 , n56912 );
not ( n72946 , n56904 );
and ( n72947 , n72946 , n31296 );
and ( n72948 , n58061 , n56904 );
or ( n72949 , n72947 , n72948 );
and ( n72950 , n72945 , n72949 );
and ( n72951 , n58061 , n56912 );
or ( n72952 , n72950 , n72951 );
and ( n72953 , n72944 , n72952 );
not ( n72954 , n56937 );
not ( n72955 , n56939 );
and ( n72956 , n72955 , n72952 );
and ( n72957 , n58085 , n56939 );
or ( n72958 , n72956 , n72957 );
and ( n72959 , n72954 , n72958 );
and ( n72960 , n58093 , n56937 );
or ( n72961 , n72959 , n72960 );
and ( n72962 , n72961 , n31452 );
or ( n72963 , n72953 , n72962 );
and ( n72964 , n72963 , n31638 );
and ( n72965 , n31296 , n47277 );
or ( n72966 , C0 , n72934 , n72943 , n72964 , n72965 );
buf ( n72967 , n72966 );
buf ( n72968 , n72967 );
buf ( n72969 , n31655 );
buf ( n72970 , RI15b472b0_293);
buf ( n72971 , n72970 );
buf ( n72972 , n30987 );
and ( n72973 , n50955 , n70040 );
xor ( n72974 , n50953 , n72973 );
and ( n72975 , n72974 , n32431 );
not ( n72976 , n50002 );
and ( n72977 , n72976 , n50953 );
and ( n72978 , n40578 , n50002 );
or ( n72979 , n72977 , n72978 );
and ( n72980 , n72979 , n32419 );
not ( n72981 , n50008 );
and ( n72982 , n72981 , n50953 );
not ( n72983 , n51594 );
and ( n72984 , n72983 , n51554 );
xor ( n72985 , n59226 , n59235 );
and ( n72986 , n72985 , n51594 );
or ( n72987 , n72984 , n72986 );
and ( n72988 , n72987 , n50008 );
or ( n72989 , n72982 , n72988 );
and ( n72990 , n72989 , n32415 );
not ( n72991 , n50067 );
and ( n72992 , n72991 , n50953 );
and ( n72993 , n60433 , n70060 );
xor ( n72994 , n60416 , n72993 );
and ( n72995 , n72994 , n50067 );
or ( n72996 , n72992 , n72995 );
and ( n72997 , n72996 , n32411 );
and ( n72998 , n50953 , n50098 );
or ( n72999 , n72975 , n72980 , n72990 , n72997 , n72998 );
and ( n73000 , n72999 , n32456 );
and ( n73001 , n50953 , n47409 );
or ( n73002 , C0 , n73000 , n73001 );
buf ( n73003 , n73002 );
buf ( n73004 , n73003 );
buf ( n73005 , n31655 );
xor ( n73006 , n54154 , n54982 );
and ( n73007 , n73006 , n33199 );
not ( n73008 , n48648 );
and ( n73009 , n73008 , n54154 );
and ( n73010 , n34439 , n48648 );
or ( n73011 , n73009 , n73010 );
and ( n73012 , n73011 , n32924 );
not ( n73013 , n48660 );
and ( n73014 , n73013 , n54154 );
and ( n73015 , n72892 , n48660 );
or ( n73016 , n73014 , n73015 );
and ( n73017 , n73016 , n33172 );
not ( n73018 , n48730 );
and ( n73019 , n73018 , n54154 );
and ( n73020 , n32723 , n55215 );
and ( n73021 , n32725 , n55217 );
and ( n73022 , n32727 , n55219 );
and ( n73023 , n32729 , n55221 );
and ( n73024 , n32731 , n55223 );
and ( n73025 , n32733 , n55225 );
and ( n73026 , n32735 , n55227 );
and ( n73027 , n32737 , n55229 );
and ( n73028 , n32739 , n55231 );
and ( n73029 , n32741 , n55233 );
and ( n73030 , n32743 , n55235 );
and ( n73031 , n32745 , n55237 );
and ( n73032 , n32747 , n55239 );
and ( n73033 , n32749 , n55241 );
and ( n73034 , n32751 , n55243 );
and ( n73035 , n32753 , n55245 );
or ( n73036 , n73020 , n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , n73035 );
and ( n73037 , n73036 , n48730 );
or ( n73038 , n73019 , n73037 );
and ( n73039 , n73038 , n33187 );
and ( n73040 , n54154 , n54713 );
or ( n73041 , n73007 , n73012 , n73017 , n73039 , n73040 );
and ( n73042 , n73041 , n33208 );
and ( n73043 , n54154 , n39805 );
or ( n73044 , C0 , n73042 , n73043 );
buf ( n73045 , n73044 );
buf ( n73046 , n73045 );
buf ( n73047 , n30987 );
buf ( n73048 , n31655 );
not ( n73049 , n41532 );
and ( n73050 , n73049 , n34439 );
and ( n73051 , n54606 , n41532 );
or ( n73052 , n73050 , n73051 );
buf ( n73053 , n73052 );
buf ( n73054 , n73053 );
buf ( n73055 , n31655 );
buf ( n73056 , n30987 );
buf ( n73057 , n31655 );
buf ( n73058 , n31655 );
buf ( n73059 , n30987 );
not ( n73060 , n46356 );
and ( n73061 , n73060 , n31210 );
not ( n73062 , n55473 );
and ( n73063 , n73062 , n31210 );
and ( n73064 , n31238 , n55473 );
or ( n73065 , n73063 , n73064 );
and ( n73066 , n73065 , n46356 );
or ( n73067 , n73061 , n73066 );
and ( n73068 , n73067 , n31649 );
not ( n73069 , n55481 );
not ( n73070 , n55473 );
and ( n73071 , n73070 , n31210 );
and ( n73072 , n49901 , n55473 );
or ( n73073 , n73071 , n73072 );
and ( n73074 , n73069 , n73073 );
and ( n73075 , n49901 , n55481 );
or ( n73076 , n73074 , n73075 );
and ( n73077 , n73076 , n31643 );
not ( n73078 , n31452 );
not ( n73079 , n55481 );
not ( n73080 , n55473 );
and ( n73081 , n73080 , n31210 );
and ( n73082 , n49901 , n55473 );
or ( n73083 , n73081 , n73082 );
and ( n73084 , n73079 , n73083 );
and ( n73085 , n49901 , n55481 );
or ( n73086 , n73084 , n73085 );
and ( n73087 , n73078 , n73086 );
not ( n73088 , n55501 );
not ( n73089 , n55503 );
and ( n73090 , n73089 , n73086 );
and ( n73091 , n49925 , n55503 );
or ( n73092 , n73090 , n73091 );
and ( n73093 , n73088 , n73092 );
and ( n73094 , n49933 , n55501 );
or ( n73095 , n73093 , n73094 );
and ( n73096 , n73095 , n31452 );
or ( n73097 , n73087 , n73096 );
and ( n73098 , n73097 , n31638 );
and ( n73099 , n31210 , n47277 );
or ( n73100 , C0 , n73068 , n73077 , n73098 , n73099 );
buf ( n73101 , n73100 );
buf ( n73102 , n73101 );
and ( n73103 , n64567 , n32494 );
not ( n73104 , n46083 );
buf ( n73105 , RI15b5f928_1126);
and ( n73106 , n73104 , n73105 );
not ( n73107 , n46290 );
and ( n73108 , n73107 , n46130 );
xor ( n73109 , n46303 , n46309 );
and ( n73110 , n73109 , n46290 );
or ( n73111 , n73108 , n73110 );
and ( n73112 , n73111 , n46083 );
or ( n73113 , n73106 , n73112 );
and ( n73114 , n73113 , n32421 );
not ( n73115 , n46326 );
and ( n73116 , n73115 , n73105 );
and ( n73117 , n73111 , n46326 );
or ( n73118 , n73116 , n73117 );
and ( n73119 , n73118 , n32417 );
and ( n73120 , n73105 , n46340 );
or ( n73121 , n73114 , n73119 , n73120 );
and ( n73122 , n73121 , n32456 );
and ( n73123 , n73105 , n46349 );
or ( n73124 , C0 , n73103 , n73122 , n73123 );
buf ( n73125 , n73124 );
buf ( n73126 , n73125 );
and ( n73127 , n58809 , n31645 );
not ( n73128 , n45274 );
buf ( n73129 , RI15b536a0_711);
and ( n73130 , n73128 , n73129 );
and ( n73131 , n58815 , n45274 );
or ( n73132 , n73130 , n73131 );
and ( n73133 , n73132 , n31373 );
not ( n73134 , n45280 );
and ( n73135 , n73134 , n73129 );
and ( n73136 , n58815 , n45280 );
or ( n73137 , n73135 , n73136 );
and ( n73138 , n73137 , n31468 );
and ( n73139 , n73129 , n45802 );
or ( n73140 , n73133 , n73138 , n73139 );
and ( n73141 , n73140 , n31557 );
and ( n73142 , n73129 , n45808 );
or ( n73143 , C0 , n73127 , n73141 , n73142 );
buf ( n73144 , n73143 );
buf ( n73145 , n73144 );
buf ( n73146 , n31655 );
buf ( n73147 , n30987 );
not ( n73148 , n40163 );
and ( n73149 , n73148 , n31784 );
not ( n73150 , n53227 );
and ( n73151 , n73150 , n31784 );
and ( n73152 , n32252 , n53227 );
or ( n73153 , n73151 , n73152 );
and ( n73154 , n73153 , n40163 );
or ( n73155 , n73149 , n73154 );
and ( n73156 , n73155 , n32498 );
not ( n73157 , n53235 );
not ( n73158 , n53227 );
and ( n73159 , n73158 , n31784 );
and ( n73160 , n40393 , n53227 );
or ( n73161 , n73159 , n73160 );
and ( n73162 , n73157 , n73161 );
and ( n73163 , n40393 , n53235 );
or ( n73164 , n73162 , n73163 );
and ( n73165 , n73164 , n32473 );
not ( n73166 , n32475 );
not ( n73167 , n53235 );
not ( n73168 , n53227 );
and ( n73169 , n73168 , n31784 );
and ( n73170 , n40393 , n53227 );
or ( n73171 , n73169 , n73170 );
and ( n73172 , n73167 , n73171 );
and ( n73173 , n40393 , n53235 );
or ( n73174 , n73172 , n73173 );
and ( n73175 , n73166 , n73174 );
not ( n73176 , n53260 );
not ( n73177 , n53262 );
and ( n73178 , n73177 , n73174 );
and ( n73179 , n40972 , n53262 );
or ( n73180 , n73178 , n73179 );
and ( n73181 , n73176 , n73180 );
and ( n73182 , n41267 , n53260 );
or ( n73183 , n73181 , n73182 );
and ( n73184 , n73183 , n32475 );
or ( n73185 , n73175 , n73184 );
and ( n73186 , n73185 , n32486 );
and ( n73187 , n31784 , n41278 );
or ( n73188 , C0 , n73156 , n73165 , n73186 , n73187 );
buf ( n73189 , n73188 );
buf ( n73190 , n73189 );
buf ( n73191 , n30987 );
buf ( n73192 , n31655 );
not ( n73193 , n34150 );
and ( n73194 , n73193 , n32735 );
not ( n73195 , n57872 );
and ( n73196 , n73195 , n32735 );
and ( n73197 , n32755 , n57872 );
or ( n73198 , n73196 , n73197 );
and ( n73199 , n73198 , n34150 );
or ( n73200 , n73194 , n73199 );
and ( n73201 , n73200 , n33381 );
not ( n73202 , n57880 );
not ( n73203 , n57872 );
and ( n73204 , n73203 , n32735 );
and ( n73205 , n35083 , n57872 );
or ( n73206 , n73204 , n73205 );
and ( n73207 , n73202 , n73206 );
and ( n73208 , n35083 , n57880 );
or ( n73209 , n73207 , n73208 );
and ( n73210 , n73209 , n33375 );
not ( n73211 , n32968 );
not ( n73212 , n57880 );
not ( n73213 , n57872 );
and ( n73214 , n73213 , n32735 );
and ( n73215 , n35083 , n57872 );
or ( n73216 , n73214 , n73215 );
and ( n73217 , n73212 , n73216 );
and ( n73218 , n35083 , n57880 );
or ( n73219 , n73217 , n73218 );
and ( n73220 , n73211 , n73219 );
not ( n73221 , n57900 );
not ( n73222 , n57902 );
and ( n73223 , n73222 , n73219 );
and ( n73224 , n35107 , n57902 );
or ( n73225 , n73223 , n73224 );
and ( n73226 , n73221 , n73225 );
and ( n73227 , n35115 , n57900 );
or ( n73228 , n73226 , n73227 );
and ( n73229 , n73228 , n32968 );
or ( n73230 , n73220 , n73229 );
and ( n73231 , n73230 , n33370 );
and ( n73232 , n32735 , n35062 );
or ( n73233 , C0 , n73201 , n73210 , n73231 , n73232 );
buf ( n73234 , n73233 );
buf ( n73235 , n73234 );
buf ( n73236 , n31655 );
buf ( n73237 , n30987 );
buf ( n73238 , n30987 );
buf ( n73239 , n31655 );
xor ( n73240 , n46237 , n49997 );
and ( n73241 , n73240 , n32431 );
not ( n73242 , n50002 );
and ( n73243 , n73242 , n46237 );
and ( n73244 , n40486 , n50002 );
or ( n73245 , n73243 , n73244 );
and ( n73246 , n73245 , n32419 );
not ( n73247 , n50008 );
and ( n73248 , n73247 , n46237 );
not ( n73249 , n47910 );
and ( n73250 , n73249 , n60901 );
and ( n73251 , n69313 , n47910 );
or ( n73252 , n73250 , n73251 );
and ( n73253 , n73252 , n50008 );
or ( n73254 , n73248 , n73253 );
and ( n73255 , n73254 , n32415 );
not ( n73256 , n50067 );
and ( n73257 , n73256 , n46237 );
and ( n73258 , n31896 , n47357 );
and ( n73259 , n31898 , n47359 );
and ( n73260 , n31900 , n47361 );
and ( n73261 , n31902 , n47363 );
and ( n73262 , n31904 , n47365 );
and ( n73263 , n31906 , n47367 );
and ( n73264 , n31908 , n47369 );
and ( n73265 , n31910 , n47371 );
and ( n73266 , n31912 , n47373 );
and ( n73267 , n31914 , n47375 );
and ( n73268 , n31916 , n47377 );
and ( n73269 , n31918 , n47379 );
and ( n73270 , n31920 , n47381 );
and ( n73271 , n31922 , n47383 );
and ( n73272 , n31924 , n47385 );
and ( n73273 , n31926 , n47387 );
or ( n73274 , n73258 , n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , n73271 , n73272 , n73273 );
and ( n73275 , n73274 , n50067 );
or ( n73276 , n73257 , n73275 );
and ( n73277 , n73276 , n32411 );
and ( n73278 , n46237 , n50098 );
or ( n73279 , n73241 , n73246 , n73255 , n73277 , n73278 );
and ( n73280 , n73279 , n32456 );
and ( n73281 , n46237 , n47409 );
or ( n73282 , C0 , n73280 , n73281 );
buf ( n73283 , n73282 );
buf ( n73284 , n73283 );
buf ( n73285 , n31655 );
not ( n73286 , n46356 );
and ( n73287 , n73286 , n31258 );
not ( n73288 , n50109 );
and ( n73289 , n73288 , n31258 );
and ( n73290 , n31272 , n50109 );
or ( n73291 , n73289 , n73290 );
and ( n73292 , n73291 , n46356 );
or ( n73293 , n73287 , n73292 );
and ( n73294 , n73293 , n31649 );
not ( n73295 , n50117 );
not ( n73296 , n50109 );
and ( n73297 , n73296 , n31258 );
and ( n73298 , n49443 , n50109 );
or ( n73299 , n73297 , n73298 );
and ( n73300 , n73295 , n73299 );
and ( n73301 , n49443 , n50117 );
or ( n73302 , n73300 , n73301 );
and ( n73303 , n73302 , n31643 );
not ( n73304 , n31452 );
not ( n73305 , n50117 );
not ( n73306 , n50109 );
and ( n73307 , n73306 , n31258 );
and ( n73308 , n49443 , n50109 );
or ( n73309 , n73307 , n73308 );
and ( n73310 , n73305 , n73309 );
and ( n73311 , n49443 , n50117 );
or ( n73312 , n73310 , n73311 );
and ( n73313 , n73304 , n73312 );
not ( n73314 , n50142 );
not ( n73315 , n50144 );
and ( n73316 , n73315 , n73312 );
and ( n73317 , n49469 , n50144 );
or ( n73318 , n73316 , n73317 );
and ( n73319 , n73314 , n73318 );
and ( n73320 , n49477 , n50142 );
or ( n73321 , n73319 , n73320 );
and ( n73322 , n73321 , n31452 );
or ( n73323 , n73313 , n73322 );
and ( n73324 , n73323 , n31638 );
and ( n73325 , n31258 , n47277 );
or ( n73326 , C0 , n73294 , n73303 , n73324 , n73325 );
buf ( n73327 , n73326 );
buf ( n73328 , n73327 );
not ( n73329 , n34150 );
and ( n73330 , n73329 , n32787 );
not ( n73331 , n56239 );
and ( n73332 , n73331 , n32787 );
and ( n73333 , n32789 , n56239 );
or ( n73334 , n73332 , n73333 );
and ( n73335 , n73334 , n34150 );
or ( n73336 , n73330 , n73335 );
and ( n73337 , n73336 , n33381 );
not ( n73338 , n56247 );
not ( n73339 , n56239 );
and ( n73340 , n73339 , n32787 );
and ( n73341 , n34301 , n56239 );
or ( n73342 , n73340 , n73341 );
and ( n73343 , n73338 , n73342 );
and ( n73344 , n34301 , n56247 );
or ( n73345 , n73343 , n73344 );
and ( n73346 , n73345 , n33375 );
not ( n73347 , n32968 );
not ( n73348 , n56247 );
not ( n73349 , n56239 );
and ( n73350 , n73349 , n32787 );
and ( n73351 , n34301 , n56239 );
or ( n73352 , n73350 , n73351 );
and ( n73353 , n73348 , n73352 );
and ( n73354 , n34301 , n56247 );
or ( n73355 , n73353 , n73354 );
and ( n73356 , n73347 , n73355 );
not ( n73357 , n56267 );
not ( n73358 , n56269 );
and ( n73359 , n73358 , n73355 );
and ( n73360 , n34761 , n56269 );
or ( n73361 , n73359 , n73360 );
and ( n73362 , n73357 , n73361 );
and ( n73363 , n35050 , n56267 );
or ( n73364 , n73362 , n73363 );
and ( n73365 , n73364 , n32968 );
or ( n73366 , n73356 , n73365 );
and ( n73367 , n73366 , n33370 );
and ( n73368 , n32787 , n35062 );
or ( n73369 , C0 , n73337 , n73346 , n73367 , n73368 );
buf ( n73370 , n73369 );
buf ( n73371 , n73370 );
buf ( n73372 , n30987 );
buf ( n73373 , n31655 );
buf ( n73374 , n31655 );
buf ( n73375 , n30987 );
not ( n73376 , n34150 );
and ( n73377 , n73376 , n32745 );
not ( n73378 , n56192 );
and ( n73379 , n73378 , n32745 );
and ( n73380 , n32755 , n56192 );
or ( n73381 , n73379 , n73380 );
and ( n73382 , n73381 , n34150 );
or ( n73383 , n73377 , n73382 );
and ( n73384 , n73383 , n33381 );
not ( n73385 , n56200 );
not ( n73386 , n56192 );
and ( n73387 , n73386 , n32745 );
and ( n73388 , n35083 , n56192 );
or ( n73389 , n73387 , n73388 );
and ( n73390 , n73385 , n73389 );
and ( n73391 , n35083 , n56200 );
or ( n73392 , n73390 , n73391 );
and ( n73393 , n73392 , n33375 );
not ( n73394 , n32968 );
not ( n73395 , n56200 );
not ( n73396 , n56192 );
and ( n73397 , n73396 , n32745 );
and ( n73398 , n35083 , n56192 );
or ( n73399 , n73397 , n73398 );
and ( n73400 , n73395 , n73399 );
and ( n73401 , n35083 , n56200 );
or ( n73402 , n73400 , n73401 );
and ( n73403 , n73394 , n73402 );
not ( n73404 , n56220 );
not ( n73405 , n56222 );
and ( n73406 , n73405 , n73402 );
and ( n73407 , n35107 , n56222 );
or ( n73408 , n73406 , n73407 );
and ( n73409 , n73404 , n73408 );
and ( n73410 , n35115 , n56220 );
or ( n73411 , n73409 , n73410 );
and ( n73412 , n73411 , n32968 );
or ( n73413 , n73403 , n73412 );
and ( n73414 , n73413 , n33370 );
and ( n73415 , n32745 , n35062 );
or ( n73416 , C0 , n73384 , n73393 , n73414 , n73415 );
buf ( n73417 , n73416 );
buf ( n73418 , n73417 );
buf ( n73419 , n31655 );
not ( n73420 , n38443 );
and ( n73421 , n73420 , n38286 );
xor ( n73422 , n53465 , n53504 );
and ( n73423 , n73422 , n38443 );
or ( n73424 , n73421 , n73423 );
and ( n73425 , n73424 , n38450 );
not ( n73426 , n39339 );
and ( n73427 , n73426 , n39186 );
xor ( n73428 , n53521 , n53560 );
and ( n73429 , n73428 , n39339 );
or ( n73430 , n73427 , n73429 );
and ( n73431 , n73430 , n39346 );
and ( n73432 , n40219 , n39359 );
or ( n73433 , n73425 , n73431 , n73432 );
buf ( n73434 , n73433 );
buf ( n73435 , n73434 );
and ( n73436 , n57515 , n48455 );
not ( n73437 , n48457 );
and ( n73438 , n73437 , n52402 );
and ( n73439 , n57515 , n48457 );
or ( n73440 , n73438 , n73439 );
and ( n73441 , n73440 , n31373 );
not ( n73442 , n44807 );
and ( n73443 , n73442 , n52402 );
and ( n73444 , n57515 , n44807 );
or ( n73445 , n73443 , n73444 );
and ( n73446 , n73445 , n31408 );
not ( n73447 , n48468 );
and ( n73448 , n73447 , n52402 );
and ( n73449 , n57515 , n48468 );
or ( n73450 , n73448 , n73449 );
and ( n73451 , n73450 , n31468 );
not ( n73452 , n44817 );
and ( n73453 , n73452 , n52402 );
and ( n73454 , n57515 , n44817 );
or ( n73455 , n73453 , n73454 );
and ( n73456 , n73455 , n31521 );
not ( n73457 , n39979 );
and ( n73458 , n73457 , n52402 );
and ( n73459 , n57503 , n39979 );
or ( n73460 , n73458 , n73459 );
and ( n73461 , n73460 , n31538 );
not ( n73462 , n45059 );
and ( n73463 , n73462 , n52402 );
and ( n73464 , n57503 , n45059 );
or ( n73465 , n73463 , n73464 );
and ( n73466 , n73465 , n31536 );
not ( n73467 , n33419 );
and ( n73468 , n73467 , n52402 );
xor ( n73469 , n57503 , n57504 );
and ( n73470 , n73469 , n33419 );
or ( n73471 , n73468 , n73470 );
and ( n73472 , n73471 , n31529 );
not ( n73473 , n33734 );
and ( n73474 , n73473 , n52402 );
not ( n73475 , n33533 );
xor ( n73476 , n57515 , n57516 );
and ( n73477 , n73475 , n73476 );
xnor ( n73478 , n57526 , n57527 );
and ( n73479 , n73478 , n33533 );
or ( n73480 , n73477 , n73479 );
and ( n73481 , n73480 , n33734 );
or ( n73482 , n73474 , n73481 );
and ( n73483 , n73482 , n31527 );
and ( n73484 , n57526 , n48513 );
or ( n73485 , n73436 , n73441 , n73446 , n73451 , n73456 , n73461 , n73466 , n73472 , n73483 , n73484 );
and ( n73486 , n73485 , n31557 );
and ( n73487 , n35390 , n33973 );
and ( n73488 , n52402 , n48524 );
or ( n73489 , C0 , n73486 , n73487 , n73488 );
buf ( n73490 , n73489 );
buf ( n73491 , n73490 );
buf ( n73492 , n30987 );
not ( n73493 , n33419 );
and ( n73494 , n73493 , n30989 );
xor ( n73495 , n33592 , n33609 );
xor ( n73496 , n73495 , n33673 );
and ( n73497 , n73496 , n33419 );
or ( n73498 , n73494 , n73497 );
and ( n73499 , n73498 , n31529 );
not ( n73500 , n33734 );
and ( n73501 , n73500 , n30989 );
not ( n73502 , n33533 );
xor ( n73503 , n33779 , n33609 );
xor ( n73504 , n73503 , n33791 );
and ( n73505 , n73502 , n73504 );
xor ( n73506 , n33872 , n33874 );
xor ( n73507 , n73506 , n33893 );
and ( n73508 , n73507 , n33533 );
or ( n73509 , n73505 , n73508 );
and ( n73510 , n73509 , n33734 );
or ( n73511 , n73501 , n73510 );
and ( n73512 , n73511 , n31527 );
and ( n73513 , n30989 , n33942 );
or ( n73514 , n73499 , n73512 , n73513 );
and ( n73515 , n73514 , n31557 );
and ( n73516 , n31621 , n31643 );
not ( n73517 , n31452 );
and ( n73518 , n73517 , n31621 );
xor ( n73519 , n30989 , n31588 );
and ( n73520 , n73519 , n31452 );
or ( n73521 , n73518 , n73520 );
and ( n73522 , n73521 , n31638 );
and ( n73523 , n31079 , n33973 );
and ( n73524 , n30989 , n33978 );
or ( n73525 , C0 , n73515 , n73516 , n73522 , n73523 , n73524 );
buf ( n73526 , n73525 );
buf ( n73527 , n73526 );
not ( n73528 , n40163 );
and ( n73529 , n73528 , n31665 );
and ( n73530 , n40188 , n40163 );
or ( n73531 , n73529 , n73530 );
and ( n73532 , n73531 , n32498 );
not ( n73533 , n55780 );
not ( n73534 , n55558 );
and ( n73535 , n73534 , n31665 );
buf ( n73536 , n73535 );
and ( n73537 , n73533 , n73536 );
buf ( n73538 , n73537 );
and ( n73539 , n73538 , n32496 );
and ( n73540 , n40430 , n32473 );
not ( n73541 , n32475 );
and ( n73542 , n73541 , n40430 );
xor ( n73543 , n40435 , n55791 );
not ( n73544 , n73543 );
buf ( n73545 , n73544 );
not ( n73546 , n73545 );
and ( n73547 , n73546 , n32475 );
or ( n73548 , n73542 , n73547 );
and ( n73549 , n73548 , n32486 );
and ( n73550 , n31665 , n55800 );
or ( n73551 , C0 , n73532 , n73539 , n73540 , n73549 , n73550 );
buf ( n73552 , n73551 );
buf ( n73553 , n73552 );
buf ( n73554 , n30987 );
not ( n73555 , n35542 );
and ( n73556 , n73555 , n41856 );
and ( n73557 , n67452 , n35542 );
or ( n73558 , n73556 , n73557 );
buf ( n73559 , n73558 );
buf ( n73560 , n73559 );
buf ( n73561 , n30987 );
buf ( n73562 , n31655 );
buf ( n73563 , n30987 );
not ( n73564 , n36587 );
and ( n73565 , n73564 , n36515 );
xor ( n73566 , n61941 , n61944 );
and ( n73567 , n73566 , n36587 );
or ( n73568 , n73565 , n73567 );
and ( n73569 , n73568 , n36596 );
not ( n73570 , n37485 );
and ( n73571 , n73570 , n37417 );
xor ( n73572 , n61957 , n61960 );
and ( n73573 , n73572 , n37485 );
or ( n73574 , n73571 , n73573 );
and ( n73575 , n73574 , n37494 );
and ( n73576 , n41864 , n37506 );
or ( n73577 , n73569 , n73575 , n73576 );
buf ( n73578 , n73577 );
buf ( n73579 , n73578 );
buf ( n73580 , n31655 );
and ( n73581 , n47657 , n50275 );
not ( n73582 , n50278 );
and ( n73583 , n73582 , n47570 );
and ( n73584 , n47657 , n50278 );
or ( n73585 , n73583 , n73584 );
and ( n73586 , n73585 , n32421 );
not ( n73587 , n50002 );
and ( n73588 , n73587 , n47570 );
and ( n73589 , n47657 , n50002 );
or ( n73590 , n73588 , n73589 );
and ( n73591 , n73590 , n32419 );
not ( n73592 , n50289 );
and ( n73593 , n73592 , n47570 );
and ( n73594 , n47657 , n50289 );
or ( n73595 , n73593 , n73594 );
and ( n73596 , n73595 , n32417 );
not ( n73597 , n50008 );
and ( n73598 , n73597 , n47570 );
and ( n73599 , n47657 , n50008 );
or ( n73600 , n73598 , n73599 );
and ( n73601 , n73600 , n32415 );
not ( n73602 , n47331 );
and ( n73603 , n73602 , n47570 );
and ( n73604 , n47602 , n47331 );
or ( n73605 , n73603 , n73604 );
and ( n73606 , n73605 , n32413 );
not ( n73607 , n50067 );
and ( n73608 , n73607 , n47570 );
and ( n73609 , n47602 , n50067 );
or ( n73610 , n73608 , n73609 );
and ( n73611 , n73610 , n32411 );
not ( n73612 , n31728 );
and ( n73613 , n73612 , n47570 );
and ( n73614 , n52083 , n31728 );
or ( n73615 , n73613 , n73614 );
and ( n73616 , n73615 , n32253 );
not ( n73617 , n32283 );
and ( n73618 , n73617 , n47570 );
and ( n73619 , n52094 , n32283 );
or ( n73620 , n73618 , n73619 );
and ( n73621 , n73620 , n32398 );
and ( n73622 , n47707 , n50334 );
or ( n73623 , n73581 , n73586 , n73591 , n73596 , n73601 , n73606 , n73611 , n73616 , n73621 , n73622 );
and ( n73624 , n73623 , n32456 );
and ( n73625 , n37547 , n32489 );
and ( n73626 , n47570 , n50345 );
or ( n73627 , C0 , n73624 , n73625 , n73626 );
buf ( n73628 , n73627 );
buf ( n73629 , n73628 );
buf ( n73630 , n31655 );
buf ( n73631 , n31655 );
buf ( n73632 , n30987 );
not ( n73633 , n35542 );
and ( n73634 , n73633 , n41862 );
buf ( n73635 , RI15b45b40_243);
and ( n73636 , n73635 , n35542 );
or ( n73637 , n73634 , n73636 );
buf ( n73638 , n73637 );
buf ( n73639 , n73638 );
not ( n73640 , n34150 );
and ( n73641 , n73640 , n32809 );
not ( n73642 , n56836 );
and ( n73643 , n73642 , n32809 );
and ( n73644 , n32823 , n56836 );
or ( n73645 , n73643 , n73644 );
and ( n73646 , n73645 , n34150 );
or ( n73647 , n73641 , n73646 );
and ( n73648 , n73647 , n33381 );
not ( n73649 , n56844 );
not ( n73650 , n56836 );
and ( n73651 , n73650 , n32809 );
and ( n73652 , n41464 , n56836 );
or ( n73653 , n73651 , n73652 );
and ( n73654 , n73649 , n73653 );
and ( n73655 , n41464 , n56844 );
or ( n73656 , n73654 , n73655 );
and ( n73657 , n73656 , n33375 );
not ( n73658 , n32968 );
not ( n73659 , n56844 );
not ( n73660 , n56836 );
and ( n73661 , n73660 , n32809 );
and ( n73662 , n41464 , n56836 );
or ( n73663 , n73661 , n73662 );
and ( n73664 , n73659 , n73663 );
and ( n73665 , n41464 , n56844 );
or ( n73666 , n73664 , n73665 );
and ( n73667 , n73658 , n73666 );
not ( n73668 , n56864 );
not ( n73669 , n56866 );
and ( n73670 , n73669 , n73666 );
and ( n73671 , n41490 , n56866 );
or ( n73672 , n73670 , n73671 );
and ( n73673 , n73668 , n73672 );
and ( n73674 , n41500 , n56864 );
or ( n73675 , n73673 , n73674 );
and ( n73676 , n73675 , n32968 );
or ( n73677 , n73667 , n73676 );
and ( n73678 , n73677 , n33370 );
and ( n73679 , n32809 , n35062 );
or ( n73680 , C0 , n73648 , n73657 , n73678 , n73679 );
buf ( n73681 , n73680 );
buf ( n73682 , n73681 );
buf ( n73683 , n30987 );
buf ( n73684 , n31655 );
buf ( n73685 , RI15b48138_324);
and ( n73686 , n73685 , n58207 );
and ( n73687 , n54736 , n44695 );
or ( n73688 , n73686 , n73687 );
buf ( n73689 , n73688 );
buf ( n73690 , n73689 );
buf ( n73691 , n31655 );
buf ( n73692 , n30987 );
buf ( n73693 , n30987 );
buf ( n73694 , n30987 );
not ( n73695 , n46356 );
and ( n73696 , n73695 , n31309 );
not ( n73697 , n47831 );
and ( n73698 , n73697 , n31309 );
and ( n73699 , n31339 , n47831 );
or ( n73700 , n73698 , n73699 );
and ( n73701 , n73700 , n46356 );
or ( n73702 , n73696 , n73701 );
and ( n73703 , n73702 , n31649 );
not ( n73704 , n47839 );
not ( n73705 , n47831 );
and ( n73706 , n73705 , n31309 );
and ( n73707 , n47449 , n47831 );
or ( n73708 , n73706 , n73707 );
and ( n73709 , n73704 , n73708 );
and ( n73710 , n47449 , n47839 );
or ( n73711 , n73709 , n73710 );
and ( n73712 , n73711 , n31643 );
not ( n73713 , n31452 );
not ( n73714 , n47839 );
not ( n73715 , n47831 );
and ( n73716 , n73715 , n31309 );
and ( n73717 , n47449 , n47831 );
or ( n73718 , n73716 , n73717 );
and ( n73719 , n73714 , n73718 );
and ( n73720 , n47449 , n47839 );
or ( n73721 , n73719 , n73720 );
and ( n73722 , n73713 , n73721 );
not ( n73723 , n47866 );
not ( n73724 , n47868 );
and ( n73725 , n73724 , n73721 );
and ( n73726 , n47485 , n47868 );
or ( n73727 , n73725 , n73726 );
and ( n73728 , n73723 , n73727 );
and ( n73729 , n47503 , n47866 );
or ( n73730 , n73728 , n73729 );
and ( n73731 , n73730 , n31452 );
or ( n73732 , n73722 , n73731 );
and ( n73733 , n73732 , n31638 );
and ( n73734 , n31309 , n47277 );
or ( n73735 , C0 , n73703 , n73712 , n73733 , n73734 );
buf ( n73736 , n73735 );
buf ( n73737 , n73736 );
buf ( n73738 , n31655 );
not ( n73739 , n35278 );
buf ( n73740 , RI15b5f400_1115);
and ( n73741 , n73739 , n73740 );
not ( n73742 , n46290 );
and ( n73743 , n73742 , n46195 );
xor ( n73744 , n46298 , n46314 );
and ( n73745 , n73744 , n46290 );
or ( n73746 , n73743 , n73745 );
and ( n73747 , n73746 , n35278 );
or ( n73748 , n73741 , n73747 );
and ( n73749 , n73748 , n32417 );
not ( n73750 , n47912 );
and ( n73751 , n73750 , n73740 );
not ( n73752 , n48101 );
and ( n73753 , n73752 , n48013 );
xor ( n73754 , n50022 , n50023 );
and ( n73755 , n73754 , n48101 );
or ( n73756 , n73753 , n73755 );
and ( n73757 , n73756 , n47912 );
or ( n73758 , n73751 , n73757 );
and ( n73759 , n73758 , n32415 );
and ( n73760 , n73740 , n48133 );
or ( n73761 , n73749 , n73759 , n73760 );
and ( n73762 , n73761 , n32456 );
and ( n73763 , n73740 , n47409 );
or ( n73764 , C0 , n73762 , n73763 );
buf ( n73765 , n73764 );
buf ( n73766 , n73765 );
buf ( n73767 , n30987 );
buf ( n73768 , RI15b46b30_277);
and ( n73769 , n73768 , n33377 );
not ( n73770 , n48545 );
and ( n73771 , n73770 , n72970 );
not ( n73772 , n39572 );
and ( n73773 , n73772 , n39477 );
xor ( n73774 , n42620 , n42633 );
and ( n73775 , n73774 , n39572 );
or ( n73776 , n73773 , n73775 );
and ( n73777 , n73776 , n48545 );
or ( n73778 , n73771 , n73777 );
and ( n73779 , n73778 , n32890 );
not ( n73780 , n48557 );
and ( n73781 , n73780 , n72970 );
and ( n73782 , n73776 , n48557 );
or ( n73783 , n73781 , n73782 );
and ( n73784 , n73783 , n33038 );
and ( n73785 , n72970 , n48571 );
or ( n73786 , n73779 , n73784 , n73785 );
and ( n73787 , n73786 , n33208 );
and ( n73788 , n72970 , n48577 );
or ( n73789 , C0 , n73769 , n73787 , n73788 );
buf ( n73790 , n73789 );
buf ( n73791 , n73790 );
buf ( n73792 , n31655 );
buf ( n73793 , n31655 );
buf ( n73794 , n30987 );
buf ( n73795 , n30987 );
buf ( n73796 , n30987 );
buf ( n73797 , n31655 );
buf ( n73798 , RI15b46608_266);
and ( n73799 , n73798 , n33377 );
not ( n73800 , n48545 );
and ( n73801 , n73800 , n65013 );
buf ( n73802 , n73801 );
and ( n73803 , n73802 , n32890 );
not ( n73804 , n48557 );
and ( n73805 , n73804 , n65013 );
not ( n73806 , n54581 );
and ( n73807 , n73806 , n54543 );
xor ( n73808 , n54543 , n54340 );
and ( n73809 , n70664 , n70665 );
xor ( n73810 , n73808 , n73809 );
and ( n73811 , n73810 , n54581 );
or ( n73812 , n73807 , n73811 );
and ( n73813 , n73812 , n48557 );
or ( n73814 , n73805 , n73813 );
and ( n73815 , n73814 , n33038 );
and ( n73816 , n65013 , n48571 );
or ( n73817 , n73803 , n73815 , n73816 );
and ( n73818 , n73817 , n33208 );
and ( n73819 , n65013 , n48577 );
or ( n73820 , C0 , n73799 , n73818 , n73819 );
buf ( n73821 , n73820 );
buf ( n73822 , n73821 );
buf ( n73823 , n31655 );
buf ( n73824 , n30987 );
buf ( n73825 , n31655 );
not ( n73826 , n31728 );
and ( n73827 , n73826 , n32464 );
xor ( n73828 , n32000 , n32033 );
xor ( n73829 , n73828 , n32069 );
and ( n73830 , n73829 , n31728 );
or ( n73831 , n73827 , n73830 );
and ( n73832 , n73831 , n32253 );
not ( n73833 , n32283 );
and ( n73834 , n73833 , n32464 );
not ( n73835 , n31823 );
xor ( n73836 , n32306 , n32033 );
xor ( n73837 , n73836 , n32308 );
and ( n73838 , n73835 , n73837 );
xor ( n73839 , n32364 , n32366 );
xor ( n73840 , n73839 , n32371 );
and ( n73841 , n73840 , n31823 );
or ( n73842 , n73838 , n73841 );
and ( n73843 , n73842 , n32283 );
or ( n73844 , n73834 , n73843 );
and ( n73845 , n73844 , n32398 );
and ( n73846 , n32464 , n32436 );
or ( n73847 , n73832 , n73845 , n73846 );
and ( n73848 , n73847 , n32456 );
and ( n73849 , n46065 , n32473 );
not ( n73850 , n32475 );
and ( n73851 , n73850 , n46065 );
and ( n73852 , n32464 , n32475 );
or ( n73853 , n73851 , n73852 );
and ( n73854 , n73853 , n32486 );
and ( n73855 , n37514 , n32489 );
and ( n73856 , n32464 , n32501 );
or ( n73857 , C0 , n73848 , n73849 , n73854 , n73855 , n73856 );
buf ( n73858 , n73857 );
buf ( n73859 , n73858 );
buf ( n73860 , n31655 );
buf ( n73861 , n30987 );
not ( n73862 , n46356 );
and ( n73863 , n73862 , n31009 );
buf ( n73864 , n73863 );
and ( n73865 , n73864 , n31649 );
not ( n73866 , n52614 );
not ( n73867 , n44702 );
and ( n73868 , n73867 , n31009 );
buf ( n73869 , n73868 );
and ( n73870 , n73866 , n73869 );
buf ( n73871 , n73870 );
and ( n73872 , n73871 , n31647 );
and ( n73873 , n31009 , n52626 );
or ( n73874 , C0 , n73865 , n73872 , C0 , C0 , n73873 );
buf ( n73875 , n73874 );
buf ( n73876 , n73875 );
not ( n73877 , n48765 );
and ( n73878 , n73877 , n33236 );
xor ( n73879 , n48866 , n48883 );
xor ( n73880 , n73879 , n48991 );
and ( n73881 , n73880 , n48765 );
or ( n73882 , n73878 , n73881 );
and ( n73883 , n73882 , n33180 );
not ( n73884 , n49054 );
and ( n73885 , n73884 , n33236 );
not ( n73886 , n48845 );
xor ( n73887 , n49083 , n48883 );
xor ( n73888 , n73887 , n49105 );
and ( n73889 , n73886 , n73888 );
xor ( n73890 , n49196 , n49198 );
xor ( n73891 , n73890 , n49231 );
and ( n73892 , n73891 , n48845 );
or ( n73893 , n73889 , n73892 );
and ( n73894 , n73893 , n49054 );
or ( n73895 , n73885 , n73894 );
and ( n73896 , n73895 , n33178 );
and ( n73897 , n33236 , n49774 );
or ( n73898 , n73883 , n73896 , n73897 );
and ( n73899 , n73898 , n33208 );
and ( n73900 , n33323 , n33375 );
not ( n73901 , n32968 );
and ( n73902 , n73901 , n33323 );
xor ( n73903 , n33236 , n49782 );
and ( n73904 , n73903 , n32968 );
or ( n73905 , n73902 , n73904 );
and ( n73906 , n73905 , n33370 );
and ( n73907 , n32999 , n35056 );
and ( n73908 , n33236 , n49794 );
or ( n73909 , C0 , n73899 , n73900 , n73906 , n73907 , n73908 );
buf ( n73910 , n73909 );
buf ( n73911 , n73910 );
buf ( n73912 , n31655 );
buf ( n73913 , n30987 );
not ( n73914 , n50828 );
not ( n73915 , n50834 );
and ( n73916 , n73915 , n40249 );
and ( n73917 , n68204 , n50834 );
or ( n73918 , n73916 , n73917 );
and ( n73919 , n73914 , n73918 );
and ( n73920 , n60218 , n50828 );
or ( n73921 , n73919 , n73920 );
buf ( n73922 , n73921 );
buf ( n73923 , n73922 );
buf ( n73924 , n30987 );
buf ( n73925 , n31655 );
buf ( n73926 , n31655 );
buf ( n73927 , n30987 );
not ( n73928 , n32953 );
and ( n73929 , n73928 , n73798 );
and ( n73930 , n73812 , n32953 );
or ( n73931 , n73929 , n73930 );
and ( n73932 , n73931 , n33038 );
not ( n73933 , n48660 );
and ( n73934 , n73933 , n73798 );
not ( n73935 , n55168 );
and ( n73936 , n73935 , n55140 );
xor ( n73937 , n55140 , n34193 );
and ( n73938 , n70676 , n70677 );
xor ( n73939 , n73937 , n73938 );
and ( n73940 , n73939 , n55168 );
or ( n73941 , n73936 , n73940 );
and ( n73942 , n73941 , n48660 );
or ( n73943 , n73934 , n73942 );
and ( n73944 , n73943 , n33172 );
and ( n73945 , n73798 , n39795 );
or ( n73946 , n73932 , n73944 , n73945 );
and ( n73947 , n73946 , n33208 );
and ( n73948 , n73798 , n39805 );
or ( n73949 , C0 , n73947 , n73948 );
buf ( n73950 , n73949 );
buf ( n73951 , n73950 );
buf ( n73952 , n30987 );
buf ( n73953 , n31655 );
buf ( n73954 , n30987 );
and ( n73955 , n49059 , n48639 );
not ( n73956 , n48642 );
and ( n73957 , n73956 , n48584 );
and ( n73958 , n49059 , n48642 );
or ( n73959 , n73957 , n73958 );
and ( n73960 , n73959 , n32890 );
not ( n73961 , n48648 );
and ( n73962 , n73961 , n48584 );
and ( n73963 , n49059 , n48648 );
or ( n73964 , n73962 , n73963 );
and ( n73965 , n73964 , n32924 );
not ( n73966 , n48654 );
and ( n73967 , n73966 , n48584 );
and ( n73968 , n49059 , n48654 );
or ( n73969 , n73967 , n73968 );
and ( n73970 , n73969 , n33038 );
not ( n73971 , n48660 );
and ( n73972 , n73971 , n48584 );
and ( n73973 , n49059 , n48660 );
or ( n73974 , n73972 , n73973 );
and ( n73975 , n73974 , n33172 );
not ( n73976 , n41576 );
and ( n73977 , n73976 , n48584 );
and ( n73978 , n48769 , n41576 );
or ( n73979 , n73977 , n73978 );
and ( n73980 , n73979 , n33189 );
not ( n73981 , n48730 );
and ( n73982 , n73981 , n48584 );
and ( n73983 , n48769 , n48730 );
or ( n73984 , n73982 , n73983 );
and ( n73985 , n73984 , n33187 );
not ( n73986 , n48765 );
and ( n73987 , n73986 , n48584 );
xor ( n73988 , n48769 , n49019 );
and ( n73989 , n73988 , n48765 );
or ( n73990 , n73987 , n73989 );
and ( n73991 , n73990 , n33180 );
not ( n73992 , n49054 );
and ( n73993 , n73992 , n48584 );
not ( n73994 , n48845 );
xor ( n73995 , n49059 , n49133 );
and ( n73996 , n73994 , n73995 );
xnor ( n73997 , n49168 , n49259 );
and ( n73998 , n73997 , n48845 );
or ( n73999 , n73996 , n73998 );
and ( n74000 , n73999 , n49054 );
or ( n74001 , n73993 , n74000 );
and ( n74002 , n74001 , n33178 );
and ( n74003 , n49168 , n49275 );
or ( n74004 , n73955 , n73960 , n73965 , n73970 , n73975 , n73980 , n73985 , n73991 , n74002 , n74003 );
and ( n74005 , n74004 , n33208 );
and ( n74006 , n32977 , n35056 );
and ( n74007 , n48584 , n49286 );
or ( n74008 , C0 , n74005 , n74006 , n74007 );
buf ( n74009 , n74008 );
buf ( n74010 , n74009 );
buf ( n74011 , n30987 );
buf ( n74012 , n31655 );
buf ( n74013 , n31655 );
buf ( n74014 , n31655 );
not ( n74015 , n33419 );
and ( n74016 , n74015 , n31568 );
and ( n74017 , n67838 , n33419 );
or ( n74018 , n74016 , n74017 );
and ( n74019 , n74018 , n31529 );
not ( n74020 , n33734 );
and ( n74021 , n74020 , n31568 );
and ( n74022 , n67849 , n33734 );
or ( n74023 , n74021 , n74022 );
and ( n74024 , n74023 , n31527 );
and ( n74025 , n31568 , n33942 );
or ( n74026 , n74019 , n74024 , n74025 );
and ( n74027 , n74026 , n31557 );
and ( n74028 , n35492 , n31643 );
not ( n74029 , n31452 );
and ( n74030 , n74029 , n35492 );
xor ( n74031 , n31568 , n42438 );
and ( n74032 , n74031 , n31452 );
or ( n74033 , n74030 , n74032 );
and ( n74034 , n74033 , n31638 );
and ( n74035 , n35394 , n33973 );
and ( n74036 , n31568 , n33978 );
or ( n74037 , C0 , n74027 , n74028 , n74034 , n74035 , n74036 );
buf ( n74038 , n74037 );
buf ( n74039 , n74038 );
buf ( n74040 , n30987 );
buf ( n74041 , n30987 );
and ( n74042 , n31576 , n31007 );
not ( n74043 , n31077 );
and ( n74044 , n74043 , n34000 );
buf ( n74045 , n74044 );
and ( n74046 , n74045 , n31373 );
not ( n74047 , n31402 );
and ( n74048 , n74047 , n34000 );
buf ( n74049 , n74048 );
and ( n74050 , n74049 , n31408 );
not ( n74051 , n31437 );
and ( n74052 , n74051 , n34000 );
not ( n74053 , n31455 );
and ( n74054 , n74053 , n34040 );
xor ( n74055 , n34000 , n34023 );
and ( n74056 , n74055 , n31455 );
or ( n74057 , n74054 , n74056 );
and ( n74058 , n74057 , n31437 );
or ( n74059 , n74052 , n74058 );
and ( n74060 , n74059 , n31468 );
not ( n74061 , n31497 );
and ( n74062 , n74061 , n34000 );
not ( n74063 , n31454 );
not ( n74064 , n31501 );
and ( n74065 , n74064 , n34040 );
xor ( n74066 , n34041 , n34075 );
and ( n74067 , n74066 , n31501 );
or ( n74068 , n74065 , n74067 );
and ( n74069 , n74063 , n74068 );
and ( n74070 , n74055 , n31454 );
or ( n74071 , n74069 , n74070 );
and ( n74072 , n74071 , n31497 );
or ( n74073 , n74062 , n74072 );
and ( n74074 , n74073 , n31521 );
and ( n74075 , n34000 , n31553 );
or ( n74076 , n74046 , n74050 , n74060 , n74074 , n74075 );
and ( n74077 , n74076 , n31557 );
not ( n74078 , n31452 );
not ( n74079 , n31619 );
and ( n74080 , n74079 , n34097 );
xor ( n74081 , n34098 , n34132 );
and ( n74082 , n74081 , n31619 );
or ( n74083 , n74080 , n74082 );
and ( n74084 , n74078 , n74083 );
and ( n74085 , n34000 , n31452 );
or ( n74086 , n74084 , n74085 );
and ( n74087 , n74086 , n31638 );
buf ( n74088 , n33973 );
and ( n74089 , n34000 , n31650 );
or ( n74090 , C0 , n74042 , n74077 , n74087 , n74088 , n74089 );
buf ( n74091 , n74090 );
buf ( n74092 , n74091 );
buf ( n74093 , n31655 );
buf ( n74094 , n30987 );
buf ( n74095 , n30987 );
buf ( n74096 , n31655 );
buf ( n74097 , n31655 );
not ( n74098 , n43755 );
and ( n74099 , n74098 , n43479 );
xor ( n74100 , n52314 , n52315 );
and ( n74101 , n74100 , n43755 );
or ( n74102 , n74099 , n74101 );
and ( n74103 , n74102 , n43774 );
not ( n74104 , n44663 );
and ( n74105 , n74104 , n44391 );
xor ( n74106 , n52352 , n52353 );
and ( n74107 , n74106 , n44663 );
or ( n74108 , n74105 , n74107 );
and ( n74109 , n74108 , n44682 );
buf ( n74110 , RI15b45690_233);
and ( n74111 , n74110 , n44695 );
or ( n74112 , n74103 , n74109 , n74111 );
buf ( n74113 , n74112 );
buf ( n74114 , n74113 );
buf ( n74115 , n30987 );
xor ( n74116 , n44764 , n44803 );
and ( n74117 , n74116 , n31548 );
not ( n74118 , n44807 );
and ( n74119 , n74118 , n44764 );
and ( n74120 , n46617 , n44807 );
or ( n74121 , n74119 , n74120 );
and ( n74122 , n74121 , n31408 );
not ( n74123 , n44817 );
and ( n74124 , n74123 , n44764 );
not ( n74125 , n44994 );
and ( n74126 , n74125 , n44966 );
xor ( n74127 , n44998 , n45022 );
and ( n74128 , n74127 , n44994 );
or ( n74129 , n74126 , n74128 );
and ( n74130 , n74129 , n44817 );
or ( n74131 , n74124 , n74130 );
and ( n74132 , n74131 , n31521 );
not ( n74133 , n45059 );
and ( n74134 , n74133 , n44764 );
xor ( n74135 , n45095 , n45134 );
and ( n74136 , n74135 , n45059 );
or ( n74137 , n74134 , n74136 );
and ( n74138 , n74137 , n31536 );
and ( n74139 , n44764 , n45148 );
or ( n74140 , n74117 , n74122 , n74132 , n74138 , n74139 );
and ( n74141 , n74140 , n31557 );
and ( n74142 , n44764 , n40154 );
or ( n74143 , C0 , n74141 , n74142 );
buf ( n74144 , n74143 );
buf ( n74145 , n74144 );
buf ( n74146 , n31655 );
not ( n74147 , n40163 );
and ( n74148 , n74147 , n31918 );
not ( n74149 , n45161 );
and ( n74150 , n74149 , n31918 );
and ( n74151 , n32200 , n45161 );
or ( n74152 , n74150 , n74151 );
and ( n74153 , n74152 , n40163 );
or ( n74154 , n74148 , n74153 );
and ( n74155 , n74154 , n32498 );
not ( n74156 , n45170 );
not ( n74157 , n45161 );
and ( n74158 , n74157 , n31918 );
and ( n74159 , n53243 , n45161 );
or ( n74160 , n74158 , n74159 );
and ( n74161 , n74156 , n74160 );
and ( n74162 , n53243 , n45170 );
or ( n74163 , n74161 , n74162 );
and ( n74164 , n74163 , n32473 );
not ( n74165 , n32475 );
not ( n74166 , n45170 );
not ( n74167 , n45161 );
and ( n74168 , n74167 , n31918 );
and ( n74169 , n53243 , n45161 );
or ( n74170 , n74168 , n74169 );
and ( n74171 , n74166 , n74170 );
and ( n74172 , n53243 , n45170 );
or ( n74173 , n74171 , n74172 );
and ( n74174 , n74165 , n74173 );
not ( n74175 , n45196 );
not ( n74176 , n45199 );
and ( n74177 , n74176 , n74173 );
and ( n74178 , n53269 , n45199 );
or ( n74179 , n74177 , n74178 );
and ( n74180 , n74175 , n74179 );
and ( n74181 , n53277 , n45196 );
or ( n74182 , n74180 , n74181 );
and ( n74183 , n74182 , n32475 );
or ( n74184 , n74174 , n74183 );
and ( n74185 , n74184 , n32486 );
and ( n74186 , n31918 , n41278 );
or ( n74187 , C0 , n74155 , n74164 , n74185 , n74186 );
buf ( n74188 , n74187 );
buf ( n74189 , n74188 );
buf ( n74190 , n30987 );
not ( n74191 , n50828 );
not ( n74192 , n50834 );
and ( n74193 , n74192 , n40505 );
buf ( n74194 , RI15b53790_713);
and ( n74195 , n74194 , n50834 );
or ( n74196 , n74193 , n74195 );
and ( n74197 , n74191 , n74196 );
buf ( n74198 , RI15b5fbf8_1132);
and ( n74199 , n74198 , n50828 );
or ( n74200 , n74197 , n74199 );
buf ( n74201 , n74200 );
buf ( n74202 , n74201 );
xor ( n74203 , n33075 , n58396 );
and ( n74204 , n74203 , n33201 );
not ( n74205 , n41576 );
and ( n74206 , n74205 , n33075 );
xor ( n74207 , n58472 , n58597 );
and ( n74208 , n74207 , n41576 );
or ( n74209 , n74206 , n74208 );
and ( n74210 , n74209 , n33189 );
and ( n74211 , n33075 , n41592 );
or ( n74212 , n74204 , n74210 , n74211 );
and ( n74213 , n74212 , n33208 );
and ( n74214 , n33075 , n39805 );
or ( n74215 , C0 , n74213 , n74214 );
buf ( n74216 , n74215 );
buf ( n74217 , n74216 );
buf ( n74218 , n30987 );
buf ( n74219 , n31655 );
buf ( n74220 , n31655 );
buf ( n74221 , n30987 );
buf ( n74222 , n30987 );
buf ( n74223 , n31655 );
buf ( n74224 , n31655 );
not ( n74225 , n50828 );
not ( n74226 , n50834 );
and ( n74227 , n74226 , n40569 );
buf ( n74228 , RI15b54078_732);
and ( n74229 , n74228 , n50834 );
or ( n74230 , n74227 , n74229 );
and ( n74231 , n74225 , n74230 );
and ( n74232 , n63558 , n50828 );
or ( n74233 , n74231 , n74232 );
buf ( n74234 , n74233 );
buf ( n74235 , n74234 );
buf ( n74236 , n30987 );
xor ( n74237 , n33113 , n52222 );
and ( n74238 , n74237 , n33201 );
not ( n74239 , n41576 );
and ( n74240 , n74239 , n33113 );
and ( n74241 , n32690 , n52252 );
and ( n74242 , n32692 , n52254 );
and ( n74243 , n32694 , n52256 );
and ( n74244 , n32696 , n52258 );
and ( n74245 , n32698 , n52260 );
and ( n74246 , n32700 , n52262 );
and ( n74247 , n32702 , n52264 );
and ( n74248 , n32704 , n52266 );
and ( n74249 , n32706 , n52268 );
and ( n74250 , n32708 , n52270 );
and ( n74251 , n32710 , n52272 );
and ( n74252 , n32712 , n52274 );
and ( n74253 , n32714 , n52276 );
and ( n74254 , n32716 , n52278 );
and ( n74255 , n32718 , n52280 );
and ( n74256 , n32720 , n52282 );
or ( n74257 , n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , n74255 , n74256 );
and ( n74258 , n74257 , n41576 );
or ( n74259 , n74240 , n74258 );
and ( n74260 , n74259 , n33189 );
and ( n74261 , n33113 , n41592 );
or ( n74262 , n74238 , n74260 , n74261 );
and ( n74263 , n74262 , n33208 );
and ( n74264 , n33113 , n39805 );
or ( n74265 , C0 , n74263 , n74264 );
buf ( n74266 , n74265 );
buf ( n74267 , n74266 );
not ( n74268 , n40163 );
and ( n74269 , n74268 , n32044 );
not ( n74270 , n54629 );
and ( n74271 , n74270 , n32044 );
and ( n74272 , n32130 , n54629 );
or ( n74273 , n74271 , n74272 );
and ( n74274 , n74273 , n40163 );
or ( n74275 , n74269 , n74274 );
and ( n74276 , n74275 , n32498 );
not ( n74277 , n54637 );
not ( n74278 , n54629 );
and ( n74279 , n74278 , n32044 );
and ( n74280 , n45833 , n54629 );
or ( n74281 , n74279 , n74280 );
and ( n74282 , n74277 , n74281 );
and ( n74283 , n45833 , n54637 );
or ( n74284 , n74282 , n74283 );
and ( n74285 , n74284 , n32473 );
not ( n74286 , n32475 );
not ( n74287 , n54637 );
not ( n74288 , n54629 );
and ( n74289 , n74288 , n32044 );
and ( n74290 , n45833 , n54629 );
or ( n74291 , n74289 , n74290 );
and ( n74292 , n74287 , n74291 );
and ( n74293 , n45833 , n54637 );
or ( n74294 , n74292 , n74293 );
and ( n74295 , n74286 , n74294 );
not ( n74296 , n54657 );
not ( n74297 , n54659 );
and ( n74298 , n74297 , n74294 );
and ( n74299 , n45857 , n54659 );
or ( n74300 , n74298 , n74299 );
and ( n74301 , n74296 , n74300 );
and ( n74302 , n45865 , n54657 );
or ( n74303 , n74301 , n74302 );
and ( n74304 , n74303 , n32475 );
or ( n74305 , n74295 , n74304 );
and ( n74306 , n74305 , n32486 );
and ( n74307 , n32044 , n41278 );
or ( n74308 , C0 , n74276 , n74285 , n74306 , n74307 );
buf ( n74309 , n74308 );
buf ( n74310 , n74309 );
buf ( n74311 , n31655 );
and ( n74312 , n53148 , n31645 );
not ( n74313 , n45274 );
and ( n74314 , n74313 , n55346 );
buf ( n74315 , n74314 );
and ( n74316 , n74315 , n31373 );
not ( n74317 , n45280 );
and ( n74318 , n74317 , n55346 );
and ( n74319 , n53154 , n45280 );
or ( n74320 , n74318 , n74319 );
and ( n74321 , n74320 , n31468 );
and ( n74322 , n55346 , n45802 );
or ( n74323 , n74316 , n74321 , n74322 );
and ( n74324 , n74323 , n31557 );
and ( n74325 , n55346 , n45808 );
or ( n74326 , C0 , n74312 , n74324 , n74325 );
buf ( n74327 , n74326 );
buf ( n74328 , n74327 );
buf ( n74329 , n30987 );
buf ( n74330 , n30987 );
buf ( n74331 , n31655 );
not ( n74332 , n32953 );
and ( n74333 , n74332 , n70129 );
not ( n74334 , n39572 );
and ( n74335 , n74334 , n39568 );
xor ( n74336 , n65461 , n65462 );
and ( n74337 , n74336 , n39572 );
or ( n74338 , n74335 , n74337 );
and ( n74339 , n74338 , n32953 );
or ( n74340 , n74333 , n74339 );
and ( n74341 , n74340 , n33038 );
not ( n74342 , n39586 );
and ( n74343 , n74342 , n70129 );
and ( n74344 , n70137 , n39586 );
or ( n74345 , n74343 , n74344 );
and ( n74346 , n74345 , n33172 );
and ( n74347 , n70129 , n39795 );
or ( n74348 , n74341 , n74346 , n74347 );
and ( n74349 , n74348 , n33208 );
and ( n74350 , n70129 , n39805 );
or ( n74351 , C0 , n74349 , n74350 );
buf ( n74352 , n74351 );
buf ( n74353 , n74352 );
buf ( n74354 , n31655 );
buf ( n74355 , n30987 );
buf ( n74356 , n30987 );
buf ( n74357 , n30987 );
buf ( n74358 , n31655 );
buf ( n74359 , n30987 );
not ( n74360 , n40163 );
and ( n74361 , n74360 , n31811 );
not ( n74362 , n57233 );
and ( n74363 , n74362 , n31811 );
and ( n74364 , n32252 , n57233 );
or ( n74365 , n74363 , n74364 );
and ( n74366 , n74365 , n40163 );
or ( n74367 , n74361 , n74366 );
and ( n74368 , n74367 , n32498 );
not ( n74369 , n57241 );
not ( n74370 , n57233 );
and ( n74371 , n74370 , n31811 );
and ( n74372 , n40393 , n57233 );
or ( n74373 , n74371 , n74372 );
and ( n74374 , n74369 , n74373 );
and ( n74375 , n40393 , n57241 );
or ( n74376 , n74374 , n74375 );
and ( n74377 , n74376 , n32473 );
not ( n74378 , n32475 );
not ( n74379 , n57241 );
not ( n74380 , n57233 );
and ( n74381 , n74380 , n31811 );
and ( n74382 , n40393 , n57233 );
or ( n74383 , n74381 , n74382 );
and ( n74384 , n74379 , n74383 );
and ( n74385 , n40393 , n57241 );
or ( n74386 , n74384 , n74385 );
and ( n74387 , n74378 , n74386 );
not ( n74388 , n57261 );
not ( n74389 , n57263 );
and ( n74390 , n74389 , n74386 );
and ( n74391 , n40972 , n57263 );
or ( n74392 , n74390 , n74391 );
and ( n74393 , n74388 , n74392 );
and ( n74394 , n41267 , n57261 );
or ( n74395 , n74393 , n74394 );
and ( n74396 , n74395 , n32475 );
or ( n74397 , n74387 , n74396 );
and ( n74398 , n74397 , n32486 );
and ( n74399 , n31811 , n41278 );
or ( n74400 , C0 , n74368 , n74377 , n74398 , n74399 );
buf ( n74401 , n74400 );
buf ( n74402 , n74401 );
xor ( n74403 , n31507 , n31509 );
and ( n74404 , n74403 , n31550 );
not ( n74405 , n39979 );
and ( n74406 , n74405 , n31507 );
buf ( n74407 , n31170 );
and ( n74408 , n74407 , n39979 );
or ( n74409 , n74406 , n74408 );
and ( n74410 , n74409 , n31538 );
and ( n74411 , n31507 , n40143 );
or ( n74412 , n74404 , n74410 , n74411 );
and ( n74413 , n74412 , n31557 );
and ( n74414 , n31507 , n40154 );
or ( n74415 , C0 , n74413 , n74414 );
buf ( n74416 , n74415 );
buf ( n74417 , n74416 );
buf ( n74418 , n30987 );
not ( n74419 , n34150 );
and ( n74420 , n74419 , n32767 );
not ( n74421 , n58762 );
and ( n74422 , n74421 , n32767 );
and ( n74423 , n32789 , n58762 );
or ( n74424 , n74422 , n74423 );
and ( n74425 , n74424 , n34150 );
or ( n74426 , n74420 , n74425 );
and ( n74427 , n74426 , n33381 );
not ( n74428 , n58770 );
not ( n74429 , n58762 );
and ( n74430 , n74429 , n32767 );
and ( n74431 , n34301 , n58762 );
or ( n74432 , n74430 , n74431 );
and ( n74433 , n74428 , n74432 );
and ( n74434 , n34301 , n58770 );
or ( n74435 , n74433 , n74434 );
and ( n74436 , n74435 , n33375 );
not ( n74437 , n32968 );
not ( n74438 , n58770 );
not ( n74439 , n58762 );
and ( n74440 , n74439 , n32767 );
and ( n74441 , n34301 , n58762 );
or ( n74442 , n74440 , n74441 );
and ( n74443 , n74438 , n74442 );
and ( n74444 , n34301 , n58770 );
or ( n74445 , n74443 , n74444 );
and ( n74446 , n74437 , n74445 );
not ( n74447 , n58790 );
not ( n74448 , n58792 );
and ( n74449 , n74448 , n74445 );
and ( n74450 , n34761 , n58792 );
or ( n74451 , n74449 , n74450 );
and ( n74452 , n74447 , n74451 );
and ( n74453 , n35050 , n58790 );
or ( n74454 , n74452 , n74453 );
and ( n74455 , n74454 , n32968 );
or ( n74456 , n74446 , n74455 );
and ( n74457 , n74456 , n33370 );
and ( n74458 , n32767 , n35062 );
or ( n74459 , C0 , n74427 , n74436 , n74457 , n74458 );
buf ( n74460 , n74459 );
buf ( n74461 , n74460 );
buf ( n74462 , n30987 );
buf ( n74463 , n31655 );
buf ( n74464 , n31655 );
buf ( n74465 , n30987 );
buf ( n74466 , n31655 );
buf ( n74467 , n31655 );
buf ( n74468 , n30987 );
and ( n74469 , n70129 , n33377 );
not ( n74470 , n48545 );
and ( n74471 , n74470 , n52669 );
and ( n74472 , n74338 , n48545 );
or ( n74473 , n74471 , n74472 );
and ( n74474 , n74473 , n32890 );
not ( n74475 , n48557 );
and ( n74476 , n74475 , n52669 );
and ( n74477 , n74338 , n48557 );
or ( n74478 , n74476 , n74477 );
and ( n74479 , n74478 , n33038 );
and ( n74480 , n52669 , n48571 );
or ( n74481 , n74474 , n74479 , n74480 );
and ( n74482 , n74481 , n33208 );
and ( n74483 , n52669 , n48577 );
or ( n74484 , C0 , n74469 , n74482 , n74483 );
buf ( n74485 , n74484 );
buf ( n74486 , n74485 );
buf ( n74487 , n30987 );
buf ( n74488 , n31655 );
not ( n74489 , n31437 );
and ( n74490 , n74489 , n56333 );
and ( n74491 , n56342 , n31437 );
or ( n74492 , n74490 , n74491 );
and ( n74493 , n74492 , n31468 );
not ( n74494 , n41837 );
and ( n74495 , n74494 , n56333 );
and ( n74496 , n62186 , n41837 );
or ( n74497 , n74495 , n74496 );
and ( n74498 , n74497 , n31521 );
and ( n74499 , n56333 , n42158 );
or ( n74500 , n74493 , n74498 , n74499 );
and ( n74501 , n74500 , n31557 );
and ( n74502 , n56333 , n40154 );
or ( n74503 , C0 , n74501 , n74502 );
buf ( n74504 , n74503 );
buf ( n74505 , n74504 );
not ( n74506 , n40163 );
and ( n74507 , n74506 , n32001 );
not ( n74508 , n56988 );
and ( n74509 , n74508 , n32001 );
and ( n74510 , n32147 , n56988 );
or ( n74511 , n74509 , n74510 );
and ( n74512 , n74511 , n40163 );
or ( n74513 , n74507 , n74512 );
and ( n74514 , n74513 , n32498 );
not ( n74515 , n56996 );
not ( n74516 , n56988 );
and ( n74517 , n74516 , n32001 );
and ( n74518 , n49314 , n56988 );
or ( n74519 , n74517 , n74518 );
and ( n74520 , n74515 , n74519 );
and ( n74521 , n49314 , n56996 );
or ( n74522 , n74520 , n74521 );
and ( n74523 , n74522 , n32473 );
not ( n74524 , n32475 );
not ( n74525 , n56996 );
not ( n74526 , n56988 );
and ( n74527 , n74526 , n32001 );
and ( n74528 , n49314 , n56988 );
or ( n74529 , n74527 , n74528 );
and ( n74530 , n74525 , n74529 );
and ( n74531 , n49314 , n56996 );
or ( n74532 , n74530 , n74531 );
and ( n74533 , n74524 , n74532 );
not ( n74534 , n57016 );
not ( n74535 , n57018 );
and ( n74536 , n74535 , n74532 );
and ( n74537 , n49340 , n57018 );
or ( n74538 , n74536 , n74537 );
and ( n74539 , n74534 , n74538 );
and ( n74540 , n49348 , n57016 );
or ( n74541 , n74539 , n74540 );
and ( n74542 , n74541 , n32475 );
or ( n74543 , n74533 , n74542 );
and ( n74544 , n74543 , n32486 );
and ( n74545 , n32001 , n41278 );
or ( n74546 , C0 , n74514 , n74523 , n74544 , n74545 );
buf ( n74547 , n74546 );
buf ( n74548 , n74547 );
buf ( n74549 , n30987 );
buf ( n74550 , n31655 );
buf ( n74551 , n31655 );
buf ( n74552 , n30987 );
not ( n74553 , n34150 );
and ( n74554 , n74553 , n32861 );
not ( n74555 , n60126 );
and ( n74556 , n74555 , n32861 );
and ( n74557 , n32889 , n60126 );
or ( n74558 , n74556 , n74557 );
and ( n74559 , n74558 , n34150 );
or ( n74560 , n74554 , n74559 );
and ( n74561 , n74560 , n33381 );
not ( n74562 , n60134 );
not ( n74563 , n60126 );
and ( n74564 , n74563 , n32861 );
and ( n74565 , n52819 , n60126 );
or ( n74566 , n74564 , n74565 );
and ( n74567 , n74562 , n74566 );
and ( n74568 , n52819 , n60134 );
or ( n74569 , n74567 , n74568 );
and ( n74570 , n74569 , n33375 );
not ( n74571 , n32968 );
not ( n74572 , n60134 );
not ( n74573 , n60126 );
and ( n74574 , n74573 , n32861 );
and ( n74575 , n52819 , n60126 );
or ( n74576 , n74574 , n74575 );
and ( n74577 , n74572 , n74576 );
and ( n74578 , n52819 , n60134 );
or ( n74579 , n74577 , n74578 );
and ( n74580 , n74571 , n74579 );
not ( n74581 , n60154 );
not ( n74582 , n60156 );
and ( n74583 , n74582 , n74579 );
and ( n74584 , n52845 , n60156 );
or ( n74585 , n74583 , n74584 );
and ( n74586 , n74581 , n74585 );
and ( n74587 , n52855 , n60154 );
or ( n74588 , n74586 , n74587 );
and ( n74589 , n74588 , n32968 );
or ( n74590 , n74580 , n74589 );
and ( n74591 , n74590 , n33370 );
and ( n74592 , n32861 , n35062 );
or ( n74593 , C0 , n74561 , n74570 , n74591 , n74592 );
buf ( n74594 , n74593 );
buf ( n74595 , n74594 );
and ( n74596 , n54688 , n33377 );
not ( n74597 , n48545 );
and ( n74598 , n74597 , n67546 );
and ( n74599 , n71468 , n48545 );
or ( n74600 , n74598 , n74599 );
and ( n74601 , n74600 , n32890 );
not ( n74602 , n48557 );
and ( n74603 , n74602 , n67546 );
and ( n74604 , n71468 , n48557 );
or ( n74605 , n74603 , n74604 );
and ( n74606 , n74605 , n33038 );
and ( n74607 , n67546 , n48571 );
or ( n74608 , n74601 , n74606 , n74607 );
and ( n74609 , n74608 , n33208 );
and ( n74610 , n67546 , n48577 );
or ( n74611 , C0 , n74596 , n74609 , n74610 );
buf ( n74612 , n74611 );
buf ( n74613 , n74612 );
buf ( n74614 , n31655 );
buf ( n74615 , n31655 );
buf ( n74616 , n30987 );
buf ( n74617 , n30987 );
buf ( n74618 , n30987 );
buf ( n74619 , n30987 );
buf ( n74620 , n31655 );
not ( n74621 , n43755 );
and ( n74622 , n74621 , n43615 );
xor ( n74623 , n52306 , n52323 );
and ( n74624 , n74623 , n43755 );
or ( n74625 , n74622 , n74624 );
and ( n74626 , n74625 , n43774 );
not ( n74627 , n44663 );
and ( n74628 , n74627 , n44527 );
xor ( n74629 , n52344 , n52361 );
and ( n74630 , n74629 , n44663 );
or ( n74631 , n74628 , n74630 );
and ( n74632 , n74631 , n44682 );
and ( n74633 , n55546 , n44695 );
or ( n74634 , n74626 , n74632 , n74633 );
buf ( n74635 , n74634 );
buf ( n74636 , n74635 );
buf ( n74637 , n31655 );
buf ( n74638 , n30987 );
buf ( n74639 , n31655 );
buf ( n74640 , n31655 );
buf ( n74641 , n30987 );
buf ( n74642 , RI15b46c98_280);
and ( n74643 , n74642 , n33377 );
not ( n74644 , n48545 );
and ( n74645 , n74644 , n57167 );
not ( n74646 , n39572 );
and ( n74647 , n74646 , n39516 );
xor ( n74648 , n42617 , n42636 );
and ( n74649 , n74648 , n39572 );
or ( n74650 , n74647 , n74649 );
and ( n74651 , n74650 , n48545 );
or ( n74652 , n74645 , n74651 );
and ( n74653 , n74652 , n32890 );
not ( n74654 , n48557 );
and ( n74655 , n74654 , n57167 );
and ( n74656 , n74650 , n48557 );
or ( n74657 , n74655 , n74656 );
and ( n74658 , n74657 , n33038 );
and ( n74659 , n57167 , n48571 );
or ( n74660 , n74653 , n74658 , n74659 );
and ( n74661 , n74660 , n33208 );
and ( n74662 , n57167 , n48577 );
or ( n74663 , C0 , n74643 , n74661 , n74662 );
buf ( n74664 , n74663 );
buf ( n74665 , n74664 );
buf ( n74666 , n30987 );
not ( n74667 , n36587 );
and ( n74668 , n74667 , n36413 );
xor ( n74669 , n50176 , n50211 );
and ( n74670 , n74669 , n36587 );
or ( n74671 , n74668 , n74670 );
and ( n74672 , n74671 , n36596 );
not ( n74673 , n37485 );
and ( n74674 , n74673 , n37315 );
xor ( n74675 , n50226 , n50261 );
and ( n74676 , n74675 , n37485 );
or ( n74677 , n74674 , n74676 );
and ( n74678 , n74677 , n37494 );
and ( n74679 , n41858 , n37506 );
or ( n74680 , n74672 , n74678 , n74679 );
buf ( n74681 , n74680 );
buf ( n74682 , n74681 );
buf ( n74683 , n31655 );
and ( n74684 , n50441 , n50275 );
not ( n74685 , n50278 );
and ( n74686 , n74685 , n50409 );
and ( n74687 , n50441 , n50278 );
or ( n74688 , n74686 , n74687 );
and ( n74689 , n74688 , n32421 );
not ( n74690 , n50002 );
and ( n74691 , n74690 , n50409 );
and ( n74692 , n50441 , n50002 );
or ( n74693 , n74691 , n74692 );
and ( n74694 , n74693 , n32419 );
not ( n74695 , n50289 );
and ( n74696 , n74695 , n50409 );
and ( n74697 , n50441 , n50289 );
or ( n74698 , n74696 , n74697 );
and ( n74699 , n74698 , n32417 );
not ( n74700 , n50008 );
and ( n74701 , n74700 , n50409 );
and ( n74702 , n50441 , n50008 );
or ( n74703 , n74701 , n74702 );
and ( n74704 , n74703 , n32415 );
not ( n74705 , n47331 );
and ( n74706 , n74705 , n50409 );
and ( n74707 , n50419 , n47331 );
or ( n74708 , n74706 , n74707 );
and ( n74709 , n74708 , n32413 );
not ( n74710 , n50067 );
and ( n74711 , n74710 , n50409 );
and ( n74712 , n50419 , n50067 );
or ( n74713 , n74711 , n74712 );
and ( n74714 , n74713 , n32411 );
not ( n74715 , n31728 );
and ( n74716 , n74715 , n50409 );
and ( n74717 , n60983 , n31728 );
or ( n74718 , n74716 , n74717 );
and ( n74719 , n74718 , n32253 );
not ( n74720 , n32283 );
and ( n74721 , n74720 , n50409 );
and ( n74722 , n60994 , n32283 );
or ( n74723 , n74721 , n74722 );
and ( n74724 , n74723 , n32398 );
and ( n74725 , n50458 , n50334 );
or ( n74726 , n74684 , n74689 , n74694 , n74699 , n74704 , n74709 , n74714 , n74719 , n74724 , n74725 );
and ( n74727 , n74726 , n32456 );
and ( n74728 , n37535 , n32489 );
and ( n74729 , n50409 , n50345 );
or ( n74730 , C0 , n74727 , n74728 , n74729 );
buf ( n74731 , n74730 );
buf ( n74732 , n74731 );
not ( n74733 , n40163 );
and ( n74734 , n74733 , n31836 );
not ( n74735 , n45227 );
and ( n74736 , n74735 , n31836 );
and ( n74737 , n32235 , n45227 );
or ( n74738 , n74736 , n74737 );
and ( n74739 , n74738 , n40163 );
or ( n74740 , n74734 , n74739 );
and ( n74741 , n74740 , n32498 );
not ( n74742 , n45235 );
not ( n74743 , n45227 );
and ( n74744 , n74743 , n31836 );
and ( n74745 , n42188 , n45227 );
or ( n74746 , n74744 , n74745 );
and ( n74747 , n74742 , n74746 );
and ( n74748 , n42188 , n45235 );
or ( n74749 , n74747 , n74748 );
and ( n74750 , n74749 , n32473 );
not ( n74751 , n32475 );
not ( n74752 , n45235 );
not ( n74753 , n45227 );
and ( n74754 , n74753 , n31836 );
and ( n74755 , n42188 , n45227 );
or ( n74756 , n74754 , n74755 );
and ( n74757 , n74752 , n74756 );
and ( n74758 , n42188 , n45235 );
or ( n74759 , n74757 , n74758 );
and ( n74760 , n74751 , n74759 );
not ( n74761 , n45255 );
not ( n74762 , n45257 );
and ( n74763 , n74762 , n74759 );
and ( n74764 , n42216 , n45257 );
or ( n74765 , n74763 , n74764 );
and ( n74766 , n74761 , n74765 );
and ( n74767 , n42224 , n45255 );
or ( n74768 , n74766 , n74767 );
and ( n74769 , n74768 , n32475 );
or ( n74770 , n74760 , n74769 );
and ( n74771 , n74770 , n32486 );
and ( n74772 , n31836 , n41278 );
or ( n74773 , C0 , n74741 , n74750 , n74771 , n74772 );
buf ( n74774 , n74773 );
buf ( n74775 , n74774 );
and ( n74776 , n60741 , n31645 );
not ( n74777 , n45274 );
buf ( n74778 , RI15b53e98_728);
and ( n74779 , n74777 , n74778 );
buf ( n74780 , n74779 );
and ( n74781 , n74780 , n31373 );
not ( n74782 , n45280 );
and ( n74783 , n74782 , n74778 );
and ( n74784 , n60747 , n45280 );
or ( n74785 , n74783 , n74784 );
and ( n74786 , n74785 , n31468 );
and ( n74787 , n74778 , n45802 );
or ( n74788 , n74781 , n74786 , n74787 );
and ( n74789 , n74788 , n31557 );
and ( n74790 , n74778 , n45808 );
or ( n74791 , C0 , n74776 , n74789 , n74790 );
buf ( n74792 , n74791 );
buf ( n74793 , n74792 );
buf ( n74794 , n31655 );
buf ( n74795 , n30987 );
buf ( n74796 , n30987 );
buf ( n74797 , n31655 );
buf ( n74798 , n31655 );
not ( n74799 , n46356 );
and ( n74800 , n74799 , n31222 );
not ( n74801 , n55263 );
and ( n74802 , n74801 , n31222 );
and ( n74803 , n31238 , n55263 );
or ( n74804 , n74802 , n74803 );
and ( n74805 , n74804 , n46356 );
or ( n74806 , n74800 , n74805 );
and ( n74807 , n74806 , n31649 );
not ( n74808 , n55271 );
not ( n74809 , n55263 );
and ( n74810 , n74809 , n31222 );
and ( n74811 , n49901 , n55263 );
or ( n74812 , n74810 , n74811 );
and ( n74813 , n74808 , n74812 );
and ( n74814 , n49901 , n55271 );
or ( n74815 , n74813 , n74814 );
and ( n74816 , n74815 , n31643 );
not ( n74817 , n31452 );
not ( n74818 , n55271 );
not ( n74819 , n55263 );
and ( n74820 , n74819 , n31222 );
and ( n74821 , n49901 , n55263 );
or ( n74822 , n74820 , n74821 );
and ( n74823 , n74818 , n74822 );
and ( n74824 , n49901 , n55271 );
or ( n74825 , n74823 , n74824 );
and ( n74826 , n74817 , n74825 );
not ( n74827 , n55291 );
not ( n74828 , n55293 );
and ( n74829 , n74828 , n74825 );
and ( n74830 , n49925 , n55293 );
or ( n74831 , n74829 , n74830 );
and ( n74832 , n74827 , n74831 );
and ( n74833 , n49933 , n55291 );
or ( n74834 , n74832 , n74833 );
and ( n74835 , n74834 , n31452 );
or ( n74836 , n74826 , n74835 );
and ( n74837 , n74836 , n31638 );
and ( n74838 , n31222 , n47277 );
or ( n74839 , C0 , n74807 , n74816 , n74837 , n74838 );
buf ( n74840 , n74839 );
buf ( n74841 , n74840 );
xor ( n74842 , n46146 , n49990 );
and ( n74843 , n74842 , n32431 );
not ( n74844 , n50002 );
and ( n74845 , n74844 , n46146 );
and ( n74846 , n40323 , n50002 );
or ( n74847 , n74845 , n74846 );
and ( n74848 , n74847 , n32419 );
not ( n74849 , n50008 );
and ( n74850 , n74849 , n46146 );
not ( n74851 , n47910 );
and ( n74852 , n74851 , n64257 );
and ( n74853 , n64273 , n47910 );
or ( n74854 , n74852 , n74853 );
and ( n74855 , n74854 , n50008 );
or ( n74856 , n74850 , n74855 );
and ( n74857 , n74856 , n32415 );
not ( n74858 , n50067 );
and ( n74859 , n74858 , n46146 );
and ( n74860 , n31893 , n50067 );
or ( n74861 , n74859 , n74860 );
and ( n74862 , n74861 , n32411 );
and ( n74863 , n46146 , n50098 );
or ( n74864 , n74843 , n74848 , n74857 , n74862 , n74863 );
and ( n74865 , n74864 , n32456 );
and ( n74866 , n46146 , n47409 );
or ( n74867 , C0 , n74865 , n74866 );
buf ( n74868 , n74867 );
buf ( n74869 , n74868 );
buf ( n74870 , n30987 );
not ( n74871 , n34150 );
and ( n74872 , n74871 , n32687 );
not ( n74873 , n56239 );
and ( n74874 , n74873 , n32687 );
and ( n74875 , n32689 , n56239 );
or ( n74876 , n74874 , n74875 );
and ( n74877 , n74876 , n34150 );
or ( n74878 , n74872 , n74877 );
and ( n74879 , n74878 , n33381 );
not ( n74880 , n56247 );
not ( n74881 , n56239 );
and ( n74882 , n74881 , n32687 );
and ( n74883 , n50682 , n56239 );
or ( n74884 , n74882 , n74883 );
and ( n74885 , n74880 , n74884 );
and ( n74886 , n50682 , n56247 );
or ( n74887 , n74885 , n74886 );
and ( n74888 , n74887 , n33375 );
not ( n74889 , n32968 );
not ( n74890 , n56247 );
not ( n74891 , n56239 );
and ( n74892 , n74891 , n32687 );
and ( n74893 , n50682 , n56239 );
or ( n74894 , n74892 , n74893 );
and ( n74895 , n74890 , n74894 );
and ( n74896 , n50682 , n56247 );
or ( n74897 , n74895 , n74896 );
and ( n74898 , n74889 , n74897 );
not ( n74899 , n56267 );
not ( n74900 , n56269 );
and ( n74901 , n74900 , n74897 );
and ( n74902 , n50706 , n56269 );
or ( n74903 , n74901 , n74902 );
and ( n74904 , n74899 , n74903 );
and ( n74905 , n50714 , n56267 );
or ( n74906 , n74904 , n74905 );
and ( n74907 , n74906 , n32968 );
or ( n74908 , n74898 , n74907 );
and ( n74909 , n74908 , n33370 );
and ( n74910 , n32687 , n35062 );
or ( n74911 , C0 , n74879 , n74888 , n74909 , n74910 );
buf ( n74912 , n74911 );
buf ( n74913 , n74912 );
buf ( n74914 , n30987 );
buf ( n74915 , n31655 );
buf ( n74916 , n31655 );
buf ( n74917 , n30987 );
not ( n74918 , n34150 );
and ( n74919 , n74918 , n32846 );
not ( n74920 , n56192 );
and ( n74921 , n74920 , n32846 );
and ( n74922 , n32856 , n56192 );
or ( n74923 , n74921 , n74922 );
and ( n74924 , n74923 , n34150 );
or ( n74925 , n74919 , n74924 );
and ( n74926 , n74925 , n33381 );
not ( n74927 , n56200 );
not ( n74928 , n56192 );
and ( n74929 , n74928 , n32846 );
and ( n74930 , n48160 , n56192 );
or ( n74931 , n74929 , n74930 );
and ( n74932 , n74927 , n74931 );
and ( n74933 , n48160 , n56200 );
or ( n74934 , n74932 , n74933 );
and ( n74935 , n74934 , n33375 );
not ( n74936 , n32968 );
not ( n74937 , n56200 );
not ( n74938 , n56192 );
and ( n74939 , n74938 , n32846 );
and ( n74940 , n48160 , n56192 );
or ( n74941 , n74939 , n74940 );
and ( n74942 , n74937 , n74941 );
and ( n74943 , n48160 , n56200 );
or ( n74944 , n74942 , n74943 );
and ( n74945 , n74936 , n74944 );
not ( n74946 , n56220 );
not ( n74947 , n56222 );
and ( n74948 , n74947 , n74944 );
and ( n74949 , n48186 , n56222 );
or ( n74950 , n74948 , n74949 );
and ( n74951 , n74946 , n74950 );
and ( n74952 , n48196 , n56220 );
or ( n74953 , n74951 , n74952 );
and ( n74954 , n74953 , n32968 );
or ( n74955 , n74945 , n74954 );
and ( n74956 , n74955 , n33370 );
and ( n74957 , n32846 , n35062 );
or ( n74958 , C0 , n74926 , n74935 , n74956 , n74957 );
buf ( n74959 , n74958 );
buf ( n74960 , n74959 );
not ( n74961 , n34150 );
and ( n74962 , n74961 , n32830 );
not ( n74963 , n59574 );
and ( n74964 , n74963 , n32830 );
and ( n74965 , n32856 , n59574 );
or ( n74966 , n74964 , n74965 );
and ( n74967 , n74966 , n34150 );
or ( n74968 , n74962 , n74967 );
and ( n74969 , n74968 , n33381 );
not ( n74970 , n59582 );
not ( n74971 , n59574 );
and ( n74972 , n74971 , n32830 );
and ( n74973 , n48160 , n59574 );
or ( n74974 , n74972 , n74973 );
and ( n74975 , n74970 , n74974 );
and ( n74976 , n48160 , n59582 );
or ( n74977 , n74975 , n74976 );
and ( n74978 , n74977 , n33375 );
not ( n74979 , n32968 );
not ( n74980 , n59582 );
not ( n74981 , n59574 );
and ( n74982 , n74981 , n32830 );
and ( n74983 , n48160 , n59574 );
or ( n74984 , n74982 , n74983 );
and ( n74985 , n74980 , n74984 );
and ( n74986 , n48160 , n59582 );
or ( n74987 , n74985 , n74986 );
and ( n74988 , n74979 , n74987 );
not ( n74989 , n59602 );
not ( n74990 , n59604 );
and ( n74991 , n74990 , n74987 );
and ( n74992 , n48186 , n59604 );
or ( n74993 , n74991 , n74992 );
and ( n74994 , n74989 , n74993 );
and ( n74995 , n48196 , n59602 );
or ( n74996 , n74994 , n74995 );
and ( n74997 , n74996 , n32968 );
or ( n74998 , n74988 , n74997 );
and ( n74999 , n74998 , n33370 );
and ( n75000 , n32830 , n35062 );
or ( n75001 , C0 , n74969 , n74978 , n74999 , n75000 );
buf ( n75002 , n75001 );
buf ( n75003 , n75002 );
buf ( n75004 , n30987 );
buf ( n75005 , n31655 );
buf ( n75006 , n31655 );
buf ( n75007 , n30987 );
buf ( n75008 , n31655 );
buf ( n75009 , n31655 );
xor ( n75010 , n46185 , n49993 );
and ( n75011 , n75010 , n32431 );
not ( n75012 , n50002 );
and ( n75013 , n75012 , n46185 );
and ( n75014 , n40514 , n50002 );
or ( n75015 , n75013 , n75014 );
and ( n75016 , n75015 , n32419 );
not ( n75017 , n50008 );
and ( n75018 , n75017 , n46185 );
not ( n75019 , n47910 );
and ( n75020 , n75019 , n73740 );
and ( n75021 , n73756 , n47910 );
or ( n75022 , n75020 , n75021 );
and ( n75023 , n75022 , n50008 );
or ( n75024 , n75018 , n75023 );
and ( n75025 , n75024 , n32415 );
not ( n75026 , n50067 );
and ( n75027 , n75026 , n46185 );
and ( n75028 , n66304 , n50067 );
or ( n75029 , n75027 , n75028 );
and ( n75030 , n75029 , n32411 );
and ( n75031 , n46185 , n50098 );
or ( n75032 , n75011 , n75016 , n75025 , n75030 , n75031 );
and ( n75033 , n75032 , n32456 );
and ( n75034 , n46185 , n47409 );
or ( n75035 , C0 , n75033 , n75034 );
buf ( n75036 , n75035 );
buf ( n75037 , n75036 );
not ( n75038 , n46356 );
and ( n75039 , n75038 , n31114 );
not ( n75040 , n55263 );
and ( n75041 , n75040 , n31114 );
and ( n75042 , n31138 , n55263 );
or ( n75043 , n75041 , n75042 );
and ( n75044 , n75043 , n46356 );
or ( n75045 , n75039 , n75044 );
and ( n75046 , n75045 , n31649 );
not ( n75047 , n55271 );
not ( n75048 , n55263 );
and ( n75049 , n75048 , n31114 );
and ( n75050 , n56920 , n55263 );
or ( n75051 , n75049 , n75050 );
and ( n75052 , n75047 , n75051 );
and ( n75053 , n56920 , n55271 );
or ( n75054 , n75052 , n75053 );
and ( n75055 , n75054 , n31643 );
not ( n75056 , n31452 );
not ( n75057 , n55271 );
not ( n75058 , n55263 );
and ( n75059 , n75058 , n31114 );
and ( n75060 , n56920 , n55263 );
or ( n75061 , n75059 , n75060 );
and ( n75062 , n75057 , n75061 );
and ( n75063 , n56920 , n55271 );
or ( n75064 , n75062 , n75063 );
and ( n75065 , n75056 , n75064 );
not ( n75066 , n55291 );
not ( n75067 , n55293 );
and ( n75068 , n75067 , n75064 );
and ( n75069 , n56946 , n55293 );
or ( n75070 , n75068 , n75069 );
and ( n75071 , n75066 , n75070 );
and ( n75072 , n56954 , n55291 );
or ( n75073 , n75071 , n75072 );
and ( n75074 , n75073 , n31452 );
or ( n75075 , n75065 , n75074 );
and ( n75076 , n75075 , n31638 );
and ( n75077 , n31114 , n47277 );
or ( n75078 , C0 , n75046 , n75055 , n75076 , n75077 );
buf ( n75079 , n75078 );
buf ( n75080 , n75079 );
buf ( n75081 , n30987 );
buf ( n75082 , n31655 );
not ( n75083 , n35542 );
and ( n75084 , n75083 , n41850 );
buf ( n75085 , RI15b455a0_231);
and ( n75086 , n75085 , n35542 );
or ( n75087 , n75084 , n75086 );
buf ( n75088 , n75087 );
buf ( n75089 , n75088 );
buf ( n75090 , n30987 );
buf ( n75091 , n30987 );
not ( n75092 , n34150 );
and ( n75093 , n75092 , n32708 );
not ( n75094 , n56836 );
and ( n75095 , n75094 , n32708 );
and ( n75096 , n32722 , n56836 );
or ( n75097 , n75095 , n75096 );
and ( n75098 , n75097 , n34150 );
or ( n75099 , n75093 , n75098 );
and ( n75100 , n75099 , n33381 );
not ( n75101 , n56844 );
not ( n75102 , n56836 );
and ( n75103 , n75102 , n32708 );
and ( n75104 , n42565 , n56836 );
or ( n75105 , n75103 , n75104 );
and ( n75106 , n75101 , n75105 );
and ( n75107 , n42565 , n56844 );
or ( n75108 , n75106 , n75107 );
and ( n75109 , n75108 , n33375 );
not ( n75110 , n32968 );
not ( n75111 , n56844 );
not ( n75112 , n56836 );
and ( n75113 , n75112 , n32708 );
and ( n75114 , n42565 , n56836 );
or ( n75115 , n75113 , n75114 );
and ( n75116 , n75111 , n75115 );
and ( n75117 , n42565 , n56844 );
or ( n75118 , n75116 , n75117 );
and ( n75119 , n75110 , n75118 );
not ( n75120 , n56864 );
not ( n75121 , n56866 );
and ( n75122 , n75121 , n75118 );
and ( n75123 , n42589 , n56866 );
or ( n75124 , n75122 , n75123 );
and ( n75125 , n75120 , n75124 );
and ( n75126 , n42597 , n56864 );
or ( n75127 , n75125 , n75126 );
and ( n75128 , n75127 , n32968 );
or ( n75129 , n75119 , n75128 );
and ( n75130 , n75129 , n33370 );
and ( n75131 , n32708 , n35062 );
or ( n75132 , C0 , n75100 , n75109 , n75130 , n75131 );
buf ( n75133 , n75132 );
buf ( n75134 , n75133 );
buf ( n75135 , n31655 );
buf ( n75136 , n31655 );
xor ( n75137 , n50971 , n64711 );
and ( n75138 , n75137 , n32431 );
not ( n75139 , n50002 );
and ( n75140 , n75139 , n50971 );
and ( n75141 , n40641 , n50002 );
or ( n75142 , n75140 , n75141 );
and ( n75143 , n75142 , n32419 );
not ( n75144 , n50008 );
and ( n75145 , n75144 , n50971 );
not ( n75146 , n51594 );
and ( n75147 , n75146 , n51446 );
xor ( n75148 , n51601 , n51605 );
and ( n75149 , n75148 , n51594 );
or ( n75150 , n75147 , n75149 );
and ( n75151 , n75150 , n50008 );
or ( n75152 , n75145 , n75151 );
and ( n75153 , n75152 , n32415 );
not ( n75154 , n50067 );
and ( n75155 , n75154 , n50971 );
and ( n75156 , n31966 , n60510 );
and ( n75157 , n31968 , n60512 );
and ( n75158 , n31970 , n60514 );
and ( n75159 , n31972 , n60516 );
and ( n75160 , n31974 , n60518 );
and ( n75161 , n31976 , n60520 );
and ( n75162 , n31978 , n60522 );
and ( n75163 , n31980 , n60524 );
and ( n75164 , n31982 , n60526 );
and ( n75165 , n31984 , n60528 );
and ( n75166 , n31986 , n60530 );
and ( n75167 , n31988 , n60532 );
and ( n75168 , n31990 , n60534 );
and ( n75169 , n31992 , n60536 );
and ( n75170 , n31994 , n60538 );
and ( n75171 , n31996 , n60540 );
or ( n75172 , n75156 , n75157 , n75158 , n75159 , n75160 , n75161 , n75162 , n75163 , n75164 , n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , n75171 );
and ( n75173 , n75172 , n50067 );
or ( n75174 , n75155 , n75173 );
and ( n75175 , n75174 , n32411 );
and ( n75176 , n50971 , n50098 );
or ( n75177 , n75138 , n75143 , n75153 , n75175 , n75176 );
and ( n75178 , n75177 , n32456 );
and ( n75179 , n50971 , n47409 );
or ( n75180 , C0 , n75178 , n75179 );
buf ( n75181 , n75180 );
buf ( n75182 , n75181 );
buf ( n75183 , n30987 );
buf ( n75184 , n31655 );
not ( n75185 , n46356 );
and ( n75186 , n75185 , n31327 );
not ( n75187 , n64746 );
and ( n75188 , n75187 , n31327 );
and ( n75189 , n31339 , n64746 );
or ( n75190 , n75188 , n75189 );
and ( n75191 , n75190 , n46356 );
or ( n75192 , n75186 , n75191 );
and ( n75193 , n75192 , n31649 );
not ( n75194 , n64754 );
not ( n75195 , n64746 );
and ( n75196 , n75195 , n31327 );
and ( n75197 , n47449 , n64746 );
or ( n75198 , n75196 , n75197 );
and ( n75199 , n75194 , n75198 );
and ( n75200 , n47449 , n64754 );
or ( n75201 , n75199 , n75200 );
and ( n75202 , n75201 , n31643 );
not ( n75203 , n31452 );
not ( n75204 , n64754 );
not ( n75205 , n64746 );
and ( n75206 , n75205 , n31327 );
and ( n75207 , n47449 , n64746 );
or ( n75208 , n75206 , n75207 );
and ( n75209 , n75204 , n75208 );
and ( n75210 , n47449 , n64754 );
or ( n75211 , n75209 , n75210 );
and ( n75212 , n75203 , n75211 );
not ( n75213 , n64774 );
not ( n75214 , n64776 );
and ( n75215 , n75214 , n75211 );
and ( n75216 , n47485 , n64776 );
or ( n75217 , n75215 , n75216 );
and ( n75218 , n75213 , n75217 );
and ( n75219 , n47503 , n64774 );
or ( n75220 , n75218 , n75219 );
and ( n75221 , n75220 , n31452 );
or ( n75222 , n75212 , n75221 );
and ( n75223 , n75222 , n31638 );
and ( n75224 , n31327 , n47277 );
or ( n75225 , C0 , n75193 , n75202 , n75223 , n75224 );
buf ( n75226 , n75225 );
buf ( n75227 , n75226 );
buf ( n75228 , n31655 );
not ( n75229 , n33419 );
and ( n75230 , n75229 , n31563 );
xor ( n75231 , n57502 , n57505 );
and ( n75232 , n75231 , n33419 );
or ( n75233 , n75230 , n75232 );
and ( n75234 , n75233 , n31529 );
not ( n75235 , n33734 );
and ( n75236 , n75235 , n31563 );
not ( n75237 , n33533 );
xor ( n75238 , n57514 , n57517 );
and ( n75239 , n75237 , n75238 );
xnor ( n75240 , n57525 , n57528 );
and ( n75241 , n75240 , n33533 );
or ( n75242 , n75239 , n75241 );
and ( n75243 , n75242 , n33734 );
or ( n75244 , n75236 , n75243 );
and ( n75245 , n75244 , n31527 );
and ( n75246 , n31563 , n33942 );
or ( n75247 , n75234 , n75245 , n75246 );
and ( n75248 , n75247 , n31557 );
and ( n75249 , n35482 , n31643 );
not ( n75250 , n31452 );
and ( n75251 , n75250 , n35482 );
xor ( n75252 , n31563 , n59437 );
and ( n75253 , n75252 , n31452 );
or ( n75254 , n75251 , n75253 );
and ( n75255 , n75254 , n31638 );
and ( n75256 , n35389 , n33973 );
and ( n75257 , n31563 , n33978 );
or ( n75258 , C0 , n75248 , n75249 , n75255 , n75256 , n75257 );
buf ( n75259 , n75258 );
buf ( n75260 , n75259 );
buf ( n75261 , n30987 );
buf ( n75262 , n30987 );
and ( n75263 , n31581 , n31007 );
not ( n75264 , n31077 );
and ( n75265 , n75264 , n34005 );
buf ( n75266 , n75265 );
and ( n75267 , n75266 , n31373 );
not ( n75268 , n31402 );
and ( n75269 , n75268 , n34005 );
buf ( n75270 , n75269 );
and ( n75271 , n75270 , n31408 );
not ( n75272 , n31437 );
and ( n75273 , n75272 , n34005 );
not ( n75274 , n31455 );
and ( n75275 , n75274 , n34050 );
xor ( n75276 , n34005 , n34018 );
and ( n75277 , n75276 , n31455 );
or ( n75278 , n75275 , n75277 );
and ( n75279 , n75278 , n31437 );
or ( n75280 , n75273 , n75279 );
and ( n75281 , n75280 , n31468 );
not ( n75282 , n31497 );
and ( n75283 , n75282 , n34005 );
not ( n75284 , n31454 );
not ( n75285 , n31501 );
and ( n75286 , n75285 , n34050 );
xor ( n75287 , n34051 , n34070 );
and ( n75288 , n75287 , n31501 );
or ( n75289 , n75286 , n75288 );
and ( n75290 , n75284 , n75289 );
and ( n75291 , n75276 , n31454 );
or ( n75292 , n75290 , n75291 );
and ( n75293 , n75292 , n31497 );
or ( n75294 , n75283 , n75293 );
and ( n75295 , n75294 , n31521 );
and ( n75296 , n34005 , n31553 );
or ( n75297 , n75267 , n75271 , n75281 , n75295 , n75296 );
and ( n75298 , n75297 , n31557 );
not ( n75299 , n31452 );
not ( n75300 , n31619 );
and ( n75301 , n75300 , n34107 );
xor ( n75302 , n34108 , n34127 );
and ( n75303 , n75302 , n31619 );
or ( n75304 , n75301 , n75303 );
and ( n75305 , n75299 , n75304 );
and ( n75306 , n34005 , n31452 );
or ( n75307 , n75305 , n75306 );
and ( n75308 , n75307 , n31638 );
buf ( n75309 , n33973 );
and ( n75310 , n34005 , n31650 );
or ( n75311 , C0 , n75263 , n75298 , n75308 , n75309 , n75310 );
buf ( n75312 , n75311 );
buf ( n75313 , n75312 );
buf ( n75314 , n31655 );
buf ( n75315 , n31655 );
buf ( n75316 , n31655 );
buf ( n75317 , n30987 );
not ( n75318 , n34150 );
and ( n75319 , n75318 , n32757 );
not ( n75320 , n56708 );
and ( n75321 , n75320 , n32757 );
and ( n75322 , n32789 , n56708 );
or ( n75323 , n75321 , n75322 );
and ( n75324 , n75323 , n34150 );
or ( n75325 , n75319 , n75324 );
and ( n75326 , n75325 , n33381 );
not ( n75327 , n56716 );
not ( n75328 , n56708 );
and ( n75329 , n75328 , n32757 );
and ( n75330 , n34301 , n56708 );
or ( n75331 , n75329 , n75330 );
and ( n75332 , n75327 , n75331 );
and ( n75333 , n34301 , n56716 );
or ( n75334 , n75332 , n75333 );
and ( n75335 , n75334 , n33375 );
not ( n75336 , n32968 );
not ( n75337 , n56716 );
not ( n75338 , n56708 );
and ( n75339 , n75338 , n32757 );
and ( n75340 , n34301 , n56708 );
or ( n75341 , n75339 , n75340 );
and ( n75342 , n75337 , n75341 );
and ( n75343 , n34301 , n56716 );
or ( n75344 , n75342 , n75343 );
and ( n75345 , n75336 , n75344 );
not ( n75346 , n56736 );
not ( n75347 , n56738 );
and ( n75348 , n75347 , n75344 );
and ( n75349 , n34761 , n56738 );
or ( n75350 , n75348 , n75349 );
and ( n75351 , n75346 , n75350 );
and ( n75352 , n35050 , n56736 );
or ( n75353 , n75351 , n75352 );
and ( n75354 , n75353 , n32968 );
or ( n75355 , n75345 , n75354 );
and ( n75356 , n75355 , n33370 );
and ( n75357 , n32757 , n35062 );
or ( n75358 , C0 , n75326 , n75335 , n75356 , n75357 );
buf ( n75359 , n75358 );
buf ( n75360 , n75359 );
buf ( n75361 , n30987 );
buf ( n75362 , n30987 );
buf ( n75363 , n31655 );
and ( n75364 , n31567 , n31007 );
not ( n75365 , n31077 );
and ( n75366 , n75365 , n35393 );
buf ( n75367 , n75366 );
and ( n75368 , n75367 , n31373 );
not ( n75369 , n31402 );
and ( n75370 , n75369 , n35393 );
buf ( n75371 , n75370 );
and ( n75372 , n75371 , n31408 );
not ( n75373 , n31437 );
and ( n75374 , n75373 , n35393 );
not ( n75375 , n31455 );
and ( n75376 , n75375 , n35435 );
xor ( n75377 , n35393 , n35405 );
and ( n75378 , n75377 , n31455 );
or ( n75379 , n75376 , n75378 );
and ( n75380 , n75379 , n31437 );
or ( n75381 , n75374 , n75380 );
and ( n75382 , n75381 , n31468 );
not ( n75383 , n31497 );
and ( n75384 , n75383 , n35393 );
not ( n75385 , n31454 );
not ( n75386 , n31501 );
and ( n75387 , n75386 , n35435 );
xor ( n75388 , n35436 , n35455 );
and ( n75389 , n75388 , n31501 );
or ( n75390 , n75387 , n75389 );
and ( n75391 , n75385 , n75390 );
and ( n75392 , n75377 , n31454 );
or ( n75393 , n75391 , n75392 );
and ( n75394 , n75393 , n31497 );
or ( n75395 , n75384 , n75394 );
and ( n75396 , n75395 , n31521 );
and ( n75397 , n35393 , n31553 );
or ( n75398 , n75368 , n75372 , n75382 , n75396 , n75397 );
and ( n75399 , n75398 , n31557 );
not ( n75400 , n31452 );
not ( n75401 , n31619 );
and ( n75402 , n75401 , n35490 );
xor ( n75403 , n35491 , n35509 );
and ( n75404 , n75403 , n31619 );
or ( n75405 , n75402 , n75404 );
and ( n75406 , n75400 , n75405 );
and ( n75407 , n35393 , n31452 );
or ( n75408 , n75406 , n75407 );
and ( n75409 , n75408 , n31638 );
and ( n75410 , n35393 , n31650 );
or ( n75411 , C0 , n75364 , n75399 , n75409 , C0 , n75410 );
buf ( n75412 , n75411 );
buf ( n75413 , n75412 );
not ( n75414 , n33419 );
and ( n75415 , n75414 , n31577 );
xor ( n75416 , n33471 , n33694 );
and ( n75417 , n75416 , n33419 );
or ( n75418 , n75415 , n75417 );
and ( n75419 , n75418 , n31529 );
not ( n75420 , n33734 );
and ( n75421 , n75420 , n31577 );
not ( n75422 , n33533 );
xor ( n75423 , n33764 , n33812 );
and ( n75424 , n75422 , n75423 );
xnor ( n75425 , n33849 , n33914 );
and ( n75426 , n75425 , n33533 );
or ( n75427 , n75424 , n75426 );
and ( n75428 , n75427 , n33734 );
or ( n75429 , n75421 , n75428 );
and ( n75430 , n75429 , n31527 );
and ( n75431 , n31577 , n33942 );
or ( n75432 , n75419 , n75430 , n75431 );
and ( n75433 , n75432 , n31557 );
and ( n75434 , n34099 , n31643 );
not ( n75435 , n31452 );
and ( n75436 , n75435 , n34099 );
xor ( n75437 , n31577 , n33960 );
and ( n75438 , n75437 , n31452 );
or ( n75439 , n75436 , n75438 );
and ( n75440 , n75439 , n31638 );
and ( n75441 , n34001 , n33973 );
and ( n75442 , n31577 , n33978 );
or ( n75443 , C0 , n75433 , n75434 , n75440 , n75441 , n75442 );
buf ( n75444 , n75443 );
buf ( n75445 , n75444 );
buf ( n75446 , n31655 );
buf ( n75447 , n30987 );
buf ( n75448 , n30987 );
buf ( n75449 , n30987 );
buf ( n75450 , n31655 );
and ( n75451 , n64914 , n33377 );
not ( n75452 , n48545 );
buf ( n75453 , RI15b47940_307);
and ( n75454 , n75452 , n75453 );
buf ( n75455 , n75454 );
and ( n75456 , n75455 , n32890 );
not ( n75457 , n48557 );
and ( n75458 , n75457 , n75453 );
and ( n75459 , n64920 , n48557 );
or ( n75460 , n75458 , n75459 );
and ( n75461 , n75460 , n33038 );
and ( n75462 , n75453 , n48571 );
or ( n75463 , n75456 , n75461 , n75462 );
and ( n75464 , n75463 , n33208 );
and ( n75465 , n75453 , n48577 );
or ( n75466 , C0 , n75451 , n75464 , n75465 );
buf ( n75467 , n75466 );
buf ( n75468 , n75467 );
buf ( n75469 , n31655 );
not ( n75470 , n33419 );
and ( n75471 , n75470 , n31628 );
and ( n75472 , n59182 , n33419 );
or ( n75473 , n75471 , n75472 );
and ( n75474 , n75473 , n31529 );
not ( n75475 , n33734 );
and ( n75476 , n75475 , n31628 );
and ( n75477 , n59193 , n33734 );
or ( n75478 , n75476 , n75477 );
and ( n75479 , n75478 , n31527 );
and ( n75480 , n31628 , n33942 );
or ( n75481 , n75474 , n75479 , n75480 );
and ( n75482 , n75481 , n31557 );
and ( n75483 , n31628 , n31643 );
buf ( n75484 , n31628 );
and ( n75485 , n75484 , n31638 );
and ( n75486 , n35687 , n33973 );
and ( n75487 , n31628 , n33978 );
or ( n75488 , C0 , n75482 , n75483 , n75485 , n75486 , n75487 );
buf ( n75489 , n75488 );
buf ( n75490 , n75489 );
not ( n75491 , n35542 );
and ( n75492 , n75491 , n41515 );
buf ( n75493 , RI15b45e10_249);
and ( n75494 , n75493 , n35542 );
or ( n75495 , n75492 , n75494 );
buf ( n75496 , n75495 );
buf ( n75497 , n75496 );
buf ( n75498 , n30987 );
buf ( n75499 , n30987 );
buf ( n75500 , n31655 );
not ( n75501 , n40163 );
and ( n75502 , n75501 , n32066 );
not ( n75503 , n40166 );
and ( n75504 , n75503 , n32066 );
and ( n75505 , n32130 , n40166 );
or ( n75506 , n75504 , n75505 );
and ( n75507 , n75506 , n40163 );
or ( n75508 , n75502 , n75507 );
and ( n75509 , n75508 , n32498 );
not ( n75510 , n40195 );
not ( n75511 , n40166 );
and ( n75512 , n75511 , n32066 );
and ( n75513 , n45833 , n40166 );
or ( n75514 , n75512 , n75513 );
and ( n75515 , n75510 , n75514 );
and ( n75516 , n45833 , n40195 );
or ( n75517 , n75515 , n75516 );
and ( n75518 , n75517 , n32473 );
not ( n75519 , n32475 );
not ( n75520 , n40195 );
not ( n75521 , n40166 );
and ( n75522 , n75521 , n32066 );
and ( n75523 , n45833 , n40166 );
or ( n75524 , n75522 , n75523 );
and ( n75525 , n75520 , n75524 );
and ( n75526 , n45833 , n40195 );
or ( n75527 , n75525 , n75526 );
and ( n75528 , n75519 , n75527 );
not ( n75529 , n40446 );
not ( n75530 , n40448 );
and ( n75531 , n75530 , n75527 );
and ( n75532 , n45857 , n40448 );
or ( n75533 , n75531 , n75532 );
and ( n75534 , n75529 , n75533 );
and ( n75535 , n45865 , n40446 );
or ( n75536 , n75534 , n75535 );
and ( n75537 , n75536 , n32475 );
or ( n75538 , n75528 , n75537 );
and ( n75539 , n75538 , n32486 );
and ( n75540 , n32066 , n41278 );
or ( n75541 , C0 , n75509 , n75518 , n75539 , n75540 );
buf ( n75542 , n75541 );
buf ( n75543 , n75542 );
not ( n75544 , n36587 );
and ( n75545 , n75544 , n36583 );
xor ( n75546 , n36583 , n36091 );
and ( n75547 , n61938 , n61947 );
xor ( n75548 , n75546 , n75547 );
and ( n75549 , n75548 , n36587 );
or ( n75550 , n75545 , n75549 );
and ( n75551 , n75550 , n36596 );
not ( n75552 , n37485 );
and ( n75553 , n75552 , n37481 );
xor ( n75554 , n37481 , n36993 );
and ( n75555 , n61954 , n61963 );
xor ( n75556 , n75554 , n75555 );
and ( n75557 , n75556 , n37485 );
or ( n75558 , n75553 , n75557 );
and ( n75559 , n75558 , n37494 );
and ( n75560 , n41515 , n37506 );
or ( n75561 , n75551 , n75559 , n75560 );
buf ( n75562 , n75561 );
buf ( n75563 , n75562 );
buf ( n75564 , n31655 );
buf ( n75565 , n30987 );
and ( n75566 , n47661 , n50275 );
not ( n75567 , n50278 );
and ( n75568 , n75567 , n47574 );
and ( n75569 , n47661 , n50278 );
or ( n75570 , n75568 , n75569 );
and ( n75571 , n75570 , n32421 );
not ( n75572 , n50002 );
and ( n75573 , n75572 , n47574 );
and ( n75574 , n47661 , n50002 );
or ( n75575 , n75573 , n75574 );
and ( n75576 , n75575 , n32419 );
not ( n75577 , n50289 );
and ( n75578 , n75577 , n47574 );
and ( n75579 , n47661 , n50289 );
or ( n75580 , n75578 , n75579 );
and ( n75581 , n75580 , n32417 );
not ( n75582 , n50008 );
and ( n75583 , n75582 , n47574 );
and ( n75584 , n47661 , n50008 );
or ( n75585 , n75583 , n75584 );
and ( n75586 , n75585 , n32415 );
not ( n75587 , n47331 );
and ( n75588 , n75587 , n47574 );
and ( n75589 , n47606 , n47331 );
or ( n75590 , n75588 , n75589 );
and ( n75591 , n75590 , n32413 );
not ( n75592 , n50067 );
and ( n75593 , n75592 , n47574 );
and ( n75594 , n47606 , n50067 );
or ( n75595 , n75593 , n75594 );
and ( n75596 , n75595 , n32411 );
not ( n75597 , n31728 );
and ( n75598 , n75597 , n47574 );
and ( n75599 , n51998 , n31728 );
or ( n75600 , n75598 , n75599 );
and ( n75601 , n75600 , n32253 );
not ( n75602 , n32283 );
and ( n75603 , n75602 , n47574 );
and ( n75604 , n52009 , n32283 );
or ( n75605 , n75603 , n75604 );
and ( n75606 , n75605 , n32398 );
and ( n75607 , n47711 , n50334 );
or ( n75608 , n75566 , n75571 , n75576 , n75581 , n75586 , n75591 , n75596 , n75601 , n75606 , n75607 );
and ( n75609 , n75608 , n32456 );
and ( n75610 , n37555 , n32489 );
and ( n75611 , n47574 , n50345 );
or ( n75612 , C0 , n75609 , n75610 , n75611 );
buf ( n75613 , n75612 );
buf ( n75614 , n75613 );
buf ( n75615 , n31655 );
and ( n75616 , n33236 , n32528 );
not ( n75617 , n32598 );
and ( n75618 , n75617 , n32999 );
and ( n75619 , n32531 , n45916 );
and ( n75620 , n75619 , n32598 );
or ( n75621 , n75618 , n75620 );
and ( n75622 , n75621 , n32890 );
not ( n75623 , n32919 );
and ( n75624 , n75623 , n32999 );
and ( n75625 , n75619 , n32919 );
or ( n75626 , n75624 , n75625 );
and ( n75627 , n75626 , n32924 );
not ( n75628 , n32953 );
and ( n75629 , n75628 , n32999 );
not ( n75630 , n32971 );
and ( n75631 , n75630 , n33123 );
xor ( n75632 , n32999 , n33006 );
and ( n75633 , n75632 , n32971 );
or ( n75634 , n75631 , n75633 );
and ( n75635 , n75634 , n32953 );
or ( n75636 , n75629 , n75635 );
and ( n75637 , n75636 , n33038 );
not ( n75638 , n33067 );
and ( n75639 , n75638 , n32999 );
not ( n75640 , n32970 );
not ( n75641 , n33071 );
and ( n75642 , n75641 , n33123 );
xor ( n75643 , n33124 , n33138 );
and ( n75644 , n75643 , n33071 );
or ( n75645 , n75642 , n75644 );
and ( n75646 , n75640 , n75645 );
and ( n75647 , n75632 , n32970 );
or ( n75648 , n75646 , n75647 );
and ( n75649 , n75648 , n33067 );
or ( n75650 , n75639 , n75649 );
and ( n75651 , n75650 , n33172 );
and ( n75652 , n32999 , n33204 );
or ( n75653 , n75622 , n75627 , n75637 , n75651 , n75652 );
and ( n75654 , n75653 , n33208 );
not ( n75655 , n32968 );
not ( n75656 , n33270 );
and ( n75657 , n75656 , n33323 );
xor ( n75658 , n33324 , n33338 );
and ( n75659 , n75658 , n33270 );
or ( n75660 , n75657 , n75659 );
and ( n75661 , n75655 , n75660 );
and ( n75662 , n32999 , n32968 );
or ( n75663 , n75661 , n75662 );
and ( n75664 , n75663 , n33370 );
buf ( n75665 , n35056 );
and ( n75666 , n32999 , n33382 );
or ( n75667 , C0 , n75616 , n75654 , n75664 , n75665 , n75666 );
buf ( n75668 , n75667 );
buf ( n75669 , n75668 );
buf ( n75670 , n30987 );
buf ( n75671 , n30987 );
and ( n75672 , n32464 , n32500 );
not ( n75673 , n35211 );
and ( n75674 , n75673 , n37514 );
and ( n75675 , n31756 , n35211 );
or ( n75676 , n75674 , n75675 );
and ( n75677 , n75676 , n32421 );
not ( n75678 , n35245 );
and ( n75679 , n75678 , n37514 );
and ( n75680 , n31756 , n35245 );
or ( n75681 , n75679 , n75680 );
and ( n75682 , n75681 , n32419 );
not ( n75683 , n35278 );
and ( n75684 , n75683 , n37514 );
not ( n75685 , n35295 );
and ( n75686 , n75685 , n45999 );
not ( n75687 , n37514 );
and ( n75688 , n75687 , n35295 );
or ( n75689 , n75686 , n75688 );
and ( n75690 , n75689 , n35278 );
or ( n75691 , n75684 , n75690 );
and ( n75692 , n75691 , n32417 );
not ( n75693 , n35331 );
and ( n75694 , n75693 , n37514 );
not ( n75695 , n35294 );
not ( n75696 , n45995 );
and ( n75697 , n75696 , n45999 );
xor ( n75698 , n46000 , n46001 );
and ( n75699 , n75698 , n45995 );
or ( n75700 , n75697 , n75699 );
and ( n75701 , n75695 , n75700 );
and ( n75702 , n75687 , n35294 );
or ( n75703 , n75701 , n75702 );
and ( n75704 , n75703 , n35331 );
or ( n75705 , n75694 , n75704 );
and ( n75706 , n75705 , n32415 );
and ( n75707 , n37514 , n35354 );
or ( n75708 , n75677 , n75682 , n75692 , n75706 , n75707 );
and ( n75709 , n75708 , n32456 );
not ( n75710 , n32475 );
not ( n75711 , n46060 );
and ( n75712 , n75711 , n46065 );
xor ( n75713 , n46066 , n46067 );
and ( n75714 , n75713 , n46060 );
or ( n75715 , n75712 , n75714 );
and ( n75716 , n75710 , n75715 );
and ( n75717 , n37514 , n32475 );
or ( n75718 , n75716 , n75717 );
and ( n75719 , n75718 , n32486 );
and ( n75720 , n37514 , n35367 );
or ( n75721 , C0 , n75672 , n75709 , n75719 , C0 , n75720 );
buf ( n75722 , n75721 );
buf ( n75723 , n75722 );
buf ( n75724 , n31655 );
buf ( n75725 , n31655 );
buf ( n75726 , n31655 );
and ( n75727 , n57416 , n32494 );
not ( n75728 , n46083 );
buf ( n75729 , RI15b5fa90_1129);
and ( n75730 , n75728 , n75729 );
not ( n75731 , n46290 );
and ( n75732 , n75731 , n46169 );
xor ( n75733 , n46300 , n46312 );
and ( n75734 , n75733 , n46290 );
or ( n75735 , n75732 , n75734 );
and ( n75736 , n75735 , n46083 );
or ( n75737 , n75730 , n75736 );
and ( n75738 , n75737 , n32421 );
not ( n75739 , n46326 );
and ( n75740 , n75739 , n75729 );
and ( n75741 , n75735 , n46326 );
or ( n75742 , n75740 , n75741 );
and ( n75743 , n75742 , n32417 );
and ( n75744 , n75729 , n46340 );
or ( n75745 , n75738 , n75743 , n75744 );
and ( n75746 , n75745 , n32456 );
and ( n75747 , n75729 , n46349 );
or ( n75748 , C0 , n75727 , n75746 , n75747 );
buf ( n75749 , n75748 );
buf ( n75750 , n75749 );
buf ( n75751 , n30987 );
not ( n75752 , n46356 );
and ( n75753 , n75752 , n31094 );
not ( n75754 , n55473 );
and ( n75755 , n75754 , n31094 );
and ( n75756 , n31138 , n55473 );
or ( n75757 , n75755 , n75756 );
and ( n75758 , n75757 , n46356 );
or ( n75759 , n75753 , n75758 );
and ( n75760 , n75759 , n31649 );
not ( n75761 , n55481 );
not ( n75762 , n55473 );
and ( n75763 , n75762 , n31094 );
and ( n75764 , n56920 , n55473 );
or ( n75765 , n75763 , n75764 );
and ( n75766 , n75761 , n75765 );
and ( n75767 , n56920 , n55481 );
or ( n75768 , n75766 , n75767 );
and ( n75769 , n75768 , n31643 );
not ( n75770 , n31452 );
not ( n75771 , n55481 );
not ( n75772 , n55473 );
and ( n75773 , n75772 , n31094 );
and ( n75774 , n56920 , n55473 );
or ( n75775 , n75773 , n75774 );
and ( n75776 , n75771 , n75775 );
and ( n75777 , n56920 , n55481 );
or ( n75778 , n75776 , n75777 );
and ( n75779 , n75770 , n75778 );
not ( n75780 , n55501 );
not ( n75781 , n55503 );
and ( n75782 , n75781 , n75778 );
and ( n75783 , n56946 , n55503 );
or ( n75784 , n75782 , n75783 );
and ( n75785 , n75780 , n75784 );
and ( n75786 , n56954 , n55501 );
or ( n75787 , n75785 , n75786 );
and ( n75788 , n75787 , n31452 );
or ( n75789 , n75779 , n75788 );
and ( n75790 , n75789 , n31638 );
and ( n75791 , n31094 , n47277 );
or ( n75792 , C0 , n75760 , n75769 , n75790 , n75791 );
buf ( n75793 , n75792 );
buf ( n75794 , n75793 );
buf ( n75795 , RI15b54348_738);
and ( n75796 , n75795 , n58921 );
and ( n75797 , n41520 , n37506 );
or ( n75798 , n75796 , n75797 );
buf ( n75799 , n75798 );
buf ( n75800 , n75799 );
and ( n75801 , n47664 , n50275 );
not ( n75802 , n50278 );
and ( n75803 , n75802 , n47577 );
and ( n75804 , n47664 , n50278 );
or ( n75805 , n75803 , n75804 );
and ( n75806 , n75805 , n32421 );
not ( n75807 , n50002 );
and ( n75808 , n75807 , n47577 );
and ( n75809 , n47664 , n50002 );
or ( n75810 , n75808 , n75809 );
and ( n75811 , n75810 , n32419 );
not ( n75812 , n50289 );
and ( n75813 , n75812 , n47577 );
and ( n75814 , n47664 , n50289 );
or ( n75815 , n75813 , n75814 );
and ( n75816 , n75815 , n32417 );
not ( n75817 , n50008 );
and ( n75818 , n75817 , n47577 );
and ( n75819 , n47664 , n50008 );
or ( n75820 , n75818 , n75819 );
and ( n75821 , n75820 , n32415 );
not ( n75822 , n47331 );
and ( n75823 , n75822 , n47577 );
and ( n75824 , n47609 , n47331 );
or ( n75825 , n75823 , n75824 );
and ( n75826 , n75825 , n32413 );
not ( n75827 , n50067 );
and ( n75828 , n75827 , n47577 );
and ( n75829 , n47609 , n50067 );
or ( n75830 , n75828 , n75829 );
and ( n75831 , n75830 , n32411 );
not ( n75832 , n31728 );
and ( n75833 , n75832 , n47577 );
xor ( n75834 , n47609 , n47620 );
and ( n75835 , n75834 , n31728 );
or ( n75836 , n75833 , n75835 );
and ( n75837 , n75836 , n32253 );
not ( n75838 , n32283 );
and ( n75839 , n75838 , n47577 );
not ( n75840 , n31823 );
xor ( n75841 , n47664 , n47675 );
and ( n75842 , n75840 , n75841 );
xnor ( n75843 , n47714 , n47725 );
and ( n75844 , n75843 , n31823 );
or ( n75845 , n75842 , n75844 );
and ( n75846 , n75845 , n32283 );
or ( n75847 , n75839 , n75846 );
and ( n75848 , n75847 , n32398 );
and ( n75849 , n47714 , n50334 );
or ( n75850 , n75801 , n75806 , n75811 , n75816 , n75821 , n75826 , n75831 , n75837 , n75848 , n75849 );
and ( n75851 , n75850 , n32456 );
and ( n75852 , n37561 , n32489 );
and ( n75853 , n47577 , n50345 );
or ( n75854 , C0 , n75851 , n75852 , n75853 );
buf ( n75855 , n75854 );
buf ( n75856 , n75855 );
buf ( n75857 , n31655 );
buf ( n75858 , n30987 );
not ( n75859 , n43755 );
and ( n75860 , n75859 , n43326 );
xor ( n75861 , n43760 , n43768 );
and ( n75862 , n75861 , n43755 );
or ( n75863 , n75860 , n75862 );
and ( n75864 , n75863 , n43774 );
not ( n75865 , n44663 );
and ( n75866 , n75865 , n44238 );
xor ( n75867 , n44668 , n44676 );
and ( n75868 , n75867 , n44663 );
or ( n75869 , n75866 , n75868 );
and ( n75870 , n75869 , n44682 );
and ( n75871 , n72666 , n44695 );
or ( n75872 , n75864 , n75870 , n75871 );
buf ( n75873 , n75872 );
buf ( n75874 , n75873 );
buf ( n75875 , n30987 );
buf ( n75876 , n31655 );
buf ( n75877 , n31655 );
buf ( n75878 , n30987 );
buf ( n75879 , RI15b60a08_1162);
and ( n75880 , n75879 , n48531 );
and ( n75881 , n50825 , n39359 );
or ( n75882 , n75880 , n75881 );
buf ( n75883 , n75882 );
buf ( n75884 , n75883 );
buf ( n75885 , n31655 );
not ( n75886 , n36587 );
and ( n75887 , n75886 , n36141 );
xor ( n75888 , n50192 , n50195 );
and ( n75889 , n75888 , n36587 );
or ( n75890 , n75887 , n75889 );
and ( n75891 , n75890 , n36596 );
not ( n75892 , n37485 );
and ( n75893 , n75892 , n37043 );
xor ( n75894 , n50242 , n50245 );
and ( n75895 , n75894 , n37485 );
or ( n75896 , n75893 , n75895 );
and ( n75897 , n75896 , n37494 );
and ( n75898 , n41842 , n37506 );
or ( n75899 , n75891 , n75897 , n75898 );
buf ( n75900 , n75899 );
buf ( n75901 , n75900 );
buf ( n75902 , n30987 );
not ( n75903 , n40163 );
and ( n75904 , n75903 , n31854 );
nor ( n75905 , n42169 , n31669 , n31665 , n31661 , n31657 );
not ( n75906 , n75905 );
and ( n75907 , n75906 , n31854 );
and ( n75908 , n32235 , n75905 );
or ( n75909 , n75907 , n75908 );
and ( n75910 , n75909 , n40163 );
or ( n75911 , n75904 , n75910 );
and ( n75912 , n75911 , n32498 );
nor ( n75913 , n42179 , n40182 , n40188 , n40194 , C0 );
not ( n75914 , n75913 );
not ( n75915 , n75905 );
and ( n75916 , n75915 , n31854 );
and ( n75917 , n42188 , n75905 );
or ( n75918 , n75916 , n75917 );
and ( n75919 , n75914 , n75918 );
and ( n75920 , n42188 , n75913 );
or ( n75921 , n75919 , n75920 );
and ( n75922 , n75921 , n32473 );
not ( n75923 , n32475 );
not ( n75924 , n75913 );
not ( n75925 , n75905 );
and ( n75926 , n75925 , n31854 );
and ( n75927 , n42188 , n75905 );
or ( n75928 , n75926 , n75927 );
and ( n75929 , n75924 , n75928 );
and ( n75930 , n42188 , n75913 );
or ( n75931 , n75929 , n75930 );
and ( n75932 , n75923 , n75931 );
nor ( n75933 , n42205 , n40425 , n40435 , n40445 , C0 );
not ( n75934 , n75933 );
nor ( n75935 , n42208 , n40421 , n40430 , n40440 , C0 );
not ( n75936 , n75935 );
and ( n75937 , n75936 , n75931 );
and ( n75938 , n42216 , n75935 );
or ( n75939 , n75937 , n75938 );
and ( n75940 , n75934 , n75939 );
and ( n75941 , n42224 , n75933 );
or ( n75942 , n75940 , n75941 );
and ( n75943 , n75942 , n32475 );
or ( n75944 , n75932 , n75943 );
and ( n75945 , n75944 , n32486 );
and ( n75946 , n31854 , n41278 );
or ( n75947 , C0 , n75912 , n75922 , n75945 , n75946 );
buf ( n75948 , n75947 );
buf ( n75949 , n75948 );
xor ( n75950 , n35447 , n39940 );
and ( n75951 , n75950 , n31550 );
not ( n75952 , n39979 );
and ( n75953 , n75952 , n35447 );
and ( n75954 , n31173 , n40095 );
and ( n75955 , n31175 , n40097 );
and ( n75956 , n31177 , n40099 );
and ( n75957 , n31179 , n40101 );
and ( n75958 , n31181 , n40103 );
and ( n75959 , n31183 , n40105 );
and ( n75960 , n31185 , n40107 );
and ( n75961 , n31187 , n40109 );
and ( n75962 , n31189 , n40111 );
and ( n75963 , n31191 , n40113 );
and ( n75964 , n31193 , n40115 );
and ( n75965 , n31195 , n40117 );
and ( n75966 , n31197 , n40119 );
and ( n75967 , n31199 , n40121 );
and ( n75968 , n31201 , n40123 );
and ( n75969 , n31203 , n40125 );
or ( n75970 , n75954 , n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , n75969 );
and ( n75971 , n75970 , n39979 );
or ( n75972 , n75953 , n75971 );
and ( n75973 , n75972 , n31538 );
and ( n75974 , n35447 , n40143 );
or ( n75975 , n75951 , n75973 , n75974 );
and ( n75976 , n75975 , n31557 );
and ( n75977 , n35447 , n40154 );
or ( n75978 , C0 , n75976 , n75977 );
buf ( n75979 , n75978 );
buf ( n75980 , n75979 );
buf ( n75981 , n31655 );
buf ( n75982 , n70838 );
buf ( n75983 , n30987 );
buf ( n75984 , n30987 );
and ( n75985 , n59412 , n48455 );
not ( n75986 , n48457 );
and ( n75987 , n75986 , n52396 );
and ( n75988 , n59412 , n48457 );
or ( n75989 , n75987 , n75988 );
and ( n75990 , n75989 , n31373 );
not ( n75991 , n44807 );
and ( n75992 , n75991 , n52396 );
and ( n75993 , n59412 , n44807 );
or ( n75994 , n75992 , n75993 );
and ( n75995 , n75994 , n31408 );
not ( n75996 , n48468 );
and ( n75997 , n75996 , n52396 );
and ( n75998 , n59412 , n48468 );
or ( n75999 , n75997 , n75998 );
and ( n76000 , n75999 , n31468 );
not ( n76001 , n44817 );
and ( n76002 , n76001 , n52396 );
and ( n76003 , n59412 , n44817 );
or ( n76004 , n76002 , n76003 );
and ( n76005 , n76004 , n31521 );
not ( n76006 , n39979 );
and ( n76007 , n76006 , n52396 );
and ( n76008 , n59399 , n39979 );
or ( n76009 , n76007 , n76008 );
and ( n76010 , n76009 , n31538 );
not ( n76011 , n45059 );
and ( n76012 , n76011 , n52396 );
and ( n76013 , n59399 , n45059 );
or ( n76014 , n76012 , n76013 );
and ( n76015 , n76014 , n31536 );
not ( n76016 , n33419 );
and ( n76017 , n76016 , n52396 );
and ( n76018 , n64224 , n33419 );
or ( n76019 , n76017 , n76018 );
and ( n76020 , n76019 , n31529 );
not ( n76021 , n33734 );
and ( n76022 , n76021 , n52396 );
and ( n76023 , n64235 , n33734 );
or ( n76024 , n76022 , n76023 );
and ( n76025 , n76024 , n31527 );
and ( n76026 , n59420 , n48513 );
or ( n76027 , n75985 , n75990 , n75995 , n76000 , n76005 , n76010 , n76015 , n76020 , n76025 , n76026 );
and ( n76028 , n76027 , n31557 );
and ( n76029 , n35387 , n33973 );
and ( n76030 , n52396 , n48524 );
or ( n76031 , C0 , n76028 , n76029 , n76030 );
buf ( n76032 , n76031 );
buf ( n76033 , n76032 );
not ( n76034 , n38443 );
and ( n76035 , n76034 , n38235 );
xor ( n76036 , n53468 , n53501 );
and ( n76037 , n76036 , n38443 );
or ( n76038 , n76035 , n76037 );
and ( n76039 , n76038 , n38450 );
not ( n76040 , n39339 );
and ( n76041 , n76040 , n39135 );
xor ( n76042 , n53524 , n53557 );
and ( n76043 , n76042 , n39339 );
or ( n76044 , n76041 , n76043 );
and ( n76045 , n76044 , n39346 );
and ( n76046 , n40216 , n39359 );
or ( n76047 , n76039 , n76045 , n76046 );
buf ( n76048 , n76047 );
buf ( n76049 , n76048 );
buf ( n76050 , n30987 );
buf ( n76051 , n31655 );
not ( n76052 , n40163 );
and ( n76053 , n76052 , n31949 );
not ( n76054 , n49298 );
and ( n76055 , n76054 , n31949 );
and ( n76056 , n32183 , n49298 );
or ( n76057 , n76055 , n76056 );
and ( n76058 , n76057 , n40163 );
or ( n76059 , n76053 , n76058 );
and ( n76060 , n76059 , n32498 );
not ( n76061 , n49306 );
not ( n76062 , n49298 );
and ( n76063 , n76062 , n31949 );
and ( n76064 , n45178 , n49298 );
or ( n76065 , n76063 , n76064 );
and ( n76066 , n76061 , n76065 );
and ( n76067 , n45178 , n49306 );
or ( n76068 , n76066 , n76067 );
and ( n76069 , n76068 , n32473 );
not ( n76070 , n32475 );
not ( n76071 , n49306 );
not ( n76072 , n49298 );
and ( n76073 , n76072 , n31949 );
and ( n76074 , n45178 , n49298 );
or ( n76075 , n76073 , n76074 );
and ( n76076 , n76071 , n76075 );
and ( n76077 , n45178 , n49306 );
or ( n76078 , n76076 , n76077 );
and ( n76079 , n76070 , n76078 );
not ( n76080 , n49331 );
not ( n76081 , n49333 );
and ( n76082 , n76081 , n76078 );
and ( n76083 , n45206 , n49333 );
or ( n76084 , n76082 , n76083 );
and ( n76085 , n76080 , n76084 );
and ( n76086 , n45214 , n49331 );
or ( n76087 , n76085 , n76086 );
and ( n76088 , n76087 , n32475 );
or ( n76089 , n76079 , n76088 );
and ( n76090 , n76089 , n32486 );
and ( n76091 , n31949 , n41278 );
or ( n76092 , C0 , n76060 , n76069 , n76090 , n76091 );
buf ( n76093 , n76092 );
buf ( n76094 , n76093 );
buf ( n76095 , n30987 );
buf ( n76096 , n30987 );
xor ( n76097 , n41769 , n44788 );
and ( n76098 , n76097 , n31548 );
not ( n76099 , n44807 );
and ( n76100 , n76099 , n41769 );
and ( n76101 , n42078 , n44807 );
or ( n76102 , n76100 , n76101 );
and ( n76103 , n76102 , n31408 );
not ( n76104 , n44817 );
and ( n76105 , n76104 , n41769 );
not ( n76106 , n41835 );
buf ( n76107 , RI15b531f0_701);
and ( n76108 , n76106 , n76107 );
not ( n76109 , n42124 );
and ( n76110 , n76109 , n42088 );
xor ( n76111 , n49375 , n49384 );
and ( n76112 , n76111 , n42124 );
or ( n76113 , n76110 , n76112 );
and ( n76114 , n76113 , n41835 );
or ( n76115 , n76108 , n76114 );
and ( n76116 , n76115 , n44817 );
or ( n76117 , n76105 , n76116 );
and ( n76118 , n76117 , n31521 );
not ( n76119 , n45059 );
and ( n76120 , n76119 , n41769 );
and ( n76121 , n31274 , n42330 );
and ( n76122 , n31276 , n42332 );
and ( n76123 , n31278 , n42334 );
and ( n76124 , n31280 , n42336 );
and ( n76125 , n31282 , n42338 );
and ( n76126 , n31284 , n42340 );
and ( n76127 , n31286 , n42342 );
and ( n76128 , n31288 , n42344 );
and ( n76129 , n31290 , n42346 );
and ( n76130 , n31292 , n42348 );
and ( n76131 , n31294 , n42350 );
and ( n76132 , n31296 , n42352 );
and ( n76133 , n31298 , n42354 );
and ( n76134 , n31300 , n42356 );
and ( n76135 , n31302 , n42358 );
and ( n76136 , n31304 , n42360 );
or ( n76137 , n76121 , n76122 , n76123 , n76124 , n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , n76135 , n76136 );
and ( n76138 , n76137 , n45059 );
or ( n76139 , n76120 , n76138 );
and ( n76140 , n76139 , n31536 );
and ( n76141 , n41769 , n45148 );
or ( n76142 , n76098 , n76103 , n76118 , n76140 , n76141 );
and ( n76143 , n76142 , n31557 );
and ( n76144 , n41769 , n40154 );
or ( n76145 , C0 , n76143 , n76144 );
buf ( n76146 , n76145 );
buf ( n76147 , n76146 );
buf ( n76148 , n31655 );
not ( n76149 , n40163 );
and ( n76150 , n76149 , n32498 );
not ( n76151 , n55780 );
and ( n76152 , n76151 , n32496 );
not ( n76153 , n35292 );
and ( n76154 , n76153 , n32439 );
buf ( n76155 , n35292 );
or ( n76156 , n76154 , n76155 );
and ( n76157 , n76156 , n32494 );
not ( n76158 , n69188 );
and ( n76159 , n76158 , n31657 );
not ( n76160 , n66481 );
and ( n76161 , n76160 , n31661 );
not ( n76162 , n64637 );
and ( n76163 , n76162 , n31665 );
not ( n76164 , n63981 );
and ( n76165 , n76164 , n31669 );
not ( n76166 , n64375 );
and ( n76167 , n76166 , n31673 );
xnor ( n76168 , n63981 , n31669 );
and ( n76169 , n76167 , n76168 );
or ( n76170 , n76165 , n76169 );
xnor ( n76171 , n64637 , n31665 );
and ( n76172 , n76170 , n76171 );
or ( n76173 , n76163 , n76172 );
xnor ( n76174 , n66481 , n31661 );
and ( n76175 , n76173 , n76174 );
or ( n76176 , n76161 , n76175 );
xnor ( n76177 , n69188 , n31657 );
and ( n76178 , n76176 , n76177 );
or ( n76179 , n76159 , n76178 );
not ( n76180 , n76179 );
not ( n76181 , n69188 );
not ( n76182 , n66481 );
buf ( n76183 , n69188 );
buf ( n76184 , n69188 );
buf ( n76185 , n69188 );
buf ( n76186 , n69188 );
buf ( n76187 , n69188 );
buf ( n76188 , n69188 );
buf ( n76189 , n69188 );
buf ( n76190 , n69188 );
buf ( n76191 , n69188 );
buf ( n76192 , n69188 );
buf ( n76193 , n69188 );
buf ( n76194 , n69188 );
buf ( n76195 , n69188 );
buf ( n76196 , n69188 );
buf ( n76197 , n69188 );
buf ( n76198 , n69188 );
buf ( n76199 , n69188 );
buf ( n76200 , n69188 );
buf ( n76201 , n69188 );
buf ( n76202 , n69188 );
buf ( n76203 , n69188 );
buf ( n76204 , n69188 );
buf ( n76205 , n69188 );
buf ( n76206 , n69188 );
buf ( n76207 , n69188 );
buf ( n76208 , n69188 );
not ( n76209 , n64637 );
or ( n76210 , n76182 , n69188 , n76183 , n76184 , n76185 , n76186 , n76187 , n76188 , n76189 , n76190 , n76191 , n76192 , n76193 , n76194 , n76195 , n76196 , n76197 , n76198 , n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , n76205 , n76206 , n76207 , n76208 , n76209 );
nand ( n76211 , n76181 , n76210 );
not ( n76212 , n50277 );
and ( n76213 , n35211 , n76212 );
and ( n76214 , n55558 , n76213 );
and ( n76215 , n76214 , n32421 );
and ( n76216 , n35245 , n35291 );
and ( n76217 , n55558 , n76216 );
and ( n76218 , n76217 , n32419 );
and ( n76219 , n35278 , n76212 );
and ( n76220 , n55558 , n76219 );
and ( n76221 , n76220 , n32417 );
and ( n76222 , n35331 , n35291 );
and ( n76223 , n55558 , n76222 );
and ( n76224 , n76223 , n32415 );
and ( n76225 , n31728 , n32253 );
and ( n76226 , n32283 , n32398 );
or ( n76227 , n76215 , n76218 , n76221 , n76224 , n76225 , n76226 , C0 );
or ( n76228 , n76211 , n76227 );
or ( n76229 , n76228 , n72237 );
or ( n76230 , n76180 , n76229 );
not ( n76231 , n76230 );
and ( n76232 , n35278 , n35295 );
not ( n76233 , n76232 );
and ( n76234 , n76233 , n32439 );
buf ( n76235 , n76234 );
and ( n76236 , n76235 , n32417 );
or ( n76237 , n46333 , n32421 );
or ( n76238 , n76237 , n32423 );
or ( n76239 , n76238 , n32425 );
or ( n76240 , n76239 , n32427 );
or ( n76241 , n76240 , n32429 );
or ( n76242 , n76241 , n32431 );
or ( n76243 , n76242 , n32433 );
or ( n76244 , n76243 , n32435 );
and ( n76245 , n32439 , n76244 );
or ( n76246 , n76236 , n76245 );
and ( n76247 , n76231 , n76246 );
buf ( n76248 , n76230 );
or ( n76249 , n76247 , n76248 );
and ( n76250 , n76249 , n32456 );
buf ( n76251 , n32473 );
not ( n76252 , n35292 );
and ( n76253 , n76252 , n32492 );
buf ( n76254 , n32486 );
and ( n76255 , n76252 , n32491 );
or ( n76256 , n32489 , n32500 );
buf ( n76257 , n76256 );
or ( n76258 , C0 , n76150 , n76152 , n76157 , n76250 , n76251 , n76253 , n76254 , n76255 , n76257 );
buf ( n76259 , n76258 );
buf ( n76260 , n76259 );
buf ( n76261 , n31655 );
not ( n76262 , n36587 );
and ( n76263 , n76262 , n36243 );
xor ( n76264 , n50186 , n50201 );
and ( n76265 , n76264 , n36587 );
or ( n76266 , n76263 , n76265 );
and ( n76267 , n76266 , n36596 );
not ( n76268 , n37485 );
and ( n76269 , n76268 , n37145 );
xor ( n76270 , n50236 , n50251 );
and ( n76271 , n76270 , n37485 );
or ( n76272 , n76269 , n76271 );
and ( n76273 , n76272 , n37494 );
and ( n76274 , n41848 , n37506 );
or ( n76275 , n76267 , n76273 , n76274 );
buf ( n76276 , n76275 );
buf ( n76277 , n76276 );
buf ( n76278 , n30987 );
and ( n76279 , n33759 , n48455 );
not ( n76280 , n48457 );
and ( n76281 , n76280 , n33424 );
and ( n76282 , n33759 , n48457 );
or ( n76283 , n76281 , n76282 );
and ( n76284 , n76283 , n31373 );
not ( n76285 , n44807 );
and ( n76286 , n76285 , n33424 );
and ( n76287 , n33759 , n44807 );
or ( n76288 , n76286 , n76287 );
and ( n76289 , n76288 , n31408 );
not ( n76290 , n48468 );
and ( n76291 , n76290 , n33424 );
and ( n76292 , n33759 , n48468 );
or ( n76293 , n76291 , n76292 );
and ( n76294 , n76293 , n31468 );
not ( n76295 , n44817 );
and ( n76296 , n76295 , n33424 );
and ( n76297 , n33759 , n44817 );
or ( n76298 , n76296 , n76297 );
and ( n76299 , n76298 , n31521 );
not ( n76300 , n39979 );
and ( n76301 , n76300 , n33424 );
and ( n76302 , n33466 , n39979 );
or ( n76303 , n76301 , n76302 );
and ( n76304 , n76303 , n31538 );
not ( n76305 , n45059 );
and ( n76306 , n76305 , n33424 );
and ( n76307 , n33466 , n45059 );
or ( n76308 , n76306 , n76307 );
and ( n76309 , n76308 , n31536 );
not ( n76310 , n33419 );
and ( n76311 , n76310 , n33424 );
xor ( n76312 , n33466 , n33699 );
and ( n76313 , n76312 , n33419 );
or ( n76314 , n76311 , n76313 );
and ( n76315 , n76314 , n31529 );
not ( n76316 , n33734 );
and ( n76317 , n76316 , n33424 );
not ( n76318 , n33533 );
xor ( n76319 , n33759 , n33817 );
and ( n76320 , n76318 , n76319 );
xnor ( n76321 , n33844 , n33919 );
and ( n76322 , n76321 , n33533 );
or ( n76323 , n76320 , n76322 );
and ( n76324 , n76323 , n33734 );
or ( n76325 , n76317 , n76324 );
and ( n76326 , n76325 , n31527 );
and ( n76327 , n33844 , n48513 );
or ( n76328 , n76279 , n76284 , n76289 , n76294 , n76299 , n76304 , n76309 , n76315 , n76326 , n76327 );
and ( n76329 , n76328 , n31557 );
and ( n76330 , n35397 , n33973 );
and ( n76331 , n33424 , n48524 );
or ( n76332 , C0 , n76329 , n76330 , n76331 );
buf ( n76333 , n76332 );
buf ( n76334 , n76333 );
buf ( n76335 , n31655 );
buf ( n76336 , n30987 );
not ( n76337 , n38443 );
and ( n76338 , n76337 , n38422 );
xor ( n76339 , n69916 , n69921 );
and ( n76340 , n76339 , n38443 );
or ( n76341 , n76338 , n76340 );
and ( n76342 , n76341 , n38450 );
not ( n76343 , n39339 );
and ( n76344 , n76343 , n39322 );
xor ( n76345 , n69930 , n69935 );
and ( n76346 , n76345 , n39339 );
or ( n76347 , n76344 , n76346 );
and ( n76348 , n76347 , n39346 );
and ( n76349 , n40226 , n39359 );
or ( n76350 , n76342 , n76348 , n76349 );
buf ( n76351 , n76350 );
buf ( n76352 , n76351 );
and ( n76353 , n33234 , n32528 );
not ( n76354 , n32598 );
and ( n76355 , n76354 , n32997 );
buf ( n76356 , n76355 );
and ( n76357 , n76356 , n32890 );
not ( n76358 , n32919 );
and ( n76359 , n76358 , n32997 );
buf ( n76360 , n76359 );
and ( n76361 , n76360 , n32924 );
not ( n76362 , n32953 );
and ( n76363 , n76362 , n32997 );
not ( n76364 , n32971 );
and ( n76365 , n76364 , n33119 );
xor ( n76366 , n32997 , n33008 );
and ( n76367 , n76366 , n32971 );
or ( n76368 , n76365 , n76367 );
and ( n76369 , n76368 , n32953 );
or ( n76370 , n76363 , n76369 );
and ( n76371 , n76370 , n33038 );
not ( n76372 , n33067 );
and ( n76373 , n76372 , n32997 );
not ( n76374 , n32970 );
not ( n76375 , n33071 );
and ( n76376 , n76375 , n33119 );
xor ( n76377 , n33120 , n33140 );
and ( n76378 , n76377 , n33071 );
or ( n76379 , n76376 , n76378 );
and ( n76380 , n76374 , n76379 );
and ( n76381 , n76366 , n32970 );
or ( n76382 , n76380 , n76381 );
and ( n76383 , n76382 , n33067 );
or ( n76384 , n76373 , n76383 );
and ( n76385 , n76384 , n33172 );
and ( n76386 , n32997 , n33204 );
or ( n76387 , n76357 , n76361 , n76371 , n76385 , n76386 );
and ( n76388 , n76387 , n33208 );
not ( n76389 , n32968 );
not ( n76390 , n33270 );
and ( n76391 , n76390 , n33319 );
xor ( n76392 , n33320 , n33340 );
and ( n76393 , n76392 , n33270 );
or ( n76394 , n76391 , n76393 );
and ( n76395 , n76389 , n76394 );
and ( n76396 , n32997 , n32968 );
or ( n76397 , n76395 , n76396 );
and ( n76398 , n76397 , n33370 );
buf ( n76399 , n35056 );
and ( n76400 , n32997 , n33382 );
or ( n76401 , C0 , n76353 , n76388 , n76398 , n76399 , n76400 );
buf ( n76402 , n76401 );
buf ( n76403 , n76402 );
buf ( n76404 , n31655 );
buf ( n76405 , n30987 );
buf ( n76406 , n30987 );
buf ( n76407 , n31655 );
not ( n76408 , n31728 );
and ( n76409 , n76408 , n46016 );
and ( n76410 , n65870 , n31728 );
or ( n76411 , n76409 , n76410 );
and ( n76412 , n76411 , n32253 );
not ( n76413 , n32283 );
and ( n76414 , n76413 , n46016 );
and ( n76415 , n65885 , n32283 );
or ( n76416 , n76414 , n76415 );
and ( n76417 , n76416 , n32398 );
and ( n76418 , n46016 , n32436 );
or ( n76419 , n76412 , n76417 , n76418 );
and ( n76420 , n76419 , n32456 );
and ( n76421 , n46060 , n32473 );
not ( n76422 , n32475 );
and ( n76423 , n76422 , n46060 );
and ( n76424 , n46017 , n50482 );
xor ( n76425 , n46016 , n76424 );
and ( n76426 , n76425 , n32475 );
or ( n76427 , n76423 , n76426 );
and ( n76428 , n76427 , n32486 );
and ( n76429 , n37512 , n32489 );
and ( n76430 , n46016 , n32501 );
or ( n76431 , C0 , n76420 , n76421 , n76428 , n76429 , n76430 );
buf ( n76432 , n76431 );
buf ( n76433 , n76432 );
buf ( n76434 , n31655 );
buf ( n76435 , n30987 );
buf ( n76436 , n30987 );
buf ( n76437 , n31655 );
xor ( n76438 , n33101 , n58383 );
and ( n76439 , n76438 , n33201 );
not ( n76440 , n41576 );
and ( n76441 , n76440 , n33101 );
and ( n76442 , n55389 , n41576 );
or ( n76443 , n76441 , n76442 );
and ( n76444 , n76443 , n33189 );
and ( n76445 , n33101 , n41592 );
or ( n76446 , n76439 , n76444 , n76445 );
and ( n76447 , n76446 , n33208 );
and ( n76448 , n33101 , n39805 );
or ( n76449 , C0 , n76447 , n76448 );
buf ( n76450 , n76449 );
buf ( n76451 , n76450 );
not ( n76452 , n50828 );
not ( n76453 , n50834 );
and ( n76454 , n76453 , n40611 );
and ( n76455 , n55346 , n50834 );
or ( n76456 , n76454 , n76455 );
and ( n76457 , n76452 , n76456 );
buf ( n76458 , RI15b60210_1145);
and ( n76459 , n76458 , n50828 );
or ( n76460 , n76457 , n76459 );
buf ( n76461 , n76460 );
buf ( n76462 , n76461 );
buf ( n76463 , n31655 );
not ( n76464 , n41532 );
and ( n76465 , n76464 , n34188 );
and ( n76466 , n66889 , n41532 );
or ( n76467 , n76465 , n76466 );
buf ( n76468 , n76467 );
buf ( n76469 , n76468 );
buf ( n76470 , n31655 );
buf ( n76471 , n30987 );
xor ( n76472 , n33121 , n52218 );
and ( n76473 , n76472 , n33201 );
not ( n76474 , n41576 );
and ( n76475 , n76474 , n33121 );
buf ( n76476 , n32854 );
and ( n76477 , n76476 , n41576 );
or ( n76478 , n76475 , n76477 );
and ( n76479 , n76478 , n33189 );
and ( n76480 , n33121 , n41592 );
or ( n76481 , n76473 , n76479 , n76480 );
and ( n76482 , n76481 , n33208 );
and ( n76483 , n33121 , n39805 );
or ( n76484 , C0 , n76482 , n76483 );
buf ( n76485 , n76484 );
buf ( n76486 , n76485 );
buf ( n76487 , n30987 );
not ( n76488 , n34150 );
and ( n76489 , n76488 , n32867 );
not ( n76490 , n58762 );
and ( n76491 , n76490 , n32867 );
and ( n76492 , n32889 , n58762 );
or ( n76493 , n76491 , n76492 );
and ( n76494 , n76493 , n34150 );
or ( n76495 , n76489 , n76494 );
and ( n76496 , n76495 , n33381 );
not ( n76497 , n58770 );
not ( n76498 , n58762 );
and ( n76499 , n76498 , n32867 );
and ( n76500 , n52819 , n58762 );
or ( n76501 , n76499 , n76500 );
and ( n76502 , n76497 , n76501 );
and ( n76503 , n52819 , n58770 );
or ( n76504 , n76502 , n76503 );
and ( n76505 , n76504 , n33375 );
not ( n76506 , n32968 );
not ( n76507 , n58770 );
not ( n76508 , n58762 );
and ( n76509 , n76508 , n32867 );
and ( n76510 , n52819 , n58762 );
or ( n76511 , n76509 , n76510 );
and ( n76512 , n76507 , n76511 );
and ( n76513 , n52819 , n58770 );
or ( n76514 , n76512 , n76513 );
and ( n76515 , n76506 , n76514 );
not ( n76516 , n58790 );
not ( n76517 , n58792 );
and ( n76518 , n76517 , n76514 );
and ( n76519 , n52845 , n58792 );
or ( n76520 , n76518 , n76519 );
and ( n76521 , n76516 , n76520 );
and ( n76522 , n52855 , n58790 );
or ( n76523 , n76521 , n76522 );
and ( n76524 , n76523 , n32968 );
or ( n76525 , n76515 , n76524 );
and ( n76526 , n76525 , n33370 );
and ( n76527 , n32867 , n35062 );
or ( n76528 , C0 , n76496 , n76505 , n76526 , n76527 );
buf ( n76529 , n76528 );
buf ( n76530 , n76529 );
buf ( n76531 , n30987 );
buf ( n76532 , n30987 );
buf ( n76533 , n31655 );
buf ( n76534 , n31655 );
xor ( n76535 , n35445 , n39941 );
and ( n76536 , n76535 , n31550 );
not ( n76537 , n39979 );
and ( n76538 , n76537 , n35445 );
and ( n76539 , n69011 , n39979 );
or ( n76540 , n76538 , n76539 );
and ( n76541 , n76540 , n31538 );
and ( n76542 , n35445 , n40143 );
or ( n76543 , n76536 , n76541 , n76542 );
and ( n76544 , n76543 , n31557 );
and ( n76545 , n35445 , n40154 );
or ( n76546 , C0 , n76544 , n76545 );
buf ( n76547 , n76546 );
buf ( n76548 , n76547 );
buf ( n76549 , RI15b478c8_306);
buf ( n76550 , n76549 );
buf ( n76551 , n31655 );
not ( n76552 , n40163 );
and ( n76553 , n76552 , n31889 );
not ( n76554 , n75905 );
and ( n76555 , n76554 , n31889 );
and ( n76556 , n32218 , n75905 );
or ( n76557 , n76555 , n76556 );
and ( n76558 , n76557 , n40163 );
or ( n76559 , n76553 , n76558 );
and ( n76560 , n76559 , n32498 );
not ( n76561 , n75913 );
not ( n76562 , n75905 );
and ( n76563 , n76562 , n31889 );
and ( n76564 , n42255 , n75905 );
or ( n76565 , n76563 , n76564 );
and ( n76566 , n76561 , n76565 );
and ( n76567 , n42255 , n75913 );
or ( n76568 , n76566 , n76567 );
and ( n76569 , n76568 , n32473 );
not ( n76570 , n32475 );
not ( n76571 , n75913 );
not ( n76572 , n75905 );
and ( n76573 , n76572 , n31889 );
and ( n76574 , n42255 , n75905 );
or ( n76575 , n76573 , n76574 );
and ( n76576 , n76571 , n76575 );
and ( n76577 , n42255 , n75913 );
or ( n76578 , n76576 , n76577 );
and ( n76579 , n76570 , n76578 );
not ( n76580 , n75933 );
not ( n76581 , n75935 );
and ( n76582 , n76581 , n76578 );
and ( n76583 , n42283 , n75935 );
or ( n76584 , n76582 , n76583 );
and ( n76585 , n76580 , n76584 );
and ( n76586 , n42291 , n75933 );
or ( n76587 , n76585 , n76586 );
and ( n76588 , n76587 , n32475 );
or ( n76589 , n76579 , n76588 );
and ( n76590 , n76589 , n32486 );
and ( n76591 , n31889 , n41278 );
or ( n76592 , C0 , n76560 , n76569 , n76590 , n76591 );
buf ( n76593 , n76592 );
buf ( n76594 , n76593 );
buf ( n76595 , n30987 );
buf ( n76596 , n30987 );
buf ( n76597 , n31655 );
buf ( n76598 , n30987 );
buf ( n76599 , n30987 );
xor ( n76600 , n34062 , n39926 );
and ( n76601 , n76600 , n31550 );
not ( n76602 , n39979 );
and ( n76603 , n76602 , n34062 );
buf ( n76604 , n31270 );
and ( n76605 , n76604 , n39979 );
or ( n76606 , n76603 , n76605 );
and ( n76607 , n76606 , n31538 );
and ( n76608 , n34062 , n40143 );
or ( n76609 , n76601 , n76607 , n76608 );
and ( n76610 , n76609 , n31557 );
and ( n76611 , n34062 , n40154 );
or ( n76612 , C0 , n76610 , n76611 );
buf ( n76613 , n76612 );
buf ( n76614 , n76613 );
not ( n76615 , n40163 );
and ( n76616 , n76615 , n31920 );
not ( n76617 , n57233 );
and ( n76618 , n76617 , n31920 );
and ( n76619 , n32200 , n57233 );
or ( n76620 , n76618 , n76619 );
and ( n76621 , n76620 , n40163 );
or ( n76622 , n76616 , n76621 );
and ( n76623 , n76622 , n32498 );
not ( n76624 , n57241 );
not ( n76625 , n57233 );
and ( n76626 , n76625 , n31920 );
and ( n76627 , n53243 , n57233 );
or ( n76628 , n76626 , n76627 );
and ( n76629 , n76624 , n76628 );
and ( n76630 , n53243 , n57241 );
or ( n76631 , n76629 , n76630 );
and ( n76632 , n76631 , n32473 );
not ( n76633 , n32475 );
not ( n76634 , n57241 );
not ( n76635 , n57233 );
and ( n76636 , n76635 , n31920 );
and ( n76637 , n53243 , n57233 );
or ( n76638 , n76636 , n76637 );
and ( n76639 , n76634 , n76638 );
and ( n76640 , n53243 , n57241 );
or ( n76641 , n76639 , n76640 );
and ( n76642 , n76633 , n76641 );
not ( n76643 , n57261 );
not ( n76644 , n57263 );
and ( n76645 , n76644 , n76641 );
and ( n76646 , n53269 , n57263 );
or ( n76647 , n76645 , n76646 );
and ( n76648 , n76643 , n76647 );
and ( n76649 , n53277 , n57261 );
or ( n76650 , n76648 , n76649 );
and ( n76651 , n76650 , n32475 );
or ( n76652 , n76642 , n76651 );
and ( n76653 , n76652 , n32486 );
and ( n76654 , n31920 , n41278 );
or ( n76655 , C0 , n76623 , n76632 , n76653 , n76654 );
buf ( n76656 , n76655 );
buf ( n76657 , n76656 );
not ( n76658 , n40163 );
and ( n76659 , n76658 , n31817 );
not ( n76660 , n75905 );
and ( n76661 , n76660 , n31817 );
and ( n76662 , n32252 , n75905 );
or ( n76663 , n76661 , n76662 );
and ( n76664 , n76663 , n40163 );
or ( n76665 , n76659 , n76664 );
and ( n76666 , n76665 , n32498 );
not ( n76667 , n75913 );
not ( n76668 , n75905 );
and ( n76669 , n76668 , n31817 );
and ( n76670 , n40393 , n75905 );
or ( n76671 , n76669 , n76670 );
and ( n76672 , n76667 , n76671 );
and ( n76673 , n40393 , n75913 );
or ( n76674 , n76672 , n76673 );
and ( n76675 , n76674 , n32473 );
not ( n76676 , n32475 );
not ( n76677 , n75913 );
not ( n76678 , n75905 );
and ( n76679 , n76678 , n31817 );
and ( n76680 , n40393 , n75905 );
or ( n76681 , n76679 , n76680 );
and ( n76682 , n76677 , n76681 );
and ( n76683 , n40393 , n75913 );
or ( n76684 , n76682 , n76683 );
and ( n76685 , n76676 , n76684 );
not ( n76686 , n75933 );
not ( n76687 , n75935 );
and ( n76688 , n76687 , n76684 );
and ( n76689 , n40972 , n75935 );
or ( n76690 , n76688 , n76689 );
and ( n76691 , n76686 , n76690 );
and ( n76692 , n41267 , n75933 );
or ( n76693 , n76691 , n76692 );
and ( n76694 , n76693 , n32475 );
or ( n76695 , n76685 , n76694 );
and ( n76696 , n76695 , n32486 );
and ( n76697 , n31817 , n41278 );
or ( n76698 , C0 , n76666 , n76675 , n76696 , n76697 );
buf ( n76699 , n76698 );
buf ( n76700 , n76699 );
buf ( n76701 , n31655 );
buf ( n76702 , RI15b47c88_314);
buf ( n76703 , n76702 );
xor ( n76704 , n33997 , n39939 );
and ( n76705 , n76704 , n31550 );
not ( n76706 , n39979 );
and ( n76707 , n76706 , n33997 );
and ( n76708 , n31140 , n40095 );
and ( n76709 , n31142 , n40097 );
and ( n76710 , n31144 , n40099 );
and ( n76711 , n31146 , n40101 );
and ( n76712 , n31148 , n40103 );
and ( n76713 , n31150 , n40105 );
and ( n76714 , n31152 , n40107 );
and ( n76715 , n31154 , n40109 );
and ( n76716 , n31156 , n40111 );
and ( n76717 , n31158 , n40113 );
and ( n76718 , n31160 , n40115 );
and ( n76719 , n31162 , n40117 );
and ( n76720 , n31164 , n40119 );
and ( n76721 , n31166 , n40121 );
and ( n76722 , n31168 , n40123 );
and ( n76723 , n31170 , n40125 );
or ( n76724 , n76708 , n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , n76721 , n76722 , n76723 );
and ( n76725 , n76724 , n39979 );
or ( n76726 , n76707 , n76725 );
and ( n76727 , n76726 , n31538 );
and ( n76728 , n33997 , n40143 );
or ( n76729 , n76705 , n76727 , n76728 );
and ( n76730 , n76729 , n31557 );
and ( n76731 , n33997 , n40154 );
or ( n76732 , C0 , n76730 , n76731 );
buf ( n76733 , n76732 );
buf ( n76734 , n76733 );
buf ( n76735 , n30987 );
buf ( n76736 , n30987 );
buf ( n76737 , n30987 );
buf ( n76738 , n30987 );
buf ( n76739 , n31655 );
buf ( n76740 , RI15b46680_267);
and ( n76741 , n76740 , n33377 );
not ( n76742 , n48545 );
and ( n76743 , n76742 , n76702 );
buf ( n76744 , n76743 );
and ( n76745 , n76744 , n32890 );
not ( n76746 , n48557 );
and ( n76747 , n76746 , n76702 );
not ( n76748 , n54581 );
and ( n76749 , n76748 , n54560 );
xor ( n76750 , n54560 , n54340 );
and ( n76751 , n73808 , n73809 );
xor ( n76752 , n76750 , n76751 );
and ( n76753 , n76752 , n54581 );
or ( n76754 , n76749 , n76753 );
and ( n76755 , n76754 , n48557 );
or ( n76756 , n76747 , n76755 );
and ( n76757 , n76756 , n33038 );
and ( n76758 , n76702 , n48571 );
or ( n76759 , n76745 , n76757 , n76758 );
and ( n76760 , n76759 , n33208 );
and ( n76761 , n76702 , n48577 );
or ( n76762 , C0 , n76741 , n76760 , n76761 );
buf ( n76763 , n76762 );
buf ( n76764 , n76763 );
buf ( n76765 , n31655 );
xor ( n76766 , n35427 , n62855 );
and ( n76767 , n76766 , n31550 );
not ( n76768 , n39979 );
and ( n76769 , n76768 , n35427 );
and ( n76770 , n45112 , n68408 );
xor ( n76771 , n45095 , n76770 );
and ( n76772 , n76771 , n39979 );
or ( n76773 , n76769 , n76772 );
and ( n76774 , n76773 , n31538 );
and ( n76775 , n35427 , n40143 );
or ( n76776 , n76767 , n76774 , n76775 );
and ( n76777 , n76776 , n31557 );
and ( n76778 , n35427 , n40154 );
or ( n76779 , C0 , n76777 , n76778 );
buf ( n76780 , n76779 );
buf ( n76781 , n76780 );
buf ( n76782 , n30987 );
buf ( n76783 , n40214 );
buf ( n76784 , n30987 );
buf ( n76785 , n31655 );
not ( n76786 , n40163 );
and ( n76787 , n76786 , n31926 );
not ( n76788 , n40166 );
and ( n76789 , n76788 , n31926 );
and ( n76790 , n32200 , n40166 );
or ( n76791 , n76789 , n76790 );
and ( n76792 , n76791 , n40163 );
or ( n76793 , n76787 , n76792 );
and ( n76794 , n76793 , n32498 );
not ( n76795 , n40195 );
not ( n76796 , n40166 );
and ( n76797 , n76796 , n31926 );
and ( n76798 , n53243 , n40166 );
or ( n76799 , n76797 , n76798 );
and ( n76800 , n76795 , n76799 );
and ( n76801 , n53243 , n40195 );
or ( n76802 , n76800 , n76801 );
and ( n76803 , n76802 , n32473 );
not ( n76804 , n32475 );
not ( n76805 , n40195 );
not ( n76806 , n40166 );
and ( n76807 , n76806 , n31926 );
and ( n76808 , n53243 , n40166 );
or ( n76809 , n76807 , n76808 );
and ( n76810 , n76805 , n76809 );
and ( n76811 , n53243 , n40195 );
or ( n76812 , n76810 , n76811 );
and ( n76813 , n76804 , n76812 );
not ( n76814 , n40446 );
not ( n76815 , n40448 );
and ( n76816 , n76815 , n76812 );
and ( n76817 , n53269 , n40448 );
or ( n76818 , n76816 , n76817 );
and ( n76819 , n76814 , n76818 );
and ( n76820 , n53277 , n40446 );
or ( n76821 , n76819 , n76820 );
and ( n76822 , n76821 , n32475 );
or ( n76823 , n76813 , n76822 );
and ( n76824 , n76823 , n32486 );
and ( n76825 , n31926 , n41278 );
or ( n76826 , C0 , n76794 , n76803 , n76824 , n76825 );
buf ( n76827 , n76826 );
buf ( n76828 , n76827 );
and ( n76829 , n33223 , n32528 );
not ( n76830 , n32598 );
and ( n76831 , n76830 , n32986 );
buf ( n76832 , n76831 );
and ( n76833 , n76832 , n32890 );
not ( n76834 , n32919 );
and ( n76835 , n76834 , n32986 );
buf ( n76836 , n76835 );
and ( n76837 , n76836 , n32924 );
not ( n76838 , n32953 );
and ( n76839 , n76838 , n32986 );
not ( n76840 , n32971 );
and ( n76841 , n76840 , n33097 );
xor ( n76842 , n32986 , n33019 );
and ( n76843 , n76842 , n32971 );
or ( n76844 , n76841 , n76843 );
and ( n76845 , n76844 , n32953 );
or ( n76846 , n76839 , n76845 );
and ( n76847 , n76846 , n33038 );
not ( n76848 , n33067 );
and ( n76849 , n76848 , n32986 );
not ( n76850 , n32970 );
not ( n76851 , n33071 );
and ( n76852 , n76851 , n33097 );
xor ( n76853 , n33098 , n33151 );
and ( n76854 , n76853 , n33071 );
or ( n76855 , n76852 , n76854 );
and ( n76856 , n76850 , n76855 );
and ( n76857 , n76842 , n32970 );
or ( n76858 , n76856 , n76857 );
and ( n76859 , n76858 , n33067 );
or ( n76860 , n76849 , n76859 );
and ( n76861 , n76860 , n33172 );
and ( n76862 , n32986 , n33204 );
or ( n76863 , n76833 , n76837 , n76847 , n76861 , n76862 );
and ( n76864 , n76863 , n33208 );
not ( n76865 , n32968 );
not ( n76866 , n33270 );
and ( n76867 , n76866 , n33297 );
xor ( n76868 , n33298 , n33351 );
and ( n76869 , n76868 , n33270 );
or ( n76870 , n76867 , n76869 );
and ( n76871 , n76865 , n76870 );
and ( n76872 , n32986 , n32968 );
or ( n76873 , n76871 , n76872 );
and ( n76874 , n76873 , n33370 );
buf ( n76875 , n35056 );
and ( n76876 , n32986 , n33382 );
or ( n76877 , C0 , n76829 , n76864 , n76874 , n76875 , n76876 );
buf ( n76878 , n76877 );
buf ( n76879 , n76878 );
buf ( n76880 , n30987 );
not ( n76881 , n31728 );
and ( n76882 , n76881 , n46027 );
xor ( n76883 , n47604 , n47625 );
and ( n76884 , n76883 , n31728 );
or ( n76885 , n76882 , n76884 );
and ( n76886 , n76885 , n32253 );
not ( n76887 , n32283 );
and ( n76888 , n76887 , n46027 );
not ( n76889 , n31823 );
xor ( n76890 , n47659 , n47680 );
and ( n76891 , n76889 , n76890 );
xnor ( n76892 , n47709 , n47730 );
and ( n76893 , n76892 , n31823 );
or ( n76894 , n76891 , n76893 );
and ( n76895 , n76894 , n32283 );
or ( n76896 , n76888 , n76895 );
and ( n76897 , n76896 , n32398 );
and ( n76898 , n46027 , n32436 );
or ( n76899 , n76886 , n76897 , n76898 );
and ( n76900 , n76899 , n32456 );
and ( n76901 , n49671 , n32473 );
not ( n76902 , n32475 );
and ( n76903 , n76902 , n49671 );
xor ( n76904 , n46027 , n47759 );
and ( n76905 , n76904 , n32475 );
or ( n76906 , n76903 , n76905 );
and ( n76907 , n76906 , n32486 );
and ( n76908 , n37551 , n32489 );
and ( n76909 , n46027 , n32501 );
or ( n76910 , C0 , n76900 , n76901 , n76907 , n76908 , n76909 );
buf ( n76911 , n76910 );
buf ( n76912 , n76911 );
buf ( n76913 , n31655 );
buf ( n76914 , n31655 );
buf ( n76915 , n30987 );
buf ( n76916 , n30987 );
buf ( n76917 , n31655 );
buf ( n76918 , n31655 );
buf ( n76919 , n30987 );
xor ( n76920 , n49573 , n60319 );
and ( n76921 , n76920 , n32433 );
not ( n76922 , n47331 );
and ( n76923 , n76922 , n49573 );
xor ( n76924 , n60467 , n60543 );
and ( n76925 , n76924 , n47331 );
or ( n76926 , n76923 , n76925 );
and ( n76927 , n76926 , n32413 );
and ( n76928 , n49573 , n47402 );
or ( n76929 , n76921 , n76927 , n76928 );
and ( n76930 , n76929 , n32456 );
and ( n76931 , n49573 , n47409 );
or ( n76932 , C0 , n76930 , n76931 );
buf ( n76933 , n76932 );
buf ( n76934 , n76933 );
not ( n76935 , n46356 );
and ( n76936 , n76935 , n31132 );
not ( n76937 , n61975 );
and ( n76938 , n76937 , n31132 );
and ( n76939 , n31138 , n61975 );
or ( n76940 , n76938 , n76939 );
and ( n76941 , n76940 , n46356 );
or ( n76942 , n76936 , n76941 );
and ( n76943 , n76942 , n31649 );
not ( n76944 , n61983 );
not ( n76945 , n61975 );
and ( n76946 , n76945 , n31132 );
and ( n76947 , n56920 , n61975 );
or ( n76948 , n76946 , n76947 );
and ( n76949 , n76944 , n76948 );
and ( n76950 , n56920 , n61983 );
or ( n76951 , n76949 , n76950 );
and ( n76952 , n76951 , n31643 );
not ( n76953 , n31452 );
not ( n76954 , n61983 );
not ( n76955 , n61975 );
and ( n76956 , n76955 , n31132 );
and ( n76957 , n56920 , n61975 );
or ( n76958 , n76956 , n76957 );
and ( n76959 , n76954 , n76958 );
and ( n76960 , n56920 , n61983 );
or ( n76961 , n76959 , n76960 );
and ( n76962 , n76953 , n76961 );
not ( n76963 , n62003 );
not ( n76964 , n62005 );
and ( n76965 , n76964 , n76961 );
and ( n76966 , n56946 , n62005 );
or ( n76967 , n76965 , n76966 );
and ( n76968 , n76963 , n76967 );
and ( n76969 , n56954 , n62003 );
or ( n76970 , n76968 , n76969 );
and ( n76971 , n76970 , n31452 );
or ( n76972 , n76962 , n76971 );
and ( n76973 , n76972 , n31638 );
and ( n76974 , n31132 , n47277 );
or ( n76975 , C0 , n76943 , n76952 , n76973 , n76974 );
buf ( n76976 , n76975 );
buf ( n76977 , n76976 );
not ( n76978 , n34150 );
and ( n76979 , n76978 , n32729 );
not ( n76980 , n59574 );
and ( n76981 , n76980 , n32729 );
and ( n76982 , n32755 , n59574 );
or ( n76983 , n76981 , n76982 );
and ( n76984 , n76983 , n34150 );
or ( n76985 , n76979 , n76984 );
and ( n76986 , n76985 , n33381 );
not ( n76987 , n59582 );
not ( n76988 , n59574 );
and ( n76989 , n76988 , n32729 );
and ( n76990 , n35083 , n59574 );
or ( n76991 , n76989 , n76990 );
and ( n76992 , n76987 , n76991 );
and ( n76993 , n35083 , n59582 );
or ( n76994 , n76992 , n76993 );
and ( n76995 , n76994 , n33375 );
not ( n76996 , n32968 );
not ( n76997 , n59582 );
not ( n76998 , n59574 );
and ( n76999 , n76998 , n32729 );
and ( n77000 , n35083 , n59574 );
or ( n77001 , n76999 , n77000 );
and ( n77002 , n76997 , n77001 );
and ( n77003 , n35083 , n59582 );
or ( n77004 , n77002 , n77003 );
and ( n77005 , n76996 , n77004 );
not ( n77006 , n59602 );
not ( n77007 , n59604 );
and ( n77008 , n77007 , n77004 );
and ( n77009 , n35107 , n59604 );
or ( n77010 , n77008 , n77009 );
and ( n77011 , n77006 , n77010 );
and ( n77012 , n35115 , n59602 );
or ( n77013 , n77011 , n77012 );
and ( n77014 , n77013 , n32968 );
or ( n77015 , n77005 , n77014 );
and ( n77016 , n77015 , n33370 );
and ( n77017 , n32729 , n35062 );
or ( n77018 , C0 , n76986 , n76995 , n77016 , n77017 );
buf ( n77019 , n77018 );
buf ( n77020 , n77019 );
buf ( n77021 , n30987 );
buf ( n77022 , n31655 );
buf ( n77023 , n31655 );
buf ( n77024 , n30987 );
buf ( n77025 , n30987 );
buf ( n77026 , n31655 );
buf ( n77027 , n31655 );
buf ( n77028 , n30987 );
and ( n77029 , n49083 , n48639 );
not ( n77030 , n48642 );
and ( n77031 , n77030 , n48606 );
and ( n77032 , n49083 , n48642 );
or ( n77033 , n77031 , n77032 );
and ( n77034 , n77033 , n32890 );
not ( n77035 , n48648 );
and ( n77036 , n77035 , n48606 );
and ( n77037 , n49083 , n48648 );
or ( n77038 , n77036 , n77037 );
and ( n77039 , n77038 , n32924 );
not ( n77040 , n48654 );
and ( n77041 , n77040 , n48606 );
and ( n77042 , n49083 , n48654 );
or ( n77043 , n77041 , n77042 );
and ( n77044 , n77043 , n33038 );
not ( n77045 , n48660 );
and ( n77046 , n77045 , n48606 );
and ( n77047 , n49083 , n48660 );
or ( n77048 , n77046 , n77047 );
and ( n77049 , n77048 , n33172 );
not ( n77050 , n41576 );
and ( n77051 , n77050 , n48606 );
and ( n77052 , n48866 , n41576 );
or ( n77053 , n77051 , n77052 );
and ( n77054 , n77053 , n33189 );
not ( n77055 , n48730 );
and ( n77056 , n77055 , n48606 );
and ( n77057 , n48866 , n48730 );
or ( n77058 , n77056 , n77057 );
and ( n77059 , n77058 , n33187 );
not ( n77060 , n48765 );
and ( n77061 , n77060 , n48606 );
and ( n77062 , n73880 , n48765 );
or ( n77063 , n77061 , n77062 );
and ( n77064 , n77063 , n33180 );
not ( n77065 , n49054 );
and ( n77066 , n77065 , n48606 );
and ( n77067 , n73893 , n49054 );
or ( n77068 , n77066 , n77067 );
and ( n77069 , n77068 , n33178 );
and ( n77070 , n49196 , n49275 );
or ( n77071 , n77029 , n77034 , n77039 , n77044 , n77049 , n77054 , n77059 , n77064 , n77069 , n77070 );
and ( n77072 , n77071 , n33208 );
and ( n77073 , n32999 , n35056 );
and ( n77074 , n48606 , n49286 );
or ( n77075 , C0 , n77072 , n77073 , n77074 );
buf ( n77076 , n77075 );
buf ( n77077 , n77076 );
not ( n77078 , n46356 );
and ( n77079 , n77078 , n31187 );
not ( n77080 , n48214 );
and ( n77081 , n77080 , n31187 );
and ( n77082 , n31205 , n48214 );
or ( n77083 , n77081 , n77082 );
and ( n77084 , n77083 , n46356 );
or ( n77085 , n77079 , n77084 );
and ( n77086 , n77085 , n31649 );
not ( n77087 , n48223 );
not ( n77088 , n48214 );
and ( n77089 , n77088 , n31187 );
and ( n77090 , n50125 , n48214 );
or ( n77091 , n77089 , n77090 );
and ( n77092 , n77087 , n77091 );
and ( n77093 , n50125 , n48223 );
or ( n77094 , n77092 , n77093 );
and ( n77095 , n77094 , n31643 );
not ( n77096 , n31452 );
not ( n77097 , n48223 );
not ( n77098 , n48214 );
and ( n77099 , n77098 , n31187 );
and ( n77100 , n50125 , n48214 );
or ( n77101 , n77099 , n77100 );
and ( n77102 , n77097 , n77101 );
and ( n77103 , n50125 , n48223 );
or ( n77104 , n77102 , n77103 );
and ( n77105 , n77096 , n77104 );
not ( n77106 , n48244 );
not ( n77107 , n48247 );
and ( n77108 , n77107 , n77104 );
and ( n77109 , n50151 , n48247 );
or ( n77110 , n77108 , n77109 );
and ( n77111 , n77106 , n77110 );
and ( n77112 , n50159 , n48244 );
or ( n77113 , n77111 , n77112 );
and ( n77114 , n77113 , n31452 );
or ( n77115 , n77105 , n77114 );
and ( n77116 , n77115 , n31638 );
and ( n77117 , n31187 , n47277 );
or ( n77118 , C0 , n77086 , n77095 , n77116 , n77117 );
buf ( n77119 , n77118 );
buf ( n77120 , n77119 );
buf ( n77121 , n31655 );
buf ( n77122 , n30987 );
buf ( n77123 , n31655 );
not ( n77124 , n48267 );
not ( n77125 , n48269 );
not ( n77126 , n48272 );
and ( n77127 , n77126 , n48276 );
buf ( n77128 , n48272 );
or ( n77129 , n77127 , n77128 );
and ( n77130 , n77125 , n77129 );
buf ( n77131 , n77130 );
and ( n77132 , n77124 , n77131 );
buf ( n77133 , n48267 );
or ( n77134 , n77132 , n77133 );
and ( n77135 , n77134 , n39358 );
and ( n77136 , n76252 , n38450 );
and ( n77137 , n48287 , n39356 );
not ( n77138 , n48297 );
not ( n77139 , n48300 );
and ( n77140 , n77139 , n48294 );
buf ( n77141 , n48300 );
or ( n77142 , n77140 , n77141 );
and ( n77143 , n77138 , n77142 );
buf ( n77144 , n48297 );
or ( n77145 , n77143 , n77144 );
and ( n77146 , n77145 , n39354 );
not ( n77147 , n48272 );
not ( n77148 , n48311 );
not ( n77149 , n48315 );
not ( n77150 , n48318 );
not ( n77151 , n48320 );
not ( n77152 , n48322 );
and ( n77153 , n77151 , n77152 );
buf ( n77154 , n77153 );
and ( n77155 , n77150 , n77154 );
buf ( n77156 , n48318 );
or ( n77157 , n77155 , n77156 );
and ( n77158 , n77149 , n77157 );
buf ( n77159 , n48315 );
or ( n77160 , n77158 , n77159 );
and ( n77161 , n77148 , n77160 );
and ( n77162 , n35282 , n48311 );
or ( n77163 , n77161 , n77162 );
and ( n77164 , n77147 , n77163 );
buf ( n77165 , n48272 );
or ( n77166 , n77164 , n77165 );
and ( n77167 , n77166 , n39352 );
buf ( n77168 , n39346 );
and ( n77169 , n48263 , n39349 );
or ( n77170 , n77135 , n77136 , n77137 , n77146 , n77167 , n77168 , n77169 , C0 );
buf ( n77171 , n77170 );
buf ( n77172 , n77171 );
and ( n77173 , n33218 , n32528 );
not ( n77174 , n32598 );
and ( n77175 , n77174 , n32981 );
buf ( n77176 , n77175 );
and ( n77177 , n77176 , n32890 );
not ( n77178 , n32919 );
and ( n77179 , n77178 , n32981 );
buf ( n77180 , n77179 );
and ( n77181 , n77180 , n32924 );
not ( n77182 , n32953 );
and ( n77183 , n77182 , n32981 );
not ( n77184 , n32971 );
and ( n77185 , n77184 , n33087 );
xor ( n77186 , n32981 , n33024 );
and ( n77187 , n77186 , n32971 );
or ( n77188 , n77185 , n77187 );
and ( n77189 , n77188 , n32953 );
or ( n77190 , n77183 , n77189 );
and ( n77191 , n77190 , n33038 );
not ( n77192 , n33067 );
and ( n77193 , n77192 , n32981 );
not ( n77194 , n32970 );
not ( n77195 , n33071 );
and ( n77196 , n77195 , n33087 );
xor ( n77197 , n33088 , n33156 );
and ( n77198 , n77197 , n33071 );
or ( n77199 , n77196 , n77198 );
and ( n77200 , n77194 , n77199 );
and ( n77201 , n77186 , n32970 );
or ( n77202 , n77200 , n77201 );
and ( n77203 , n77202 , n33067 );
or ( n77204 , n77193 , n77203 );
and ( n77205 , n77204 , n33172 );
and ( n77206 , n32981 , n33204 );
or ( n77207 , n77177 , n77181 , n77191 , n77205 , n77206 );
and ( n77208 , n77207 , n33208 );
not ( n77209 , n32968 );
not ( n77210 , n33270 );
and ( n77211 , n77210 , n33287 );
xor ( n77212 , n33288 , n33356 );
and ( n77213 , n77212 , n33270 );
or ( n77214 , n77211 , n77213 );
and ( n77215 , n77209 , n77214 );
and ( n77216 , n32981 , n32968 );
or ( n77217 , n77215 , n77216 );
and ( n77218 , n77217 , n33370 );
and ( n77219 , n32981 , n33382 );
or ( n77220 , C0 , n77173 , n77208 , n77218 , C0 , n77219 );
buf ( n77221 , n77220 );
buf ( n77222 , n77221 );
buf ( n77223 , n30987 );
buf ( n77224 , n31655 );
not ( n77225 , n31728 );
and ( n77226 , n77225 , n46032 );
and ( n77227 , n75834 , n31728 );
or ( n77228 , n77226 , n77227 );
and ( n77229 , n77228 , n32253 );
not ( n77230 , n32283 );
and ( n77231 , n77230 , n46032 );
and ( n77232 , n75845 , n32283 );
or ( n77233 , n77231 , n77232 );
and ( n77234 , n77233 , n32398 );
and ( n77235 , n46032 , n32436 );
or ( n77236 , n77229 , n77234 , n77235 );
and ( n77237 , n77236 , n32456 );
and ( n77238 , n49681 , n32473 );
not ( n77239 , n32475 );
and ( n77240 , n77239 , n49681 );
xor ( n77241 , n46032 , n47754 );
and ( n77242 , n77241 , n32475 );
or ( n77243 , n77240 , n77242 );
and ( n77244 , n77243 , n32486 );
and ( n77245 , n37561 , n32489 );
and ( n77246 , n46032 , n32501 );
or ( n77247 , C0 , n77237 , n77238 , n77244 , n77245 , n77246 );
buf ( n77248 , n77247 );
buf ( n77249 , n77248 );
buf ( n77250 , n31655 );
buf ( n77251 , n30987 );
buf ( n77252 , n31655 );
xor ( n77253 , n44770 , n44797 );
and ( n77254 , n77253 , n31548 );
not ( n77255 , n44807 );
and ( n77256 , n77255 , n44770 );
and ( n77257 , n46647 , n44807 );
or ( n77258 , n77256 , n77257 );
and ( n77259 , n77258 , n31408 );
not ( n77260 , n44817 );
and ( n77261 , n77260 , n44770 );
and ( n77262 , n53164 , n44817 );
or ( n77263 , n77261 , n77262 );
and ( n77264 , n77263 , n31521 );
not ( n77265 , n45059 );
and ( n77266 , n77265 , n44770 );
and ( n77267 , n31307 , n40095 );
and ( n77268 , n31309 , n40097 );
and ( n77269 , n31311 , n40099 );
and ( n77270 , n31313 , n40101 );
and ( n77271 , n31315 , n40103 );
and ( n77272 , n31317 , n40105 );
and ( n77273 , n31319 , n40107 );
and ( n77274 , n31321 , n40109 );
and ( n77275 , n31323 , n40111 );
and ( n77276 , n31325 , n40113 );
and ( n77277 , n31327 , n40115 );
and ( n77278 , n31329 , n40117 );
and ( n77279 , n31331 , n40119 );
and ( n77280 , n31333 , n40121 );
and ( n77281 , n31335 , n40123 );
and ( n77282 , n31337 , n40125 );
or ( n77283 , n77267 , n77268 , n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , n77281 , n77282 );
and ( n77284 , n77283 , n45059 );
or ( n77285 , n77266 , n77284 );
and ( n77286 , n77285 , n31536 );
and ( n77287 , n44770 , n45148 );
or ( n77288 , n77254 , n77259 , n77264 , n77286 , n77287 );
and ( n77289 , n77288 , n31557 );
and ( n77290 , n44770 , n40154 );
or ( n77291 , C0 , n77289 , n77290 );
buf ( n77292 , n77291 );
buf ( n77293 , n77292 );
not ( n77294 , n40163 );
and ( n77295 , n77294 , n31986 );
not ( n77296 , n55888 );
and ( n77297 , n77296 , n31986 );
and ( n77298 , n32165 , n55888 );
or ( n77299 , n77297 , n77298 );
and ( n77300 , n77299 , n40163 );
or ( n77301 , n77295 , n77300 );
and ( n77302 , n77301 , n32498 );
not ( n77303 , n55896 );
not ( n77304 , n55888 );
and ( n77305 , n77304 , n31986 );
and ( n77306 , n59005 , n55888 );
or ( n77307 , n77305 , n77306 );
and ( n77308 , n77303 , n77307 );
and ( n77309 , n59005 , n55896 );
or ( n77310 , n77308 , n77309 );
and ( n77311 , n77310 , n32473 );
not ( n77312 , n32475 );
not ( n77313 , n55896 );
not ( n77314 , n55888 );
and ( n77315 , n77314 , n31986 );
and ( n77316 , n59005 , n55888 );
or ( n77317 , n77315 , n77316 );
and ( n77318 , n77313 , n77317 );
and ( n77319 , n59005 , n55896 );
or ( n77320 , n77318 , n77319 );
and ( n77321 , n77312 , n77320 );
not ( n77322 , n55916 );
not ( n77323 , n55918 );
and ( n77324 , n77323 , n77320 );
and ( n77325 , n59029 , n55918 );
or ( n77326 , n77324 , n77325 );
and ( n77327 , n77322 , n77326 );
and ( n77328 , n59037 , n55916 );
or ( n77329 , n77327 , n77328 );
and ( n77330 , n77329 , n32475 );
or ( n77331 , n77321 , n77330 );
and ( n77332 , n77331 , n32486 );
and ( n77333 , n31986 , n41278 );
or ( n77334 , C0 , n77302 , n77311 , n77332 , n77333 );
buf ( n77335 , n77334 );
buf ( n77336 , n77335 );
buf ( n77337 , n30987 );
buf ( n77338 , n30987 );
buf ( n77339 , n31655 );
and ( n77340 , n51725 , n31645 );
not ( n77341 , n45274 );
and ( n77342 , n77341 , n69688 );
buf ( n77343 , n77342 );
and ( n77344 , n77343 , n31373 );
not ( n77345 , n45280 );
and ( n77346 , n77345 , n69688 );
and ( n77347 , n51731 , n45280 );
or ( n77348 , n77346 , n77347 );
and ( n77349 , n77348 , n31468 );
and ( n77350 , n69688 , n45802 );
or ( n77351 , n77344 , n77349 , n77350 );
and ( n77352 , n77351 , n31557 );
and ( n77353 , n69688 , n45808 );
or ( n77354 , C0 , n77340 , n77352 , n77353 );
buf ( n77355 , n77354 );
buf ( n77356 , n77355 );
buf ( n77357 , n30987 );
not ( n77358 , n40163 );
and ( n77359 , n77358 , n31974 );
not ( n77360 , n54629 );
and ( n77361 , n77360 , n31974 );
and ( n77362 , n32165 , n54629 );
or ( n77363 , n77361 , n77362 );
and ( n77364 , n77363 , n40163 );
or ( n77365 , n77359 , n77364 );
and ( n77366 , n77365 , n32498 );
not ( n77367 , n54637 );
not ( n77368 , n54629 );
and ( n77369 , n77368 , n31974 );
and ( n77370 , n59005 , n54629 );
or ( n77371 , n77369 , n77370 );
and ( n77372 , n77367 , n77371 );
and ( n77373 , n59005 , n54637 );
or ( n77374 , n77372 , n77373 );
and ( n77375 , n77374 , n32473 );
not ( n77376 , n32475 );
not ( n77377 , n54637 );
not ( n77378 , n54629 );
and ( n77379 , n77378 , n31974 );
and ( n77380 , n59005 , n54629 );
or ( n77381 , n77379 , n77380 );
and ( n77382 , n77377 , n77381 );
and ( n77383 , n59005 , n54637 );
or ( n77384 , n77382 , n77383 );
and ( n77385 , n77376 , n77384 );
not ( n77386 , n54657 );
not ( n77387 , n54659 );
and ( n77388 , n77387 , n77384 );
and ( n77389 , n59029 , n54659 );
or ( n77390 , n77388 , n77389 );
and ( n77391 , n77386 , n77390 );
and ( n77392 , n59037 , n54657 );
or ( n77393 , n77391 , n77392 );
and ( n77394 , n77393 , n32475 );
or ( n77395 , n77385 , n77394 );
and ( n77396 , n77395 , n32486 );
and ( n77397 , n31974 , n41278 );
or ( n77398 , C0 , n77366 , n77375 , n77396 , n77397 );
buf ( n77399 , n77398 );
buf ( n77400 , n77399 );
buf ( n77401 , n31655 );
buf ( n77402 , n30987 );
and ( n77403 , n46031 , n32500 );
not ( n77404 , n35211 );
and ( n77405 , n77404 , n37559 );
buf ( n77406 , n77405 );
and ( n77407 , n77406 , n32421 );
not ( n77408 , n35245 );
and ( n77409 , n77408 , n37559 );
buf ( n77410 , n77409 );
and ( n77411 , n77410 , n32419 );
not ( n77412 , n35278 );
and ( n77413 , n77412 , n37559 );
not ( n77414 , n35295 );
and ( n77415 , n77414 , n49589 );
xor ( n77416 , n37559 , n49536 );
and ( n77417 , n77416 , n35295 );
or ( n77418 , n77415 , n77417 );
and ( n77419 , n77418 , n35278 );
or ( n77420 , n77413 , n77419 );
and ( n77421 , n77420 , n32417 );
not ( n77422 , n35331 );
and ( n77423 , n77422 , n37559 );
not ( n77424 , n35294 );
not ( n77425 , n45995 );
and ( n77426 , n77425 , n49589 );
xor ( n77427 , n49590 , n49622 );
and ( n77428 , n77427 , n45995 );
or ( n77429 , n77426 , n77428 );
and ( n77430 , n77424 , n77429 );
and ( n77431 , n77416 , n35294 );
or ( n77432 , n77430 , n77431 );
and ( n77433 , n77432 , n35331 );
or ( n77434 , n77423 , n77433 );
and ( n77435 , n77434 , n32415 );
and ( n77436 , n37559 , n35354 );
or ( n77437 , n77407 , n77411 , n77421 , n77435 , n77436 );
and ( n77438 , n77437 , n32456 );
not ( n77439 , n32475 );
not ( n77440 , n46060 );
and ( n77441 , n77440 , n49679 );
xor ( n77442 , n49680 , n49716 );
and ( n77443 , n77442 , n46060 );
or ( n77444 , n77441 , n77443 );
and ( n77445 , n77439 , n77444 );
and ( n77446 , n37559 , n32475 );
or ( n77447 , n77445 , n77446 );
and ( n77448 , n77447 , n32486 );
buf ( n77449 , n32489 );
and ( n77450 , n37559 , n35367 );
or ( n77451 , C0 , n77403 , n77438 , n77448 , n77449 , n77450 );
buf ( n77452 , n77451 );
buf ( n77453 , n77452 );
buf ( n77454 , n40219 );
buf ( n77455 , n30987 );
buf ( n77456 , n31655 );
not ( n77457 , n48765 );
and ( n77458 , n77457 , n33219 );
xor ( n77459 , n48774 , n49014 );
and ( n77460 , n77459 , n48765 );
or ( n77461 , n77458 , n77460 );
and ( n77462 , n77461 , n33180 );
not ( n77463 , n49054 );
and ( n77464 , n77463 , n33219 );
not ( n77465 , n48845 );
xor ( n77466 , n49064 , n49128 );
and ( n77467 , n77465 , n77466 );
xnor ( n77468 , n49173 , n49254 );
and ( n77469 , n77468 , n48845 );
or ( n77470 , n77467 , n77469 );
and ( n77471 , n77470 , n49054 );
or ( n77472 , n77464 , n77471 );
and ( n77473 , n77472 , n33178 );
and ( n77474 , n33219 , n49774 );
or ( n77475 , n77462 , n77473 , n77474 );
and ( n77476 , n77475 , n33208 );
and ( n77477 , n33289 , n33375 );
not ( n77478 , n32968 );
and ( n77479 , n77478 , n33289 );
xor ( n77480 , n33219 , n59699 );
and ( n77481 , n77480 , n32968 );
or ( n77482 , n77479 , n77481 );
and ( n77483 , n77482 , n33370 );
and ( n77484 , n32982 , n35056 );
and ( n77485 , n33219 , n49794 );
or ( n77486 , C0 , n77476 , n77477 , n77483 , n77484 , n77485 );
buf ( n77487 , n77486 );
buf ( n77488 , n77487 );
not ( n77489 , n40163 );
and ( n77490 , n77489 , n32060 );
not ( n77491 , n57233 );
and ( n77492 , n77491 , n32060 );
and ( n77493 , n32130 , n57233 );
or ( n77494 , n77492 , n77493 );
and ( n77495 , n77494 , n40163 );
or ( n77496 , n77490 , n77495 );
and ( n77497 , n77496 , n32498 );
not ( n77498 , n57241 );
not ( n77499 , n57233 );
and ( n77500 , n77499 , n32060 );
and ( n77501 , n45833 , n57233 );
or ( n77502 , n77500 , n77501 );
and ( n77503 , n77498 , n77502 );
and ( n77504 , n45833 , n57241 );
or ( n77505 , n77503 , n77504 );
and ( n77506 , n77505 , n32473 );
not ( n77507 , n32475 );
not ( n77508 , n57241 );
not ( n77509 , n57233 );
and ( n77510 , n77509 , n32060 );
and ( n77511 , n45833 , n57233 );
or ( n77512 , n77510 , n77511 );
and ( n77513 , n77508 , n77512 );
and ( n77514 , n45833 , n57241 );
or ( n77515 , n77513 , n77514 );
and ( n77516 , n77507 , n77515 );
not ( n77517 , n57261 );
not ( n77518 , n57263 );
and ( n77519 , n77518 , n77515 );
and ( n77520 , n45857 , n57263 );
or ( n77521 , n77519 , n77520 );
and ( n77522 , n77517 , n77521 );
and ( n77523 , n45865 , n57261 );
or ( n77524 , n77522 , n77523 );
and ( n77525 , n77524 , n32475 );
or ( n77526 , n77516 , n77525 );
and ( n77527 , n77526 , n32486 );
and ( n77528 , n32060 , n41278 );
or ( n77529 , C0 , n77497 , n77506 , n77527 , n77528 );
buf ( n77530 , n77529 );
buf ( n77531 , n77530 );
buf ( n77532 , n30987 );
buf ( n77533 , n31655 );
buf ( n77534 , n30987 );
xor ( n77535 , n34054 , n39930 );
and ( n77536 , n77535 , n31550 );
not ( n77537 , n39979 );
and ( n77538 , n77537 , n34054 );
and ( n77539 , n31086 , n42330 );
and ( n77540 , n31090 , n42332 );
and ( n77541 , n31094 , n42334 );
and ( n77542 , n31098 , n42336 );
and ( n77543 , n31101 , n42338 );
and ( n77544 , n31105 , n42340 );
and ( n77545 , n31108 , n42342 );
and ( n77546 , n31111 , n42344 );
and ( n77547 , n31114 , n42346 );
and ( n77548 , n31117 , n42348 );
and ( n77549 , n31120 , n42350 );
and ( n77550 , n31123 , n42352 );
and ( n77551 , n31126 , n42354 );
and ( n77552 , n31129 , n42356 );
and ( n77553 , n31132 , n42358 );
and ( n77554 , n31135 , n42360 );
or ( n77555 , n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , n77551 , n77552 , n77553 , n77554 );
and ( n77556 , n77555 , n39979 );
or ( n77557 , n77538 , n77556 );
and ( n77558 , n77557 , n31538 );
and ( n77559 , n34054 , n40143 );
or ( n77560 , n77536 , n77558 , n77559 );
and ( n77561 , n77560 , n31557 );
and ( n77562 , n34054 , n40154 );
or ( n77563 , C0 , n77561 , n77562 );
buf ( n77564 , n77563 );
buf ( n77565 , n77564 );
buf ( n77566 , n31655 );
buf ( n77567 , n48547 );
buf ( n77568 , n30987 );
and ( n77569 , n50953 , n72973 );
xor ( n77570 , n50951 , n77569 );
and ( n77571 , n77570 , n32431 );
not ( n77572 , n50002 );
and ( n77573 , n77572 , n50951 );
and ( n77574 , n40571 , n50002 );
or ( n77575 , n77573 , n77574 );
and ( n77576 , n77575 , n32419 );
not ( n77577 , n50008 );
and ( n77578 , n77577 , n50951 );
not ( n77579 , n51594 );
and ( n77580 , n77579 , n51566 );
xor ( n77581 , n59225 , n59236 );
and ( n77582 , n77581 , n51594 );
or ( n77583 , n77580 , n77582 );
and ( n77584 , n77583 , n50008 );
or ( n77585 , n77578 , n77584 );
and ( n77586 , n77585 , n32415 );
not ( n77587 , n50067 );
and ( n77588 , n77587 , n50951 );
and ( n77589 , n60416 , n72993 );
xor ( n77590 , n60399 , n77589 );
and ( n77591 , n77590 , n50067 );
or ( n77592 , n77588 , n77591 );
and ( n77593 , n77592 , n32411 );
and ( n77594 , n50951 , n50098 );
or ( n77595 , n77571 , n77576 , n77586 , n77593 , n77594 );
and ( n77596 , n77595 , n32456 );
and ( n77597 , n50951 , n47409 );
or ( n77598 , C0 , n77596 , n77597 );
buf ( n77599 , n77598 );
buf ( n77600 , n77599 );
buf ( n77601 , n31655 );
not ( n77602 , n46356 );
and ( n77603 , n77602 , n31262 );
not ( n77604 , n56904 );
and ( n77605 , n77604 , n31262 );
and ( n77606 , n31272 , n56904 );
or ( n77607 , n77605 , n77606 );
and ( n77608 , n77607 , n46356 );
or ( n77609 , n77603 , n77608 );
and ( n77610 , n77609 , n31649 );
not ( n77611 , n56912 );
not ( n77612 , n56904 );
and ( n77613 , n77612 , n31262 );
and ( n77614 , n49443 , n56904 );
or ( n77615 , n77613 , n77614 );
and ( n77616 , n77611 , n77615 );
and ( n77617 , n49443 , n56912 );
or ( n77618 , n77616 , n77617 );
and ( n77619 , n77618 , n31643 );
not ( n77620 , n31452 );
not ( n77621 , n56912 );
not ( n77622 , n56904 );
and ( n77623 , n77622 , n31262 );
and ( n77624 , n49443 , n56904 );
or ( n77625 , n77623 , n77624 );
and ( n77626 , n77621 , n77625 );
and ( n77627 , n49443 , n56912 );
or ( n77628 , n77626 , n77627 );
and ( n77629 , n77620 , n77628 );
not ( n77630 , n56937 );
not ( n77631 , n56939 );
and ( n77632 , n77631 , n77628 );
and ( n77633 , n49469 , n56939 );
or ( n77634 , n77632 , n77633 );
and ( n77635 , n77630 , n77634 );
and ( n77636 , n49477 , n56937 );
or ( n77637 , n77635 , n77636 );
and ( n77638 , n77637 , n31452 );
or ( n77639 , n77629 , n77638 );
and ( n77640 , n77639 , n31638 );
and ( n77641 , n31262 , n47277 );
or ( n77642 , C0 , n77610 , n77619 , n77640 , n77641 );
buf ( n77643 , n77642 );
buf ( n77644 , n77643 );
buf ( n77645 , n31655 );
buf ( n77646 , n30987 );
not ( n77647 , n32953 );
buf ( n77648 , RI15b46158_256);
and ( n77649 , n77647 , n77648 );
not ( n77650 , n54581 );
and ( n77651 , n77650 , n54373 );
xor ( n77652 , n64020 , n64021 );
and ( n77653 , n77652 , n54581 );
or ( n77654 , n77651 , n77653 );
and ( n77655 , n77654 , n32953 );
or ( n77656 , n77649 , n77655 );
and ( n77657 , n77656 , n33038 );
not ( n77658 , n48660 );
and ( n77659 , n77658 , n77648 );
not ( n77660 , n55168 );
and ( n77661 , n77660 , n55020 );
xor ( n77662 , n55174 , n55178 );
and ( n77663 , n77662 , n55168 );
or ( n77664 , n77661 , n77663 );
and ( n77665 , n77664 , n48660 );
or ( n77666 , n77659 , n77665 );
and ( n77667 , n77666 , n33172 );
and ( n77668 , n77648 , n39795 );
or ( n77669 , n77657 , n77667 , n77668 );
and ( n77670 , n77669 , n33208 );
and ( n77671 , n77648 , n39805 );
or ( n77672 , C0 , n77670 , n77671 );
buf ( n77673 , n77672 );
buf ( n77674 , n77673 );
buf ( n77675 , n30987 );
buf ( n77676 , n31655 );
and ( n77677 , n69733 , n32494 );
not ( n77678 , n46083 );
buf ( n77679 , RI15b5fc70_1133);
and ( n77680 , n77678 , n77679 );
and ( n77681 , n69739 , n46083 );
or ( n77682 , n77680 , n77681 );
and ( n77683 , n77682 , n32421 );
not ( n77684 , n46326 );
and ( n77685 , n77684 , n77679 );
and ( n77686 , n69739 , n46326 );
or ( n77687 , n77685 , n77686 );
and ( n77688 , n77687 , n32417 );
and ( n77689 , n77679 , n46340 );
or ( n77690 , n77683 , n77688 , n77689 );
and ( n77691 , n77690 , n32456 );
and ( n77692 , n77679 , n46349 );
or ( n77693 , C0 , n77677 , n77691 , n77692 );
buf ( n77694 , n77693 );
buf ( n77695 , n77694 );
buf ( n77696 , n31655 );
buf ( n77697 , n30987 );
not ( n77698 , n46356 );
and ( n77699 , n77698 , n31246 );
not ( n77700 , n46362 );
and ( n77701 , n77700 , n31246 );
and ( n77702 , n31272 , n46362 );
or ( n77703 , n77701 , n77702 );
and ( n77704 , n77703 , n46356 );
or ( n77705 , n77699 , n77704 );
and ( n77706 , n77705 , n31649 );
not ( n77707 , n46393 );
not ( n77708 , n46362 );
and ( n77709 , n77708 , n31246 );
and ( n77710 , n49443 , n46362 );
or ( n77711 , n77709 , n77710 );
and ( n77712 , n77707 , n77711 );
and ( n77713 , n49443 , n46393 );
or ( n77714 , n77712 , n77713 );
and ( n77715 , n77714 , n31643 );
not ( n77716 , n31452 );
not ( n77717 , n46393 );
not ( n77718 , n46362 );
and ( n77719 , n77718 , n31246 );
and ( n77720 , n49443 , n46362 );
or ( n77721 , n77719 , n77720 );
and ( n77722 , n77717 , n77721 );
and ( n77723 , n49443 , n46393 );
or ( n77724 , n77722 , n77723 );
and ( n77725 , n77716 , n77724 );
not ( n77726 , n46550 );
not ( n77727 , n46554 );
and ( n77728 , n77727 , n77724 );
and ( n77729 , n49469 , n46554 );
or ( n77730 , n77728 , n77729 );
and ( n77731 , n77726 , n77730 );
and ( n77732 , n49477 , n46550 );
or ( n77733 , n77731 , n77732 );
and ( n77734 , n77733 , n31452 );
or ( n77735 , n77725 , n77734 );
and ( n77736 , n77735 , n31638 );
and ( n77737 , n31246 , n47277 );
or ( n77738 , C0 , n77706 , n77715 , n77736 , n77737 );
buf ( n77739 , n77738 );
buf ( n77740 , n77739 );
buf ( n77741 , n31655 );
not ( n77742 , n31077 );
and ( n77743 , n58919 , n77742 );
and ( n77744 , n77743 , n31373 );
not ( n77745 , n31402 );
and ( n77746 , n58919 , n77745 );
and ( n77747 , n77746 , n31408 );
not ( n77748 , n31437 );
and ( n77749 , n58919 , n77748 );
and ( n77750 , n77749 , n31468 );
not ( n77751 , n31497 );
and ( n77752 , n58919 , n77751 );
and ( n77753 , n77752 , n31521 );
and ( n77754 , n58919 , n31553 );
or ( n77755 , n77744 , n77747 , n77750 , n77753 , n77754 );
and ( n77756 , n77755 , n31557 );
buf ( n77757 , n31640 );
or ( n77758 , n33973 , n31638 );
or ( n77759 , n77758 , n31641 );
or ( n77760 , n77759 , n31643 );
or ( n77761 , n77760 , n31645 );
or ( n77762 , n77761 , n31647 );
or ( n77763 , n77762 , n31649 );
or ( n77764 , n77763 , n31007 );
and ( n77765 , n58919 , n77764 );
or ( n77766 , C0 , n77756 , n77757 , n77765 );
buf ( n77767 , n77766 );
buf ( n77768 , n77767 );
buf ( n77769 , n30987 );
buf ( n77770 , n30987 );
not ( n77771 , n40163 );
and ( n77772 , n77771 , n31943 );
not ( n77773 , n52903 );
and ( n77774 , n77773 , n31943 );
and ( n77775 , n32183 , n52903 );
or ( n77776 , n77774 , n77775 );
and ( n77777 , n77776 , n40163 );
or ( n77778 , n77772 , n77777 );
and ( n77779 , n77778 , n32498 );
not ( n77780 , n52911 );
not ( n77781 , n52903 );
and ( n77782 , n77781 , n31943 );
and ( n77783 , n45178 , n52903 );
or ( n77784 , n77782 , n77783 );
and ( n77785 , n77780 , n77784 );
and ( n77786 , n45178 , n52911 );
or ( n77787 , n77785 , n77786 );
and ( n77788 , n77787 , n32473 );
not ( n77789 , n32475 );
not ( n77790 , n52911 );
not ( n77791 , n52903 );
and ( n77792 , n77791 , n31943 );
and ( n77793 , n45178 , n52903 );
or ( n77794 , n77792 , n77793 );
and ( n77795 , n77790 , n77794 );
and ( n77796 , n45178 , n52911 );
or ( n77797 , n77795 , n77796 );
and ( n77798 , n77789 , n77797 );
not ( n77799 , n52931 );
not ( n77800 , n52933 );
and ( n77801 , n77800 , n77797 );
and ( n77802 , n45206 , n52933 );
or ( n77803 , n77801 , n77802 );
and ( n77804 , n77799 , n77803 );
and ( n77805 , n45214 , n52931 );
or ( n77806 , n77804 , n77805 );
and ( n77807 , n77806 , n32475 );
or ( n77808 , n77798 , n77807 );
and ( n77809 , n77808 , n32486 );
and ( n77810 , n31943 , n41278 );
or ( n77811 , C0 , n77779 , n77788 , n77809 , n77810 );
buf ( n77812 , n77811 );
buf ( n77813 , n77812 );
buf ( n77814 , n31655 );
buf ( n77815 , n31655 );
buf ( n77816 , n30987 );
not ( n77817 , n32598 );
and ( n77818 , n69147 , n77817 );
and ( n77819 , n77818 , n32890 );
not ( n77820 , n32919 );
and ( n77821 , n69147 , n77820 );
and ( n77822 , n77821 , n32924 );
not ( n77823 , n32953 );
and ( n77824 , n69147 , n77823 );
and ( n77825 , n77824 , n33038 );
not ( n77826 , n33067 );
and ( n77827 , n69147 , n77826 );
and ( n77828 , n77827 , n33172 );
and ( n77829 , n69147 , n33204 );
or ( n77830 , n77819 , n77822 , n77825 , n77828 , n77829 );
and ( n77831 , n77830 , n33208 );
buf ( n77832 , n33372 );
or ( n77833 , n35056 , n33370 );
or ( n77834 , n77833 , n33373 );
or ( n77835 , n77834 , n33375 );
or ( n77836 , n77835 , n33377 );
or ( n77837 , n77836 , n33379 );
or ( n77838 , n77837 , n33381 );
or ( n77839 , n77838 , n32528 );
and ( n77840 , n69147 , n77839 );
or ( n77841 , C0 , n77831 , n77832 , n77840 );
buf ( n77842 , n77841 );
buf ( n77843 , n77842 );
buf ( n77844 , n30987 );
buf ( n77845 , n31655 );
not ( n77846 , n46356 );
and ( n77847 , n77846 , n31331 );
not ( n77848 , n49427 );
and ( n77849 , n77848 , n31331 );
and ( n77850 , n31339 , n49427 );
or ( n77851 , n77849 , n77850 );
and ( n77852 , n77851 , n46356 );
or ( n77853 , n77847 , n77852 );
and ( n77854 , n77853 , n31649 );
not ( n77855 , n49435 );
not ( n77856 , n49427 );
and ( n77857 , n77856 , n31331 );
and ( n77858 , n47449 , n49427 );
or ( n77859 , n77857 , n77858 );
and ( n77860 , n77855 , n77859 );
and ( n77861 , n47449 , n49435 );
or ( n77862 , n77860 , n77861 );
and ( n77863 , n77862 , n31643 );
not ( n77864 , n31452 );
not ( n77865 , n49435 );
not ( n77866 , n49427 );
and ( n77867 , n77866 , n31331 );
and ( n77868 , n47449 , n49427 );
or ( n77869 , n77867 , n77868 );
and ( n77870 , n77865 , n77869 );
and ( n77871 , n47449 , n49435 );
or ( n77872 , n77870 , n77871 );
and ( n77873 , n77864 , n77872 );
not ( n77874 , n49460 );
not ( n77875 , n49462 );
and ( n77876 , n77875 , n77872 );
and ( n77877 , n47485 , n49462 );
or ( n77878 , n77876 , n77877 );
and ( n77879 , n77874 , n77878 );
and ( n77880 , n47503 , n49460 );
or ( n77881 , n77879 , n77880 );
and ( n77882 , n77881 , n31452 );
or ( n77883 , n77873 , n77882 );
and ( n77884 , n77883 , n31638 );
and ( n77885 , n31331 , n47277 );
or ( n77886 , C0 , n77854 , n77863 , n77884 , n77885 );
buf ( n77887 , n77886 );
buf ( n77888 , n77887 );
buf ( n77889 , n40209 );
buf ( n77890 , n31655 );
xor ( n77891 , n45984 , n47291 );
and ( n77892 , n77891 , n32433 );
not ( n77893 , n47331 );
and ( n77894 , n77893 , n45984 );
buf ( n77895 , n31996 );
and ( n77896 , n77895 , n47331 );
or ( n77897 , n77894 , n77896 );
and ( n77898 , n77897 , n32413 );
and ( n77899 , n45984 , n47402 );
or ( n77900 , n77892 , n77898 , n77899 );
and ( n77901 , n77900 , n32456 );
and ( n77902 , n45984 , n47409 );
or ( n77903 , C0 , n77901 , n77902 );
buf ( n77904 , n77903 );
buf ( n77905 , n77904 );
buf ( n77906 , n31655 );
buf ( n77907 , n30987 );
buf ( n77908 , n30987 );
buf ( n77909 , n30987 );
xor ( n77910 , n41704 , n44783 );
and ( n77911 , n77910 , n31548 );
not ( n77912 , n44807 );
and ( n77913 , n77912 , n41704 );
and ( n77914 , n41998 , n44807 );
or ( n77915 , n77913 , n77914 );
and ( n77916 , n77915 , n31408 );
not ( n77917 , n44817 );
and ( n77918 , n77917 , n41704 );
not ( n77919 , n41835 );
and ( n77920 , n77919 , n41604 );
and ( n77921 , n42146 , n41835 );
or ( n77922 , n77920 , n77921 );
and ( n77923 , n77922 , n44817 );
or ( n77924 , n77918 , n77923 );
and ( n77925 , n77924 , n31521 );
not ( n77926 , n45059 );
and ( n77927 , n77926 , n41704 );
and ( n77928 , n77555 , n45059 );
or ( n77929 , n77927 , n77928 );
and ( n77930 , n77929 , n31536 );
and ( n77931 , n41704 , n45148 );
or ( n77932 , n77911 , n77916 , n77925 , n77930 , n77931 );
and ( n77933 , n77932 , n31557 );
and ( n77934 , n41704 , n40154 );
or ( n77935 , C0 , n77933 , n77934 );
buf ( n77936 , n77935 );
buf ( n77937 , n77936 );
buf ( n77938 , n31655 );
not ( n77939 , n40163 );
and ( n77940 , n77939 , n32052 );
not ( n77941 , n50540 );
and ( n77942 , n77941 , n32052 );
and ( n77943 , n32130 , n50540 );
or ( n77944 , n77942 , n77943 );
and ( n77945 , n77944 , n40163 );
or ( n77946 , n77940 , n77945 );
and ( n77947 , n77946 , n32498 );
not ( n77948 , n50548 );
not ( n77949 , n50540 );
and ( n77950 , n77949 , n32052 );
and ( n77951 , n45833 , n50540 );
or ( n77952 , n77950 , n77951 );
and ( n77953 , n77948 , n77952 );
and ( n77954 , n45833 , n50548 );
or ( n77955 , n77953 , n77954 );
and ( n77956 , n77955 , n32473 );
not ( n77957 , n32475 );
not ( n77958 , n50548 );
not ( n77959 , n50540 );
and ( n77960 , n77959 , n32052 );
and ( n77961 , n45833 , n50540 );
or ( n77962 , n77960 , n77961 );
and ( n77963 , n77958 , n77962 );
and ( n77964 , n45833 , n50548 );
or ( n77965 , n77963 , n77964 );
and ( n77966 , n77957 , n77965 );
not ( n77967 , n50568 );
not ( n77968 , n50570 );
and ( n77969 , n77968 , n77965 );
and ( n77970 , n45857 , n50570 );
or ( n77971 , n77969 , n77970 );
and ( n77972 , n77967 , n77971 );
and ( n77973 , n45865 , n50568 );
or ( n77974 , n77972 , n77973 );
and ( n77975 , n77974 , n32475 );
or ( n77976 , n77966 , n77975 );
and ( n77977 , n77976 , n32486 );
and ( n77978 , n32052 , n41278 );
or ( n77979 , C0 , n77947 , n77956 , n77977 , n77978 );
buf ( n77980 , n77979 );
buf ( n77981 , n77980 );
xor ( n77982 , n35443 , n39942 );
and ( n77983 , n77982 , n31550 );
not ( n77984 , n39979 );
and ( n77985 , n77984 , n35443 );
and ( n77986 , n31240 , n40095 );
and ( n77987 , n31242 , n40097 );
and ( n77988 , n31244 , n40099 );
and ( n77989 , n31246 , n40101 );
and ( n77990 , n31248 , n40103 );
and ( n77991 , n31250 , n40105 );
and ( n77992 , n31252 , n40107 );
and ( n77993 , n31254 , n40109 );
and ( n77994 , n31256 , n40111 );
and ( n77995 , n31258 , n40113 );
and ( n77996 , n31260 , n40115 );
and ( n77997 , n31262 , n40117 );
and ( n77998 , n31264 , n40119 );
and ( n77999 , n31266 , n40121 );
and ( n78000 , n31268 , n40123 );
and ( n78001 , n31270 , n40125 );
or ( n78002 , n77986 , n77987 , n77988 , n77989 , n77990 , n77991 , n77992 , n77993 , n77994 , n77995 , n77996 , n77997 , n77998 , n77999 , n78000 , n78001 );
and ( n78003 , n78002 , n39979 );
or ( n78004 , n77985 , n78003 );
and ( n78005 , n78004 , n31538 );
and ( n78006 , n35443 , n40143 );
or ( n78007 , n77983 , n78005 , n78006 );
and ( n78008 , n78007 , n31557 );
and ( n78009 , n35443 , n40154 );
or ( n78010 , C0 , n78008 , n78009 );
buf ( n78011 , n78010 );
buf ( n78012 , n78011 );
buf ( n78013 , n54078 );
buf ( n78014 , n31655 );
not ( n78015 , n40163 );
and ( n78016 , n78015 , n31924 );
not ( n78017 , n75905 );
and ( n78018 , n78017 , n31924 );
and ( n78019 , n32200 , n75905 );
or ( n78020 , n78018 , n78019 );
and ( n78021 , n78020 , n40163 );
or ( n78022 , n78016 , n78021 );
and ( n78023 , n78022 , n32498 );
not ( n78024 , n75913 );
not ( n78025 , n75905 );
and ( n78026 , n78025 , n31924 );
and ( n78027 , n53243 , n75905 );
or ( n78028 , n78026 , n78027 );
and ( n78029 , n78024 , n78028 );
and ( n78030 , n53243 , n75913 );
or ( n78031 , n78029 , n78030 );
and ( n78032 , n78031 , n32473 );
not ( n78033 , n32475 );
not ( n78034 , n75913 );
not ( n78035 , n75905 );
and ( n78036 , n78035 , n31924 );
and ( n78037 , n53243 , n75905 );
or ( n78038 , n78036 , n78037 );
and ( n78039 , n78034 , n78038 );
and ( n78040 , n53243 , n75913 );
or ( n78041 , n78039 , n78040 );
and ( n78042 , n78033 , n78041 );
not ( n78043 , n75933 );
not ( n78044 , n75935 );
and ( n78045 , n78044 , n78041 );
and ( n78046 , n53269 , n75935 );
or ( n78047 , n78045 , n78046 );
and ( n78048 , n78043 , n78047 );
and ( n78049 , n53277 , n75933 );
or ( n78050 , n78048 , n78049 );
and ( n78051 , n78050 , n32475 );
or ( n78052 , n78042 , n78051 );
and ( n78053 , n78052 , n32486 );
and ( n78054 , n31924 , n41278 );
or ( n78055 , C0 , n78023 , n78032 , n78053 , n78054 );
buf ( n78056 , n78055 );
buf ( n78057 , n78056 );
buf ( n78058 , n30987 );
buf ( n78059 , n30987 );
buf ( n78060 , n31655 );
buf ( n78061 , n30987 );
not ( n78062 , n35278 );
and ( n78063 , n78062 , n64567 );
and ( n78064 , n73111 , n35278 );
or ( n78065 , n78063 , n78064 );
and ( n78066 , n78065 , n32417 );
not ( n78067 , n47912 );
and ( n78068 , n78067 , n64567 );
and ( n78069 , n64573 , n47912 );
or ( n78070 , n78068 , n78069 );
and ( n78071 , n78070 , n32415 );
and ( n78072 , n64567 , n48133 );
or ( n78073 , n78066 , n78071 , n78072 );
and ( n78074 , n78073 , n32456 );
and ( n78075 , n64567 , n47409 );
or ( n78076 , C0 , n78074 , n78075 );
buf ( n78077 , n78076 );
buf ( n78078 , n78077 );
not ( n78079 , n46356 );
and ( n78080 , n78079 , n31206 );
not ( n78081 , n63024 );
and ( n78082 , n78081 , n31206 );
and ( n78083 , n31238 , n63024 );
or ( n78084 , n78082 , n78083 );
and ( n78085 , n78084 , n46356 );
or ( n78086 , n78080 , n78085 );
and ( n78087 , n78086 , n31649 );
not ( n78088 , n63032 );
not ( n78089 , n63024 );
and ( n78090 , n78089 , n31206 );
and ( n78091 , n49901 , n63024 );
or ( n78092 , n78090 , n78091 );
and ( n78093 , n78088 , n78092 );
and ( n78094 , n49901 , n63032 );
or ( n78095 , n78093 , n78094 );
and ( n78096 , n78095 , n31643 );
not ( n78097 , n31452 );
not ( n78098 , n63032 );
not ( n78099 , n63024 );
and ( n78100 , n78099 , n31206 );
and ( n78101 , n49901 , n63024 );
or ( n78102 , n78100 , n78101 );
and ( n78103 , n78098 , n78102 );
and ( n78104 , n49901 , n63032 );
or ( n78105 , n78103 , n78104 );
and ( n78106 , n78097 , n78105 );
not ( n78107 , n63052 );
not ( n78108 , n63054 );
and ( n78109 , n78108 , n78105 );
and ( n78110 , n49925 , n63054 );
or ( n78111 , n78109 , n78110 );
and ( n78112 , n78107 , n78111 );
and ( n78113 , n49933 , n63052 );
or ( n78114 , n78112 , n78113 );
and ( n78115 , n78114 , n31452 );
or ( n78116 , n78106 , n78115 );
and ( n78117 , n78116 , n31638 );
and ( n78118 , n31206 , n47277 );
or ( n78119 , C0 , n78087 , n78096 , n78117 , n78118 );
buf ( n78120 , n78119 );
buf ( n78121 , n78120 );
not ( n78122 , n40163 );
and ( n78123 , n78122 , n32062 );
not ( n78124 , n42238 );
and ( n78125 , n78124 , n32062 );
and ( n78126 , n32130 , n42238 );
or ( n78127 , n78125 , n78126 );
and ( n78128 , n78127 , n40163 );
or ( n78129 , n78123 , n78128 );
and ( n78130 , n78129 , n32498 );
not ( n78131 , n42247 );
not ( n78132 , n42238 );
and ( n78133 , n78132 , n32062 );
and ( n78134 , n45833 , n42238 );
or ( n78135 , n78133 , n78134 );
and ( n78136 , n78131 , n78135 );
and ( n78137 , n45833 , n42247 );
or ( n78138 , n78136 , n78137 );
and ( n78139 , n78138 , n32473 );
not ( n78140 , n32475 );
not ( n78141 , n42247 );
not ( n78142 , n42238 );
and ( n78143 , n78142 , n32062 );
and ( n78144 , n45833 , n42238 );
or ( n78145 , n78143 , n78144 );
and ( n78146 , n78141 , n78145 );
and ( n78147 , n45833 , n42247 );
or ( n78148 , n78146 , n78147 );
and ( n78149 , n78140 , n78148 );
not ( n78150 , n42273 );
not ( n78151 , n42276 );
and ( n78152 , n78151 , n78148 );
and ( n78153 , n45857 , n42276 );
or ( n78154 , n78152 , n78153 );
and ( n78155 , n78150 , n78154 );
and ( n78156 , n45865 , n42273 );
or ( n78157 , n78155 , n78156 );
and ( n78158 , n78157 , n32475 );
or ( n78159 , n78149 , n78158 );
and ( n78160 , n78159 , n32486 );
and ( n78161 , n32062 , n41278 );
or ( n78162 , C0 , n78130 , n78139 , n78160 , n78161 );
buf ( n78163 , n78162 );
buf ( n78164 , n78163 );
buf ( n78165 , n31655 );
xor ( n78166 , n34038 , n39938 );
and ( n78167 , n78166 , n31550 );
not ( n78168 , n39979 );
and ( n78169 , n78168 , n34038 );
and ( n78170 , n68670 , n39979 );
or ( n78171 , n78169 , n78170 );
and ( n78172 , n78171 , n31538 );
and ( n78173 , n34038 , n40143 );
or ( n78174 , n78167 , n78172 , n78173 );
and ( n78175 , n78174 , n31557 );
and ( n78176 , n34038 , n40154 );
or ( n78177 , C0 , n78175 , n78176 );
buf ( n78178 , n78177 );
buf ( n78179 , n78178 );
buf ( n78180 , n30987 );
buf ( n78181 , n30987 );
buf ( n78182 , n31655 );
and ( n78183 , n49369 , n31645 );
not ( n78184 , n45274 );
buf ( n78185 , RI15b53a60_719);
and ( n78186 , n78184 , n78185 );
not ( n78187 , n41809 );
and ( n78188 , n78187 , n41805 );
xor ( n78189 , n41805 , n41611 );
and ( n78190 , n62432 , n62439 );
xor ( n78191 , n78189 , n78190 );
and ( n78192 , n78191 , n41809 );
or ( n78193 , n78188 , n78192 );
and ( n78194 , n78193 , n45274 );
or ( n78195 , n78186 , n78194 );
and ( n78196 , n78195 , n31373 );
not ( n78197 , n45280 );
and ( n78198 , n78197 , n78185 );
and ( n78199 , n78193 , n45280 );
or ( n78200 , n78198 , n78199 );
and ( n78201 , n78200 , n31468 );
and ( n78202 , n78185 , n45802 );
or ( n78203 , n78196 , n78201 , n78202 );
and ( n78204 , n78203 , n31557 );
and ( n78205 , n78185 , n45808 );
or ( n78206 , C0 , n78183 , n78204 , n78205 );
buf ( n78207 , n78206 );
buf ( n78208 , n78207 );
not ( n78209 , n40163 );
and ( n78210 , n78209 , n31787 );
not ( n78211 , n54629 );
and ( n78212 , n78211 , n31787 );
and ( n78213 , n32252 , n54629 );
or ( n78214 , n78212 , n78213 );
and ( n78215 , n78214 , n40163 );
or ( n78216 , n78210 , n78215 );
and ( n78217 , n78216 , n32498 );
not ( n78218 , n54637 );
not ( n78219 , n54629 );
and ( n78220 , n78219 , n31787 );
and ( n78221 , n40393 , n54629 );
or ( n78222 , n78220 , n78221 );
and ( n78223 , n78218 , n78222 );
and ( n78224 , n40393 , n54637 );
or ( n78225 , n78223 , n78224 );
and ( n78226 , n78225 , n32473 );
not ( n78227 , n32475 );
not ( n78228 , n54637 );
not ( n78229 , n54629 );
and ( n78230 , n78229 , n31787 );
and ( n78231 , n40393 , n54629 );
or ( n78232 , n78230 , n78231 );
and ( n78233 , n78228 , n78232 );
and ( n78234 , n40393 , n54637 );
or ( n78235 , n78233 , n78234 );
and ( n78236 , n78227 , n78235 );
not ( n78237 , n54657 );
not ( n78238 , n54659 );
and ( n78239 , n78238 , n78235 );
and ( n78240 , n40972 , n54659 );
or ( n78241 , n78239 , n78240 );
and ( n78242 , n78237 , n78241 );
and ( n78243 , n41267 , n54657 );
or ( n78244 , n78242 , n78243 );
and ( n78245 , n78244 , n32475 );
or ( n78246 , n78236 , n78245 );
and ( n78247 , n78246 , n32486 );
and ( n78248 , n31787 , n41278 );
or ( n78249 , C0 , n78217 , n78226 , n78247 , n78248 );
buf ( n78250 , n78249 );
buf ( n78251 , n78250 );
buf ( n78252 , n30987 );
and ( n78253 , n48793 , n34150 );
buf ( n78254 , n78253 );
and ( n78255 , n78254 , n33381 );
and ( n78256 , n56667 , n33379 );
and ( n78257 , n57739 , n33208 );
and ( n78258 , n32547 , n61311 );
or ( n78259 , C0 , n78255 , n78256 , n78257 , n78258 );
buf ( n78260 , n78259 );
buf ( n78261 , n78260 );
buf ( n78262 , n31655 );
buf ( n78263 , n30987 );
buf ( n78264 , n30987 );
buf ( n78265 , n31655 );
not ( n78266 , n50828 );
not ( n78267 , n50834 );
and ( n78268 , n78267 , n40484 );
buf ( n78269 , RI15b538f8_716);
and ( n78270 , n78269 , n50834 );
or ( n78271 , n78268 , n78270 );
and ( n78272 , n78266 , n78271 );
and ( n78273 , n60904 , n50828 );
or ( n78274 , n78272 , n78273 );
buf ( n78275 , n78274 );
buf ( n78276 , n78275 );
buf ( n78277 , n30987 );
xor ( n78278 , n33081 , n58393 );
and ( n78279 , n78278 , n33201 );
not ( n78280 , n41576 );
and ( n78281 , n78280 , n33081 );
xor ( n78282 , n58523 , n58594 );
and ( n78283 , n78282 , n41576 );
or ( n78284 , n78281 , n78283 );
and ( n78285 , n78284 , n33189 );
and ( n78286 , n33081 , n41592 );
or ( n78287 , n78279 , n78285 , n78286 );
and ( n78288 , n78287 , n33208 );
and ( n78289 , n33081 , n39805 );
or ( n78290 , C0 , n78288 , n78289 );
buf ( n78291 , n78290 );
buf ( n78292 , n78291 );
buf ( n78293 , n31655 );
buf ( n78294 , n31655 );
buf ( n78295 , n30987 );
buf ( n78296 , RI15b5eb18_1096);
and ( n78297 , n78296 , n32494 );
not ( n78298 , n46083 );
and ( n78299 , n78298 , n69692 );
buf ( n78300 , n78299 );
and ( n78301 , n78300 , n32421 );
not ( n78302 , n46326 );
and ( n78303 , n78302 , n69692 );
not ( n78304 , n51396 );
and ( n78305 , n78304 , n51222 );
xor ( n78306 , n51401 , n51409 );
and ( n78307 , n78306 , n51396 );
or ( n78308 , n78305 , n78307 );
and ( n78309 , n78308 , n46326 );
or ( n78310 , n78303 , n78309 );
and ( n78311 , n78310 , n32417 );
and ( n78312 , n69692 , n46340 );
or ( n78313 , n78301 , n78311 , n78312 );
and ( n78314 , n78313 , n32456 );
and ( n78315 , n69692 , n46349 );
or ( n78316 , n78297 , n78314 , n78315 );
buf ( n78317 , n78316 );
buf ( n78318 , n78317 );
buf ( n78319 , n31655 );
buf ( n78320 , n30987 );
buf ( n78321 , n31655 );
not ( n78322 , n46356 );
and ( n78323 , n78322 , n31181 );
and ( n78324 , n31025 , n31021 , n48213 , n31013 , n46361 );
not ( n78325 , n78324 );
and ( n78326 , n78325 , n31181 );
and ( n78327 , n31205 , n78324 );
or ( n78328 , n78326 , n78327 );
and ( n78329 , n78328 , n46356 );
or ( n78330 , n78323 , n78329 );
and ( n78331 , n78330 , n31649 );
and ( n78332 , n46373 , n46379 , n48222 , n46392 );
not ( n78333 , n78332 );
not ( n78334 , n78324 );
and ( n78335 , n78334 , n31181 );
and ( n78336 , n50125 , n78324 );
or ( n78337 , n78335 , n78336 );
and ( n78338 , n78333 , n78337 );
and ( n78339 , n50125 , n78332 );
or ( n78340 , n78338 , n78339 );
and ( n78341 , n78340 , n31643 );
not ( n78342 , n31452 );
not ( n78343 , n78332 );
not ( n78344 , n78324 );
and ( n78345 , n78344 , n31181 );
and ( n78346 , n50125 , n78324 );
or ( n78347 , n78345 , n78346 );
and ( n78348 , n78343 , n78347 );
and ( n78349 , n50125 , n78332 );
or ( n78350 , n78348 , n78349 );
and ( n78351 , n78342 , n78350 );
and ( n78352 , n46519 , n46528 , n48243 , n46549 );
not ( n78353 , n78352 );
and ( n78354 , n46515 , n46524 , n48246 , n46544 );
not ( n78355 , n78354 );
and ( n78356 , n78355 , n78350 );
and ( n78357 , n50151 , n78354 );
or ( n78358 , n78356 , n78357 );
and ( n78359 , n78353 , n78358 );
and ( n78360 , n50159 , n78352 );
or ( n78361 , n78359 , n78360 );
and ( n78362 , n78361 , n31452 );
or ( n78363 , n78351 , n78362 );
and ( n78364 , n78363 , n31638 );
and ( n78365 , n31181 , n47277 );
or ( n78366 , n78331 , n78341 , n78364 , n78365 );
buf ( n78367 , n78366 );
buf ( n78368 , n78367 );
not ( n78369 , n41532 );
and ( n78370 , n78369 , n34375 );
and ( n78371 , n53290 , n41532 );
or ( n78372 , n78370 , n78371 );
buf ( n78373 , n78372 );
buf ( n78374 , n78373 );
buf ( n78375 , n31655 );
buf ( n78376 , n31655 );
buf ( n78377 , n30987 );
buf ( n78378 , n30987 );
and ( n78379 , n54150 , n54984 );
and ( n78380 , n54148 , n78379 );
and ( n78381 , n54146 , n78380 );
and ( n78382 , n54144 , n78381 );
and ( n78383 , n54142 , n78382 );
and ( n78384 , n54140 , n78383 );
and ( n78385 , n54138 , n78384 );
xor ( n78386 , n54136 , n78385 );
and ( n78387 , n78386 , n33199 );
not ( n78388 , n48648 );
and ( n78389 , n78388 , n54136 );
and ( n78390 , n34421 , n48648 );
or ( n78391 , n78389 , n78390 );
and ( n78392 , n78391 , n32924 );
not ( n78393 , n48660 );
and ( n78394 , n78393 , n54136 );
and ( n78395 , n73941 , n48660 );
or ( n78396 , n78394 , n78395 );
and ( n78397 , n78396 , n33172 );
not ( n78398 , n48730 );
and ( n78399 , n78398 , n54136 );
and ( n78400 , n58574 , n58591 );
and ( n78401 , n58557 , n78400 );
and ( n78402 , n58540 , n78401 );
and ( n78403 , n58523 , n78402 );
and ( n78404 , n58506 , n78403 );
xor ( n78405 , n58489 , n78404 );
and ( n78406 , n78405 , n48730 );
or ( n78407 , n78399 , n78406 );
and ( n78408 , n78407 , n33187 );
and ( n78409 , n54136 , n54713 );
or ( n78410 , n78387 , n78392 , n78397 , n78408 , n78409 );
and ( n78411 , n78410 , n33208 );
and ( n78412 , n54136 , n39805 );
or ( n78413 , C0 , n78411 , n78412 );
buf ( n78414 , n78413 );
buf ( n78415 , n78414 );
and ( n78416 , n49063 , n48639 );
not ( n78417 , n48642 );
and ( n78418 , n78417 , n48588 );
and ( n78419 , n49063 , n48642 );
or ( n78420 , n78418 , n78419 );
and ( n78421 , n78420 , n32890 );
not ( n78422 , n48648 );
and ( n78423 , n78422 , n48588 );
and ( n78424 , n49063 , n48648 );
or ( n78425 , n78423 , n78424 );
and ( n78426 , n78425 , n32924 );
not ( n78427 , n48654 );
and ( n78428 , n78427 , n48588 );
and ( n78429 , n49063 , n48654 );
or ( n78430 , n78428 , n78429 );
and ( n78431 , n78430 , n33038 );
not ( n78432 , n48660 );
and ( n78433 , n78432 , n48588 );
and ( n78434 , n49063 , n48660 );
or ( n78435 , n78433 , n78434 );
and ( n78436 , n78435 , n33172 );
not ( n78437 , n41576 );
and ( n78438 , n78437 , n48588 );
and ( n78439 , n48773 , n41576 );
or ( n78440 , n78438 , n78439 );
and ( n78441 , n78440 , n33189 );
not ( n78442 , n48730 );
and ( n78443 , n78442 , n48588 );
and ( n78444 , n48773 , n48730 );
or ( n78445 , n78443 , n78444 );
and ( n78446 , n78445 , n33187 );
not ( n78447 , n48765 );
and ( n78448 , n78447 , n48588 );
xor ( n78449 , n48773 , n49015 );
and ( n78450 , n78449 , n48765 );
or ( n78451 , n78448 , n78450 );
and ( n78452 , n78451 , n33180 );
not ( n78453 , n49054 );
and ( n78454 , n78453 , n48588 );
not ( n78455 , n48845 );
xor ( n78456 , n49063 , n49129 );
and ( n78457 , n78455 , n78456 );
xnor ( n78458 , n49172 , n49255 );
and ( n78459 , n78458 , n48845 );
or ( n78460 , n78457 , n78459 );
and ( n78461 , n78460 , n49054 );
or ( n78462 , n78454 , n78461 );
and ( n78463 , n78462 , n33178 );
and ( n78464 , n49172 , n49275 );
or ( n78465 , n78416 , n78421 , n78426 , n78431 , n78436 , n78441 , n78446 , n78452 , n78463 , n78464 );
and ( n78466 , n78465 , n33208 );
and ( n78467 , n32981 , n35056 );
and ( n78468 , n48588 , n49286 );
or ( n78469 , C0 , n78466 , n78467 , n78468 );
buf ( n78470 , n78469 );
buf ( n78471 , n78470 );
buf ( n78472 , n30987 );
buf ( n78473 , n31655 );
buf ( n78474 , n31655 );
buf ( n78475 , n30987 );
buf ( n78476 , n31655 );
not ( n78477 , n46356 );
and ( n78478 , n78477 , n31111 );
not ( n78479 , n48214 );
and ( n78480 , n78479 , n31111 );
and ( n78481 , n31138 , n48214 );
or ( n78482 , n78480 , n78481 );
and ( n78483 , n78482 , n46356 );
or ( n78484 , n78478 , n78483 );
and ( n78485 , n78484 , n31649 );
not ( n78486 , n48223 );
not ( n78487 , n48214 );
and ( n78488 , n78487 , n31111 );
and ( n78489 , n56920 , n48214 );
or ( n78490 , n78488 , n78489 );
and ( n78491 , n78486 , n78490 );
and ( n78492 , n56920 , n48223 );
or ( n78493 , n78491 , n78492 );
and ( n78494 , n78493 , n31643 );
not ( n78495 , n31452 );
not ( n78496 , n48223 );
not ( n78497 , n48214 );
and ( n78498 , n78497 , n31111 );
and ( n78499 , n56920 , n48214 );
or ( n78500 , n78498 , n78499 );
and ( n78501 , n78496 , n78500 );
and ( n78502 , n56920 , n48223 );
or ( n78503 , n78501 , n78502 );
and ( n78504 , n78495 , n78503 );
not ( n78505 , n48244 );
not ( n78506 , n48247 );
and ( n78507 , n78506 , n78503 );
and ( n78508 , n56946 , n48247 );
or ( n78509 , n78507 , n78508 );
and ( n78510 , n78505 , n78509 );
and ( n78511 , n56954 , n48244 );
or ( n78512 , n78510 , n78511 );
and ( n78513 , n78512 , n31452 );
or ( n78514 , n78504 , n78513 );
and ( n78515 , n78514 , n31638 );
and ( n78516 , n31111 , n47277 );
or ( n78517 , C0 , n78485 , n78494 , n78515 , n78516 );
buf ( n78518 , n78517 );
buf ( n78519 , n78518 );
buf ( n78520 , n30987 );
not ( n78521 , n46087 );
and ( n78522 , n78521 , n32431 );
not ( n78523 , n50002 );
and ( n78524 , n78523 , n46087 );
and ( n78525 , n40234 , n50002 );
or ( n78526 , n78524 , n78525 );
and ( n78527 , n78526 , n32419 );
not ( n78528 , n50008 );
and ( n78529 , n78528 , n46087 );
not ( n78530 , n47910 );
buf ( n78531 , RI15b5f040_1107);
and ( n78532 , n78530 , n78531 );
not ( n78533 , n48101 );
and ( n78534 , n78533 , n47918 );
xor ( n78535 , n48111 , n40244 );
and ( n78536 , n78535 , n48101 );
or ( n78537 , n78534 , n78536 );
and ( n78538 , n78537 , n47910 );
or ( n78539 , n78532 , n78538 );
and ( n78540 , n78539 , n50008 );
or ( n78541 , n78529 , n78540 );
and ( n78542 , n78541 , n32415 );
not ( n78543 , n50067 );
and ( n78544 , n78543 , n46087 );
and ( n78545 , n32068 , n50067 );
or ( n78546 , n78544 , n78545 );
and ( n78547 , n78546 , n32411 );
and ( n78548 , n46087 , n50098 );
or ( n78549 , n78522 , n78527 , n78542 , n78547 , n78548 );
and ( n78550 , n78549 , n32456 );
and ( n78551 , n46087 , n47409 );
or ( n78552 , C0 , n78550 , n78551 );
buf ( n78553 , n78552 );
buf ( n78554 , n78553 );
buf ( n78555 , n31655 );
not ( n78556 , n48765 );
and ( n78557 , n78556 , n33333 );
and ( n78558 , n61384 , n48765 );
or ( n78559 , n78557 , n78558 );
and ( n78560 , n78559 , n33180 );
not ( n78561 , n49054 );
and ( n78562 , n78561 , n33333 );
and ( n78563 , n61395 , n49054 );
or ( n78564 , n78562 , n78563 );
and ( n78565 , n78564 , n33178 );
and ( n78566 , n33333 , n49774 );
or ( n78567 , n78560 , n78565 , n78566 );
and ( n78568 , n78567 , n33208 );
and ( n78569 , n33333 , n33375 );
buf ( n78570 , n33333 );
and ( n78571 , n78570 , n33370 );
and ( n78572 , n42695 , n35056 );
and ( n78573 , n33333 , n49794 );
or ( n78574 , C0 , n78568 , n78569 , n78571 , n78572 , n78573 );
buf ( n78575 , n78574 );
buf ( n78576 , n78575 );
buf ( n78577 , n30987 );
not ( n78578 , n50828 );
not ( n78579 , n50834 );
and ( n78580 , n78579 , n40339 );
and ( n78581 , n65190 , n50834 );
or ( n78582 , n78580 , n78581 );
and ( n78583 , n78578 , n78582 );
and ( n78584 , n75729 , n50828 );
or ( n78585 , n78583 , n78584 );
buf ( n78586 , n78585 );
buf ( n78587 , n78586 );
buf ( n78588 , n31655 );
buf ( n78589 , n31655 );
buf ( n78590 , n30987 );
buf ( n78591 , n31655 );
buf ( n78592 , n30987 );
and ( n78593 , n54136 , n78385 );
xor ( n78594 , n54134 , n78593 );
and ( n78595 , n78594 , n33199 );
not ( n78596 , n48648 );
and ( n78597 , n78596 , n54134 );
and ( n78598 , n34419 , n48648 );
or ( n78599 , n78597 , n78598 );
and ( n78600 , n78599 , n32924 );
not ( n78601 , n48660 );
and ( n78602 , n78601 , n54134 );
not ( n78603 , n55168 );
and ( n78604 , n78603 , n55152 );
xor ( n78605 , n55152 , n34193 );
and ( n78606 , n73937 , n73938 );
xor ( n78607 , n78605 , n78606 );
and ( n78608 , n78607 , n55168 );
or ( n78609 , n78604 , n78608 );
and ( n78610 , n78609 , n48660 );
or ( n78611 , n78602 , n78610 );
and ( n78612 , n78611 , n33172 );
not ( n78613 , n48730 );
and ( n78614 , n78613 , n54134 );
and ( n78615 , n58489 , n78404 );
xor ( n78616 , n58472 , n78615 );
and ( n78617 , n78616 , n48730 );
or ( n78618 , n78614 , n78617 );
and ( n78619 , n78618 , n33187 );
and ( n78620 , n54134 , n54713 );
or ( n78621 , n78595 , n78600 , n78612 , n78619 , n78620 );
and ( n78622 , n78621 , n33208 );
and ( n78623 , n54134 , n39805 );
or ( n78624 , C0 , n78622 , n78623 );
buf ( n78625 , n78624 );
buf ( n78626 , n78625 );
not ( n78627 , n41532 );
and ( n78628 , n78627 , n34377 );
and ( n78629 , n74194 , n41532 );
or ( n78630 , n78628 , n78629 );
buf ( n78631 , n78630 );
buf ( n78632 , n78631 );
buf ( n78633 , n30987 );
buf ( n78634 , n31655 );
and ( n78635 , n32293 , n50275 );
not ( n78636 , n50278 );
and ( n78637 , n78636 , n31732 );
and ( n78638 , n32293 , n50278 );
or ( n78639 , n78637 , n78638 );
and ( n78640 , n78639 , n32421 );
not ( n78641 , n50002 );
and ( n78642 , n78641 , n31732 );
and ( n78643 , n32293 , n50002 );
or ( n78644 , n78642 , n78643 );
and ( n78645 , n78644 , n32419 );
not ( n78646 , n50289 );
and ( n78647 , n78646 , n31732 );
and ( n78648 , n32293 , n50289 );
or ( n78649 , n78647 , n78648 );
and ( n78650 , n78649 , n32417 );
not ( n78651 , n50008 );
and ( n78652 , n78651 , n31732 );
and ( n78653 , n32293 , n50008 );
or ( n78654 , n78652 , n78653 );
and ( n78655 , n78654 , n32415 );
not ( n78656 , n47331 );
and ( n78657 , n78656 , n31732 );
and ( n78658 , n31748 , n47331 );
or ( n78659 , n78657 , n78658 );
and ( n78660 , n78659 , n32413 );
not ( n78661 , n50067 );
and ( n78662 , n78661 , n31732 );
and ( n78663 , n31748 , n50067 );
or ( n78664 , n78662 , n78663 );
and ( n78665 , n78664 , n32411 );
not ( n78666 , n31728 );
and ( n78667 , n78666 , n31732 );
and ( n78668 , n32091 , n31728 );
or ( n78669 , n78667 , n78668 );
and ( n78670 , n78669 , n32253 );
not ( n78671 , n32283 );
and ( n78672 , n78671 , n31732 );
and ( n78673 , n32395 , n32283 );
or ( n78674 , n78672 , n78673 );
and ( n78675 , n78674 , n32398 );
and ( n78676 , n32339 , n50334 );
or ( n78677 , n78635 , n78640 , n78645 , n78650 , n78655 , n78660 , n78665 , n78670 , n78675 , n78676 );
and ( n78678 , n78677 , n32456 );
and ( n78679 , n32488 , n32489 );
and ( n78680 , n31732 , n50345 );
or ( n78681 , C0 , n78678 , n78679 , n78680 );
buf ( n78682 , n78681 );
buf ( n78683 , n78682 );
buf ( n78684 , n30987 );
not ( n78685 , n31437 );
buf ( n78686 , RI15b52728_678);
and ( n78687 , n78685 , n78686 );
not ( n78688 , n45766 );
and ( n78689 , n78688 , n45609 );
xor ( n78690 , n45773 , n45783 );
and ( n78691 , n78690 , n45766 );
or ( n78692 , n78689 , n78691 );
and ( n78693 , n78692 , n31437 );
or ( n78694 , n78687 , n78693 );
and ( n78695 , n78694 , n31468 );
not ( n78696 , n44817 );
and ( n78697 , n78696 , n78686 );
and ( n78698 , n55853 , n44817 );
or ( n78699 , n78697 , n78698 );
and ( n78700 , n78699 , n31521 );
and ( n78701 , n78686 , n42158 );
or ( n78702 , n78695 , n78700 , n78701 );
and ( n78703 , n78702 , n31557 );
and ( n78704 , n78686 , n40154 );
or ( n78705 , C0 , n78703 , n78704 );
buf ( n78706 , n78705 );
buf ( n78707 , n78706 );
buf ( n78708 , n31655 );
buf ( n78709 , n31655 );
buf ( n78710 , n30987 );
not ( n78711 , n46356 );
and ( n78712 , n78711 , n31214 );
not ( n78713 , n78324 );
and ( n78714 , n78713 , n31214 );
and ( n78715 , n31238 , n78324 );
or ( n78716 , n78714 , n78715 );
and ( n78717 , n78716 , n46356 );
or ( n78718 , n78712 , n78717 );
and ( n78719 , n78718 , n31649 );
not ( n78720 , n78332 );
not ( n78721 , n78324 );
and ( n78722 , n78721 , n31214 );
and ( n78723 , n49901 , n78324 );
or ( n78724 , n78722 , n78723 );
and ( n78725 , n78720 , n78724 );
and ( n78726 , n49901 , n78332 );
or ( n78727 , n78725 , n78726 );
and ( n78728 , n78727 , n31643 );
not ( n78729 , n31452 );
not ( n78730 , n78332 );
not ( n78731 , n78324 );
and ( n78732 , n78731 , n31214 );
and ( n78733 , n49901 , n78324 );
or ( n78734 , n78732 , n78733 );
and ( n78735 , n78730 , n78734 );
and ( n78736 , n49901 , n78332 );
or ( n78737 , n78735 , n78736 );
and ( n78738 , n78729 , n78737 );
not ( n78739 , n78352 );
not ( n78740 , n78354 );
and ( n78741 , n78740 , n78737 );
and ( n78742 , n49925 , n78354 );
or ( n78743 , n78741 , n78742 );
and ( n78744 , n78739 , n78743 );
and ( n78745 , n49933 , n78352 );
or ( n78746 , n78744 , n78745 );
and ( n78747 , n78746 , n31452 );
or ( n78748 , n78738 , n78747 );
and ( n78749 , n78748 , n31638 );
and ( n78750 , n31214 , n47277 );
or ( n78751 , C0 , n78719 , n78728 , n78749 , n78750 );
buf ( n78752 , n78751 );
buf ( n78753 , n78752 );
buf ( n78754 , n31655 );
buf ( n78755 , RI15b5eaa0_1095);
and ( n78756 , n78755 , n32494 );
not ( n78757 , n46083 );
buf ( n78758 , RI15b600a8_1142);
and ( n78759 , n78757 , n78758 );
buf ( n78760 , n78759 );
and ( n78761 , n78760 , n32421 );
not ( n78762 , n46326 );
and ( n78763 , n78762 , n78758 );
not ( n78764 , n51396 );
and ( n78765 , n78764 , n51205 );
xor ( n78766 , n51402 , n51408 );
and ( n78767 , n78766 , n51396 );
or ( n78768 , n78765 , n78767 );
and ( n78769 , n78768 , n46326 );
or ( n78770 , n78763 , n78769 );
and ( n78771 , n78770 , n32417 );
and ( n78772 , n78758 , n46340 );
or ( n78773 , n78761 , n78771 , n78772 );
and ( n78774 , n78773 , n32456 );
and ( n78775 , n78758 , n46349 );
or ( n78776 , C0 , n78756 , n78774 , n78775 );
buf ( n78777 , n78776 );
buf ( n78778 , n78777 );
not ( n78779 , n35278 );
buf ( n78780 , RI15b5ede8_1102);
and ( n78781 , n78779 , n78780 );
not ( n78782 , n51396 );
and ( n78783 , n78782 , n51324 );
xor ( n78784 , n53328 , n53335 );
and ( n78785 , n78784 , n51396 );
or ( n78786 , n78783 , n78785 );
and ( n78787 , n78786 , n35278 );
or ( n78788 , n78781 , n78787 );
and ( n78789 , n78788 , n32417 );
not ( n78790 , n50008 );
and ( n78791 , n78790 , n78780 );
and ( n78792 , n70054 , n50008 );
or ( n78793 , n78791 , n78792 );
and ( n78794 , n78793 , n32415 );
and ( n78795 , n78780 , n48133 );
or ( n78796 , n78789 , n78794 , n78795 );
and ( n78797 , n78796 , n32456 );
and ( n78798 , n78780 , n47409 );
or ( n78799 , C0 , n78797 , n78798 );
buf ( n78800 , n78799 );
buf ( n78801 , n78800 );
buf ( n78802 , n30987 );
buf ( n78803 , n31655 );
and ( n78804 , n33779 , n48455 );
not ( n78805 , n48457 );
and ( n78806 , n78805 , n33440 );
and ( n78807 , n33779 , n48457 );
or ( n78808 , n78806 , n78807 );
and ( n78809 , n78808 , n31373 );
not ( n78810 , n44807 );
and ( n78811 , n78810 , n33440 );
and ( n78812 , n33779 , n44807 );
or ( n78813 , n78811 , n78812 );
and ( n78814 , n78813 , n31408 );
not ( n78815 , n48468 );
and ( n78816 , n78815 , n33440 );
and ( n78817 , n33779 , n48468 );
or ( n78818 , n78816 , n78817 );
and ( n78819 , n78818 , n31468 );
not ( n78820 , n44817 );
and ( n78821 , n78820 , n33440 );
and ( n78822 , n33779 , n44817 );
or ( n78823 , n78821 , n78822 );
and ( n78824 , n78823 , n31521 );
not ( n78825 , n39979 );
and ( n78826 , n78825 , n33440 );
and ( n78827 , n33592 , n39979 );
or ( n78828 , n78826 , n78827 );
and ( n78829 , n78828 , n31538 );
not ( n78830 , n45059 );
and ( n78831 , n78830 , n33440 );
and ( n78832 , n33592 , n45059 );
or ( n78833 , n78831 , n78832 );
and ( n78834 , n78833 , n31536 );
not ( n78835 , n33419 );
and ( n78836 , n78835 , n33440 );
and ( n78837 , n73496 , n33419 );
or ( n78838 , n78836 , n78837 );
and ( n78839 , n78838 , n31529 );
not ( n78840 , n33734 );
and ( n78841 , n78840 , n33440 );
and ( n78842 , n73509 , n33734 );
or ( n78843 , n78841 , n78842 );
and ( n78844 , n78843 , n31527 );
and ( n78845 , n33872 , n48513 );
or ( n78846 , n78804 , n78809 , n78814 , n78819 , n78824 , n78829 , n78834 , n78839 , n78844 , n78845 );
and ( n78847 , n78846 , n31557 );
and ( n78848 , n31079 , n33973 );
and ( n78849 , n33440 , n48524 );
or ( n78850 , C0 , n78847 , n78848 , n78849 );
buf ( n78851 , n78850 );
buf ( n78852 , n78851 );
buf ( n78853 , n30987 );
buf ( n78854 , n31655 );
not ( n78855 , n46356 );
and ( n78856 , n78855 , n31311 );
not ( n78857 , n55473 );
and ( n78858 , n78857 , n31311 );
and ( n78859 , n31339 , n55473 );
or ( n78860 , n78858 , n78859 );
and ( n78861 , n78860 , n46356 );
or ( n78862 , n78856 , n78861 );
and ( n78863 , n78862 , n31649 );
not ( n78864 , n55481 );
not ( n78865 , n55473 );
and ( n78866 , n78865 , n31311 );
and ( n78867 , n47449 , n55473 );
or ( n78868 , n78866 , n78867 );
and ( n78869 , n78864 , n78868 );
and ( n78870 , n47449 , n55481 );
or ( n78871 , n78869 , n78870 );
and ( n78872 , n78871 , n31643 );
not ( n78873 , n31452 );
not ( n78874 , n55481 );
not ( n78875 , n55473 );
and ( n78876 , n78875 , n31311 );
and ( n78877 , n47449 , n55473 );
or ( n78878 , n78876 , n78877 );
and ( n78879 , n78874 , n78878 );
and ( n78880 , n47449 , n55481 );
or ( n78881 , n78879 , n78880 );
and ( n78882 , n78873 , n78881 );
not ( n78883 , n55501 );
not ( n78884 , n55503 );
and ( n78885 , n78884 , n78881 );
and ( n78886 , n47485 , n55503 );
or ( n78887 , n78885 , n78886 );
and ( n78888 , n78883 , n78887 );
and ( n78889 , n47503 , n55501 );
or ( n78890 , n78888 , n78889 );
and ( n78891 , n78890 , n31452 );
or ( n78892 , n78882 , n78891 );
and ( n78893 , n78892 , n31638 );
and ( n78894 , n31311 , n47277 );
or ( n78895 , C0 , n78863 , n78872 , n78893 , n78894 );
buf ( n78896 , n78895 );
buf ( n78897 , n78896 );
and ( n78898 , n78531 , n32494 );
not ( n78899 , n46083 );
and ( n78900 , n78899 , n66893 );
not ( n78901 , n46290 );
and ( n78902 , n78901 , n46091 );
xor ( n78903 , n46306 , n46092 );
and ( n78904 , n78903 , n46290 );
or ( n78905 , n78902 , n78904 );
and ( n78906 , n78905 , n46083 );
or ( n78907 , n78900 , n78906 );
and ( n78908 , n78907 , n32421 );
not ( n78909 , n46326 );
and ( n78910 , n78909 , n66893 );
and ( n78911 , n78905 , n46326 );
or ( n78912 , n78910 , n78911 );
and ( n78913 , n78912 , n32417 );
and ( n78914 , n66893 , n46340 );
or ( n78915 , n78908 , n78913 , n78914 );
and ( n78916 , n78915 , n32456 );
and ( n78917 , n66893 , n46349 );
or ( n78918 , C0 , n78898 , n78916 , n78917 );
buf ( n78919 , n78918 );
buf ( n78920 , n78919 );
buf ( n78921 , n31655 );
buf ( n78922 , n31655 );
buf ( n78923 , n30987 );
not ( n78924 , n58883 );
and ( n78925 , n78924 , n58207 );
and ( n78926 , n54731 , n44695 );
or ( n78927 , n78925 , n78926 );
buf ( n78928 , n78927 );
buf ( n78929 , n78928 );
buf ( n78930 , n30987 );
buf ( n78931 , n31655 );
buf ( n78932 , n30987 );
not ( n78933 , n40163 );
and ( n78934 , n78933 , n31840 );
not ( n78935 , n52120 );
and ( n78936 , n78935 , n31840 );
and ( n78937 , n32235 , n52120 );
or ( n78938 , n78936 , n78937 );
and ( n78939 , n78938 , n40163 );
or ( n78940 , n78934 , n78939 );
and ( n78941 , n78940 , n32498 );
not ( n78942 , n52128 );
not ( n78943 , n52120 );
and ( n78944 , n78943 , n31840 );
and ( n78945 , n42188 , n52120 );
or ( n78946 , n78944 , n78945 );
and ( n78947 , n78942 , n78946 );
and ( n78948 , n42188 , n52128 );
or ( n78949 , n78947 , n78948 );
and ( n78950 , n78949 , n32473 );
not ( n78951 , n32475 );
not ( n78952 , n52128 );
not ( n78953 , n52120 );
and ( n78954 , n78953 , n31840 );
and ( n78955 , n42188 , n52120 );
or ( n78956 , n78954 , n78955 );
and ( n78957 , n78952 , n78956 );
and ( n78958 , n42188 , n52128 );
or ( n78959 , n78957 , n78958 );
and ( n78960 , n78951 , n78959 );
not ( n78961 , n52148 );
not ( n78962 , n52150 );
and ( n78963 , n78962 , n78959 );
and ( n78964 , n42216 , n52150 );
or ( n78965 , n78963 , n78964 );
and ( n78966 , n78961 , n78965 );
and ( n78967 , n42224 , n52148 );
or ( n78968 , n78966 , n78967 );
and ( n78969 , n78968 , n32475 );
or ( n78970 , n78960 , n78969 );
and ( n78971 , n78970 , n32486 );
and ( n78972 , n31840 , n41278 );
or ( n78973 , C0 , n78941 , n78950 , n78971 , n78972 );
buf ( n78974 , n78973 );
buf ( n78975 , n78974 );
buf ( n78976 , n31655 );
not ( n78977 , n72565 );
and ( n78978 , n78977 , n72566 );
and ( n78979 , n53761 , n67908 );
or ( n78980 , n78978 , C0 , n78979 );
buf ( n78981 , n78980 );
buf ( n78982 , n78981 );
buf ( n78983 , n30987 );
buf ( n78984 , n31655 );
buf ( n78985 , n30987 );
not ( n78986 , n32953 );
and ( n78987 , n78986 , n76740 );
and ( n78988 , n76754 , n32953 );
or ( n78989 , n78987 , n78988 );
and ( n78990 , n78989 , n33038 );
not ( n78991 , n48660 );
and ( n78992 , n78991 , n76740 );
and ( n78993 , n78609 , n48660 );
or ( n78994 , n78992 , n78993 );
and ( n78995 , n78994 , n33172 );
and ( n78996 , n76740 , n39795 );
or ( n78997 , n78990 , n78995 , n78996 );
and ( n78998 , n78997 , n33208 );
and ( n78999 , n76740 , n39805 );
or ( n79000 , C0 , n78998 , n78999 );
buf ( n79001 , n79000 );
buf ( n79002 , n79001 );
buf ( n79003 , n30987 );
buf ( n79004 , n31655 );
not ( n79005 , n68284 );
not ( n79006 , n68286 );
not ( n79007 , n68289 );
and ( n79008 , n79006 , n79007 );
buf ( n79009 , n68286 );
or ( n79010 , n79008 , n79009 );
and ( n79011 , n79005 , n79010 );
buf ( n79012 , n79011 );
and ( n79013 , n79012 , n44694 );
not ( n79014 , n68304 );
and ( n79015 , n79014 , n44692 );
not ( n79016 , n68313 );
not ( n79017 , n68316 );
and ( n79018 , n79017 , n48294 );
buf ( n79019 , n68316 );
or ( n79020 , n79018 , n79019 );
and ( n79021 , n79016 , n79020 );
buf ( n79022 , n79021 );
and ( n79023 , n79022 , n44690 );
not ( n79024 , n68289 );
not ( n79025 , n68327 );
not ( n79026 , n68331 );
not ( n79027 , n68334 );
and ( n79028 , n79026 , n79027 );
buf ( n79029 , n68331 );
or ( n79030 , n79028 , n79029 );
and ( n79031 , n79025 , n79030 );
and ( n79032 , n32956 , n68327 );
or ( n79033 , n79031 , n79032 );
and ( n79034 , n79024 , n79033 );
buf ( n79035 , n79034 );
and ( n79036 , n79035 , n44688 );
buf ( n79037 , n44682 );
not ( n79038 , n68281 );
and ( n79039 , n79038 , n44685 );
buf ( n79040 , n44686 );
or ( n79041 , n79013 , C0 , n79015 , n79023 , n79036 , n79037 , n79039 , n79040 );
buf ( n79042 , n79041 );
buf ( n79043 , n79042 );
buf ( n79044 , n30987 );
buf ( n79045 , n30987 );
buf ( n79046 , n31655 );
buf ( n79047 , n31655 );
buf ( n79048 , n31655 );
buf ( n79049 , n31655 );
buf ( n79050 , n30987 );
not ( n79051 , n34150 );
and ( n79052 , n79051 , n32747 );
not ( n79053 , n56093 );
and ( n79054 , n79053 , n32747 );
and ( n79055 , n32755 , n56093 );
or ( n79056 , n79054 , n79055 );
and ( n79057 , n79056 , n34150 );
or ( n79058 , n79052 , n79057 );
and ( n79059 , n79058 , n33381 );
not ( n79060 , n56101 );
not ( n79061 , n56093 );
and ( n79062 , n79061 , n32747 );
and ( n79063 , n35083 , n56093 );
or ( n79064 , n79062 , n79063 );
and ( n79065 , n79060 , n79064 );
and ( n79066 , n35083 , n56101 );
or ( n79067 , n79065 , n79066 );
and ( n79068 , n79067 , n33375 );
not ( n79069 , n32968 );
not ( n79070 , n56101 );
not ( n79071 , n56093 );
and ( n79072 , n79071 , n32747 );
and ( n79073 , n35083 , n56093 );
or ( n79074 , n79072 , n79073 );
and ( n79075 , n79070 , n79074 );
and ( n79076 , n35083 , n56101 );
or ( n79077 , n79075 , n79076 );
and ( n79078 , n79069 , n79077 );
not ( n79079 , n56121 );
not ( n79080 , n56123 );
and ( n79081 , n79080 , n79077 );
and ( n79082 , n35107 , n56123 );
or ( n79083 , n79081 , n79082 );
and ( n79084 , n79079 , n79083 );
and ( n79085 , n35115 , n56121 );
or ( n79086 , n79084 , n79085 );
and ( n79087 , n79086 , n32968 );
or ( n79088 , n79078 , n79087 );
and ( n79089 , n79088 , n33370 );
and ( n79090 , n32747 , n35062 );
or ( n79091 , C0 , n79059 , n79068 , n79089 , n79090 );
buf ( n79092 , n79091 );
buf ( n79093 , n79092 );
not ( n79094 , n34150 );
and ( n79095 , n79094 , n32785 );
not ( n79096 , n56140 );
and ( n79097 , n79096 , n32785 );
and ( n79098 , n32789 , n56140 );
or ( n79099 , n79097 , n79098 );
and ( n79100 , n79099 , n34150 );
or ( n79101 , n79095 , n79100 );
and ( n79102 , n79101 , n33381 );
not ( n79103 , n56148 );
not ( n79104 , n56140 );
and ( n79105 , n79104 , n32785 );
and ( n79106 , n34301 , n56140 );
or ( n79107 , n79105 , n79106 );
and ( n79108 , n79103 , n79107 );
and ( n79109 , n34301 , n56148 );
or ( n79110 , n79108 , n79109 );
and ( n79111 , n79110 , n33375 );
not ( n79112 , n32968 );
not ( n79113 , n56148 );
not ( n79114 , n56140 );
and ( n79115 , n79114 , n32785 );
and ( n79116 , n34301 , n56140 );
or ( n79117 , n79115 , n79116 );
and ( n79118 , n79113 , n79117 );
and ( n79119 , n34301 , n56148 );
or ( n79120 , n79118 , n79119 );
and ( n79121 , n79112 , n79120 );
not ( n79122 , n56168 );
not ( n79123 , n56170 );
and ( n79124 , n79123 , n79120 );
and ( n79125 , n34761 , n56170 );
or ( n79126 , n79124 , n79125 );
and ( n79127 , n79122 , n79126 );
and ( n79128 , n35050 , n56168 );
or ( n79129 , n79127 , n79128 );
and ( n79130 , n79129 , n32968 );
or ( n79131 , n79121 , n79130 );
and ( n79132 , n79131 , n33370 );
and ( n79133 , n32785 , n35062 );
or ( n79134 , C0 , n79102 , n79111 , n79132 , n79133 );
buf ( n79135 , n79134 );
buf ( n79136 , n79135 );
buf ( n79137 , n30987 );
not ( n79138 , n38443 );
and ( n79139 , n79138 , n38337 );
xor ( n79140 , n53462 , n53507 );
and ( n79141 , n79140 , n38443 );
or ( n79142 , n79139 , n79141 );
and ( n79143 , n79142 , n38450 );
not ( n79144 , n39339 );
and ( n79145 , n79144 , n39237 );
xor ( n79146 , n53518 , n53563 );
and ( n79147 , n79146 , n39339 );
or ( n79148 , n79145 , n79147 );
and ( n79149 , n79148 , n39346 );
and ( n79150 , n40222 , n39359 );
or ( n79151 , n79143 , n79149 , n79150 );
buf ( n79152 , n79151 );
buf ( n79153 , n79152 );
and ( n79154 , n42404 , n48455 );
not ( n79155 , n48457 );
and ( n79156 , n79155 , n42377 );
and ( n79157 , n42404 , n48457 );
or ( n79158 , n79156 , n79157 );
and ( n79159 , n79158 , n31373 );
not ( n79160 , n44807 );
and ( n79161 , n79160 , n42377 );
and ( n79162 , n42404 , n44807 );
or ( n79163 , n79161 , n79162 );
and ( n79164 , n79163 , n31408 );
not ( n79165 , n48468 );
and ( n79166 , n79165 , n42377 );
and ( n79167 , n42404 , n48468 );
or ( n79168 , n79166 , n79167 );
and ( n79169 , n79168 , n31468 );
not ( n79170 , n44817 );
and ( n79171 , n79170 , n42377 );
and ( n79172 , n42404 , n44817 );
or ( n79173 , n79171 , n79172 );
and ( n79174 , n79173 , n31521 );
not ( n79175 , n39979 );
and ( n79176 , n79175 , n42377 );
and ( n79177 , n42385 , n39979 );
or ( n79178 , n79176 , n79177 );
and ( n79179 , n79178 , n31538 );
not ( n79180 , n45059 );
and ( n79181 , n79180 , n42377 );
and ( n79182 , n42385 , n45059 );
or ( n79183 , n79181 , n79182 );
and ( n79184 , n79183 , n31536 );
not ( n79185 , n33419 );
and ( n79186 , n79185 , n42377 );
and ( n79187 , n62990 , n33419 );
or ( n79188 , n79186 , n79187 );
and ( n79189 , n79188 , n31529 );
not ( n79190 , n33734 );
and ( n79191 , n79190 , n42377 );
and ( n79192 , n63001 , n33734 );
or ( n79193 , n79191 , n79192 );
and ( n79194 , n79193 , n31527 );
and ( n79195 , n42418 , n48513 );
or ( n79196 , n79154 , n79159 , n79164 , n79169 , n79174 , n79179 , n79184 , n79189 , n79194 , n79195 );
and ( n79197 , n79196 , n31557 );
and ( n79198 , n35393 , n33973 );
and ( n79199 , n42377 , n48524 );
or ( n79200 , C0 , n79197 , n79198 , n79199 );
buf ( n79201 , n79200 );
buf ( n79202 , n79201 );
buf ( n79203 , n30987 );
buf ( n79204 , n31655 );
buf ( n79205 , RI15b5eb90_1097);
and ( n79206 , n79205 , n32494 );
not ( n79207 , n46083 );
buf ( n79208 , RI15b60198_1144);
and ( n79209 , n79207 , n79208 );
buf ( n79210 , n79209 );
and ( n79211 , n79210 , n32421 );
not ( n79212 , n46326 );
and ( n79213 , n79212 , n79208 );
not ( n79214 , n51396 );
and ( n79215 , n79214 , n51239 );
xor ( n79216 , n51400 , n51410 );
and ( n79217 , n79216 , n51396 );
or ( n79218 , n79215 , n79217 );
and ( n79219 , n79218 , n46326 );
or ( n79220 , n79213 , n79219 );
and ( n79221 , n79220 , n32417 );
and ( n79222 , n79208 , n46340 );
or ( n79223 , n79211 , n79221 , n79222 );
and ( n79224 , n79223 , n32456 );
and ( n79225 , n79208 , n46349 );
or ( n79226 , C0 , n79206 , n79224 , n79225 );
buf ( n79227 , n79226 );
buf ( n79228 , n79227 );
buf ( n79229 , n31655 );
not ( n79230 , n46356 );
and ( n79231 , n79230 , n31148 );
not ( n79232 , n78324 );
and ( n79233 , n79232 , n31148 );
and ( n79234 , n31172 , n78324 );
or ( n79235 , n79233 , n79234 );
and ( n79236 , n79235 , n46356 );
or ( n79237 , n79231 , n79236 );
and ( n79238 , n79237 , n31649 );
not ( n79239 , n78332 );
not ( n79240 , n78324 );
and ( n79241 , n79240 , n31148 );
and ( n79242 , n46495 , n78324 );
or ( n79243 , n79241 , n79242 );
and ( n79244 , n79239 , n79243 );
and ( n79245 , n46495 , n78332 );
or ( n79246 , n79244 , n79245 );
and ( n79247 , n79246 , n31643 );
not ( n79248 , n31452 );
not ( n79249 , n78332 );
not ( n79250 , n78324 );
and ( n79251 , n79250 , n31148 );
and ( n79252 , n46495 , n78324 );
or ( n79253 , n79251 , n79252 );
and ( n79254 , n79249 , n79253 );
and ( n79255 , n46495 , n78332 );
or ( n79256 , n79254 , n79255 );
and ( n79257 , n79248 , n79256 );
not ( n79258 , n78352 );
not ( n79259 , n78354 );
and ( n79260 , n79259 , n79256 );
and ( n79261 , n46984 , n78354 );
or ( n79262 , n79260 , n79261 );
and ( n79263 , n79258 , n79262 );
and ( n79264 , n47267 , n78352 );
or ( n79265 , n79263 , n79264 );
and ( n79266 , n79265 , n31452 );
or ( n79267 , n79257 , n79266 );
and ( n79268 , n79267 , n31638 );
and ( n79269 , n31148 , n47277 );
or ( n79270 , C0 , n79238 , n79247 , n79268 , n79269 );
buf ( n79271 , n79270 );
buf ( n79272 , n79271 );
buf ( n79273 , n30987 );
buf ( n79274 , n31655 );
buf ( n79275 , n67631 );
nor ( n79276 , n67617 , n67626 , n67630 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
buf ( n79277 , n79276 );
buf ( n79278 , n67704 );
or ( n79279 , n79275 , n79277 , n79278 , C0 );
and ( n79280 , n79279 , n67665 );
buf ( n79281 , n67631 );
buf ( n79282 , n79276 );
buf ( n79283 , n67704 );
or ( n79284 , C0 , n79281 , n79282 , n79283 , C0 );
and ( n79285 , n79284 , n67701 );
buf ( n79286 , n67631 );
buf ( n79287 , n79276 );
buf ( n79288 , n67704 );
or ( n79289 , C0 , n79286 , n79287 , n79288 , C0 );
and ( n79290 , n79289 , n67737 );
or ( n79291 , C0 , n79280 , n79285 , n79290 );
buf ( n79292 , n79291 );
buf ( n79293 , n79292 );
not ( n79294 , n46356 );
and ( n79295 , n79294 , n31152 );
not ( n79296 , n52734 );
and ( n79297 , n79296 , n31152 );
and ( n79298 , n31172 , n52734 );
or ( n79299 , n79297 , n79298 );
and ( n79300 , n79299 , n46356 );
or ( n79301 , n79295 , n79300 );
and ( n79302 , n79301 , n31649 );
not ( n79303 , n52742 );
not ( n79304 , n52734 );
and ( n79305 , n79304 , n31152 );
and ( n79306 , n46495 , n52734 );
or ( n79307 , n79305 , n79306 );
and ( n79308 , n79303 , n79307 );
and ( n79309 , n46495 , n52742 );
or ( n79310 , n79308 , n79309 );
and ( n79311 , n79310 , n31643 );
not ( n79312 , n31452 );
not ( n79313 , n52742 );
not ( n79314 , n52734 );
and ( n79315 , n79314 , n31152 );
and ( n79316 , n46495 , n52734 );
or ( n79317 , n79315 , n79316 );
and ( n79318 , n79313 , n79317 );
and ( n79319 , n46495 , n52742 );
or ( n79320 , n79318 , n79319 );
and ( n79321 , n79312 , n79320 );
not ( n79322 , n52762 );
not ( n79323 , n52764 );
and ( n79324 , n79323 , n79320 );
and ( n79325 , n46984 , n52764 );
or ( n79326 , n79324 , n79325 );
and ( n79327 , n79322 , n79326 );
and ( n79328 , n47267 , n52762 );
or ( n79329 , n79327 , n79328 );
and ( n79330 , n79329 , n31452 );
or ( n79331 , n79321 , n79330 );
and ( n79332 , n79331 , n31638 );
and ( n79333 , n31152 , n47277 );
or ( n79334 , C0 , n79302 , n79311 , n79332 , n79333 );
buf ( n79335 , n79334 );
buf ( n79336 , n79335 );
buf ( n79337 , n30987 );
buf ( n79338 , n31655 );
buf ( n79339 , n31655 );
not ( n79340 , n41532 );
and ( n79341 , n79340 , n34373 );
and ( n79342 , n60249 , n41532 );
or ( n79343 , n79341 , n79342 );
buf ( n79344 , n79343 );
buf ( n79345 , n79344 );
buf ( n79346 , n31655 );
buf ( n79347 , n30987 );
xor ( n79348 , n54138 , n78384 );
and ( n79349 , n79348 , n33199 );
not ( n79350 , n48648 );
and ( n79351 , n79350 , n54138 );
and ( n79352 , n34423 , n48648 );
or ( n79353 , n79351 , n79352 );
and ( n79354 , n79353 , n32924 );
not ( n79355 , n48660 );
and ( n79356 , n79355 , n54138 );
and ( n79357 , n70680 , n48660 );
or ( n79358 , n79356 , n79357 );
and ( n79359 , n79358 , n33172 );
not ( n79360 , n48730 );
and ( n79361 , n79360 , n54138 );
xor ( n79362 , n58506 , n78403 );
and ( n79363 , n79362 , n48730 );
or ( n79364 , n79361 , n79363 );
and ( n79365 , n79364 , n33187 );
and ( n79366 , n54138 , n54713 );
or ( n79367 , n79349 , n79354 , n79359 , n79365 , n79366 );
and ( n79368 , n79367 , n33208 );
and ( n79369 , n54138 , n39805 );
or ( n79370 , C0 , n79368 , n79369 );
buf ( n79371 , n79370 );
buf ( n79372 , n79371 );
buf ( n79373 , n30987 );
buf ( n79374 , n31655 );
buf ( n79375 , n30987 );
buf ( n79376 , n31655 );
buf ( n79377 , n31655 );
buf ( n79378 , n30987 );
and ( n79379 , n49078 , n48639 );
not ( n79380 , n48642 );
and ( n79381 , n79380 , n48603 );
and ( n79382 , n49078 , n48642 );
or ( n79383 , n79381 , n79382 );
and ( n79384 , n79383 , n32890 );
not ( n79385 , n48648 );
and ( n79386 , n79385 , n48603 );
and ( n79387 , n49078 , n48648 );
or ( n79388 , n79386 , n79387 );
and ( n79389 , n79388 , n32924 );
not ( n79390 , n48654 );
and ( n79391 , n79390 , n48603 );
and ( n79392 , n49078 , n48654 );
or ( n79393 , n79391 , n79392 );
and ( n79394 , n79393 , n33038 );
not ( n79395 , n48660 );
and ( n79396 , n79395 , n48603 );
and ( n79397 , n49078 , n48660 );
or ( n79398 , n79396 , n79397 );
and ( n79399 , n79398 , n33172 );
not ( n79400 , n41576 );
and ( n79401 , n79400 , n48603 );
and ( n79402 , n48788 , n41576 );
or ( n79403 , n79401 , n79402 );
and ( n79404 , n79403 , n33189 );
not ( n79405 , n48730 );
and ( n79406 , n79405 , n48603 );
and ( n79407 , n48788 , n48730 );
or ( n79408 , n79406 , n79407 );
and ( n79409 , n79408 , n33187 );
not ( n79410 , n48765 );
and ( n79411 , n79410 , n48603 );
and ( n79412 , n49745 , n48765 );
or ( n79413 , n79411 , n79412 );
and ( n79414 , n79413 , n33180 );
not ( n79415 , n49054 );
and ( n79416 , n79415 , n48603 );
and ( n79417 , n49756 , n49054 );
or ( n79418 , n79416 , n79417 );
and ( n79419 , n79418 , n33178 );
and ( n79420 , n49187 , n49275 );
or ( n79421 , n79379 , n79384 , n79389 , n79394 , n79399 , n79404 , n79409 , n79414 , n79419 , n79420 );
and ( n79422 , n79421 , n33208 );
and ( n79423 , n32996 , n35056 );
and ( n79424 , n48603 , n49286 );
or ( n79425 , C0 , n79422 , n79423 , n79424 );
buf ( n79426 , n79425 );
buf ( n79427 , n79426 );
buf ( n79428 , n54728 );
buf ( n79429 , n31655 );
and ( n79430 , n33238 , n32528 );
not ( n79431 , n32598 );
and ( n79432 , n79431 , n33001 );
and ( n79433 , n48807 , n32598 );
or ( n79434 , n79432 , n79433 );
and ( n79435 , n79434 , n32890 );
not ( n79436 , n32919 );
and ( n79437 , n79436 , n33001 );
and ( n79438 , n48807 , n32919 );
or ( n79439 , n79437 , n79438 );
and ( n79440 , n79439 , n32924 );
not ( n79441 , n32953 );
and ( n79442 , n79441 , n33001 );
not ( n79443 , n32971 );
and ( n79444 , n79443 , n33127 );
xor ( n79445 , n33001 , n33004 );
and ( n79446 , n79445 , n32971 );
or ( n79447 , n79444 , n79446 );
and ( n79448 , n79447 , n32953 );
or ( n79449 , n79442 , n79448 );
and ( n79450 , n79449 , n33038 );
not ( n79451 , n33067 );
and ( n79452 , n79451 , n33001 );
not ( n79453 , n32970 );
not ( n79454 , n33071 );
and ( n79455 , n79454 , n33127 );
xor ( n79456 , n33128 , n33136 );
and ( n79457 , n79456 , n33071 );
or ( n79458 , n79455 , n79457 );
and ( n79459 , n79453 , n79458 );
and ( n79460 , n79445 , n32970 );
or ( n79461 , n79459 , n79460 );
and ( n79462 , n79461 , n33067 );
or ( n79463 , n79452 , n79462 );
and ( n79464 , n79463 , n33172 );
and ( n79465 , n33001 , n33204 );
or ( n79466 , n79435 , n79440 , n79450 , n79464 , n79465 );
and ( n79467 , n79466 , n33208 );
not ( n79468 , n32968 );
not ( n79469 , n33270 );
and ( n79470 , n79469 , n33327 );
xor ( n79471 , n33328 , n33336 );
and ( n79472 , n79471 , n33270 );
or ( n79473 , n79470 , n79472 );
and ( n79474 , n79468 , n79473 );
and ( n79475 , n33001 , n32968 );
or ( n79476 , n79474 , n79475 );
and ( n79477 , n79476 , n33370 );
and ( n79478 , n33001 , n33382 );
or ( n79479 , C0 , n79430 , n79467 , n79477 , C0 , n79478 );
buf ( n79480 , n79479 );
buf ( n79481 , n79480 );
buf ( n79482 , n30987 );
buf ( n79483 , n30987 );
and ( n79484 , n32462 , n32500 );
not ( n79485 , n35211 );
and ( n79486 , n79485 , n37583 );
and ( n79487 , n31770 , n35211 );
or ( n79488 , n79486 , n79487 );
and ( n79489 , n79488 , n32421 );
not ( n79490 , n35245 );
and ( n79491 , n79490 , n37583 );
and ( n79492 , n31770 , n35245 );
or ( n79493 , n79491 , n79492 );
and ( n79494 , n79493 , n32419 );
not ( n79495 , n35278 );
and ( n79496 , n79495 , n37583 );
not ( n79497 , n35295 );
and ( n79498 , n79497 , n47290 );
xor ( n79499 , n37583 , n49523 );
and ( n79500 , n79499 , n35295 );
or ( n79501 , n79498 , n79500 );
and ( n79502 , n79501 , n35278 );
or ( n79503 , n79496 , n79502 );
and ( n79504 , n79503 , n32417 );
not ( n79505 , n35331 );
and ( n79506 , n79505 , n37583 );
not ( n79507 , n35294 );
not ( n79508 , n45995 );
and ( n79509 , n79508 , n47290 );
xor ( n79510 , n49608 , n49609 );
and ( n79511 , n79510 , n45995 );
or ( n79512 , n79509 , n79511 );
and ( n79513 , n79507 , n79512 );
and ( n79514 , n79499 , n35294 );
or ( n79515 , n79513 , n79514 );
and ( n79516 , n79515 , n35331 );
or ( n79517 , n79506 , n79516 );
and ( n79518 , n79517 , n32415 );
and ( n79519 , n37583 , n35354 );
or ( n79520 , n79489 , n79494 , n79504 , n79518 , n79519 );
and ( n79521 , n79520 , n32456 );
not ( n79522 , n32475 );
not ( n79523 , n46060 );
and ( n79524 , n79523 , n49701 );
xor ( n79525 , n49702 , n49703 );
and ( n79526 , n79525 , n46060 );
or ( n79527 , n79524 , n79526 );
and ( n79528 , n79522 , n79527 );
and ( n79529 , n37583 , n32475 );
or ( n79530 , n79528 , n79529 );
and ( n79531 , n79530 , n32486 );
and ( n79532 , n37583 , n35367 );
or ( n79533 , C0 , n79484 , n79521 , n79531 , C0 , n79532 );
buf ( n79534 , n79533 );
buf ( n79535 , n79534 );
buf ( n79536 , n31655 );
buf ( n79537 , n30987 );
buf ( n79538 , n31655 );
and ( n79539 , n66940 , n33377 );
not ( n79540 , n48545 );
and ( n79541 , n79540 , n76549 );
buf ( n79542 , n79541 );
and ( n79543 , n79542 , n32890 );
not ( n79544 , n48557 );
and ( n79545 , n79544 , n76549 );
and ( n79546 , n66946 , n48557 );
or ( n79547 , n79545 , n79546 );
and ( n79548 , n79547 , n33038 );
and ( n79549 , n76549 , n48571 );
or ( n79550 , n79543 , n79548 , n79549 );
and ( n79551 , n79550 , n33208 );
and ( n79552 , n76549 , n48577 );
or ( n79553 , C0 , n79539 , n79551 , n79552 );
buf ( n79554 , n79553 );
buf ( n79555 , n79554 );
buf ( n79556 , n31655 );
buf ( n79557 , n30987 );
buf ( n79558 , n30987 );
buf ( n79559 , n66430 );
buf ( n79560 , n42810 );
or ( n79561 , C0 , C0 , C0 , n79559 , n79560 );
and ( n79562 , n79561 , n42806 );
buf ( n79563 , n42736 );
buf ( n79564 , n66430 );
buf ( n79565 , n42810 );
or ( n79566 , C0 , C0 , n79563 , n79564 , n79565 );
and ( n79567 , n79566 , n42842 );
or ( n79568 , C0 , C0 , n79562 , n79567 );
buf ( n79569 , n79568 );
buf ( n79570 , n79569 );
buf ( n79571 , n30987 );
buf ( n79572 , n31655 );
buf ( n79573 , n31655 );
buf ( n79574 , n31655 );
buf ( n79575 , n30987 );
buf ( n79576 , n30987 );
buf ( n79577 , n31655 );
buf ( n79578 , RI15b481b0_325);
and ( n79579 , n79578 , n58207 );
and ( n79580 , n54737 , n44695 );
or ( n79581 , n79579 , n79580 );
buf ( n79582 , n79581 );
buf ( n79583 , n79582 );
buf ( n79584 , n31655 );
buf ( n79585 , n40224 );
not ( n79586 , n34150 );
and ( n79587 , n79586 , n32807 );
not ( n79588 , n57038 );
and ( n79589 , n79588 , n32807 );
and ( n79590 , n32823 , n57038 );
or ( n79591 , n79589 , n79590 );
and ( n79592 , n79591 , n34150 );
or ( n79593 , n79587 , n79592 );
and ( n79594 , n79593 , n33381 );
not ( n79595 , n57046 );
not ( n79596 , n57038 );
and ( n79597 , n79596 , n32807 );
and ( n79598 , n41464 , n57038 );
or ( n79599 , n79597 , n79598 );
and ( n79600 , n79595 , n79599 );
and ( n79601 , n41464 , n57046 );
or ( n79602 , n79600 , n79601 );
and ( n79603 , n79602 , n33375 );
not ( n79604 , n32968 );
not ( n79605 , n57046 );
not ( n79606 , n57038 );
and ( n79607 , n79606 , n32807 );
and ( n79608 , n41464 , n57038 );
or ( n79609 , n79607 , n79608 );
and ( n79610 , n79605 , n79609 );
and ( n79611 , n41464 , n57046 );
or ( n79612 , n79610 , n79611 );
and ( n79613 , n79604 , n79612 );
not ( n79614 , n57066 );
not ( n79615 , n57068 );
and ( n79616 , n79615 , n79612 );
and ( n79617 , n41490 , n57068 );
or ( n79618 , n79616 , n79617 );
and ( n79619 , n79614 , n79618 );
and ( n79620 , n41500 , n57066 );
or ( n79621 , n79619 , n79620 );
and ( n79622 , n79621 , n32968 );
or ( n79623 , n79613 , n79622 );
and ( n79624 , n79623 , n33370 );
and ( n79625 , n32807 , n35062 );
or ( n79626 , C0 , n79594 , n79603 , n79624 , n79625 );
buf ( n79627 , n79626 );
buf ( n79628 , n79627 );
buf ( n79629 , n31655 );
buf ( n79630 , n30987 );
buf ( n79631 , n30987 );
buf ( n79632 , n31655 );
buf ( n79633 , RI15b545a0_743);
and ( n79634 , n79633 , n58921 );
and ( n79635 , n41530 , n37506 );
or ( n79636 , n79634 , n79635 );
buf ( n79637 , n79636 );
buf ( n79638 , n79637 );
not ( n79639 , n38443 );
and ( n79640 , n79639 , n37980 );
xor ( n79641 , n53483 , n53486 );
and ( n79642 , n79641 , n38443 );
or ( n79643 , n79640 , n79642 );
and ( n79644 , n79643 , n38450 );
not ( n79645 , n39339 );
and ( n79646 , n79645 , n38880 );
xor ( n79647 , n53539 , n53542 );
and ( n79648 , n79647 , n39339 );
or ( n79649 , n79646 , n79648 );
and ( n79650 , n79649 , n39346 );
and ( n79651 , n40201 , n39359 );
or ( n79652 , n79644 , n79650 , n79651 );
buf ( n79653 , n79652 );
buf ( n79654 , n79653 );
buf ( n79655 , n30987 );
not ( n79656 , n35542 );
and ( n79657 , n79656 , n41844 );
buf ( n79658 , RI15b452d0_225);
and ( n79659 , n79658 , n35542 );
or ( n79660 , n79657 , n79659 );
buf ( n79661 , n79660 );
buf ( n79662 , n79661 );
buf ( n79663 , n31655 );
buf ( n79664 , n30987 );
not ( n79665 , n33419 );
and ( n79666 , n79665 , n31585 );
and ( n79667 , n59315 , n33419 );
or ( n79668 , n79666 , n79667 );
and ( n79669 , n79668 , n31529 );
not ( n79670 , n33734 );
and ( n79671 , n79670 , n31585 );
and ( n79672 , n59328 , n33734 );
or ( n79673 , n79671 , n79672 );
and ( n79674 , n79673 , n31527 );
and ( n79675 , n31585 , n33942 );
or ( n79676 , n79669 , n79674 , n79675 );
and ( n79677 , n79676 , n31557 );
and ( n79678 , n34115 , n31643 );
not ( n79679 , n31452 );
and ( n79680 , n79679 , n34115 );
xor ( n79681 , n31585 , n33952 );
and ( n79682 , n79681 , n31452 );
or ( n79683 , n79680 , n79682 );
and ( n79684 , n79683 , n31638 );
and ( n79685 , n34009 , n33973 );
and ( n79686 , n31585 , n33978 );
or ( n79687 , C0 , n79677 , n79678 , n79684 , n79685 , n79686 );
buf ( n79688 , n79687 );
buf ( n79689 , n79688 );
and ( n79690 , n76227 , n32456 );
and ( n79691 , n55558 , n47409 );
or ( n79692 , C0 , n79690 , n79691 );
buf ( n79693 , n79692 );
buf ( n79694 , n79693 );
buf ( n79695 , n30987 );
not ( n79696 , n46356 );
and ( n79697 , n79696 , n31254 );
not ( n79698 , n48214 );
and ( n79699 , n79698 , n31254 );
and ( n79700 , n31272 , n48214 );
or ( n79701 , n79699 , n79700 );
and ( n79702 , n79701 , n46356 );
or ( n79703 , n79697 , n79702 );
and ( n79704 , n79703 , n31649 );
not ( n79705 , n48223 );
not ( n79706 , n48214 );
and ( n79707 , n79706 , n31254 );
and ( n79708 , n49443 , n48214 );
or ( n79709 , n79707 , n79708 );
and ( n79710 , n79705 , n79709 );
and ( n79711 , n49443 , n48223 );
or ( n79712 , n79710 , n79711 );
and ( n79713 , n79712 , n31643 );
not ( n79714 , n31452 );
not ( n79715 , n48223 );
not ( n79716 , n48214 );
and ( n79717 , n79716 , n31254 );
and ( n79718 , n49443 , n48214 );
or ( n79719 , n79717 , n79718 );
and ( n79720 , n79715 , n79719 );
and ( n79721 , n49443 , n48223 );
or ( n79722 , n79720 , n79721 );
and ( n79723 , n79714 , n79722 );
not ( n79724 , n48244 );
not ( n79725 , n48247 );
and ( n79726 , n79725 , n79722 );
and ( n79727 , n49469 , n48247 );
or ( n79728 , n79726 , n79727 );
and ( n79729 , n79724 , n79728 );
and ( n79730 , n49477 , n48244 );
or ( n79731 , n79729 , n79730 );
and ( n79732 , n79731 , n31452 );
or ( n79733 , n79723 , n79732 );
and ( n79734 , n79733 , n31638 );
and ( n79735 , n31254 , n47277 );
or ( n79736 , C0 , n79704 , n79713 , n79734 , n79735 );
buf ( n79737 , n79736 );
buf ( n79738 , n79737 );
buf ( n79739 , n31655 );
buf ( n79740 , n30987 );
buf ( n79741 , n31655 );
and ( n79742 , n67635 , n52726 );
buf ( n79743 , n79742 );
buf ( n79744 , n79743 );
buf ( n79745 , n30987 );
buf ( n79746 , n31655 );
buf ( n79747 , n31655 );
buf ( n79748 , n30987 );
not ( n79749 , n46356 );
and ( n79750 , n79749 , n31234 );
not ( n79751 , n61975 );
and ( n79752 , n79751 , n31234 );
and ( n79753 , n31238 , n61975 );
or ( n79754 , n79752 , n79753 );
and ( n79755 , n79754 , n46356 );
or ( n79756 , n79750 , n79755 );
and ( n79757 , n79756 , n31649 );
not ( n79758 , n61983 );
not ( n79759 , n61975 );
and ( n79760 , n79759 , n31234 );
and ( n79761 , n49901 , n61975 );
or ( n79762 , n79760 , n79761 );
and ( n79763 , n79758 , n79762 );
and ( n79764 , n49901 , n61983 );
or ( n79765 , n79763 , n79764 );
and ( n79766 , n79765 , n31643 );
not ( n79767 , n31452 );
not ( n79768 , n61983 );
not ( n79769 , n61975 );
and ( n79770 , n79769 , n31234 );
and ( n79771 , n49901 , n61975 );
or ( n79772 , n79770 , n79771 );
and ( n79773 , n79768 , n79772 );
and ( n79774 , n49901 , n61983 );
or ( n79775 , n79773 , n79774 );
and ( n79776 , n79767 , n79775 );
not ( n79777 , n62003 );
not ( n79778 , n62005 );
and ( n79779 , n79778 , n79775 );
and ( n79780 , n49925 , n62005 );
or ( n79781 , n79779 , n79780 );
and ( n79782 , n79777 , n79781 );
and ( n79783 , n49933 , n62003 );
or ( n79784 , n79782 , n79783 );
and ( n79785 , n79784 , n31452 );
or ( n79786 , n79776 , n79785 );
and ( n79787 , n79786 , n31638 );
and ( n79788 , n31234 , n47277 );
or ( n79789 , C0 , n79757 , n79766 , n79787 , n79788 );
buf ( n79790 , n79789 );
buf ( n79791 , n79790 );
xor ( n79792 , n49579 , n60316 );
and ( n79793 , n79792 , n32433 );
not ( n79794 , n47331 );
and ( n79795 , n79794 , n49579 );
and ( n79796 , n66696 , n47331 );
or ( n79797 , n79795 , n79796 );
and ( n79798 , n79797 , n32413 );
and ( n79799 , n49579 , n47402 );
or ( n79800 , n79793 , n79798 , n79799 );
and ( n79801 , n79800 , n32456 );
and ( n79802 , n49579 , n47409 );
or ( n79803 , C0 , n79801 , n79802 );
buf ( n79804 , n79803 );
buf ( n79805 , n79804 );
buf ( n79806 , n31655 );
buf ( n79807 , n30987 );
and ( n79808 , n54134 , n78593 );
xor ( n79809 , n54132 , n79808 );
and ( n79810 , n79809 , n33199 );
not ( n79811 , n48648 );
and ( n79812 , n79811 , n54132 );
and ( n79813 , n34417 , n48648 );
or ( n79814 , n79812 , n79813 );
and ( n79815 , n79814 , n32924 );
not ( n79816 , n48660 );
and ( n79817 , n79816 , n54132 );
not ( n79818 , n55168 );
and ( n79819 , n79818 , n55164 );
xor ( n79820 , n55164 , n34193 );
and ( n79821 , n78605 , n78606 );
xor ( n79822 , n79820 , n79821 );
and ( n79823 , n79822 , n55168 );
or ( n79824 , n79819 , n79823 );
and ( n79825 , n79824 , n48660 );
or ( n79826 , n79817 , n79825 );
and ( n79827 , n79826 , n33172 );
not ( n79828 , n48730 );
and ( n79829 , n79828 , n54132 );
and ( n79830 , n58472 , n78615 );
xor ( n79831 , n58455 , n79830 );
and ( n79832 , n79831 , n48730 );
or ( n79833 , n79829 , n79832 );
and ( n79834 , n79833 , n33187 );
and ( n79835 , n54132 , n54713 );
or ( n79836 , n79810 , n79815 , n79827 , n79834 , n79835 );
and ( n79837 , n79836 , n33208 );
and ( n79838 , n54132 , n39805 );
or ( n79839 , C0 , n79837 , n79838 );
buf ( n79840 , n79839 );
buf ( n79841 , n79840 );
buf ( n79842 , n30987 );
buf ( n79843 , n31655 );
not ( n79844 , n41532 );
and ( n79845 , n79844 , n34379 );
and ( n79846 , n58614 , n41532 );
or ( n79847 , n79845 , n79846 );
buf ( n79848 , n79847 );
buf ( n79849 , n79848 );
and ( n79850 , n69611 , n31645 );
not ( n79851 , n45274 );
and ( n79852 , n79851 , n52207 );
buf ( n79853 , n79852 );
and ( n79854 , n79853 , n31373 );
not ( n79855 , n45280 );
and ( n79856 , n79855 , n52207 );
and ( n79857 , n69617 , n45280 );
or ( n79858 , n79856 , n79857 );
and ( n79859 , n79858 , n31468 );
and ( n79860 , n52207 , n45802 );
or ( n79861 , n79854 , n79859 , n79860 );
and ( n79862 , n79861 , n31557 );
and ( n79863 , n52207 , n45808 );
or ( n79864 , C0 , n79850 , n79862 , n79863 );
buf ( n79865 , n79864 );
buf ( n79866 , n79865 );
buf ( n79867 , n31655 );
buf ( n79868 , n30987 );
buf ( n79869 , n30987 );
not ( n79870 , n40163 );
and ( n79871 , n79870 , n31906 );
not ( n79872 , n45227 );
and ( n79873 , n79872 , n31906 );
and ( n79874 , n32200 , n45227 );
or ( n79875 , n79873 , n79874 );
and ( n79876 , n79875 , n40163 );
or ( n79877 , n79871 , n79876 );
and ( n79878 , n79877 , n32498 );
not ( n79879 , n45235 );
not ( n79880 , n45227 );
and ( n79881 , n79880 , n31906 );
and ( n79882 , n53243 , n45227 );
or ( n79883 , n79881 , n79882 );
and ( n79884 , n79879 , n79883 );
and ( n79885 , n53243 , n45235 );
or ( n79886 , n79884 , n79885 );
and ( n79887 , n79886 , n32473 );
not ( n79888 , n32475 );
not ( n79889 , n45235 );
not ( n79890 , n45227 );
and ( n79891 , n79890 , n31906 );
and ( n79892 , n53243 , n45227 );
or ( n79893 , n79891 , n79892 );
and ( n79894 , n79889 , n79893 );
and ( n79895 , n53243 , n45235 );
or ( n79896 , n79894 , n79895 );
and ( n79897 , n79888 , n79896 );
not ( n79898 , n45255 );
not ( n79899 , n45257 );
and ( n79900 , n79899 , n79896 );
and ( n79901 , n53269 , n45257 );
or ( n79902 , n79900 , n79901 );
and ( n79903 , n79898 , n79902 );
and ( n79904 , n53277 , n45255 );
or ( n79905 , n79903 , n79904 );
and ( n79906 , n79905 , n32475 );
or ( n79907 , n79897 , n79906 );
and ( n79908 , n79907 , n32486 );
and ( n79909 , n31906 , n41278 );
or ( n79910 , C0 , n79878 , n79887 , n79908 , n79909 );
buf ( n79911 , n79910 );
buf ( n79912 , n79911 );
and ( n79913 , n47669 , n50275 );
not ( n79914 , n50278 );
and ( n79915 , n79914 , n47582 );
and ( n79916 , n47669 , n50278 );
or ( n79917 , n79915 , n79916 );
and ( n79918 , n79917 , n32421 );
not ( n79919 , n50002 );
and ( n79920 , n79919 , n47582 );
and ( n79921 , n47669 , n50002 );
or ( n79922 , n79920 , n79921 );
and ( n79923 , n79922 , n32419 );
not ( n79924 , n50289 );
and ( n79925 , n79924 , n47582 );
and ( n79926 , n47669 , n50289 );
or ( n79927 , n79925 , n79926 );
and ( n79928 , n79927 , n32417 );
not ( n79929 , n50008 );
and ( n79930 , n79929 , n47582 );
and ( n79931 , n47669 , n50008 );
or ( n79932 , n79930 , n79931 );
and ( n79933 , n79932 , n32415 );
not ( n79934 , n47331 );
and ( n79935 , n79934 , n47582 );
and ( n79936 , n47614 , n47331 );
or ( n79937 , n79935 , n79936 );
and ( n79938 , n79937 , n32413 );
not ( n79939 , n50067 );
and ( n79940 , n79939 , n47582 );
and ( n79941 , n47614 , n50067 );
or ( n79942 , n79940 , n79941 );
and ( n79943 , n79942 , n32411 );
not ( n79944 , n31728 );
and ( n79945 , n79944 , n47582 );
and ( n79946 , n49801 , n31728 );
or ( n79947 , n79945 , n79946 );
and ( n79948 , n79947 , n32253 );
not ( n79949 , n32283 );
and ( n79950 , n79949 , n47582 );
and ( n79951 , n49812 , n32283 );
or ( n79952 , n79950 , n79951 );
and ( n79953 , n79952 , n32398 );
and ( n79954 , n47719 , n50334 );
or ( n79955 , n79913 , n79918 , n79923 , n79928 , n79933 , n79938 , n79943 , n79948 , n79953 , n79954 );
and ( n79956 , n79955 , n32456 );
and ( n79957 , n37571 , n32489 );
and ( n79958 , n47582 , n50345 );
or ( n79959 , C0 , n79956 , n79957 , n79958 );
buf ( n79960 , n79959 );
buf ( n79961 , n79960 );
buf ( n79962 , n30987 );
buf ( n79963 , n31655 );
not ( n79964 , n31437 );
and ( n79965 , n79964 , n54603 );
and ( n79966 , n54616 , n31437 );
or ( n79967 , n79965 , n79966 );
and ( n79968 , n79967 , n31468 );
not ( n79969 , n44817 );
and ( n79970 , n79969 , n54603 );
and ( n79971 , n68989 , n44817 );
or ( n79972 , n79970 , n79971 );
and ( n79973 , n79972 , n31521 );
and ( n79974 , n54603 , n42158 );
or ( n79975 , n79968 , n79973 , n79974 );
and ( n79976 , n79975 , n31557 );
and ( n79977 , n54603 , n40154 );
or ( n79978 , C0 , n79976 , n79977 );
buf ( n79979 , n79978 );
buf ( n79980 , n79979 );
buf ( n79981 , n31655 );
buf ( n79982 , n30987 );
buf ( n79983 , n30987 );
buf ( n79984 , n31655 );
not ( n79985 , n32953 );
buf ( n79986 , RI15b46d88_282);
and ( n79987 , n79985 , n79986 );
not ( n79988 , n39572 );
and ( n79989 , n79988 , n39542 );
xor ( n79990 , n42615 , n42638 );
and ( n79991 , n79990 , n39572 );
or ( n79992 , n79989 , n79991 );
and ( n79993 , n79992 , n32953 );
or ( n79994 , n79987 , n79993 );
and ( n79995 , n79994 , n33038 );
not ( n79996 , n39586 );
and ( n79997 , n79996 , n79986 );
not ( n79998 , n39775 );
and ( n79999 , n79998 , n39747 );
xor ( n80000 , n42651 , n42674 );
and ( n80001 , n80000 , n39775 );
or ( n80002 , n79999 , n80001 );
and ( n80003 , n80002 , n39586 );
or ( n80004 , n79997 , n80003 );
and ( n80005 , n80004 , n33172 );
and ( n80006 , n79986 , n39795 );
or ( n80007 , n79995 , n80005 , n80006 );
and ( n80008 , n80007 , n33208 );
and ( n80009 , n79986 , n39805 );
or ( n80010 , C0 , n80008 , n80009 );
buf ( n80011 , n80010 );
buf ( n80012 , n80011 );
buf ( n80013 , n31655 );
not ( n80014 , n34150 );
and ( n80015 , n80014 , n32769 );
not ( n80016 , n57872 );
and ( n80017 , n80016 , n32769 );
and ( n80018 , n32789 , n57872 );
or ( n80019 , n80017 , n80018 );
and ( n80020 , n80019 , n34150 );
or ( n80021 , n80015 , n80020 );
and ( n80022 , n80021 , n33381 );
not ( n80023 , n57880 );
not ( n80024 , n57872 );
and ( n80025 , n80024 , n32769 );
and ( n80026 , n34301 , n57872 );
or ( n80027 , n80025 , n80026 );
and ( n80028 , n80023 , n80027 );
and ( n80029 , n34301 , n57880 );
or ( n80030 , n80028 , n80029 );
and ( n80031 , n80030 , n33375 );
not ( n80032 , n32968 );
not ( n80033 , n57880 );
not ( n80034 , n57872 );
and ( n80035 , n80034 , n32769 );
and ( n80036 , n34301 , n57872 );
or ( n80037 , n80035 , n80036 );
and ( n80038 , n80033 , n80037 );
and ( n80039 , n34301 , n57880 );
or ( n80040 , n80038 , n80039 );
and ( n80041 , n80032 , n80040 );
not ( n80042 , n57900 );
not ( n80043 , n57902 );
and ( n80044 , n80043 , n80040 );
and ( n80045 , n34761 , n57902 );
or ( n80046 , n80044 , n80045 );
and ( n80047 , n80042 , n80046 );
and ( n80048 , n35050 , n57900 );
or ( n80049 , n80047 , n80048 );
and ( n80050 , n80049 , n32968 );
or ( n80051 , n80041 , n80050 );
and ( n80052 , n80051 , n33370 );
and ( n80053 , n32769 , n35062 );
or ( n80054 , C0 , n80022 , n80031 , n80052 , n80053 );
buf ( n80055 , n80054 );
buf ( n80056 , n80055 );
buf ( n80057 , n31655 );
buf ( n80058 , n30987 );
buf ( n80059 , n30987 );
buf ( n80060 , n30987 );
buf ( n80061 , n31655 );
buf ( n80062 , n31655 );
buf ( n80063 , n30987 );
not ( n80064 , n34150 );
and ( n80065 , n80064 , n32640 );
not ( n80066 , n56192 );
and ( n80067 , n80066 , n32640 );
and ( n80068 , n32655 , n56192 );
or ( n80069 , n80067 , n80068 );
and ( n80070 , n80069 , n34150 );
or ( n80071 , n80065 , n80070 );
and ( n80072 , n80071 , n33381 );
not ( n80073 , n56200 );
not ( n80074 , n56192 );
and ( n80075 , n80074 , n32640 );
and ( n80076 , n56044 , n56192 );
or ( n80077 , n80075 , n80076 );
and ( n80078 , n80073 , n80077 );
and ( n80079 , n56044 , n56200 );
or ( n80080 , n80078 , n80079 );
and ( n80081 , n80080 , n33375 );
not ( n80082 , n32968 );
not ( n80083 , n56200 );
not ( n80084 , n56192 );
and ( n80085 , n80084 , n32640 );
and ( n80086 , n56044 , n56192 );
or ( n80087 , n80085 , n80086 );
and ( n80088 , n80083 , n80087 );
and ( n80089 , n56044 , n56200 );
or ( n80090 , n80088 , n80089 );
and ( n80091 , n80082 , n80090 );
not ( n80092 , n56220 );
not ( n80093 , n56222 );
and ( n80094 , n80093 , n80090 );
and ( n80095 , n56068 , n56222 );
or ( n80096 , n80094 , n80095 );
and ( n80097 , n80092 , n80096 );
and ( n80098 , n56076 , n56220 );
or ( n80099 , n80097 , n80098 );
and ( n80100 , n80099 , n32968 );
or ( n80101 , n80091 , n80100 );
and ( n80102 , n80101 , n33370 );
and ( n80103 , n32640 , n35062 );
or ( n80104 , C0 , n80072 , n80081 , n80102 , n80103 );
buf ( n80105 , n80104 );
buf ( n80106 , n80105 );
not ( n80107 , n34150 );
and ( n80108 , n80107 , n32887 );
not ( n80109 , n56239 );
and ( n80110 , n80109 , n32887 );
and ( n80111 , n32889 , n56239 );
or ( n80112 , n80110 , n80111 );
and ( n80113 , n80112 , n34150 );
or ( n80114 , n80108 , n80113 );
and ( n80115 , n80114 , n33381 );
not ( n80116 , n56247 );
not ( n80117 , n56239 );
and ( n80118 , n80117 , n32887 );
and ( n80119 , n52819 , n56239 );
or ( n80120 , n80118 , n80119 );
and ( n80121 , n80116 , n80120 );
and ( n80122 , n52819 , n56247 );
or ( n80123 , n80121 , n80122 );
and ( n80124 , n80123 , n33375 );
not ( n80125 , n32968 );
not ( n80126 , n56247 );
not ( n80127 , n56239 );
and ( n80128 , n80127 , n32887 );
and ( n80129 , n52819 , n56239 );
or ( n80130 , n80128 , n80129 );
and ( n80131 , n80126 , n80130 );
and ( n80132 , n52819 , n56247 );
or ( n80133 , n80131 , n80132 );
and ( n80134 , n80125 , n80133 );
not ( n80135 , n56267 );
not ( n80136 , n56269 );
and ( n80137 , n80136 , n80133 );
and ( n80138 , n52845 , n56269 );
or ( n80139 , n80137 , n80138 );
and ( n80140 , n80135 , n80139 );
and ( n80141 , n52855 , n56267 );
or ( n80142 , n80140 , n80141 );
and ( n80143 , n80142 , n32968 );
or ( n80144 , n80134 , n80143 );
and ( n80145 , n80144 , n33370 );
and ( n80146 , n32887 , n35062 );
or ( n80147 , C0 , n80115 , n80124 , n80145 , n80146 );
buf ( n80148 , n80147 );
buf ( n80149 , n80148 );
buf ( n80150 , n31655 );
buf ( n80151 , n30987 );
not ( n80152 , n46356 );
and ( n80153 , n80152 , n31248 );
not ( n80154 , n78324 );
and ( n80155 , n80154 , n31248 );
and ( n80156 , n31272 , n78324 );
or ( n80157 , n80155 , n80156 );
and ( n80158 , n80157 , n46356 );
or ( n80159 , n80153 , n80158 );
and ( n80160 , n80159 , n31649 );
not ( n80161 , n78332 );
not ( n80162 , n78324 );
and ( n80163 , n80162 , n31248 );
and ( n80164 , n49443 , n78324 );
or ( n80165 , n80163 , n80164 );
and ( n80166 , n80161 , n80165 );
and ( n80167 , n49443 , n78332 );
or ( n80168 , n80166 , n80167 );
and ( n80169 , n80168 , n31643 );
not ( n80170 , n31452 );
not ( n80171 , n78332 );
not ( n80172 , n78324 );
and ( n80173 , n80172 , n31248 );
and ( n80174 , n49443 , n78324 );
or ( n80175 , n80173 , n80174 );
and ( n80176 , n80171 , n80175 );
and ( n80177 , n49443 , n78332 );
or ( n80178 , n80176 , n80177 );
and ( n80179 , n80170 , n80178 );
not ( n80180 , n78352 );
not ( n80181 , n78354 );
and ( n80182 , n80181 , n80178 );
and ( n80183 , n49469 , n78354 );
or ( n80184 , n80182 , n80183 );
and ( n80185 , n80180 , n80184 );
and ( n80186 , n49477 , n78352 );
or ( n80187 , n80185 , n80186 );
and ( n80188 , n80187 , n31452 );
or ( n80189 , n80179 , n80188 );
and ( n80190 , n80189 , n31638 );
and ( n80191 , n31248 , n47277 );
or ( n80192 , C0 , n80160 , n80169 , n80190 , n80191 );
buf ( n80193 , n80192 );
buf ( n80194 , n80193 );
buf ( n80195 , n31655 );
buf ( n80196 , RI15b5ea28_1094);
and ( n80197 , n80196 , n32494 );
not ( n80198 , n46083 );
and ( n80199 , n80198 , n66178 );
buf ( n80200 , n80199 );
and ( n80201 , n80200 , n32421 );
not ( n80202 , n46326 );
and ( n80203 , n80202 , n66178 );
not ( n80204 , n51396 );
and ( n80205 , n80204 , n51188 );
xor ( n80206 , n51403 , n51407 );
and ( n80207 , n80206 , n51396 );
or ( n80208 , n80205 , n80207 );
and ( n80209 , n80208 , n46326 );
or ( n80210 , n80203 , n80209 );
and ( n80211 , n80210 , n32417 );
and ( n80212 , n66178 , n46340 );
or ( n80213 , n80201 , n80211 , n80212 );
and ( n80214 , n80213 , n32456 );
and ( n80215 , n66178 , n46349 );
or ( n80216 , C0 , n80197 , n80214 , n80215 );
buf ( n80217 , n80216 );
buf ( n80218 , n80217 );
xor ( n80219 , n39415 , n54967 );
and ( n80220 , n80219 , n33199 );
not ( n80221 , n48648 );
and ( n80222 , n80221 , n39415 );
and ( n80223 , n34234 , n48648 );
or ( n80224 , n80222 , n80223 );
and ( n80225 , n80224 , n32924 );
not ( n80226 , n48660 );
and ( n80227 , n80226 , n39415 );
not ( n80228 , n39584 );
and ( n80229 , n80228 , n48543 );
not ( n80230 , n39775 );
and ( n80231 , n80230 , n39639 );
xor ( n80232 , n42660 , n42665 );
and ( n80233 , n80232 , n39775 );
or ( n80234 , n80231 , n80233 );
and ( n80235 , n80234 , n39584 );
or ( n80236 , n80229 , n80235 );
and ( n80237 , n80236 , n48660 );
or ( n80238 , n80227 , n80237 );
and ( n80239 , n80238 , n33172 );
not ( n80240 , n48730 );
and ( n80241 , n80240 , n39415 );
and ( n80242 , n48902 , n48730 );
or ( n80243 , n80241 , n80242 );
and ( n80244 , n80243 , n33187 );
and ( n80245 , n39415 , n54713 );
or ( n80246 , n80220 , n80225 , n80239 , n80244 , n80245 );
and ( n80247 , n80246 , n33208 );
and ( n80248 , n39415 , n39805 );
or ( n80249 , C0 , n80247 , n80248 );
buf ( n80250 , n80249 );
buf ( n80251 , n80250 );
buf ( n80252 , n31655 );
buf ( n80253 , n30987 );
buf ( n80254 , n30987 );
buf ( n80255 , n31655 );
not ( n80256 , n41532 );
buf ( n80257 , n80256 );
buf ( n80258 , n80257 );
buf ( n80259 , n30987 );
and ( n80260 , n49066 , n48639 );
not ( n80261 , n48642 );
and ( n80262 , n80261 , n48591 );
and ( n80263 , n49066 , n48642 );
or ( n80264 , n80262 , n80263 );
and ( n80265 , n80264 , n32890 );
not ( n80266 , n48648 );
and ( n80267 , n80266 , n48591 );
and ( n80268 , n49066 , n48648 );
or ( n80269 , n80267 , n80268 );
and ( n80270 , n80269 , n32924 );
not ( n80271 , n48654 );
and ( n80272 , n80271 , n48591 );
and ( n80273 , n49066 , n48654 );
or ( n80274 , n80272 , n80273 );
and ( n80275 , n80274 , n33038 );
not ( n80276 , n48660 );
and ( n80277 , n80276 , n48591 );
and ( n80278 , n49066 , n48660 );
or ( n80279 , n80277 , n80278 );
and ( n80280 , n80279 , n33172 );
not ( n80281 , n41576 );
and ( n80282 , n80281 , n48591 );
and ( n80283 , n48776 , n41576 );
or ( n80284 , n80282 , n80283 );
and ( n80285 , n80284 , n33189 );
not ( n80286 , n48730 );
and ( n80287 , n80286 , n48591 );
and ( n80288 , n48776 , n48730 );
or ( n80289 , n80287 , n80288 );
and ( n80290 , n80289 , n33187 );
not ( n80291 , n48765 );
and ( n80292 , n80291 , n48591 );
and ( n80293 , n62511 , n48765 );
or ( n80294 , n80292 , n80293 );
and ( n80295 , n80294 , n33180 );
not ( n80296 , n49054 );
and ( n80297 , n80296 , n48591 );
and ( n80298 , n62522 , n49054 );
or ( n80299 , n80297 , n80298 );
and ( n80300 , n80299 , n33178 );
and ( n80301 , n49175 , n49275 );
or ( n80302 , n80260 , n80265 , n80270 , n80275 , n80280 , n80285 , n80290 , n80295 , n80300 , n80301 );
and ( n80303 , n80302 , n33208 );
and ( n80304 , n32984 , n35056 );
and ( n80305 , n48591 , n49286 );
or ( n80306 , C0 , n80303 , n80304 , n80305 );
buf ( n80307 , n80306 );
buf ( n80308 , n80307 );
buf ( n80309 , n31655 );
buf ( n80310 , n31655 );
buf ( n80311 , n30987 );
buf ( n80312 , n30987 );
not ( n80313 , n36587 );
and ( n80314 , n80313 , n36430 );
xor ( n80315 , n50175 , n50212 );
and ( n80316 , n80315 , n36587 );
or ( n80317 , n80314 , n80316 );
and ( n80318 , n80317 , n36596 );
not ( n80319 , n37485 );
and ( n80320 , n80319 , n37332 );
xor ( n80321 , n50225 , n50262 );
and ( n80322 , n80321 , n37485 );
or ( n80323 , n80320 , n80322 );
and ( n80324 , n80323 , n37494 );
and ( n80325 , n41859 , n37506 );
or ( n80326 , n80318 , n80324 , n80325 );
buf ( n80327 , n80326 );
buf ( n80328 , n80327 );
buf ( n80329 , n31655 );
and ( n80330 , n50442 , n50275 );
not ( n80331 , n50278 );
and ( n80332 , n80331 , n50410 );
and ( n80333 , n50442 , n50278 );
or ( n80334 , n80332 , n80333 );
and ( n80335 , n80334 , n32421 );
not ( n80336 , n50002 );
and ( n80337 , n80336 , n50410 );
and ( n80338 , n50442 , n50002 );
or ( n80339 , n80337 , n80338 );
and ( n80340 , n80339 , n32419 );
not ( n80341 , n50289 );
and ( n80342 , n80341 , n50410 );
and ( n80343 , n50442 , n50289 );
or ( n80344 , n80342 , n80343 );
and ( n80345 , n80344 , n32417 );
not ( n80346 , n50008 );
and ( n80347 , n80346 , n50410 );
and ( n80348 , n50442 , n50008 );
or ( n80349 , n80347 , n80348 );
and ( n80350 , n80349 , n32415 );
not ( n80351 , n47331 );
and ( n80352 , n80351 , n50410 );
and ( n80353 , n50420 , n47331 );
or ( n80354 , n80352 , n80353 );
and ( n80355 , n80354 , n32413 );
not ( n80356 , n50067 );
and ( n80357 , n80356 , n50410 );
and ( n80358 , n50420 , n50067 );
or ( n80359 , n80357 , n80358 );
and ( n80360 , n80359 , n32411 );
not ( n80361 , n31728 );
and ( n80362 , n80361 , n50410 );
xor ( n80363 , n50420 , n50423 );
and ( n80364 , n80363 , n31728 );
or ( n80365 , n80362 , n80364 );
and ( n80366 , n80365 , n32253 );
not ( n80367 , n32283 );
and ( n80368 , n80367 , n50410 );
not ( n80369 , n31823 );
xor ( n80370 , n50442 , n50445 );
and ( n80371 , n80369 , n80370 );
xnor ( n80372 , n50459 , n50462 );
and ( n80373 , n80372 , n31823 );
or ( n80374 , n80371 , n80373 );
and ( n80375 , n80374 , n32283 );
or ( n80376 , n80368 , n80375 );
and ( n80377 , n80376 , n32398 );
and ( n80378 , n50459 , n50334 );
or ( n80379 , n80330 , n80335 , n80340 , n80345 , n80350 , n80355 , n80360 , n80366 , n80377 , n80378 );
and ( n80380 , n80379 , n32456 );
and ( n80381 , n37537 , n32489 );
and ( n80382 , n50410 , n50345 );
or ( n80383 , C0 , n80380 , n80381 , n80382 );
buf ( n80384 , n80383 );
buf ( n80385 , n80384 );
buf ( n80386 , n30987 );
buf ( n80387 , n40204 );
not ( n80388 , n34150 );
and ( n80389 , n80388 , n32631 );
not ( n80390 , n57038 );
and ( n80391 , n80390 , n32631 );
and ( n80392 , n32655 , n57038 );
or ( n80393 , n80391 , n80392 );
and ( n80394 , n80393 , n34150 );
or ( n80395 , n80389 , n80394 );
and ( n80396 , n80395 , n33381 );
not ( n80397 , n57046 );
not ( n80398 , n57038 );
and ( n80399 , n80398 , n32631 );
and ( n80400 , n56044 , n57038 );
or ( n80401 , n80399 , n80400 );
and ( n80402 , n80397 , n80401 );
and ( n80403 , n56044 , n57046 );
or ( n80404 , n80402 , n80403 );
and ( n80405 , n80404 , n33375 );
not ( n80406 , n32968 );
not ( n80407 , n57046 );
not ( n80408 , n57038 );
and ( n80409 , n80408 , n32631 );
and ( n80410 , n56044 , n57038 );
or ( n80411 , n80409 , n80410 );
and ( n80412 , n80407 , n80411 );
and ( n80413 , n56044 , n57046 );
or ( n80414 , n80412 , n80413 );
and ( n80415 , n80406 , n80414 );
not ( n80416 , n57066 );
not ( n80417 , n57068 );
and ( n80418 , n80417 , n80414 );
and ( n80419 , n56068 , n57068 );
or ( n80420 , n80418 , n80419 );
and ( n80421 , n80416 , n80420 );
and ( n80422 , n56076 , n57066 );
or ( n80423 , n80421 , n80422 );
and ( n80424 , n80423 , n32968 );
or ( n80425 , n80415 , n80424 );
and ( n80426 , n80425 , n33370 );
and ( n80427 , n32631 , n35062 );
or ( n80428 , C0 , n80396 , n80405 , n80426 , n80427 );
buf ( n80429 , n80428 );
buf ( n80430 , n80429 );
buf ( n80431 , n30987 );
buf ( n80432 , n31655 );
buf ( n80433 , n31655 );
buf ( n80434 , n31655 );
not ( n80435 , n38443 );
and ( n80436 , n80435 , n38031 );
xor ( n80437 , n53480 , n53489 );
and ( n80438 , n80437 , n38443 );
or ( n80439 , n80436 , n80438 );
and ( n80440 , n80439 , n38450 );
not ( n80441 , n39339 );
and ( n80442 , n80441 , n38931 );
xor ( n80443 , n53536 , n53545 );
and ( n80444 , n80443 , n39339 );
or ( n80445 , n80442 , n80444 );
and ( n80446 , n80445 , n39346 );
and ( n80447 , n40204 , n39359 );
or ( n80448 , n80440 , n80446 , n80447 );
buf ( n80449 , n80448 );
buf ( n80450 , n80449 );
buf ( n80451 , RI15b54438_740);
and ( n80452 , n80451 , n58921 );
and ( n80453 , n41527 , n37506 );
or ( n80454 , n80452 , n80453 );
buf ( n80455 , n80454 );
buf ( n80456 , n80455 );
buf ( n80457 , n30987 );
xor ( n80458 , n35441 , n39943 );
and ( n80459 , n80458 , n31550 );
not ( n80460 , n39979 );
and ( n80461 , n80460 , n35441 );
and ( n80462 , n55875 , n39979 );
or ( n80463 , n80461 , n80462 );
and ( n80464 , n80463 , n31538 );
and ( n80465 , n35441 , n40143 );
or ( n80466 , n80459 , n80464 , n80465 );
and ( n80467 , n80466 , n31557 );
and ( n80468 , n35441 , n40154 );
or ( n80469 , C0 , n80467 , n80468 );
buf ( n80470 , n80469 );
buf ( n80471 , n80470 );
buf ( n80472 , RI15b47508_298);
buf ( n80473 , n80472 );
buf ( n80474 , n31655 );
not ( n80475 , n40163 );
and ( n80476 , n80475 , n31959 );
not ( n80477 , n75905 );
and ( n80478 , n80477 , n31959 );
and ( n80479 , n32183 , n75905 );
or ( n80480 , n80478 , n80479 );
and ( n80481 , n80480 , n40163 );
or ( n80482 , n80476 , n80481 );
and ( n80483 , n80482 , n32498 );
not ( n80484 , n75913 );
not ( n80485 , n75905 );
and ( n80486 , n80485 , n31959 );
and ( n80487 , n45178 , n75905 );
or ( n80488 , n80486 , n80487 );
and ( n80489 , n80484 , n80488 );
and ( n80490 , n45178 , n75913 );
or ( n80491 , n80489 , n80490 );
and ( n80492 , n80491 , n32473 );
not ( n80493 , n32475 );
not ( n80494 , n75913 );
not ( n80495 , n75905 );
and ( n80496 , n80495 , n31959 );
and ( n80497 , n45178 , n75905 );
or ( n80498 , n80496 , n80497 );
and ( n80499 , n80494 , n80498 );
and ( n80500 , n45178 , n75913 );
or ( n80501 , n80499 , n80500 );
and ( n80502 , n80493 , n80501 );
not ( n80503 , n75933 );
not ( n80504 , n75935 );
and ( n80505 , n80504 , n80501 );
and ( n80506 , n45206 , n75935 );
or ( n80507 , n80505 , n80506 );
and ( n80508 , n80503 , n80507 );
and ( n80509 , n45214 , n75933 );
or ( n80510 , n80508 , n80509 );
and ( n80511 , n80510 , n32475 );
or ( n80512 , n80502 , n80511 );
and ( n80513 , n80512 , n32486 );
and ( n80514 , n31959 , n41278 );
or ( n80515 , C0 , n80483 , n80492 , n80513 , n80514 );
buf ( n80516 , n80515 );
buf ( n80517 , n80516 );
buf ( n80518 , n30987 );
buf ( n80519 , n30987 );
buf ( n80520 , n30987 );
buf ( n80521 , n31655 );
not ( n80522 , n46356 );
and ( n80523 , n80522 , n31360 );
not ( n80524 , n64746 );
and ( n80525 , n80524 , n31360 );
and ( n80526 , n31372 , n64746 );
or ( n80527 , n80525 , n80526 );
and ( n80528 , n80527 , n46356 );
or ( n80529 , n80523 , n80528 );
and ( n80530 , n80529 , n31649 );
not ( n80531 , n64754 );
not ( n80532 , n64746 );
and ( n80533 , n80532 , n31360 );
and ( n80534 , n47849 , n64746 );
or ( n80535 , n80533 , n80534 );
and ( n80536 , n80531 , n80535 );
and ( n80537 , n47849 , n64754 );
or ( n80538 , n80536 , n80537 );
and ( n80539 , n80538 , n31643 );
not ( n80540 , n31452 );
not ( n80541 , n64754 );
not ( n80542 , n64746 );
and ( n80543 , n80542 , n31360 );
and ( n80544 , n47849 , n64746 );
or ( n80545 , n80543 , n80544 );
and ( n80546 , n80541 , n80545 );
and ( n80547 , n47849 , n64754 );
or ( n80548 , n80546 , n80547 );
and ( n80549 , n80540 , n80548 );
not ( n80550 , n64774 );
not ( n80551 , n64776 );
and ( n80552 , n80551 , n80548 );
and ( n80553 , n47877 , n64776 );
or ( n80554 , n80552 , n80553 );
and ( n80555 , n80550 , n80554 );
and ( n80556 , n47887 , n64774 );
or ( n80557 , n80555 , n80556 );
and ( n80558 , n80557 , n31452 );
or ( n80559 , n80549 , n80558 );
and ( n80560 , n80559 , n31638 );
and ( n80561 , n31360 , n47277 );
or ( n80562 , C0 , n80530 , n80539 , n80560 , n80561 );
buf ( n80563 , n80562 );
buf ( n80564 , n80563 );
buf ( n80565 , n31655 );
xor ( n80566 , n50973 , n64710 );
and ( n80567 , n80566 , n32431 );
not ( n80568 , n50002 );
and ( n80569 , n80568 , n50973 );
and ( n80570 , n40648 , n50002 );
or ( n80571 , n80569 , n80570 );
and ( n80572 , n80571 , n32419 );
not ( n80573 , n50008 );
and ( n80574 , n80573 , n50973 );
not ( n80575 , n51594 );
and ( n80576 , n80575 , n51434 );
xor ( n80577 , n51602 , n51604 );
and ( n80578 , n80577 , n51594 );
or ( n80579 , n80576 , n80578 );
and ( n80580 , n80579 , n50008 );
or ( n80581 , n80574 , n80580 );
and ( n80582 , n80581 , n32415 );
not ( n80583 , n50067 );
and ( n80584 , n80583 , n50973 );
and ( n80585 , n65687 , n50067 );
or ( n80586 , n80584 , n80585 );
and ( n80587 , n80586 , n32411 );
and ( n80588 , n50973 , n50098 );
or ( n80589 , n80567 , n80572 , n80582 , n80587 , n80588 );
and ( n80590 , n80589 , n32456 );
and ( n80591 , n50973 , n47409 );
or ( n80592 , C0 , n80590 , n80591 );
buf ( n80593 , n80592 );
buf ( n80594 , n80593 );
not ( n80595 , n40163 );
and ( n80596 , n80595 , n32027 );
not ( n80597 , n42238 );
and ( n80598 , n80597 , n32027 );
and ( n80599 , n32147 , n42238 );
or ( n80600 , n80598 , n80599 );
and ( n80601 , n80600 , n40163 );
or ( n80602 , n80596 , n80601 );
and ( n80603 , n80602 , n32498 );
not ( n80604 , n42247 );
not ( n80605 , n42238 );
and ( n80606 , n80605 , n32027 );
and ( n80607 , n49314 , n42238 );
or ( n80608 , n80606 , n80607 );
and ( n80609 , n80604 , n80608 );
and ( n80610 , n49314 , n42247 );
or ( n80611 , n80609 , n80610 );
and ( n80612 , n80611 , n32473 );
not ( n80613 , n32475 );
not ( n80614 , n42247 );
not ( n80615 , n42238 );
and ( n80616 , n80615 , n32027 );
and ( n80617 , n49314 , n42238 );
or ( n80618 , n80616 , n80617 );
and ( n80619 , n80614 , n80618 );
and ( n80620 , n49314 , n42247 );
or ( n80621 , n80619 , n80620 );
and ( n80622 , n80613 , n80621 );
not ( n80623 , n42273 );
not ( n80624 , n42276 );
and ( n80625 , n80624 , n80621 );
and ( n80626 , n49340 , n42276 );
or ( n80627 , n80625 , n80626 );
and ( n80628 , n80623 , n80627 );
and ( n80629 , n49348 , n42273 );
or ( n80630 , n80628 , n80629 );
and ( n80631 , n80630 , n32475 );
or ( n80632 , n80622 , n80631 );
and ( n80633 , n80632 , n32486 );
and ( n80634 , n32027 , n41278 );
or ( n80635 , C0 , n80603 , n80612 , n80633 , n80634 );
buf ( n80636 , n80635 );
buf ( n80637 , n80636 );
buf ( n80638 , n31655 );
xor ( n80639 , n34040 , n39937 );
and ( n80640 , n80639 , n31550 );
not ( n80641 , n39979 );
and ( n80642 , n80641 , n34040 );
and ( n80643 , n49413 , n39979 );
or ( n80644 , n80642 , n80643 );
and ( n80645 , n80644 , n31538 );
and ( n80646 , n34040 , n40143 );
or ( n80647 , n80640 , n80645 , n80646 );
and ( n80648 , n80647 , n31557 );
and ( n80649 , n34040 , n40154 );
or ( n80650 , C0 , n80648 , n80649 );
buf ( n80651 , n80650 );
buf ( n80652 , n80651 );
buf ( n80653 , n30987 );
buf ( n80654 , n30987 );
and ( n80655 , n33232 , n32528 );
not ( n80656 , n32598 );
and ( n80657 , n80656 , n32995 );
buf ( n80658 , n80657 );
and ( n80659 , n80658 , n32890 );
not ( n80660 , n32919 );
and ( n80661 , n80660 , n32995 );
buf ( n80662 , n80661 );
and ( n80663 , n80662 , n32924 );
not ( n80664 , n32953 );
and ( n80665 , n80664 , n32995 );
not ( n80666 , n32971 );
and ( n80667 , n80666 , n33115 );
xor ( n80668 , n32995 , n33010 );
and ( n80669 , n80668 , n32971 );
or ( n80670 , n80667 , n80669 );
and ( n80671 , n80670 , n32953 );
or ( n80672 , n80665 , n80671 );
and ( n80673 , n80672 , n33038 );
not ( n80674 , n33067 );
and ( n80675 , n80674 , n32995 );
not ( n80676 , n32970 );
not ( n80677 , n33071 );
and ( n80678 , n80677 , n33115 );
xor ( n80679 , n33116 , n33142 );
and ( n80680 , n80679 , n33071 );
or ( n80681 , n80678 , n80680 );
and ( n80682 , n80676 , n80681 );
and ( n80683 , n80668 , n32970 );
or ( n80684 , n80682 , n80683 );
and ( n80685 , n80684 , n33067 );
or ( n80686 , n80675 , n80685 );
and ( n80687 , n80686 , n33172 );
and ( n80688 , n32995 , n33204 );
or ( n80689 , n80659 , n80663 , n80673 , n80687 , n80688 );
and ( n80690 , n80689 , n33208 );
not ( n80691 , n32968 );
not ( n80692 , n33270 );
and ( n80693 , n80692 , n33315 );
xor ( n80694 , n33316 , n33342 );
and ( n80695 , n80694 , n33270 );
or ( n80696 , n80693 , n80695 );
and ( n80697 , n80691 , n80696 );
and ( n80698 , n32995 , n32968 );
or ( n80699 , n80697 , n80698 );
and ( n80700 , n80699 , n33370 );
buf ( n80701 , n35056 );
and ( n80702 , n32995 , n33382 );
or ( n80703 , C0 , n80655 , n80690 , n80700 , n80701 , n80702 );
buf ( n80704 , n80703 );
buf ( n80705 , n80704 );
buf ( n80706 , n31655 );
buf ( n80707 , n30987 );
buf ( n80708 , n30987 );
buf ( n80709 , n31655 );
not ( n80710 , n31728 );
and ( n80711 , n80710 , n46018 );
and ( n80712 , n71537 , n31728 );
or ( n80713 , n80711 , n80712 );
and ( n80714 , n80713 , n32253 );
not ( n80715 , n32283 );
and ( n80716 , n80715 , n46018 );
and ( n80717 , n71548 , n32283 );
or ( n80718 , n80716 , n80717 );
and ( n80719 , n80718 , n32398 );
and ( n80720 , n46018 , n32436 );
or ( n80721 , n80714 , n80719 , n80720 );
and ( n80722 , n80721 , n32456 );
and ( n80723 , n49654 , n32473 );
not ( n80724 , n32475 );
and ( n80725 , n80724 , n49654 );
xor ( n80726 , n46018 , n50481 );
and ( n80727 , n80726 , n32475 );
or ( n80728 , n80725 , n80727 );
and ( n80729 , n80728 , n32486 );
and ( n80730 , n37533 , n32489 );
and ( n80731 , n46018 , n32501 );
or ( n80732 , C0 , n80722 , n80723 , n80729 , n80730 , n80731 );
buf ( n80733 , n80732 );
buf ( n80734 , n80733 );
and ( n80735 , n50897 , n32494 );
not ( n80736 , n46083 );
and ( n80737 , n80736 , n76458 );
buf ( n80738 , n80737 );
and ( n80739 , n80738 , n32421 );
not ( n80740 , n46326 );
and ( n80741 , n80740 , n76458 );
and ( n80742 , n51414 , n46326 );
or ( n80743 , n80741 , n80742 );
and ( n80744 , n80743 , n32417 );
and ( n80745 , n76458 , n46340 );
or ( n80746 , n80739 , n80744 , n80745 );
and ( n80747 , n80746 , n32456 );
and ( n80748 , n76458 , n46349 );
or ( n80749 , C0 , n80735 , n80747 , n80748 );
buf ( n80750 , n80749 );
buf ( n80751 , n80750 );
buf ( n80752 , n31655 );
not ( n80753 , n46356 );
and ( n80754 , n80753 , n31101 );
not ( n80755 , n78324 );
and ( n80756 , n80755 , n31101 );
and ( n80757 , n31138 , n78324 );
or ( n80758 , n80756 , n80757 );
and ( n80759 , n80758 , n46356 );
or ( n80760 , n80754 , n80759 );
and ( n80761 , n80760 , n31649 );
not ( n80762 , n78332 );
not ( n80763 , n78324 );
and ( n80764 , n80763 , n31101 );
and ( n80765 , n56920 , n78324 );
or ( n80766 , n80764 , n80765 );
and ( n80767 , n80762 , n80766 );
and ( n80768 , n56920 , n78332 );
or ( n80769 , n80767 , n80768 );
and ( n80770 , n80769 , n31643 );
not ( n80771 , n31452 );
not ( n80772 , n78332 );
not ( n80773 , n78324 );
and ( n80774 , n80773 , n31101 );
and ( n80775 , n56920 , n78324 );
or ( n80776 , n80774 , n80775 );
and ( n80777 , n80772 , n80776 );
and ( n80778 , n56920 , n78332 );
or ( n80779 , n80777 , n80778 );
and ( n80780 , n80771 , n80779 );
not ( n80781 , n78352 );
not ( n80782 , n78354 );
and ( n80783 , n80782 , n80779 );
and ( n80784 , n56946 , n78354 );
or ( n80785 , n80783 , n80784 );
and ( n80786 , n80781 , n80785 );
and ( n80787 , n56954 , n78352 );
or ( n80788 , n80786 , n80787 );
and ( n80789 , n80788 , n31452 );
or ( n80790 , n80780 , n80789 );
and ( n80791 , n80790 , n31638 );
and ( n80792 , n31101 , n47277 );
or ( n80793 , C0 , n80761 , n80770 , n80791 , n80792 );
buf ( n80794 , n80793 );
buf ( n80795 , n80794 );
buf ( n80796 , n30987 );
buf ( n80797 , n31655 );
buf ( n80798 , n30987 );
buf ( n80799 , n31655 );
buf ( n80800 , RI15b466f8_268);
and ( n80801 , n80800 , n33377 );
not ( n80802 , n48545 );
and ( n80803 , n80802 , n35538 );
buf ( n80804 , n80803 );
and ( n80805 , n80804 , n32890 );
not ( n80806 , n48557 );
and ( n80807 , n80806 , n35538 );
not ( n80808 , n54581 );
and ( n80809 , n80808 , n54577 );
xor ( n80810 , n54577 , n54340 );
and ( n80811 , n76750 , n76751 );
xor ( n80812 , n80810 , n80811 );
and ( n80813 , n80812 , n54581 );
or ( n80814 , n80809 , n80813 );
and ( n80815 , n80814 , n48557 );
or ( n80816 , n80807 , n80815 );
and ( n80817 , n80816 , n33038 );
and ( n80818 , n35538 , n48571 );
or ( n80819 , n80805 , n80817 , n80818 );
and ( n80820 , n80819 , n33208 );
and ( n80821 , n35538 , n48577 );
or ( n80822 , C0 , n80801 , n80820 , n80821 );
buf ( n80823 , n80822 );
buf ( n80824 , n80823 );
buf ( n80825 , n31655 );
buf ( n80826 , n30987 );
buf ( n80827 , n31655 );
buf ( n80828 , n30987 );
not ( n80829 , n40163 );
and ( n80830 , n80829 , n31988 );
not ( n80831 , n45161 );
and ( n80832 , n80831 , n31988 );
and ( n80833 , n32165 , n45161 );
or ( n80834 , n80832 , n80833 );
and ( n80835 , n80834 , n40163 );
or ( n80836 , n80830 , n80835 );
and ( n80837 , n80836 , n32498 );
not ( n80838 , n45170 );
not ( n80839 , n45161 );
and ( n80840 , n80839 , n31988 );
and ( n80841 , n59005 , n45161 );
or ( n80842 , n80840 , n80841 );
and ( n80843 , n80838 , n80842 );
and ( n80844 , n59005 , n45170 );
or ( n80845 , n80843 , n80844 );
and ( n80846 , n80845 , n32473 );
not ( n80847 , n32475 );
not ( n80848 , n45170 );
not ( n80849 , n45161 );
and ( n80850 , n80849 , n31988 );
and ( n80851 , n59005 , n45161 );
or ( n80852 , n80850 , n80851 );
and ( n80853 , n80848 , n80852 );
and ( n80854 , n59005 , n45170 );
or ( n80855 , n80853 , n80854 );
and ( n80856 , n80847 , n80855 );
not ( n80857 , n45196 );
not ( n80858 , n45199 );
and ( n80859 , n80858 , n80855 );
and ( n80860 , n59029 , n45199 );
or ( n80861 , n80859 , n80860 );
and ( n80862 , n80857 , n80861 );
and ( n80863 , n59037 , n45196 );
or ( n80864 , n80862 , n80863 );
and ( n80865 , n80864 , n32475 );
or ( n80866 , n80856 , n80865 );
and ( n80867 , n80866 , n32486 );
and ( n80868 , n31988 , n41278 );
or ( n80869 , C0 , n80837 , n80846 , n80867 , n80868 );
buf ( n80870 , n80869 );
buf ( n80871 , n80870 );
xor ( n80872 , n45330 , n61852 );
and ( n80873 , n80872 , n31548 );
not ( n80874 , n44807 );
and ( n80875 , n80874 , n45330 );
and ( n80876 , n46611 , n44807 );
or ( n80877 , n80875 , n80876 );
and ( n80878 , n80877 , n31408 );
not ( n80879 , n44817 );
and ( n80880 , n80879 , n45330 );
not ( n80881 , n44994 );
and ( n80882 , n80881 , n44990 );
xor ( n80883 , n44990 , n41881 );
and ( n80884 , n44997 , n45023 );
xor ( n80885 , n80883 , n80884 );
and ( n80886 , n80885 , n44994 );
or ( n80887 , n80882 , n80886 );
and ( n80888 , n80887 , n44817 );
or ( n80889 , n80880 , n80888 );
and ( n80890 , n80889 , n31521 );
not ( n80891 , n45059 );
and ( n80892 , n80891 , n45330 );
and ( n80893 , n31340 , n40003 );
and ( n80894 , n31342 , n40005 );
and ( n80895 , n31344 , n40007 );
and ( n80896 , n31346 , n40009 );
and ( n80897 , n31348 , n40011 );
and ( n80898 , n31350 , n40013 );
and ( n80899 , n31352 , n40015 );
and ( n80900 , n31354 , n40017 );
and ( n80901 , n31356 , n40019 );
and ( n80902 , n31358 , n40021 );
and ( n80903 , n31360 , n40023 );
and ( n80904 , n31362 , n40025 );
and ( n80905 , n31364 , n40027 );
and ( n80906 , n31366 , n40029 );
and ( n80907 , n31368 , n40031 );
and ( n80908 , n31370 , n40033 );
or ( n80909 , n80893 , n80894 , n80895 , n80896 , n80897 , n80898 , n80899 , n80900 , n80901 , n80902 , n80903 , n80904 , n80905 , n80906 , n80907 , n80908 );
and ( n80910 , n45078 , n45135 );
xor ( n80911 , n80909 , n80910 );
and ( n80912 , n80911 , n45059 );
or ( n80913 , n80892 , n80912 );
and ( n80914 , n80913 , n31536 );
and ( n80915 , n45330 , n45148 );
or ( n80916 , n80873 , n80878 , n80890 , n80914 , n80915 );
and ( n80917 , n80916 , n31557 );
and ( n80918 , n45330 , n40154 );
or ( n80919 , C0 , n80917 , n80918 );
buf ( n80920 , n80919 );
buf ( n80921 , n80920 );
buf ( n80922 , n30987 );
not ( n80923 , n31728 );
and ( n80924 , n80923 , n35182 );
and ( n80925 , n65789 , n31728 );
or ( n80926 , n80924 , n80925 );
and ( n80927 , n80926 , n32253 );
not ( n80928 , n32283 );
and ( n80929 , n80928 , n35182 );
and ( n80930 , n65800 , n32283 );
or ( n80931 , n80929 , n80930 );
and ( n80932 , n80931 , n32398 );
and ( n80933 , n35182 , n32436 );
or ( n80934 , n80927 , n80932 , n80933 );
and ( n80935 , n80934 , n32456 );
and ( n80936 , n35182 , n32473 );
buf ( n80937 , n35182 );
and ( n80938 , n80937 , n32486 );
and ( n80939 , n35213 , n32489 );
and ( n80940 , n35182 , n32501 );
or ( n80941 , C0 , n80935 , n80936 , n80938 , n80939 , n80940 );
buf ( n80942 , n80941 );
buf ( n80943 , n80942 );
buf ( n80944 , n31655 );
buf ( n80945 , n30987 );
not ( n80946 , n46356 );
and ( n80947 , n80946 , n31135 );
not ( n80948 , n60564 );
and ( n80949 , n80948 , n31135 );
and ( n80950 , n31138 , n60564 );
or ( n80951 , n80949 , n80950 );
and ( n80952 , n80951 , n46356 );
or ( n80953 , n80947 , n80952 );
and ( n80954 , n80953 , n31649 );
not ( n80955 , n60572 );
not ( n80956 , n60564 );
and ( n80957 , n80956 , n31135 );
and ( n80958 , n56920 , n60564 );
or ( n80959 , n80957 , n80958 );
and ( n80960 , n80955 , n80959 );
and ( n80961 , n56920 , n60572 );
or ( n80962 , n80960 , n80961 );
and ( n80963 , n80962 , n31643 );
not ( n80964 , n31452 );
not ( n80965 , n60572 );
not ( n80966 , n60564 );
and ( n80967 , n80966 , n31135 );
and ( n80968 , n56920 , n60564 );
or ( n80969 , n80967 , n80968 );
and ( n80970 , n80965 , n80969 );
and ( n80971 , n56920 , n60572 );
or ( n80972 , n80970 , n80971 );
and ( n80973 , n80964 , n80972 );
not ( n80974 , n60592 );
not ( n80975 , n60594 );
and ( n80976 , n80975 , n80972 );
and ( n80977 , n56946 , n60594 );
or ( n80978 , n80976 , n80977 );
and ( n80979 , n80974 , n80978 );
and ( n80980 , n56954 , n60592 );
or ( n80981 , n80979 , n80980 );
and ( n80982 , n80981 , n31452 );
or ( n80983 , n80973 , n80982 );
and ( n80984 , n80983 , n31638 );
and ( n80985 , n31135 , n47277 );
or ( n80986 , C0 , n80954 , n80963 , n80984 , n80985 );
buf ( n80987 , n80986 );
buf ( n80988 , n80987 );
buf ( n80989 , n30987 );
buf ( n80990 , n31655 );
buf ( n80991 , n30987 );
not ( n80992 , n33419 );
and ( n80993 , n80992 , n31572 );
and ( n80994 , n76312 , n33419 );
or ( n80995 , n80993 , n80994 );
and ( n80996 , n80995 , n31529 );
not ( n80997 , n33734 );
and ( n80998 , n80997 , n31572 );
and ( n80999 , n76323 , n33734 );
or ( n81000 , n80998 , n80999 );
and ( n81001 , n81000 , n31527 );
and ( n81002 , n31572 , n33942 );
or ( n81003 , n80996 , n81001 , n81002 );
and ( n81004 , n81003 , n31557 );
and ( n81005 , n35499 , n31643 );
not ( n81006 , n31452 );
and ( n81007 , n81006 , n35499 );
xor ( n81008 , n31572 , n33965 );
and ( n81009 , n81008 , n31452 );
or ( n81010 , n81007 , n81009 );
and ( n81011 , n81010 , n31638 );
and ( n81012 , n35397 , n33973 );
and ( n81013 , n31572 , n33978 );
or ( n81014 , C0 , n81004 , n81005 , n81011 , n81012 , n81013 );
buf ( n81015 , n81014 );
buf ( n81016 , n81015 );
and ( n81017 , n31572 , n31007 );
not ( n81018 , n31077 );
and ( n81019 , n81018 , n35397 );
buf ( n81020 , n81019 );
and ( n81021 , n81020 , n31373 );
not ( n81022 , n31402 );
and ( n81023 , n81022 , n35397 );
buf ( n81024 , n81023 );
and ( n81025 , n81024 , n31408 );
not ( n81026 , n31437 );
and ( n81027 , n81026 , n35397 );
not ( n81028 , n31455 );
and ( n81029 , n81028 , n35445 );
xor ( n81030 , n35397 , n35400 );
and ( n81031 , n81030 , n31455 );
or ( n81032 , n81029 , n81031 );
and ( n81033 , n81032 , n31437 );
or ( n81034 , n81027 , n81033 );
and ( n81035 , n81034 , n31468 );
not ( n81036 , n31497 );
and ( n81037 , n81036 , n35397 );
not ( n81038 , n31454 );
not ( n81039 , n31501 );
and ( n81040 , n81039 , n35445 );
xor ( n81041 , n35446 , n35450 );
and ( n81042 , n81041 , n31501 );
or ( n81043 , n81040 , n81042 );
and ( n81044 , n81038 , n81043 );
and ( n81045 , n81030 , n31454 );
or ( n81046 , n81044 , n81045 );
and ( n81047 , n81046 , n31497 );
or ( n81048 , n81037 , n81047 );
and ( n81049 , n81048 , n31521 );
and ( n81050 , n35397 , n31553 );
or ( n81051 , n81021 , n81025 , n81035 , n81049 , n81050 );
and ( n81052 , n81051 , n31557 );
not ( n81053 , n31452 );
not ( n81054 , n31619 );
and ( n81055 , n81054 , n35499 );
xor ( n81056 , n35500 , n35504 );
and ( n81057 , n81056 , n31619 );
or ( n81058 , n81055 , n81057 );
and ( n81059 , n81053 , n81058 );
and ( n81060 , n35397 , n31452 );
or ( n81061 , n81059 , n81060 );
and ( n81062 , n81061 , n31638 );
buf ( n81063 , n33973 );
and ( n81064 , n35397 , n31650 );
or ( n81065 , C0 , n81017 , n81052 , n81062 , n81063 , n81064 );
buf ( n81066 , n81065 );
buf ( n81067 , n81066 );
buf ( n81068 , n30987 );
buf ( n81069 , n31655 );
buf ( n81070 , n31655 );
buf ( n81071 , n31655 );
not ( n81072 , n40163 );
and ( n81073 , n81072 , n31972 );
not ( n81074 , n53227 );
and ( n81075 , n81074 , n31972 );
and ( n81076 , n32165 , n53227 );
or ( n81077 , n81075 , n81076 );
and ( n81078 , n81077 , n40163 );
or ( n81079 , n81073 , n81078 );
and ( n81080 , n81079 , n32498 );
not ( n81081 , n53235 );
not ( n81082 , n53227 );
and ( n81083 , n81082 , n31972 );
and ( n81084 , n59005 , n53227 );
or ( n81085 , n81083 , n81084 );
and ( n81086 , n81081 , n81085 );
and ( n81087 , n59005 , n53235 );
or ( n81088 , n81086 , n81087 );
and ( n81089 , n81088 , n32473 );
not ( n81090 , n32475 );
not ( n81091 , n53235 );
not ( n81092 , n53227 );
and ( n81093 , n81092 , n31972 );
and ( n81094 , n59005 , n53227 );
or ( n81095 , n81093 , n81094 );
and ( n81096 , n81091 , n81095 );
and ( n81097 , n59005 , n53235 );
or ( n81098 , n81096 , n81097 );
and ( n81099 , n81090 , n81098 );
not ( n81100 , n53260 );
not ( n81101 , n53262 );
and ( n81102 , n81101 , n81098 );
and ( n81103 , n59029 , n53262 );
or ( n81104 , n81102 , n81103 );
and ( n81105 , n81100 , n81104 );
and ( n81106 , n59037 , n53260 );
or ( n81107 , n81105 , n81106 );
and ( n81108 , n81107 , n32475 );
or ( n81109 , n81099 , n81108 );
and ( n81110 , n81109 , n32486 );
and ( n81111 , n31972 , n41278 );
or ( n81112 , C0 , n81080 , n81089 , n81110 , n81111 );
buf ( n81113 , n81112 );
buf ( n81114 , n81113 );
and ( n81115 , n65626 , n31645 );
not ( n81116 , n45274 );
and ( n81117 , n81116 , n78269 );
not ( n81118 , n41809 );
and ( n81119 , n81118 , n41766 );
xor ( n81120 , n62434 , n62437 );
and ( n81121 , n81120 , n41809 );
or ( n81122 , n81119 , n81121 );
and ( n81123 , n81122 , n45274 );
or ( n81124 , n81117 , n81123 );
and ( n81125 , n81124 , n31373 );
not ( n81126 , n45280 );
and ( n81127 , n81126 , n78269 );
and ( n81128 , n81122 , n45280 );
or ( n81129 , n81127 , n81128 );
and ( n81130 , n81129 , n31468 );
and ( n81131 , n78269 , n45802 );
or ( n81132 , n81125 , n81130 , n81131 );
and ( n81133 , n81132 , n31557 );
and ( n81134 , n78269 , n45808 );
or ( n81135 , C0 , n81115 , n81133 , n81134 );
buf ( n81136 , n81135 );
buf ( n81137 , n81136 );
buf ( n81138 , n30987 );
buf ( n81139 , n31655 );
buf ( n81140 , n30987 );
buf ( n81141 , n30987 );
and ( n81142 , n55411 , n33377 );
not ( n81143 , n48545 );
buf ( n81144 , RI15b47148_290);
and ( n81145 , n81143 , n81144 );
not ( n81146 , n39572 );
and ( n81147 , n81146 , n39438 );
xor ( n81148 , n42623 , n42630 );
and ( n81149 , n81148 , n39572 );
or ( n81150 , n81147 , n81149 );
and ( n81151 , n81150 , n48545 );
or ( n81152 , n81145 , n81151 );
and ( n81153 , n81152 , n32890 );
not ( n81154 , n48557 );
and ( n81155 , n81154 , n81144 );
and ( n81156 , n81150 , n48557 );
or ( n81157 , n81155 , n81156 );
and ( n81158 , n81157 , n33038 );
and ( n81159 , n81144 , n48571 );
or ( n81160 , n81153 , n81158 , n81159 );
and ( n81161 , n81160 , n33208 );
and ( n81162 , n81144 , n48577 );
or ( n81163 , C0 , n81142 , n81161 , n81162 );
buf ( n81164 , n81163 );
buf ( n81165 , n81164 );
buf ( n81166 , n31655 );
not ( n81167 , n41532 );
and ( n81168 , n81167 , n34371 );
and ( n81169 , n78269 , n41532 );
or ( n81170 , n81168 , n81169 );
buf ( n81171 , n81170 );
buf ( n81172 , n81171 );
buf ( n81173 , n31655 );
buf ( n81174 , n30987 );
xor ( n81175 , n54140 , n78383 );
and ( n81176 , n81175 , n33199 );
not ( n81177 , n48648 );
and ( n81178 , n81177 , n54140 );
and ( n81179 , n34425 , n48648 );
or ( n81180 , n81178 , n81179 );
and ( n81181 , n81180 , n32924 );
not ( n81182 , n48660 );
and ( n81183 , n81182 , n54140 );
and ( n81184 , n67530 , n48660 );
or ( n81185 , n81183 , n81184 );
and ( n81186 , n81185 , n33172 );
not ( n81187 , n48730 );
and ( n81188 , n81187 , n54140 );
xor ( n81189 , n58523 , n78402 );
and ( n81190 , n81189 , n48730 );
or ( n81191 , n81188 , n81190 );
and ( n81192 , n81191 , n33187 );
and ( n81193 , n54140 , n54713 );
or ( n81194 , n81176 , n81181 , n81186 , n81192 , n81193 );
and ( n81195 , n81194 , n33208 );
and ( n81196 , n54140 , n39805 );
or ( n81197 , C0 , n81195 , n81196 );
buf ( n81198 , n81197 );
buf ( n81199 , n81198 );
buf ( n81200 , n30987 );
buf ( n81201 , n31655 );
not ( n81202 , n35211 );
and ( n81203 , n63293 , n81202 );
and ( n81204 , n81203 , n32421 );
not ( n81205 , n35245 );
and ( n81206 , n81205 , n63293 );
buf ( n81207 , n35245 );
or ( n81208 , n81206 , n81207 );
and ( n81209 , n81208 , n32419 );
not ( n81210 , n35278 );
and ( n81211 , n63293 , n81210 );
and ( n81212 , n81211 , n32417 );
not ( n81213 , n35331 );
and ( n81214 , n81213 , n63293 );
buf ( n81215 , n35331 );
or ( n81216 , n81214 , n81215 );
and ( n81217 , n81216 , n32415 );
and ( n81218 , n63293 , n35354 );
or ( n81219 , n81204 , n81209 , n81212 , n81217 , n81218 );
and ( n81220 , n81219 , n32456 );
or ( n81221 , n32486 , n32492 );
or ( n81222 , n81221 , n32473 );
or ( n81223 , n81222 , n32494 );
or ( n81224 , n81223 , n32496 );
or ( n81225 , n81224 , n32498 );
or ( n81226 , n81225 , n32500 );
and ( n81227 , n63293 , n81226 );
buf ( n81228 , n68574 );
or ( n81229 , C0 , n81220 , n81227 , n81228 );
buf ( n81230 , n81229 );
buf ( n81231 , n81230 );
buf ( n81232 , n30987 );
buf ( n81233 , n31655 );
buf ( n81234 , n31655 );
not ( n81235 , n46356 );
and ( n81236 , n81235 , n31252 );
not ( n81237 , n52734 );
and ( n81238 , n81237 , n31252 );
and ( n81239 , n31272 , n52734 );
or ( n81240 , n81238 , n81239 );
and ( n81241 , n81240 , n46356 );
or ( n81242 , n81236 , n81241 );
and ( n81243 , n81242 , n31649 );
not ( n81244 , n52742 );
not ( n81245 , n52734 );
and ( n81246 , n81245 , n31252 );
and ( n81247 , n49443 , n52734 );
or ( n81248 , n81246 , n81247 );
and ( n81249 , n81244 , n81248 );
and ( n81250 , n49443 , n52742 );
or ( n81251 , n81249 , n81250 );
and ( n81252 , n81251 , n31643 );
not ( n81253 , n31452 );
not ( n81254 , n52742 );
not ( n81255 , n52734 );
and ( n81256 , n81255 , n31252 );
and ( n81257 , n49443 , n52734 );
or ( n81258 , n81256 , n81257 );
and ( n81259 , n81254 , n81258 );
and ( n81260 , n49443 , n52742 );
or ( n81261 , n81259 , n81260 );
and ( n81262 , n81253 , n81261 );
not ( n81263 , n52762 );
not ( n81264 , n52764 );
and ( n81265 , n81264 , n81261 );
and ( n81266 , n49469 , n52764 );
or ( n81267 , n81265 , n81266 );
and ( n81268 , n81263 , n81267 );
and ( n81269 , n49477 , n52762 );
or ( n81270 , n81268 , n81269 );
and ( n81271 , n81270 , n31452 );
or ( n81272 , n81262 , n81271 );
and ( n81273 , n81272 , n31638 );
and ( n81274 , n31252 , n47277 );
or ( n81275 , C0 , n81243 , n81252 , n81273 , n81274 );
buf ( n81276 , n81275 );
buf ( n81277 , n81276 );
not ( n81278 , n34150 );
and ( n81279 , n81278 , n32667 );
not ( n81280 , n58762 );
and ( n81281 , n81280 , n32667 );
and ( n81282 , n32689 , n58762 );
or ( n81283 , n81281 , n81282 );
and ( n81284 , n81283 , n34150 );
or ( n81285 , n81279 , n81284 );
and ( n81286 , n81285 , n33381 );
not ( n81287 , n58770 );
not ( n81288 , n58762 );
and ( n81289 , n81288 , n32667 );
and ( n81290 , n50682 , n58762 );
or ( n81291 , n81289 , n81290 );
and ( n81292 , n81287 , n81291 );
and ( n81293 , n50682 , n58770 );
or ( n81294 , n81292 , n81293 );
and ( n81295 , n81294 , n33375 );
not ( n81296 , n32968 );
not ( n81297 , n58770 );
not ( n81298 , n58762 );
and ( n81299 , n81298 , n32667 );
and ( n81300 , n50682 , n58762 );
or ( n81301 , n81299 , n81300 );
and ( n81302 , n81297 , n81301 );
and ( n81303 , n50682 , n58770 );
or ( n81304 , n81302 , n81303 );
and ( n81305 , n81296 , n81304 );
not ( n81306 , n58790 );
not ( n81307 , n58792 );
and ( n81308 , n81307 , n81304 );
and ( n81309 , n50706 , n58792 );
or ( n81310 , n81308 , n81309 );
and ( n81311 , n81306 , n81310 );
and ( n81312 , n50714 , n58790 );
or ( n81313 , n81311 , n81312 );
and ( n81314 , n81313 , n32968 );
or ( n81315 , n81305 , n81314 );
and ( n81316 , n81315 , n33370 );
and ( n81317 , n32667 , n35062 );
or ( n81318 , C0 , n81286 , n81295 , n81316 , n81317 );
buf ( n81319 , n81318 );
buf ( n81320 , n81319 );
buf ( n81321 , n30987 );
buf ( n81322 , n31655 );
buf ( n81323 , n31655 );
buf ( n81324 , n30987 );
buf ( n81325 , n31655 );
not ( n81326 , n35542 );
and ( n81327 , n81326 , n41857 );
buf ( n81328 , RI15b458e8_238);
and ( n81329 , n81328 , n35542 );
or ( n81330 , n81327 , n81329 );
buf ( n81331 , n81330 );
buf ( n81332 , n81331 );
buf ( n81333 , n31655 );
not ( n81334 , n48765 );
and ( n81335 , n81334 , n32510 );
and ( n81336 , n48582 , n48696 );
xor ( n81337 , n56473 , n81336 );
and ( n81338 , n48697 , n49021 );
xor ( n81339 , n81337 , n81338 );
and ( n81340 , n81339 , n48765 );
or ( n81341 , n81335 , n81340 );
and ( n81342 , n81341 , n33180 );
not ( n81343 , n49054 );
and ( n81344 , n81343 , n32510 );
not ( n81345 , n48845 );
and ( n81346 , n48582 , n48637 );
xor ( n81347 , n56473 , n81346 );
and ( n81348 , n48638 , n49135 );
xor ( n81349 , n81347 , n81348 );
and ( n81350 , n81345 , n81349 );
and ( n81351 , n48582 , n49165 );
xor ( n81352 , n56473 , n81351 );
or ( n81353 , n49166 , n49261 );
xnor ( n81354 , n81352 , n81353 );
and ( n81355 , n81354 , n48845 );
or ( n81356 , n81350 , n81355 );
and ( n81357 , n81356 , n49054 );
or ( n81358 , n81344 , n81357 );
and ( n81359 , n81358 , n33178 );
and ( n81360 , n32510 , n49774 );
or ( n81361 , n81342 , n81359 , n81360 );
and ( n81362 , n81361 , n33208 );
and ( n81363 , n33272 , n33375 );
not ( n81364 , n32968 );
and ( n81365 , n81364 , n33272 );
and ( n81366 , n33212 , n66023 );
xor ( n81367 , n32510 , n81366 );
and ( n81368 , n81367 , n32968 );
or ( n81369 , n81365 , n81368 );
and ( n81370 , n81369 , n33370 );
and ( n81371 , n32600 , n35056 );
and ( n81372 , n32510 , n49794 );
or ( n81373 , C0 , n81362 , n81363 , n81370 , n81371 , n81372 );
buf ( n81374 , n81373 );
buf ( n81375 , n81374 );
and ( n81376 , n31730 , n32500 );
not ( n81377 , n35211 );
and ( n81378 , n81377 , n32488 );
buf ( n81379 , n81378 );
and ( n81380 , n81379 , n32421 );
not ( n81381 , n35245 );
and ( n81382 , n81381 , n32488 );
buf ( n81383 , n81382 );
and ( n81384 , n81383 , n32419 );
not ( n81385 , n35278 );
and ( n81386 , n81385 , n32488 );
not ( n81387 , n35295 );
and ( n81388 , n81387 , n47285 );
xor ( n81389 , n32488 , n49528 );
and ( n81390 , n81389 , n35295 );
or ( n81391 , n81388 , n81390 );
and ( n81392 , n81391 , n35278 );
or ( n81393 , n81386 , n81392 );
and ( n81394 , n81393 , n32417 );
not ( n81395 , n35331 );
and ( n81396 , n81395 , n32488 );
not ( n81397 , n35294 );
not ( n81398 , n45995 );
and ( n81399 , n81398 , n47285 );
xor ( n81400 , n49603 , n49614 );
and ( n81401 , n81400 , n45995 );
or ( n81402 , n81399 , n81401 );
and ( n81403 , n81397 , n81402 );
and ( n81404 , n81389 , n35294 );
or ( n81405 , n81403 , n81404 );
and ( n81406 , n81405 , n35331 );
or ( n81407 , n81396 , n81406 );
and ( n81408 , n81407 , n32415 );
and ( n81409 , n32488 , n35354 );
or ( n81410 , n81380 , n81384 , n81394 , n81408 , n81409 );
and ( n81411 , n81410 , n32456 );
not ( n81412 , n32475 );
not ( n81413 , n46060 );
and ( n81414 , n81413 , n32471 );
xor ( n81415 , n49694 , n49708 );
and ( n81416 , n81415 , n46060 );
or ( n81417 , n81414 , n81416 );
and ( n81418 , n81412 , n81417 );
and ( n81419 , n32488 , n32475 );
or ( n81420 , n81418 , n81419 );
and ( n81421 , n81420 , n32486 );
buf ( n81422 , n32489 );
and ( n81423 , n32488 , n35367 );
or ( n81424 , C0 , n81376 , n81411 , n81421 , n81422 , n81423 );
buf ( n81425 , n81424 );
buf ( n81426 , n81425 );
buf ( n81427 , n30987 );
buf ( n81428 , n30987 );
buf ( n81429 , n31655 );
and ( n81430 , n71254 , n32494 );
not ( n81431 , n46083 );
and ( n81432 , n81431 , n35529 );
buf ( n81433 , n81432 );
and ( n81434 , n81433 , n32421 );
not ( n81435 , n46326 );
and ( n81436 , n81435 , n35529 );
and ( n81437 , n71262 , n46326 );
or ( n81438 , n81436 , n81437 );
and ( n81439 , n81438 , n32417 );
and ( n81440 , n35529 , n46340 );
or ( n81441 , n81434 , n81439 , n81440 );
and ( n81442 , n81441 , n32456 );
and ( n81443 , n35529 , n46349 );
or ( n81444 , C0 , n81430 , n81442 , n81443 );
buf ( n81445 , n81444 );
buf ( n81446 , n81445 );
buf ( n81447 , n31655 );
not ( n81448 , n46356 );
and ( n81449 , n81448 , n31105 );
not ( n81450 , n53353 );
and ( n81451 , n81450 , n31105 );
and ( n81452 , n31138 , n53353 );
or ( n81453 , n81451 , n81452 );
and ( n81454 , n81453 , n46356 );
or ( n81455 , n81449 , n81454 );
and ( n81456 , n81455 , n31649 );
not ( n81457 , n53361 );
not ( n81458 , n53353 );
and ( n81459 , n81458 , n31105 );
and ( n81460 , n56920 , n53353 );
or ( n81461 , n81459 , n81460 );
and ( n81462 , n81457 , n81461 );
and ( n81463 , n56920 , n53361 );
or ( n81464 , n81462 , n81463 );
and ( n81465 , n81464 , n31643 );
not ( n81466 , n31452 );
not ( n81467 , n53361 );
not ( n81468 , n53353 );
and ( n81469 , n81468 , n31105 );
and ( n81470 , n56920 , n53353 );
or ( n81471 , n81469 , n81470 );
and ( n81472 , n81467 , n81471 );
and ( n81473 , n56920 , n53361 );
or ( n81474 , n81472 , n81473 );
and ( n81475 , n81466 , n81474 );
not ( n81476 , n53381 );
not ( n81477 , n53383 );
and ( n81478 , n81477 , n81474 );
and ( n81479 , n56946 , n53383 );
or ( n81480 , n81478 , n81479 );
and ( n81481 , n81476 , n81480 );
and ( n81482 , n56954 , n53381 );
or ( n81483 , n81481 , n81482 );
and ( n81484 , n81483 , n31452 );
or ( n81485 , n81475 , n81484 );
and ( n81486 , n81485 , n31638 );
and ( n81487 , n31105 , n47277 );
or ( n81488 , C0 , n81456 , n81465 , n81486 , n81487 );
buf ( n81489 , n81488 );
buf ( n81490 , n81489 );
buf ( n81491 , n30987 );
buf ( n81492 , n30987 );
buf ( n81493 , n31655 );
buf ( n81494 , n31655 );
buf ( n81495 , n30987 );
not ( n81496 , n41532 );
and ( n81497 , n81496 , n34423 );
and ( n81498 , n59978 , n41532 );
or ( n81499 , n81497 , n81498 );
buf ( n81500 , n81499 );
buf ( n81501 , n81500 );
xor ( n81502 , n39506 , n54974 );
and ( n81503 , n81502 , n33199 );
not ( n81504 , n48648 );
and ( n81505 , n81504 , n39506 );
and ( n81506 , n34373 , n48648 );
or ( n81507 , n81505 , n81506 );
and ( n81508 , n81507 , n32924 );
not ( n81509 , n48660 );
and ( n81510 , n81509 , n39506 );
not ( n81511 , n39584 );
and ( n81512 , n81511 , n74642 );
not ( n81513 , n39775 );
and ( n81514 , n81513 , n39723 );
xor ( n81515 , n42653 , n42672 );
and ( n81516 , n81515 , n39775 );
or ( n81517 , n81514 , n81516 );
and ( n81518 , n81517 , n39584 );
or ( n81519 , n81512 , n81518 );
and ( n81520 , n81519 , n48660 );
or ( n81521 , n81510 , n81520 );
and ( n81522 , n81521 , n33172 );
not ( n81523 , n48730 );
and ( n81524 , n81523 , n39506 );
and ( n81525 , n32723 , n52252 );
and ( n81526 , n32725 , n52254 );
and ( n81527 , n32727 , n52256 );
and ( n81528 , n32729 , n52258 );
and ( n81529 , n32731 , n52260 );
and ( n81530 , n32733 , n52262 );
and ( n81531 , n32735 , n52264 );
and ( n81532 , n32737 , n52266 );
and ( n81533 , n32739 , n52268 );
and ( n81534 , n32741 , n52270 );
and ( n81535 , n32743 , n52272 );
and ( n81536 , n32745 , n52274 );
and ( n81537 , n32747 , n52276 );
and ( n81538 , n32749 , n52278 );
and ( n81539 , n32751 , n52280 );
and ( n81540 , n32753 , n52282 );
or ( n81541 , n81525 , n81526 , n81527 , n81528 , n81529 , n81530 , n81531 , n81532 , n81533 , n81534 , n81535 , n81536 , n81537 , n81538 , n81539 , n81540 );
and ( n81542 , n81541 , n48730 );
or ( n81543 , n81524 , n81542 );
and ( n81544 , n81543 , n33187 );
and ( n81545 , n39506 , n54713 );
or ( n81546 , n81503 , n81508 , n81522 , n81544 , n81545 );
and ( n81547 , n81546 , n33208 );
and ( n81548 , n39506 , n39805 );
or ( n81549 , C0 , n81547 , n81548 );
buf ( n81550 , n81549 );
buf ( n81551 , n81550 );
buf ( n81552 , n30987 );
buf ( n81553 , n31655 );
buf ( n81554 , n31655 );
buf ( n81555 , n30987 );
not ( n81556 , n43755 );
and ( n81557 , n81556 , n43394 );
xor ( n81558 , n50501 , n50504 );
and ( n81559 , n81558 , n43755 );
or ( n81560 , n81557 , n81559 );
and ( n81561 , n81560 , n43774 );
not ( n81562 , n44663 );
and ( n81563 , n81562 , n44306 );
xor ( n81564 , n50519 , n50522 );
and ( n81565 , n81564 , n44663 );
or ( n81566 , n81563 , n81565 );
and ( n81567 , n81566 , n44682 );
and ( n81568 , n47416 , n44695 );
or ( n81569 , n81561 , n81567 , n81568 );
buf ( n81570 , n81569 );
buf ( n81571 , n81570 );
buf ( n81572 , n30987 );
and ( n81573 , n32306 , n50275 );
not ( n81574 , n50278 );
and ( n81575 , n81574 , n31739 );
and ( n81576 , n32306 , n50278 );
or ( n81577 , n81575 , n81576 );
and ( n81578 , n81577 , n32421 );
not ( n81579 , n50002 );
and ( n81580 , n81579 , n31739 );
and ( n81581 , n32306 , n50002 );
or ( n81582 , n81580 , n81581 );
and ( n81583 , n81582 , n32419 );
not ( n81584 , n50289 );
and ( n81585 , n81584 , n31739 );
and ( n81586 , n32306 , n50289 );
or ( n81587 , n81585 , n81586 );
and ( n81588 , n81587 , n32417 );
not ( n81589 , n50008 );
and ( n81590 , n81589 , n31739 );
and ( n81591 , n32306 , n50008 );
or ( n81592 , n81590 , n81591 );
and ( n81593 , n81592 , n32415 );
not ( n81594 , n47331 );
and ( n81595 , n81594 , n31739 );
and ( n81596 , n32000 , n47331 );
or ( n81597 , n81595 , n81596 );
and ( n81598 , n81597 , n32413 );
not ( n81599 , n50067 );
and ( n81600 , n81599 , n31739 );
and ( n81601 , n32000 , n50067 );
or ( n81602 , n81600 , n81601 );
and ( n81603 , n81602 , n32411 );
not ( n81604 , n31728 );
and ( n81605 , n81604 , n31739 );
and ( n81606 , n73829 , n31728 );
or ( n81607 , n81605 , n81606 );
and ( n81608 , n81607 , n32253 );
not ( n81609 , n32283 );
and ( n81610 , n81609 , n31739 );
and ( n81611 , n73842 , n32283 );
or ( n81612 , n81610 , n81611 );
and ( n81613 , n81612 , n32398 );
and ( n81614 , n32364 , n50334 );
or ( n81615 , n81573 , n81578 , n81583 , n81588 , n81593 , n81598 , n81603 , n81608 , n81613 , n81614 );
and ( n81616 , n81615 , n32456 );
and ( n81617 , n37514 , n32489 );
and ( n81618 , n31739 , n50345 );
or ( n81619 , C0 , n81616 , n81617 , n81618 );
buf ( n81620 , n81619 );
buf ( n81621 , n81620 );
not ( n81622 , n31437 );
buf ( n81623 , RI15b52a70_685);
and ( n81624 , n81622 , n81623 );
not ( n81625 , n45766 );
and ( n81626 , n81625 , n45728 );
xor ( n81627 , n45887 , n45892 );
and ( n81628 , n81627 , n45766 );
or ( n81629 , n81626 , n81628 );
and ( n81630 , n81629 , n31437 );
or ( n81631 , n81624 , n81630 );
and ( n81632 , n81631 , n31468 );
not ( n81633 , n44817 );
and ( n81634 , n81633 , n81623 );
and ( n81635 , n74129 , n44817 );
or ( n81636 , n81634 , n81635 );
and ( n81637 , n81636 , n31521 );
and ( n81638 , n81623 , n42158 );
or ( n81639 , n81632 , n81637 , n81638 );
and ( n81640 , n81639 , n31557 );
and ( n81641 , n81623 , n40154 );
or ( n81642 , C0 , n81640 , n81641 );
buf ( n81643 , n81642 );
buf ( n81644 , n81643 );
buf ( n81645 , n31655 );
and ( n81646 , n32296 , n50275 );
not ( n81647 , n50278 );
and ( n81648 , n81647 , n31734 );
and ( n81649 , n32296 , n50278 );
or ( n81650 , n81648 , n81649 );
and ( n81651 , n81650 , n32421 );
not ( n81652 , n50002 );
and ( n81653 , n81652 , n31734 );
and ( n81654 , n32296 , n50002 );
or ( n81655 , n81653 , n81654 );
and ( n81656 , n81655 , n32419 );
not ( n81657 , n50289 );
and ( n81658 , n81657 , n31734 );
and ( n81659 , n32296 , n50289 );
or ( n81660 , n81658 , n81659 );
and ( n81661 , n81660 , n32417 );
not ( n81662 , n50008 );
and ( n81663 , n81662 , n31734 );
and ( n81664 , n32296 , n50008 );
or ( n81665 , n81663 , n81664 );
and ( n81666 , n81665 , n32415 );
not ( n81667 , n47331 );
and ( n81668 , n81667 , n31734 );
and ( n81669 , n31825 , n47331 );
or ( n81670 , n81668 , n81669 );
and ( n81671 , n81670 , n32413 );
not ( n81672 , n50067 );
and ( n81673 , n81672 , n31734 );
and ( n81674 , n31825 , n50067 );
or ( n81675 , n81673 , n81674 );
and ( n81676 , n81675 , n32411 );
not ( n81677 , n31728 );
and ( n81678 , n81677 , n31734 );
and ( n81679 , n44730 , n31728 );
or ( n81680 , n81678 , n81679 );
and ( n81681 , n81680 , n32253 );
not ( n81682 , n32283 );
and ( n81683 , n81682 , n31734 );
and ( n81684 , n44743 , n32283 );
or ( n81685 , n81683 , n81684 );
and ( n81686 , n81685 , n32398 );
and ( n81687 , n32344 , n50334 );
or ( n81688 , n81646 , n81651 , n81656 , n81661 , n81666 , n81671 , n81676 , n81681 , n81686 , n81687 );
and ( n81689 , n81688 , n32456 );
and ( n81690 , n37577 , n32489 );
and ( n81691 , n31734 , n50345 );
or ( n81692 , C0 , n81689 , n81690 , n81691 );
buf ( n81693 , n81692 );
buf ( n81694 , n81693 );
buf ( n81695 , n30987 );
not ( n81696 , n31437 );
buf ( n81697 , RI15b52818_680);
and ( n81698 , n81696 , n81697 );
not ( n81699 , n45766 );
and ( n81700 , n81699 , n45643 );
xor ( n81701 , n45771 , n45785 );
and ( n81702 , n81701 , n45766 );
or ( n81703 , n81700 , n81702 );
and ( n81704 , n81703 , n31437 );
or ( n81705 , n81698 , n81704 );
and ( n81706 , n81705 , n31468 );
not ( n81707 , n44817 );
and ( n81708 , n81707 , n81697 );
not ( n81709 , n44994 );
and ( n81710 , n81709 , n44906 );
xor ( n81711 , n45003 , n45017 );
and ( n81712 , n81711 , n44994 );
or ( n81713 , n81710 , n81712 );
and ( n81714 , n81713 , n44817 );
or ( n81715 , n81708 , n81714 );
and ( n81716 , n81715 , n31521 );
and ( n81717 , n81697 , n42158 );
or ( n81718 , n81706 , n81716 , n81717 );
and ( n81719 , n81718 , n31557 );
and ( n81720 , n81697 , n40154 );
or ( n81721 , C0 , n81719 , n81720 );
buf ( n81722 , n81721 );
buf ( n81723 , n81722 );
buf ( n81724 , n31655 );
buf ( n81725 , n31655 );
buf ( n81726 , n30987 );
not ( n81727 , n34150 );
and ( n81728 , n81727 , n32828 );
not ( n81729 , n60126 );
and ( n81730 , n81729 , n32828 );
and ( n81731 , n32856 , n60126 );
or ( n81732 , n81730 , n81731 );
and ( n81733 , n81732 , n34150 );
or ( n81734 , n81728 , n81733 );
and ( n81735 , n81734 , n33381 );
not ( n81736 , n60134 );
not ( n81737 , n60126 );
and ( n81738 , n81737 , n32828 );
and ( n81739 , n48160 , n60126 );
or ( n81740 , n81738 , n81739 );
and ( n81741 , n81736 , n81740 );
and ( n81742 , n48160 , n60134 );
or ( n81743 , n81741 , n81742 );
and ( n81744 , n81743 , n33375 );
not ( n81745 , n32968 );
not ( n81746 , n60134 );
not ( n81747 , n60126 );
and ( n81748 , n81747 , n32828 );
and ( n81749 , n48160 , n60126 );
or ( n81750 , n81748 , n81749 );
and ( n81751 , n81746 , n81750 );
and ( n81752 , n48160 , n60134 );
or ( n81753 , n81751 , n81752 );
and ( n81754 , n81745 , n81753 );
not ( n81755 , n60154 );
not ( n81756 , n60156 );
and ( n81757 , n81756 , n81753 );
and ( n81758 , n48186 , n60156 );
or ( n81759 , n81757 , n81758 );
and ( n81760 , n81755 , n81759 );
and ( n81761 , n48196 , n60154 );
or ( n81762 , n81760 , n81761 );
and ( n81763 , n81762 , n32968 );
or ( n81764 , n81754 , n81763 );
and ( n81765 , n81764 , n33370 );
and ( n81766 , n32828 , n35062 );
or ( n81767 , C0 , n81735 , n81744 , n81765 , n81766 );
buf ( n81768 , n81767 );
buf ( n81769 , n81768 );
buf ( n81770 , n30987 );
buf ( n81771 , n31655 );
not ( n81772 , n32953 );
and ( n81773 , n81772 , n48543 );
and ( n81774 , n48553 , n32953 );
or ( n81775 , n81773 , n81774 );
and ( n81776 , n81775 , n33038 );
not ( n81777 , n39586 );
and ( n81778 , n81777 , n48543 );
and ( n81779 , n80234 , n39586 );
or ( n81780 , n81778 , n81779 );
and ( n81781 , n81780 , n33172 );
and ( n81782 , n48543 , n39795 );
or ( n81783 , n81776 , n81781 , n81782 );
and ( n81784 , n81783 , n33208 );
and ( n81785 , n48543 , n39805 );
or ( n81786 , C0 , n81784 , n81785 );
buf ( n81787 , n81786 );
buf ( n81788 , n81787 );
buf ( n81789 , n30987 );
buf ( n81790 , n31655 );
buf ( n81791 , n31655 );
buf ( n81792 , n30987 );
not ( n81793 , n46356 );
and ( n81794 , n81793 , n31197 );
not ( n81795 , n49427 );
and ( n81796 , n81795 , n31197 );
and ( n81797 , n31205 , n49427 );
or ( n81798 , n81796 , n81797 );
and ( n81799 , n81798 , n46356 );
or ( n81800 , n81794 , n81799 );
and ( n81801 , n81800 , n31649 );
not ( n81802 , n49435 );
not ( n81803 , n49427 );
and ( n81804 , n81803 , n31197 );
and ( n81805 , n50125 , n49427 );
or ( n81806 , n81804 , n81805 );
and ( n81807 , n81802 , n81806 );
and ( n81808 , n50125 , n49435 );
or ( n81809 , n81807 , n81808 );
and ( n81810 , n81809 , n31643 );
not ( n81811 , n31452 );
not ( n81812 , n49435 );
not ( n81813 , n49427 );
and ( n81814 , n81813 , n31197 );
and ( n81815 , n50125 , n49427 );
or ( n81816 , n81814 , n81815 );
and ( n81817 , n81812 , n81816 );
and ( n81818 , n50125 , n49435 );
or ( n81819 , n81817 , n81818 );
and ( n81820 , n81811 , n81819 );
not ( n81821 , n49460 );
not ( n81822 , n49462 );
and ( n81823 , n81822 , n81819 );
and ( n81824 , n50151 , n49462 );
or ( n81825 , n81823 , n81824 );
and ( n81826 , n81821 , n81825 );
and ( n81827 , n50159 , n49460 );
or ( n81828 , n81826 , n81827 );
and ( n81829 , n81828 , n31452 );
or ( n81830 , n81820 , n81829 );
and ( n81831 , n81830 , n31638 );
and ( n81832 , n31197 , n47277 );
or ( n81833 , C0 , n81801 , n81810 , n81831 , n81832 );
buf ( n81834 , n81833 );
buf ( n81835 , n81834 );
not ( n81836 , n35542 );
and ( n81837 , n81836 , n41863 );
and ( n81838 , n68176 , n35542 );
or ( n81839 , n81837 , n81838 );
buf ( n81840 , n81839 );
buf ( n81841 , n81840 );
xor ( n81842 , n47287 , n47295 );
and ( n81843 , n81842 , n32433 );
not ( n81844 , n47331 );
and ( n81845 , n81844 , n47287 );
buf ( n81846 , n31856 );
and ( n81847 , n81846 , n47331 );
or ( n81848 , n81845 , n81847 );
and ( n81849 , n81848 , n32413 );
and ( n81850 , n47287 , n47402 );
or ( n81851 , n81843 , n81849 , n81850 );
and ( n81852 , n81851 , n32456 );
and ( n81853 , n47287 , n47409 );
or ( n81854 , C0 , n81852 , n81853 );
buf ( n81855 , n81854 );
buf ( n81856 , n81855 );
buf ( n81857 , n31655 );
buf ( n81858 , n31655 );
buf ( n81859 , n30987 );
xor ( n81860 , n39389 , n54676 );
and ( n81861 , n81860 , n33199 );
not ( n81862 , n48648 );
and ( n81863 , n81862 , n39389 );
and ( n81864 , n34208 , n48648 );
or ( n81865 , n81863 , n81864 );
and ( n81866 , n81865 , n32924 );
not ( n81867 , n48660 );
and ( n81868 , n81867 , n39389 );
not ( n81869 , n39584 );
and ( n81870 , n81869 , n61232 );
and ( n81871 , n61248 , n39584 );
or ( n81872 , n81870 , n81871 );
and ( n81873 , n81872 , n48660 );
or ( n81874 , n81868 , n81873 );
and ( n81875 , n81874 , n33172 );
not ( n81876 , n48730 );
and ( n81877 , n81876 , n39389 );
and ( n81878 , n48940 , n48730 );
or ( n81879 , n81877 , n81878 );
and ( n81880 , n81879 , n33187 );
and ( n81881 , n39389 , n54713 );
or ( n81882 , n81861 , n81866 , n81875 , n81880 , n81881 );
and ( n81883 , n81882 , n33208 );
and ( n81884 , n39389 , n39805 );
or ( n81885 , C0 , n81883 , n81884 );
buf ( n81886 , n81885 );
buf ( n81887 , n81886 );
buf ( n81888 , n30987 );
buf ( n81889 , n30987 );
buf ( n81890 , n31655 );
buf ( n81891 , n31655 );
buf ( n81892 , n31655 );
not ( n81893 , n36587 );
and ( n81894 , n81893 , n36226 );
xor ( n81895 , n50187 , n50200 );
and ( n81896 , n81895 , n36587 );
or ( n81897 , n81894 , n81896 );
and ( n81898 , n81897 , n36596 );
not ( n81899 , n37485 );
and ( n81900 , n81899 , n37128 );
xor ( n81901 , n50237 , n50250 );
and ( n81902 , n81901 , n37485 );
or ( n81903 , n81900 , n81902 );
and ( n81904 , n81903 , n37494 );
and ( n81905 , n41847 , n37506 );
or ( n81906 , n81898 , n81904 , n81905 );
buf ( n81907 , n81906 );
buf ( n81908 , n81907 );
buf ( n81909 , n30987 );
not ( n81910 , n35292 );
and ( n81911 , n81910 , n32441 );
buf ( n81912 , n81911 );
and ( n81913 , n81912 , n32494 );
not ( n81914 , n76230 );
not ( n81915 , n76232 );
and ( n81916 , n81915 , n32441 );
buf ( n81917 , n76232 );
or ( n81918 , n81916 , n81917 );
and ( n81919 , n81918 , n32417 );
and ( n81920 , n32441 , n76244 );
or ( n81921 , n81919 , n81920 );
and ( n81922 , n81914 , n81921 );
buf ( n81923 , n76230 );
or ( n81924 , n81922 , n81923 );
and ( n81925 , n81924 , n32456 );
and ( n81926 , n76252 , n32492 );
not ( n81927 , n32475 );
and ( n81928 , n81927 , n32486 );
not ( n81929 , n76252 );
and ( n81930 , n81929 , n32491 );
or ( n81931 , C0 , C0 , C0 , n81913 , n81925 , C0 , n81926 , n81928 , n81930 , C0 );
buf ( n81932 , n81931 );
buf ( n81933 , n81932 );
buf ( n81934 , n31655 );
buf ( n81935 , n30987 );
and ( n81936 , n54132 , n79808 );
xor ( n81937 , n39374 , n81936 );
and ( n81938 , n81937 , n33199 );
not ( n81939 , n48648 );
and ( n81940 , n81939 , n39374 );
and ( n81941 , n34193 , n48648 );
or ( n81942 , n81940 , n81941 );
and ( n81943 , n81942 , n32924 );
not ( n81944 , n48660 );
and ( n81945 , n81944 , n39374 );
buf ( n81946 , n81945 );
and ( n81947 , n81946 , n33172 );
not ( n81948 , n48730 );
and ( n81949 , n81948 , n39374 );
buf ( n81950 , n81949 );
and ( n81951 , n81950 , n33187 );
and ( n81952 , n39374 , n54713 );
or ( n81953 , n81938 , n81943 , n81947 , n81951 , n81952 );
and ( n81954 , n81953 , n33208 );
and ( n81955 , n39374 , n39805 );
or ( n81956 , C0 , n81954 , n81955 );
buf ( n81957 , n81956 );
buf ( n81958 , n81957 );
buf ( n81959 , n30987 );
buf ( n81960 , n31655 );
not ( n81961 , n41532 );
and ( n81962 , n81961 , n34273 );
and ( n81963 , n73129 , n41532 );
or ( n81964 , n81962 , n81963 );
buf ( n81965 , n81964 );
buf ( n81966 , n81965 );
buf ( n81967 , n31655 );
buf ( n81968 , n30987 );
not ( n81969 , n35278 );
and ( n81970 , n81969 , n57416 );
and ( n81971 , n75735 , n35278 );
or ( n81972 , n81970 , n81971 );
and ( n81973 , n81972 , n32417 );
not ( n81974 , n47912 );
and ( n81975 , n81974 , n57416 );
and ( n81976 , n57422 , n47912 );
or ( n81977 , n81975 , n81976 );
and ( n81978 , n81977 , n32415 );
and ( n81979 , n57416 , n48133 );
or ( n81980 , n81973 , n81978 , n81979 );
and ( n81981 , n81980 , n32456 );
and ( n81982 , n57416 , n47409 );
or ( n81983 , C0 , n81981 , n81982 );
buf ( n81984 , n81983 );
buf ( n81985 , n81984 );
not ( n81986 , n46356 );
and ( n81987 , n81986 , n31086 );
not ( n81988 , n63024 );
and ( n81989 , n81988 , n31086 );
and ( n81990 , n31138 , n63024 );
or ( n81991 , n81989 , n81990 );
and ( n81992 , n81991 , n46356 );
or ( n81993 , n81987 , n81992 );
and ( n81994 , n81993 , n31649 );
not ( n81995 , n63032 );
not ( n81996 , n63024 );
and ( n81997 , n81996 , n31086 );
and ( n81998 , n56920 , n63024 );
or ( n81999 , n81997 , n81998 );
and ( n82000 , n81995 , n81999 );
and ( n82001 , n56920 , n63032 );
or ( n82002 , n82000 , n82001 );
and ( n82003 , n82002 , n31643 );
not ( n82004 , n31452 );
not ( n82005 , n63032 );
not ( n82006 , n63024 );
and ( n82007 , n82006 , n31086 );
and ( n82008 , n56920 , n63024 );
or ( n82009 , n82007 , n82008 );
and ( n82010 , n82005 , n82009 );
and ( n82011 , n56920 , n63032 );
or ( n82012 , n82010 , n82011 );
and ( n82013 , n82004 , n82012 );
not ( n82014 , n63052 );
not ( n82015 , n63054 );
and ( n82016 , n82015 , n82012 );
and ( n82017 , n56946 , n63054 );
or ( n82018 , n82016 , n82017 );
and ( n82019 , n82014 , n82018 );
and ( n82020 , n56954 , n63052 );
or ( n82021 , n82019 , n82020 );
and ( n82022 , n82021 , n31452 );
or ( n82023 , n82013 , n82022 );
and ( n82024 , n82023 , n31638 );
and ( n82025 , n31086 , n47277 );
or ( n82026 , C0 , n81994 , n82003 , n82024 , n82025 );
buf ( n82027 , n82026 );
buf ( n82028 , n82027 );
buf ( n82029 , n30987 );
buf ( n82030 , n30987 );
buf ( n82031 , n31655 );
not ( n82032 , n34150 );
and ( n82033 , n82032 , n32743 );
not ( n82034 , n56413 );
and ( n82035 , n82034 , n32743 );
and ( n82036 , n32755 , n56413 );
or ( n82037 , n82035 , n82036 );
and ( n82038 , n82037 , n34150 );
or ( n82039 , n82033 , n82038 );
and ( n82040 , n82039 , n33381 );
not ( n82041 , n56421 );
not ( n82042 , n56413 );
and ( n82043 , n82042 , n32743 );
and ( n82044 , n35083 , n56413 );
or ( n82045 , n82043 , n82044 );
and ( n82046 , n82041 , n82045 );
and ( n82047 , n35083 , n56421 );
or ( n82048 , n82046 , n82047 );
and ( n82049 , n82048 , n33375 );
not ( n82050 , n32968 );
not ( n82051 , n56421 );
not ( n82052 , n56413 );
and ( n82053 , n82052 , n32743 );
and ( n82054 , n35083 , n56413 );
or ( n82055 , n82053 , n82054 );
and ( n82056 , n82051 , n82055 );
and ( n82057 , n35083 , n56421 );
or ( n82058 , n82056 , n82057 );
and ( n82059 , n82050 , n82058 );
not ( n82060 , n56441 );
not ( n82061 , n56443 );
and ( n82062 , n82061 , n82058 );
and ( n82063 , n35107 , n56443 );
or ( n82064 , n82062 , n82063 );
and ( n82065 , n82060 , n82064 );
and ( n82066 , n35115 , n56441 );
or ( n82067 , n82065 , n82066 );
and ( n82068 , n82067 , n32968 );
or ( n82069 , n82059 , n82068 );
and ( n82070 , n82069 , n33370 );
and ( n82071 , n32743 , n35062 );
or ( n82072 , C0 , n82040 , n82049 , n82070 , n82071 );
buf ( n82073 , n82072 );
buf ( n82074 , n82073 );
not ( n82075 , n34150 );
and ( n82076 , n82075 , n32542 );
and ( n82077 , n34170 , n34150 );
or ( n82078 , n82076 , n82077 );
and ( n82079 , n82078 , n33381 );
not ( n82080 , n56687 );
not ( n82081 , n56464 );
and ( n82082 , n82081 , n32542 );
buf ( n82083 , n82082 );
and ( n82084 , n82080 , n82083 );
buf ( n82085 , n82084 );
and ( n82086 , n82085 , n33379 );
and ( n82087 , n34329 , n33375 );
not ( n82088 , n32968 );
and ( n82089 , n82088 , n34329 );
xor ( n82090 , n34333 , n34325 );
not ( n82091 , n82090 );
buf ( n82092 , n82091 );
not ( n82093 , n82092 );
and ( n82094 , n82093 , n32968 );
or ( n82095 , n82089 , n82094 );
and ( n82096 , n82095 , n33370 );
and ( n82097 , n32542 , n56699 );
or ( n82098 , C0 , n82079 , n82086 , n82087 , n82096 , n82097 );
buf ( n82099 , n82098 );
buf ( n82100 , n82099 );
buf ( n82101 , n31655 );
buf ( n82102 , n30987 );
buf ( n82103 , n30987 );
not ( n82104 , n34150 );
and ( n82105 , n82104 , n32811 );
not ( n82106 , n56413 );
and ( n82107 , n82106 , n32811 );
and ( n82108 , n32823 , n56413 );
or ( n82109 , n82107 , n82108 );
and ( n82110 , n82109 , n34150 );
or ( n82111 , n82105 , n82110 );
and ( n82112 , n82111 , n33381 );
not ( n82113 , n56421 );
not ( n82114 , n56413 );
and ( n82115 , n82114 , n32811 );
and ( n82116 , n41464 , n56413 );
or ( n82117 , n82115 , n82116 );
and ( n82118 , n82113 , n82117 );
and ( n82119 , n41464 , n56421 );
or ( n82120 , n82118 , n82119 );
and ( n82121 , n82120 , n33375 );
not ( n82122 , n32968 );
not ( n82123 , n56421 );
not ( n82124 , n56413 );
and ( n82125 , n82124 , n32811 );
and ( n82126 , n41464 , n56413 );
or ( n82127 , n82125 , n82126 );
and ( n82128 , n82123 , n82127 );
and ( n82129 , n41464 , n56421 );
or ( n82130 , n82128 , n82129 );
and ( n82131 , n82122 , n82130 );
not ( n82132 , n56441 );
not ( n82133 , n56443 );
and ( n82134 , n82133 , n82130 );
and ( n82135 , n41490 , n56443 );
or ( n82136 , n82134 , n82135 );
and ( n82137 , n82132 , n82136 );
and ( n82138 , n41500 , n56441 );
or ( n82139 , n82137 , n82138 );
and ( n82140 , n82139 , n32968 );
or ( n82141 , n82131 , n82140 );
and ( n82142 , n82141 , n33370 );
and ( n82143 , n32811 , n35062 );
or ( n82144 , C0 , n82112 , n82121 , n82142 , n82143 );
buf ( n82145 , n82144 );
buf ( n82146 , n82145 );
buf ( n82147 , n31655 );
buf ( n82148 , n31655 );
and ( n82149 , n57801 , n33208 );
and ( n82150 , n56464 , n39805 );
or ( n82151 , C0 , n82149 , n82150 );
buf ( n82152 , n82151 );
buf ( n82153 , n82152 );
buf ( n82154 , n30987 );
not ( n82155 , n40163 );
and ( n82156 , n82155 , n32038 );
not ( n82157 , n42171 );
and ( n82158 , n82157 , n32038 );
and ( n82159 , n32130 , n42171 );
or ( n82160 , n82158 , n82159 );
and ( n82161 , n82160 , n40163 );
or ( n82162 , n82156 , n82161 );
and ( n82163 , n82162 , n32498 );
not ( n82164 , n42180 );
not ( n82165 , n42171 );
and ( n82166 , n82165 , n32038 );
and ( n82167 , n45833 , n42171 );
or ( n82168 , n82166 , n82167 );
and ( n82169 , n82164 , n82168 );
and ( n82170 , n45833 , n42180 );
or ( n82171 , n82169 , n82170 );
and ( n82172 , n82171 , n32473 );
not ( n82173 , n32475 );
not ( n82174 , n42180 );
not ( n82175 , n42171 );
and ( n82176 , n82175 , n32038 );
and ( n82177 , n45833 , n42171 );
or ( n82178 , n82176 , n82177 );
and ( n82179 , n82174 , n82178 );
and ( n82180 , n45833 , n42180 );
or ( n82181 , n82179 , n82180 );
and ( n82182 , n82173 , n82181 );
not ( n82183 , n42206 );
not ( n82184 , n42209 );
and ( n82185 , n82184 , n82181 );
and ( n82186 , n45857 , n42209 );
or ( n82187 , n82185 , n82186 );
and ( n82188 , n82183 , n82187 );
and ( n82189 , n45865 , n42206 );
or ( n82190 , n82188 , n82189 );
and ( n82191 , n82190 , n32475 );
or ( n82192 , n82182 , n82191 );
and ( n82193 , n82192 , n32486 );
and ( n82194 , n32038 , n41278 );
or ( n82195 , C0 , n82163 , n82172 , n82193 , n82194 );
buf ( n82196 , n82195 );
buf ( n82197 , n82196 );
not ( n82198 , n31437 );
and ( n82199 , n82198 , n62425 );
and ( n82200 , n62442 , n31437 );
or ( n82201 , n82199 , n82200 );
and ( n82202 , n82201 , n31468 );
not ( n82203 , n41837 );
and ( n82204 , n82203 , n62425 );
not ( n82205 , n42124 );
and ( n82206 , n82205 , n42104 );
xor ( n82207 , n49374 , n49385 );
and ( n82208 , n82207 , n42124 );
or ( n82209 , n82206 , n82208 );
and ( n82210 , n82209 , n41837 );
or ( n82211 , n82204 , n82210 );
and ( n82212 , n82211 , n31521 );
and ( n82213 , n62425 , n42158 );
or ( n82214 , n82202 , n82212 , n82213 );
and ( n82215 , n82214 , n31557 );
and ( n82216 , n62425 , n40154 );
or ( n82217 , C0 , n82215 , n82216 );
buf ( n82218 , n82217 );
buf ( n82219 , n82218 );
buf ( n82220 , n31655 );
buf ( n82221 , n31655 );
buf ( n82222 , n30987 );
not ( n82223 , n34150 );
and ( n82224 , n82223 , n32661 );
not ( n82225 , n60126 );
and ( n82226 , n82225 , n32661 );
and ( n82227 , n32689 , n60126 );
or ( n82228 , n82226 , n82227 );
and ( n82229 , n82228 , n34150 );
or ( n82230 , n82224 , n82229 );
and ( n82231 , n82230 , n33381 );
not ( n82232 , n60134 );
not ( n82233 , n60126 );
and ( n82234 , n82233 , n32661 );
and ( n82235 , n50682 , n60126 );
or ( n82236 , n82234 , n82235 );
and ( n82237 , n82232 , n82236 );
and ( n82238 , n50682 , n60134 );
or ( n82239 , n82237 , n82238 );
and ( n82240 , n82239 , n33375 );
not ( n82241 , n32968 );
not ( n82242 , n60134 );
not ( n82243 , n60126 );
and ( n82244 , n82243 , n32661 );
and ( n82245 , n50682 , n60126 );
or ( n82246 , n82244 , n82245 );
and ( n82247 , n82242 , n82246 );
and ( n82248 , n50682 , n60134 );
or ( n82249 , n82247 , n82248 );
and ( n82250 , n82241 , n82249 );
not ( n82251 , n60154 );
not ( n82252 , n60156 );
and ( n82253 , n82252 , n82249 );
and ( n82254 , n50706 , n60156 );
or ( n82255 , n82253 , n82254 );
and ( n82256 , n82251 , n82255 );
and ( n82257 , n50714 , n60154 );
or ( n82258 , n82256 , n82257 );
and ( n82259 , n82258 , n32968 );
or ( n82260 , n82250 , n82259 );
and ( n82261 , n82260 , n33370 );
and ( n82262 , n32661 , n35062 );
or ( n82263 , C0 , n82231 , n82240 , n82261 , n82262 );
buf ( n82264 , n82263 );
buf ( n82265 , n82264 );
buf ( n82266 , n30987 );
buf ( n82267 , n31655 );
buf ( n82268 , n30987 );
buf ( n82269 , n31655 );
not ( n82270 , n40163 );
and ( n82271 , n82270 , n31832 );
not ( n82272 , n53227 );
and ( n82273 , n82272 , n31832 );
and ( n82274 , n32235 , n53227 );
or ( n82275 , n82273 , n82274 );
and ( n82276 , n82275 , n40163 );
or ( n82277 , n82271 , n82276 );
and ( n82278 , n82277 , n32498 );
not ( n82279 , n53235 );
not ( n82280 , n53227 );
and ( n82281 , n82280 , n31832 );
and ( n82282 , n42188 , n53227 );
or ( n82283 , n82281 , n82282 );
and ( n82284 , n82279 , n82283 );
and ( n82285 , n42188 , n53235 );
or ( n82286 , n82284 , n82285 );
and ( n82287 , n82286 , n32473 );
not ( n82288 , n32475 );
not ( n82289 , n53235 );
not ( n82290 , n53227 );
and ( n82291 , n82290 , n31832 );
and ( n82292 , n42188 , n53227 );
or ( n82293 , n82291 , n82292 );
and ( n82294 , n82289 , n82293 );
and ( n82295 , n42188 , n53235 );
or ( n82296 , n82294 , n82295 );
and ( n82297 , n82288 , n82296 );
not ( n82298 , n53260 );
not ( n82299 , n53262 );
and ( n82300 , n82299 , n82296 );
and ( n82301 , n42216 , n53262 );
or ( n82302 , n82300 , n82301 );
and ( n82303 , n82298 , n82302 );
and ( n82304 , n42224 , n53260 );
or ( n82305 , n82303 , n82304 );
and ( n82306 , n82305 , n32475 );
or ( n82307 , n82297 , n82306 );
and ( n82308 , n82307 , n32486 );
and ( n82309 , n31832 , n41278 );
or ( n82310 , C0 , n82278 , n82287 , n82308 , n82309 );
buf ( n82311 , n82310 );
buf ( n82312 , n82311 );
and ( n82313 , n41604 , n31645 );
not ( n82314 , n45274 );
and ( n82315 , n82314 , n58614 );
and ( n82316 , n41831 , n45274 );
or ( n82317 , n82315 , n82316 );
and ( n82318 , n82317 , n31373 );
not ( n82319 , n45280 );
and ( n82320 , n82319 , n58614 );
and ( n82321 , n41831 , n45280 );
or ( n82322 , n82320 , n82321 );
and ( n82323 , n82322 , n31468 );
and ( n82324 , n58614 , n45802 );
or ( n82325 , n82318 , n82323 , n82324 );
and ( n82326 , n82325 , n31557 );
and ( n82327 , n58614 , n45808 );
or ( n82328 , C0 , n82313 , n82326 , n82327 );
buf ( n82329 , n82328 );
buf ( n82330 , n82329 );
buf ( n82331 , n31655 );
buf ( n82332 , n30987 );
not ( n82333 , n46356 );
and ( n82334 , n82333 , n31282 );
not ( n82335 , n78324 );
and ( n82336 , n82335 , n31282 );
and ( n82337 , n31306 , n78324 );
or ( n82338 , n82336 , n82337 );
and ( n82339 , n82338 , n46356 );
or ( n82340 , n82334 , n82339 );
and ( n82341 , n82340 , n31649 );
not ( n82342 , n78332 );
not ( n82343 , n78324 );
and ( n82344 , n82343 , n31282 );
and ( n82345 , n58061 , n78324 );
or ( n82346 , n82344 , n82345 );
and ( n82347 , n82342 , n82346 );
and ( n82348 , n58061 , n78332 );
or ( n82349 , n82347 , n82348 );
and ( n82350 , n82349 , n31643 );
not ( n82351 , n31452 );
not ( n82352 , n78332 );
not ( n82353 , n78324 );
and ( n82354 , n82353 , n31282 );
and ( n82355 , n58061 , n78324 );
or ( n82356 , n82354 , n82355 );
and ( n82357 , n82352 , n82356 );
and ( n82358 , n58061 , n78332 );
or ( n82359 , n82357 , n82358 );
and ( n82360 , n82351 , n82359 );
not ( n82361 , n78352 );
not ( n82362 , n78354 );
and ( n82363 , n82362 , n82359 );
and ( n82364 , n58085 , n78354 );
or ( n82365 , n82363 , n82364 );
and ( n82366 , n82361 , n82365 );
and ( n82367 , n58093 , n78352 );
or ( n82368 , n82366 , n82367 );
and ( n82369 , n82368 , n31452 );
or ( n82370 , n82360 , n82369 );
and ( n82371 , n82370 , n31638 );
and ( n82372 , n31282 , n47277 );
or ( n82373 , C0 , n82341 , n82350 , n82371 , n82372 );
buf ( n82374 , n82373 );
buf ( n82375 , n82374 );
buf ( n82376 , n31655 );
buf ( n82377 , RI15b5e9b0_1093);
and ( n82378 , n82377 , n32494 );
not ( n82379 , n46083 );
buf ( n82380 , RI15b5ffb8_1140);
and ( n82381 , n82379 , n82380 );
buf ( n82382 , n82381 );
and ( n82383 , n82382 , n32421 );
not ( n82384 , n46326 );
and ( n82385 , n82384 , n82380 );
not ( n82386 , n51396 );
and ( n82387 , n82386 , n51171 );
xor ( n82388 , n51404 , n51406 );
and ( n82389 , n82388 , n51396 );
or ( n82390 , n82387 , n82389 );
and ( n82391 , n82390 , n46326 );
or ( n82392 , n82385 , n82391 );
and ( n82393 , n82392 , n32417 );
and ( n82394 , n82380 , n46340 );
or ( n82395 , n82383 , n82393 , n82394 );
and ( n82396 , n82395 , n32456 );
and ( n82397 , n82380 , n46349 );
or ( n82398 , C0 , n82378 , n82396 , n82397 );
buf ( n82399 , n82398 );
buf ( n82400 , n82399 );
buf ( n82401 , n31655 );
buf ( n82402 , n30987 );
not ( n82403 , n50828 );
not ( n82404 , n50834 );
and ( n82405 , n82404 , n40267 );
and ( n82406 , n59536 , n50834 );
or ( n82407 , n82405 , n82406 );
and ( n82408 , n82403 , n82407 );
buf ( n82409 , RI15b5f8b0_1125);
and ( n82410 , n82409 , n50828 );
or ( n82411 , n82408 , n82410 );
buf ( n82412 , n82411 );
buf ( n82413 , n82412 );
buf ( n82414 , n30987 );
buf ( n82415 , n31655 );
not ( n82416 , n48765 );
and ( n82417 , n82416 , n33237 );
and ( n82418 , n62630 , n48765 );
or ( n82419 , n82417 , n82418 );
and ( n82420 , n82419 , n33180 );
not ( n82421 , n49054 );
and ( n82422 , n82421 , n33237 );
and ( n82423 , n62643 , n49054 );
or ( n82424 , n82422 , n82423 );
and ( n82425 , n82424 , n33178 );
and ( n82426 , n33237 , n49774 );
or ( n82427 , n82420 , n82425 , n82426 );
and ( n82428 , n82427 , n33208 );
and ( n82429 , n33325 , n33375 );
not ( n82430 , n32968 );
and ( n82431 , n82430 , n33325 );
xor ( n82432 , n33237 , n49781 );
and ( n82433 , n82432 , n32968 );
or ( n82434 , n82431 , n82433 );
and ( n82435 , n82434 , n33370 );
and ( n82436 , n33000 , n35056 );
and ( n82437 , n33237 , n49794 );
or ( n82438 , C0 , n82428 , n82429 , n82435 , n82436 , n82437 );
buf ( n82439 , n82438 );
buf ( n82440 , n82439 );
buf ( n82441 , n31655 );
buf ( n82442 , n30987 );
buf ( n82443 , n30987 );
buf ( n82444 , n31655 );
not ( n82445 , n50828 );
buf ( n82446 , n82445 );
buf ( n82447 , n82446 );
xor ( n82448 , n39441 , n54969 );
and ( n82449 , n82448 , n33199 );
not ( n82450 , n48648 );
and ( n82451 , n82450 , n39441 );
and ( n82452 , n34260 , n48648 );
or ( n82453 , n82451 , n82452 );
and ( n82454 , n82453 , n32924 );
not ( n82455 , n48660 );
and ( n82456 , n82455 , n39441 );
not ( n82457 , n39584 );
and ( n82458 , n82457 , n58018 );
and ( n82459 , n58034 , n39584 );
or ( n82460 , n82458 , n82459 );
and ( n82461 , n82460 , n48660 );
or ( n82462 , n82456 , n82461 );
and ( n82463 , n82462 , n33172 );
not ( n82464 , n48730 );
and ( n82465 , n82464 , n39441 );
and ( n82466 , n48864 , n48730 );
or ( n82467 , n82465 , n82466 );
and ( n82468 , n82467 , n33187 );
and ( n82469 , n39441 , n54713 );
or ( n82470 , n82449 , n82454 , n82463 , n82468 , n82469 );
and ( n82471 , n82470 , n33208 );
and ( n82472 , n39441 , n39805 );
or ( n82473 , C0 , n82471 , n82472 );
buf ( n82474 , n82473 );
buf ( n82475 , n82474 );
buf ( n82476 , n31655 );
buf ( n82477 , n30987 );
not ( n82478 , n34150 );
and ( n82479 , n82478 , n32791 );
not ( n82480 , n56708 );
and ( n82481 , n82480 , n32791 );
and ( n82482 , n32823 , n56708 );
or ( n82483 , n82481 , n82482 );
and ( n82484 , n82483 , n34150 );
or ( n82485 , n82479 , n82484 );
and ( n82486 , n82485 , n33381 );
not ( n82487 , n56716 );
not ( n82488 , n56708 );
and ( n82489 , n82488 , n32791 );
and ( n82490 , n41464 , n56708 );
or ( n82491 , n82489 , n82490 );
and ( n82492 , n82487 , n82491 );
and ( n82493 , n41464 , n56716 );
or ( n82494 , n82492 , n82493 );
and ( n82495 , n82494 , n33375 );
not ( n82496 , n32968 );
not ( n82497 , n56716 );
not ( n82498 , n56708 );
and ( n82499 , n82498 , n32791 );
and ( n82500 , n41464 , n56708 );
or ( n82501 , n82499 , n82500 );
and ( n82502 , n82497 , n82501 );
and ( n82503 , n41464 , n56716 );
or ( n82504 , n82502 , n82503 );
and ( n82505 , n82496 , n82504 );
not ( n82506 , n56736 );
not ( n82507 , n56738 );
and ( n82508 , n82507 , n82504 );
and ( n82509 , n41490 , n56738 );
or ( n82510 , n82508 , n82509 );
and ( n82511 , n82506 , n82510 );
and ( n82512 , n41500 , n56736 );
or ( n82513 , n82511 , n82512 );
and ( n82514 , n82513 , n32968 );
or ( n82515 , n82505 , n82514 );
and ( n82516 , n82515 , n33370 );
and ( n82517 , n32791 , n35062 );
or ( n82518 , C0 , n82486 , n82495 , n82516 , n82517 );
buf ( n82519 , n82518 );
buf ( n82520 , n82519 );
buf ( n82521 , n30987 );
buf ( n82522 , n31655 );
not ( n82523 , n41532 );
and ( n82524 , n82523 , n34437 );
and ( n82525 , n69688 , n41532 );
or ( n82526 , n82524 , n82525 );
buf ( n82527 , n82526 );
buf ( n82528 , n82527 );
buf ( n82529 , n31655 );
buf ( n82530 , n30987 );
xor ( n82531 , n54156 , n54981 );
and ( n82532 , n82531 , n33199 );
not ( n82533 , n48648 );
and ( n82534 , n82533 , n54156 );
and ( n82535 , n34441 , n48648 );
or ( n82536 , n82534 , n82535 );
and ( n82537 , n82536 , n32924 );
not ( n82538 , n48660 );
and ( n82539 , n82538 , n54156 );
and ( n82540 , n77664 , n48660 );
or ( n82541 , n82539 , n82540 );
and ( n82542 , n82541 , n33172 );
not ( n82543 , n48730 );
and ( n82544 , n82543 , n54156 );
and ( n82545 , n69721 , n48730 );
or ( n82546 , n82544 , n82545 );
and ( n82547 , n82546 , n33187 );
and ( n82548 , n54156 , n54713 );
or ( n82549 , n82532 , n82537 , n82542 , n82547 , n82548 );
and ( n82550 , n82549 , n33208 );
and ( n82551 , n54156 , n39805 );
or ( n82552 , C0 , n82550 , n82551 );
buf ( n82553 , n82552 );
buf ( n82554 , n82553 );
buf ( n82555 , n30987 );
buf ( n82556 , n31655 );
buf ( n82557 , n30987 );
not ( n82558 , n31437 );
and ( n82559 , n82558 , n49369 );
and ( n82560 , n78193 , n31437 );
or ( n82561 , n82559 , n82560 );
and ( n82562 , n82561 , n31468 );
not ( n82563 , n41837 );
and ( n82564 , n82563 , n49369 );
and ( n82565 , n49389 , n41837 );
or ( n82566 , n82564 , n82565 );
and ( n82567 , n82566 , n31521 );
and ( n82568 , n49369 , n42158 );
or ( n82569 , n82562 , n82567 , n82568 );
and ( n82570 , n82569 , n31557 );
and ( n82571 , n49369 , n40154 );
or ( n82572 , C0 , n82570 , n82571 );
buf ( n82573 , n82572 );
buf ( n82574 , n82573 );
buf ( n82575 , n31655 );
not ( n82576 , n40163 );
and ( n82577 , n82576 , n31781 );
not ( n82578 , n56287 );
and ( n82579 , n82578 , n31781 );
and ( n82580 , n32252 , n56287 );
or ( n82581 , n82579 , n82580 );
and ( n82582 , n82581 , n40163 );
or ( n82583 , n82577 , n82582 );
and ( n82584 , n82583 , n32498 );
not ( n82585 , n56295 );
not ( n82586 , n56287 );
and ( n82587 , n82586 , n31781 );
and ( n82588 , n40393 , n56287 );
or ( n82589 , n82587 , n82588 );
and ( n82590 , n82585 , n82589 );
and ( n82591 , n40393 , n56295 );
or ( n82592 , n82590 , n82591 );
and ( n82593 , n82592 , n32473 );
not ( n82594 , n32475 );
not ( n82595 , n56295 );
not ( n82596 , n56287 );
and ( n82597 , n82596 , n31781 );
and ( n82598 , n40393 , n56287 );
or ( n82599 , n82597 , n82598 );
and ( n82600 , n82595 , n82599 );
and ( n82601 , n40393 , n56295 );
or ( n82602 , n82600 , n82601 );
and ( n82603 , n82594 , n82602 );
not ( n82604 , n56315 );
not ( n82605 , n56317 );
and ( n82606 , n82605 , n82602 );
and ( n82607 , n40972 , n56317 );
or ( n82608 , n82606 , n82607 );
and ( n82609 , n82604 , n82608 );
and ( n82610 , n41267 , n56315 );
or ( n82611 , n82609 , n82610 );
and ( n82612 , n82611 , n32475 );
or ( n82613 , n82603 , n82612 );
and ( n82614 , n82613 , n32486 );
and ( n82615 , n31781 , n41278 );
or ( n82616 , C0 , n82584 , n82593 , n82614 , n82615 );
buf ( n82617 , n82616 );
buf ( n82618 , n82617 );
buf ( n82619 , n30987 );
not ( n82620 , n40163 );
and ( n82621 , n82620 , n32003 );
not ( n82622 , n42171 );
and ( n82623 , n82622 , n32003 );
and ( n82624 , n32147 , n42171 );
or ( n82625 , n82623 , n82624 );
and ( n82626 , n82625 , n40163 );
or ( n82627 , n82621 , n82626 );
and ( n82628 , n82627 , n32498 );
not ( n82629 , n42180 );
not ( n82630 , n42171 );
and ( n82631 , n82630 , n32003 );
and ( n82632 , n49314 , n42171 );
or ( n82633 , n82631 , n82632 );
and ( n82634 , n82629 , n82633 );
and ( n82635 , n49314 , n42180 );
or ( n82636 , n82634 , n82635 );
and ( n82637 , n82636 , n32473 );
not ( n82638 , n32475 );
not ( n82639 , n42180 );
not ( n82640 , n42171 );
and ( n82641 , n82640 , n32003 );
and ( n82642 , n49314 , n42171 );
or ( n82643 , n82641 , n82642 );
and ( n82644 , n82639 , n82643 );
and ( n82645 , n49314 , n42180 );
or ( n82646 , n82644 , n82645 );
and ( n82647 , n82638 , n82646 );
not ( n82648 , n42206 );
not ( n82649 , n42209 );
and ( n82650 , n82649 , n82646 );
and ( n82651 , n49340 , n42209 );
or ( n82652 , n82650 , n82651 );
and ( n82653 , n82648 , n82652 );
and ( n82654 , n49348 , n42206 );
or ( n82655 , n82653 , n82654 );
and ( n82656 , n82655 , n32475 );
or ( n82657 , n82647 , n82656 );
and ( n82658 , n82657 , n32486 );
and ( n82659 , n32003 , n41278 );
or ( n82660 , C0 , n82628 , n82637 , n82658 , n82659 );
buf ( n82661 , n82660 );
buf ( n82662 , n82661 );
buf ( n82663 , n31655 );
not ( n82664 , n31437 );
and ( n82665 , n82664 , n76107 );
not ( n82666 , n41809 );
and ( n82667 , n82666 , n41779 );
xor ( n82668 , n62433 , n62438 );
and ( n82669 , n82668 , n41809 );
or ( n82670 , n82667 , n82669 );
and ( n82671 , n82670 , n31437 );
or ( n82672 , n82665 , n82671 );
and ( n82673 , n82672 , n31468 );
not ( n82674 , n41837 );
and ( n82675 , n82674 , n76107 );
and ( n82676 , n76113 , n41837 );
or ( n82677 , n82675 , n82676 );
and ( n82678 , n82677 , n31521 );
and ( n82679 , n76107 , n42158 );
or ( n82680 , n82673 , n82678 , n82679 );
and ( n82681 , n82680 , n31557 );
and ( n82682 , n76107 , n40154 );
or ( n82683 , C0 , n82681 , n82682 );
buf ( n82684 , n82683 );
buf ( n82685 , n82684 );
buf ( n82686 , n30987 );
and ( n82687 , n31580 , n31007 );
not ( n82688 , n31077 );
and ( n82689 , n82688 , n34004 );
buf ( n82690 , n82689 );
and ( n82691 , n82690 , n31373 );
not ( n82692 , n31402 );
and ( n82693 , n82692 , n34004 );
buf ( n82694 , n82693 );
and ( n82695 , n82694 , n31408 );
not ( n82696 , n31437 );
and ( n82697 , n82696 , n34004 );
not ( n82698 , n31455 );
and ( n82699 , n82698 , n34048 );
xor ( n82700 , n34004 , n34019 );
and ( n82701 , n82700 , n31455 );
or ( n82702 , n82699 , n82701 );
and ( n82703 , n82702 , n31437 );
or ( n82704 , n82697 , n82703 );
and ( n82705 , n82704 , n31468 );
not ( n82706 , n31497 );
and ( n82707 , n82706 , n34004 );
not ( n82708 , n31454 );
not ( n82709 , n31501 );
and ( n82710 , n82709 , n34048 );
xor ( n82711 , n34049 , n34071 );
and ( n82712 , n82711 , n31501 );
or ( n82713 , n82710 , n82712 );
and ( n82714 , n82708 , n82713 );
and ( n82715 , n82700 , n31454 );
or ( n82716 , n82714 , n82715 );
and ( n82717 , n82716 , n31497 );
or ( n82718 , n82707 , n82717 );
and ( n82719 , n82718 , n31521 );
and ( n82720 , n34004 , n31553 );
or ( n82721 , n82691 , n82695 , n82705 , n82719 , n82720 );
and ( n82722 , n82721 , n31557 );
not ( n82723 , n31452 );
not ( n82724 , n31619 );
and ( n82725 , n82724 , n34105 );
xor ( n82726 , n34106 , n34128 );
and ( n82727 , n82726 , n31619 );
or ( n82728 , n82725 , n82727 );
and ( n82729 , n82723 , n82728 );
and ( n82730 , n34004 , n31452 );
or ( n82731 , n82729 , n82730 );
and ( n82732 , n82731 , n31638 );
buf ( n82733 , n33973 );
and ( n82734 , n34004 , n31650 );
or ( n82735 , C0 , n82687 , n82722 , n82732 , n82733 , n82734 );
buf ( n82736 , n82735 );
buf ( n82737 , n82736 );
buf ( n82738 , n31655 );
buf ( n82739 , n31655 );
not ( n82740 , n33419 );
and ( n82741 , n82740 , n31564 );
and ( n82742 , n73469 , n33419 );
or ( n82743 , n82741 , n82742 );
and ( n82744 , n82743 , n31529 );
not ( n82745 , n33734 );
and ( n82746 , n82745 , n31564 );
and ( n82747 , n73480 , n33734 );
or ( n82748 , n82746 , n82747 );
and ( n82749 , n82748 , n31527 );
and ( n82750 , n31564 , n33942 );
or ( n82751 , n82744 , n82749 , n82750 );
and ( n82752 , n82751 , n31557 );
and ( n82753 , n35484 , n31643 );
not ( n82754 , n31452 );
and ( n82755 , n82754 , n35484 );
xor ( n82756 , n31564 , n59436 );
and ( n82757 , n82756 , n31452 );
or ( n82758 , n82755 , n82757 );
and ( n82759 , n82758 , n31638 );
and ( n82760 , n35390 , n33973 );
and ( n82761 , n31564 , n33978 );
or ( n82762 , C0 , n82752 , n82753 , n82759 , n82760 , n82761 );
buf ( n82763 , n82762 );
buf ( n82764 , n82763 );
buf ( n82765 , n30987 );
buf ( n82766 , n31655 );
buf ( n82767 , n31655 );
buf ( n82768 , n30987 );
xor ( n82769 , n39545 , n54977 );
and ( n82770 , n82769 , n33199 );
not ( n82771 , n48648 );
and ( n82772 , n82771 , n39545 );
and ( n82773 , n34367 , n48648 );
or ( n82774 , n82772 , n82773 );
and ( n82775 , n82774 , n32924 );
not ( n82776 , n48660 );
and ( n82777 , n82776 , n39545 );
not ( n82778 , n39584 );
and ( n82779 , n82778 , n42610 );
and ( n82780 , n42678 , n39584 );
or ( n82781 , n82779 , n82780 );
and ( n82782 , n82781 , n48660 );
or ( n82783 , n82777 , n82782 );
and ( n82784 , n82783 , n33172 );
not ( n82785 , n48730 );
and ( n82786 , n82785 , n39545 );
and ( n82787 , n32824 , n52252 );
and ( n82788 , n32826 , n52254 );
and ( n82789 , n32828 , n52256 );
and ( n82790 , n32830 , n52258 );
and ( n82791 , n32832 , n52260 );
and ( n82792 , n32834 , n52262 );
and ( n82793 , n32836 , n52264 );
and ( n82794 , n32838 , n52266 );
and ( n82795 , n32840 , n52268 );
and ( n82796 , n32842 , n52270 );
and ( n82797 , n32844 , n52272 );
and ( n82798 , n32846 , n52274 );
and ( n82799 , n32848 , n52276 );
and ( n82800 , n32850 , n52278 );
and ( n82801 , n32852 , n52280 );
and ( n82802 , n32854 , n52282 );
or ( n82803 , n82787 , n82788 , n82789 , n82790 , n82791 , n82792 , n82793 , n82794 , n82795 , n82796 , n82797 , n82798 , n82799 , n82800 , n82801 , n82802 );
and ( n82804 , n82803 , n48730 );
or ( n82805 , n82786 , n82804 );
and ( n82806 , n82805 , n33187 );
and ( n82807 , n39545 , n54713 );
or ( n82808 , n82770 , n82775 , n82784 , n82806 , n82807 );
and ( n82809 , n82808 , n33208 );
and ( n82810 , n39545 , n39805 );
or ( n82811 , C0 , n82809 , n82810 );
buf ( n82812 , n82811 );
buf ( n82813 , n82812 );
not ( n82814 , n41532 );
and ( n82815 , n82814 , n34429 );
and ( n82816 , n74778 , n41532 );
or ( n82817 , n82815 , n82816 );
buf ( n82818 , n82817 );
buf ( n82819 , n82818 );
buf ( n82820 , n30987 );
not ( n82821 , n46356 );
and ( n82822 , n82821 , n31366 );
not ( n82823 , n47423 );
and ( n82824 , n82823 , n31366 );
and ( n82825 , n31372 , n47423 );
or ( n82826 , n82824 , n82825 );
and ( n82827 , n82826 , n46356 );
or ( n82828 , n82822 , n82827 );
and ( n82829 , n82828 , n31649 );
not ( n82830 , n47431 );
not ( n82831 , n47423 );
and ( n82832 , n82831 , n31366 );
and ( n82833 , n47849 , n47423 );
or ( n82834 , n82832 , n82833 );
and ( n82835 , n82830 , n82834 );
and ( n82836 , n47849 , n47431 );
or ( n82837 , n82835 , n82836 );
and ( n82838 , n82837 , n31643 );
not ( n82839 , n31452 );
not ( n82840 , n47431 );
not ( n82841 , n47423 );
and ( n82842 , n82841 , n31366 );
and ( n82843 , n47849 , n47423 );
or ( n82844 , n82842 , n82843 );
and ( n82845 , n82840 , n82844 );
and ( n82846 , n47849 , n47431 );
or ( n82847 , n82845 , n82846 );
and ( n82848 , n82839 , n82847 );
not ( n82849 , n47466 );
not ( n82850 , n47468 );
and ( n82851 , n82850 , n82847 );
and ( n82852 , n47877 , n47468 );
or ( n82853 , n82851 , n82852 );
and ( n82854 , n82849 , n82853 );
and ( n82855 , n47887 , n47466 );
or ( n82856 , n82854 , n82855 );
and ( n82857 , n82856 , n31452 );
or ( n82858 , n82848 , n82857 );
and ( n82859 , n82858 , n31638 );
and ( n82860 , n31366 , n47277 );
or ( n82861 , C0 , n82829 , n82838 , n82859 , n82860 );
buf ( n82862 , n82861 );
buf ( n82863 , n82862 );
buf ( n82864 , n31655 );
buf ( n82865 , n31655 );
buf ( n82866 , n30987 );
xor ( n82867 , n47284 , n47298 );
and ( n82868 , n82867 , n32433 );
not ( n82869 , n47331 );
and ( n82870 , n82869 , n47284 );
and ( n82871 , n61496 , n47331 );
or ( n82872 , n82870 , n82871 );
and ( n82873 , n82872 , n32413 );
and ( n82874 , n47284 , n47402 );
or ( n82875 , n82868 , n82873 , n82874 );
and ( n82876 , n82875 , n32456 );
and ( n82877 , n47284 , n47409 );
or ( n82878 , C0 , n82876 , n82877 );
buf ( n82879 , n82878 );
buf ( n82880 , n82879 );
not ( n82881 , n35542 );
and ( n82882 , n82881 , n41851 );
and ( n82883 , n50531 , n35542 );
or ( n82884 , n82882 , n82883 );
buf ( n82885 , n82884 );
buf ( n82886 , n82885 );
not ( n82887 , n40163 );
and ( n82888 , n82887 , n31805 );
not ( n82889 , n55888 );
and ( n82890 , n82889 , n31805 );
and ( n82891 , n32252 , n55888 );
or ( n82892 , n82890 , n82891 );
and ( n82893 , n82892 , n40163 );
or ( n82894 , n82888 , n82893 );
and ( n82895 , n82894 , n32498 );
not ( n82896 , n55896 );
not ( n82897 , n55888 );
and ( n82898 , n82897 , n31805 );
and ( n82899 , n40393 , n55888 );
or ( n82900 , n82898 , n82899 );
and ( n82901 , n82896 , n82900 );
and ( n82902 , n40393 , n55896 );
or ( n82903 , n82901 , n82902 );
and ( n82904 , n82903 , n32473 );
not ( n82905 , n32475 );
not ( n82906 , n55896 );
not ( n82907 , n55888 );
and ( n82908 , n82907 , n31805 );
and ( n82909 , n40393 , n55888 );
or ( n82910 , n82908 , n82909 );
and ( n82911 , n82906 , n82910 );
and ( n82912 , n40393 , n55896 );
or ( n82913 , n82911 , n82912 );
and ( n82914 , n82905 , n82913 );
not ( n82915 , n55916 );
not ( n82916 , n55918 );
and ( n82917 , n82916 , n82913 );
and ( n82918 , n40972 , n55918 );
or ( n82919 , n82917 , n82918 );
and ( n82920 , n82915 , n82919 );
and ( n82921 , n41267 , n55916 );
or ( n82922 , n82920 , n82921 );
and ( n82923 , n82922 , n32475 );
or ( n82924 , n82914 , n82923 );
and ( n82925 , n82924 , n32486 );
and ( n82926 , n31805 , n41278 );
or ( n82927 , C0 , n82895 , n82904 , n82925 , n82926 );
buf ( n82928 , n82927 );
buf ( n82929 , n82928 );
xor ( n82930 , n44775 , n44792 );
and ( n82931 , n82930 , n31548 );
not ( n82932 , n44807 );
and ( n82933 , n82932 , n44775 );
and ( n82934 , n46672 , n44807 );
or ( n82935 , n82933 , n82934 );
and ( n82936 , n82935 , n31408 );
not ( n82937 , n44817 );
and ( n82938 , n82937 , n44775 );
not ( n82939 , n44994 );
and ( n82940 , n82939 , n44834 );
xor ( n82941 , n45009 , n45011 );
and ( n82942 , n82941 , n44994 );
or ( n82943 , n82940 , n82942 );
and ( n82944 , n82943 , n44817 );
or ( n82945 , n82938 , n82944 );
and ( n82946 , n82945 , n31521 );
not ( n82947 , n45059 );
and ( n82948 , n82947 , n44775 );
and ( n82949 , n76724 , n45059 );
or ( n82950 , n82948 , n82949 );
and ( n82951 , n82950 , n31536 );
and ( n82952 , n44775 , n45148 );
or ( n82953 , n82931 , n82936 , n82946 , n82951 , n82952 );
and ( n82954 , n82953 , n31557 );
and ( n82955 , n44775 , n40154 );
or ( n82956 , C0 , n82954 , n82955 );
buf ( n82957 , n82956 );
buf ( n82958 , n82957 );
buf ( n82959 , n30987 );
buf ( n82960 , n31655 );
buf ( n82961 , n30987 );
buf ( n82962 , n31655 );
buf ( n82963 , n30987 );
not ( n82964 , n46356 );
and ( n82965 , n82964 , n31307 );
not ( n82966 , n63024 );
and ( n82967 , n82966 , n31307 );
and ( n82968 , n31339 , n63024 );
or ( n82969 , n82967 , n82968 );
and ( n82970 , n82969 , n46356 );
or ( n82971 , n82965 , n82970 );
and ( n82972 , n82971 , n31649 );
not ( n82973 , n63032 );
not ( n82974 , n63024 );
and ( n82975 , n82974 , n31307 );
and ( n82976 , n47449 , n63024 );
or ( n82977 , n82975 , n82976 );
and ( n82978 , n82973 , n82977 );
and ( n82979 , n47449 , n63032 );
or ( n82980 , n82978 , n82979 );
and ( n82981 , n82980 , n31643 );
not ( n82982 , n31452 );
not ( n82983 , n63032 );
not ( n82984 , n63024 );
and ( n82985 , n82984 , n31307 );
and ( n82986 , n47449 , n63024 );
or ( n82987 , n82985 , n82986 );
and ( n82988 , n82983 , n82987 );
and ( n82989 , n47449 , n63032 );
or ( n82990 , n82988 , n82989 );
and ( n82991 , n82982 , n82990 );
not ( n82992 , n63052 );
not ( n82993 , n63054 );
and ( n82994 , n82993 , n82990 );
and ( n82995 , n47485 , n63054 );
or ( n82996 , n82994 , n82995 );
and ( n82997 , n82992 , n82996 );
and ( n82998 , n47503 , n63052 );
or ( n82999 , n82997 , n82998 );
and ( n83000 , n82999 , n31452 );
or ( n83001 , n82991 , n83000 );
and ( n83002 , n83001 , n31638 );
and ( n83003 , n31307 , n47277 );
or ( n83004 , C0 , n82972 , n82981 , n83002 , n83003 );
buf ( n83005 , n83004 );
buf ( n83006 , n83005 );
not ( n83007 , n35278 );
and ( n83008 , n83007 , n78531 );
and ( n83009 , n78905 , n35278 );
or ( n83010 , n83008 , n83009 );
and ( n83011 , n83010 , n32417 );
not ( n83012 , n47912 );
and ( n83013 , n83012 , n78531 );
and ( n83014 , n78537 , n47912 );
or ( n83015 , n83013 , n83014 );
and ( n83016 , n83015 , n32415 );
and ( n83017 , n78531 , n48133 );
or ( n83018 , n83011 , n83016 , n83017 );
and ( n83019 , n83018 , n32456 );
and ( n83020 , n78531 , n47409 );
or ( n83021 , C0 , n83019 , n83020 );
buf ( n83022 , n83021 );
buf ( n83023 , n83022 );
buf ( n83024 , n31655 );
xor ( n83025 , n49567 , n60322 );
and ( n83026 , n83025 , n32433 );
not ( n83027 , n47331 );
and ( n83028 , n83027 , n49567 );
xor ( n83029 , n60416 , n60546 );
and ( n83030 , n83029 , n47331 );
or ( n83031 , n83028 , n83030 );
and ( n83032 , n83031 , n32413 );
and ( n83033 , n49567 , n47402 );
or ( n83034 , n83026 , n83032 , n83033 );
and ( n83035 , n83034 , n32456 );
and ( n83036 , n49567 , n47409 );
or ( n83037 , C0 , n83035 , n83036 );
buf ( n83038 , n83037 );
buf ( n83039 , n83038 );
buf ( n83040 , n30987 );
not ( n83041 , n46356 );
and ( n83042 , n83041 , n31304 );
not ( n83043 , n60564 );
and ( n83044 , n83043 , n31304 );
and ( n83045 , n31306 , n60564 );
or ( n83046 , n83044 , n83045 );
and ( n83047 , n83046 , n46356 );
or ( n83048 , n83042 , n83047 );
and ( n83049 , n83048 , n31649 );
not ( n83050 , n60572 );
not ( n83051 , n60564 );
and ( n83052 , n83051 , n31304 );
and ( n83053 , n58061 , n60564 );
or ( n83054 , n83052 , n83053 );
and ( n83055 , n83050 , n83054 );
and ( n83056 , n58061 , n60572 );
or ( n83057 , n83055 , n83056 );
and ( n83058 , n83057 , n31643 );
not ( n83059 , n31452 );
not ( n83060 , n60572 );
not ( n83061 , n60564 );
and ( n83062 , n83061 , n31304 );
and ( n83063 , n58061 , n60564 );
or ( n83064 , n83062 , n83063 );
and ( n83065 , n83060 , n83064 );
and ( n83066 , n58061 , n60572 );
or ( n83067 , n83065 , n83066 );
and ( n83068 , n83059 , n83067 );
not ( n83069 , n60592 );
not ( n83070 , n60594 );
and ( n83071 , n83070 , n83067 );
and ( n83072 , n58085 , n60594 );
or ( n83073 , n83071 , n83072 );
and ( n83074 , n83069 , n83073 );
and ( n83075 , n58093 , n60592 );
or ( n83076 , n83074 , n83075 );
and ( n83077 , n83076 , n31452 );
or ( n83078 , n83068 , n83077 );
and ( n83079 , n83078 , n31638 );
and ( n83080 , n31304 , n47277 );
or ( n83081 , C0 , n83049 , n83058 , n83079 , n83080 );
buf ( n83082 , n83081 );
buf ( n83083 , n83082 );
buf ( n83084 , n30987 );
buf ( n83085 , n31655 );
buf ( n83086 , RI15b46ef0_285);
buf ( n83087 , n83086 );
buf ( n83088 , n30987 );
and ( n83089 , n50951 , n77569 );
xor ( n83090 , n50949 , n83089 );
and ( n83091 , n83090 , n32431 );
not ( n83092 , n50002 );
and ( n83093 , n83092 , n50949 );
and ( n83094 , n40564 , n50002 );
or ( n83095 , n83093 , n83094 );
and ( n83096 , n83095 , n32419 );
not ( n83097 , n50008 );
and ( n83098 , n83097 , n50949 );
and ( n83099 , n59240 , n50008 );
or ( n83100 , n83098 , n83099 );
and ( n83101 , n83100 , n32415 );
not ( n83102 , n50067 );
and ( n83103 , n83102 , n50949 );
and ( n83104 , n60399 , n77589 );
xor ( n83105 , n60382 , n83104 );
and ( n83106 , n83105 , n50067 );
or ( n83107 , n83103 , n83106 );
and ( n83108 , n83107 , n32411 );
and ( n83109 , n50949 , n50098 );
or ( n83110 , n83091 , n83096 , n83101 , n83108 , n83109 );
and ( n83111 , n83110 , n32456 );
and ( n83112 , n50949 , n47409 );
or ( n83113 , C0 , n83111 , n83112 );
buf ( n83114 , n83113 );
buf ( n83115 , n83114 );
buf ( n83116 , n31655 );
not ( n83117 , n46356 );
and ( n83118 , n83117 , n31228 );
not ( n83119 , n56904 );
and ( n83120 , n83119 , n31228 );
and ( n83121 , n31238 , n56904 );
or ( n83122 , n83120 , n83121 );
and ( n83123 , n83122 , n46356 );
or ( n83124 , n83118 , n83123 );
and ( n83125 , n83124 , n31649 );
not ( n83126 , n56912 );
not ( n83127 , n56904 );
and ( n83128 , n83127 , n31228 );
and ( n83129 , n49901 , n56904 );
or ( n83130 , n83128 , n83129 );
and ( n83131 , n83126 , n83130 );
and ( n83132 , n49901 , n56912 );
or ( n83133 , n83131 , n83132 );
and ( n83134 , n83133 , n31643 );
not ( n83135 , n31452 );
not ( n83136 , n56912 );
not ( n83137 , n56904 );
and ( n83138 , n83137 , n31228 );
and ( n83139 , n49901 , n56904 );
or ( n83140 , n83138 , n83139 );
and ( n83141 , n83136 , n83140 );
and ( n83142 , n49901 , n56912 );
or ( n83143 , n83141 , n83142 );
and ( n83144 , n83135 , n83143 );
not ( n83145 , n56937 );
not ( n83146 , n56939 );
and ( n83147 , n83146 , n83143 );
and ( n83148 , n49925 , n56939 );
or ( n83149 , n83147 , n83148 );
and ( n83150 , n83145 , n83149 );
and ( n83151 , n49933 , n56937 );
or ( n83152 , n83150 , n83151 );
and ( n83153 , n83152 , n31452 );
or ( n83154 , n83144 , n83153 );
and ( n83155 , n83154 , n31638 );
and ( n83156 , n31228 , n47277 );
or ( n83157 , C0 , n83125 , n83134 , n83155 , n83156 );
buf ( n83158 , n83157 );
buf ( n83159 , n83158 );
buf ( n83160 , n31655 );
not ( n83161 , n43755 );
and ( n83162 , n83161 , n43700 );
xor ( n83163 , n52301 , n52328 );
and ( n83164 , n83163 , n43755 );
or ( n83165 , n83162 , n83164 );
and ( n83166 , n83165 , n43774 );
not ( n83167 , n44663 );
and ( n83168 , n83167 , n44612 );
xor ( n83169 , n52339 , n52366 );
and ( n83170 , n83169 , n44663 );
or ( n83171 , n83168 , n83170 );
and ( n83172 , n83171 , n44682 );
buf ( n83173 , RI15b45ca8_246);
and ( n83174 , n83173 , n44695 );
or ( n83175 , n83166 , n83172 , n83174 );
buf ( n83176 , n83175 );
buf ( n83177 , n83176 );
buf ( n83178 , n30987 );
buf ( n83179 , n31655 );
buf ( n83180 , n31655 );
buf ( n83181 , n30987 );
buf ( n83182 , n30987 );
not ( n83183 , n32953 );
and ( n83184 , n83183 , n54075 );
and ( n83185 , n54589 , n32953 );
or ( n83186 , n83184 , n83185 );
and ( n83187 , n83186 , n33038 );
not ( n83188 , n48660 );
and ( n83189 , n83188 , n54075 );
not ( n83190 , n55168 );
and ( n83191 , n83190 , n55008 );
xor ( n83192 , n55175 , n55177 );
and ( n83193 , n83192 , n55168 );
or ( n83194 , n83191 , n83193 );
and ( n83195 , n83194 , n48660 );
or ( n83196 , n83189 , n83195 );
and ( n83197 , n83196 , n33172 );
and ( n83198 , n54075 , n39795 );
or ( n83199 , n83187 , n83197 , n83198 );
and ( n83200 , n83199 , n33208 );
and ( n83201 , n54075 , n39805 );
or ( n83202 , C0 , n83200 , n83201 );
buf ( n83203 , n83202 );
buf ( n83204 , n83203 );
buf ( n83205 , n30987 );
buf ( n83206 , n31655 );
buf ( n83207 , n31655 );
and ( n83208 , n59253 , n32494 );
not ( n83209 , n46083 );
and ( n83210 , n83209 , n56401 );
buf ( n83211 , n83210 );
and ( n83212 , n83211 , n32421 );
not ( n83213 , n46326 );
and ( n83214 , n83213 , n56401 );
and ( n83215 , n59259 , n46326 );
or ( n83216 , n83214 , n83215 );
and ( n83217 , n83216 , n32417 );
and ( n83218 , n56401 , n46340 );
or ( n83219 , n83212 , n83217 , n83218 );
and ( n83220 , n83219 , n32456 );
and ( n83221 , n56401 , n46349 );
or ( n83222 , C0 , n83208 , n83220 , n83221 );
buf ( n83223 , n83222 );
buf ( n83224 , n83223 );
buf ( n83225 , n31655 );
not ( n83226 , n46356 );
and ( n83227 , n83226 , n31350 );
not ( n83228 , n53353 );
and ( n83229 , n83228 , n31350 );
and ( n83230 , n31372 , n53353 );
or ( n83231 , n83229 , n83230 );
and ( n83232 , n83231 , n46356 );
or ( n83233 , n83227 , n83232 );
and ( n83234 , n83233 , n31649 );
not ( n83235 , n53361 );
not ( n83236 , n53353 );
and ( n83237 , n83236 , n31350 );
and ( n83238 , n47849 , n53353 );
or ( n83239 , n83237 , n83238 );
and ( n83240 , n83235 , n83239 );
and ( n83241 , n47849 , n53361 );
or ( n83242 , n83240 , n83241 );
and ( n83243 , n83242 , n31643 );
not ( n83244 , n31452 );
not ( n83245 , n53361 );
not ( n83246 , n53353 );
and ( n83247 , n83246 , n31350 );
and ( n83248 , n47849 , n53353 );
or ( n83249 , n83247 , n83248 );
and ( n83250 , n83245 , n83249 );
and ( n83251 , n47849 , n53361 );
or ( n83252 , n83250 , n83251 );
and ( n83253 , n83244 , n83252 );
not ( n83254 , n53381 );
not ( n83255 , n53383 );
and ( n83256 , n83255 , n83252 );
and ( n83257 , n47877 , n53383 );
or ( n83258 , n83256 , n83257 );
and ( n83259 , n83254 , n83258 );
and ( n83260 , n47887 , n53381 );
or ( n83261 , n83259 , n83260 );
and ( n83262 , n83261 , n31452 );
or ( n83263 , n83253 , n83262 );
and ( n83264 , n83263 , n31638 );
and ( n83265 , n31350 , n47277 );
or ( n83266 , C0 , n83234 , n83243 , n83264 , n83265 );
buf ( n83267 , n83266 );
buf ( n83268 , n83267 );
buf ( n83269 , n30987 );
buf ( n83270 , n31655 );
not ( n83271 , n31437 );
and ( n83272 , n83271 , n52176 );
not ( n83273 , n41809 );
and ( n83274 , n83273 , n41610 );
xor ( n83275 , n41820 , n41611 );
and ( n83276 , n83275 , n41809 );
or ( n83277 , n83274 , n83276 );
and ( n83278 , n83277 , n31437 );
or ( n83279 , n83272 , n83278 );
and ( n83280 , n83279 , n31468 );
not ( n83281 , n41837 );
and ( n83282 , n83281 , n52176 );
and ( n83283 , n52182 , n41837 );
or ( n83284 , n83282 , n83283 );
and ( n83285 , n83284 , n31521 );
and ( n83286 , n52176 , n42158 );
or ( n83287 , n83280 , n83285 , n83286 );
and ( n83288 , n83287 , n31557 );
and ( n83289 , n52176 , n40154 );
or ( n83290 , C0 , n83288 , n83289 );
buf ( n83291 , n83290 );
buf ( n83292 , n83291 );
not ( n83293 , n40163 );
and ( n83294 , n83293 , n31826 );
not ( n83295 , n56988 );
and ( n83296 , n83295 , n31826 );
and ( n83297 , n32235 , n56988 );
or ( n83298 , n83296 , n83297 );
and ( n83299 , n83298 , n40163 );
or ( n83300 , n83294 , n83299 );
and ( n83301 , n83300 , n32498 );
not ( n83302 , n56996 );
not ( n83303 , n56988 );
and ( n83304 , n83303 , n31826 );
and ( n83305 , n42188 , n56988 );
or ( n83306 , n83304 , n83305 );
and ( n83307 , n83302 , n83306 );
and ( n83308 , n42188 , n56996 );
or ( n83309 , n83307 , n83308 );
and ( n83310 , n83309 , n32473 );
not ( n83311 , n32475 );
not ( n83312 , n56996 );
not ( n83313 , n56988 );
and ( n83314 , n83313 , n31826 );
and ( n83315 , n42188 , n56988 );
or ( n83316 , n83314 , n83315 );
and ( n83317 , n83312 , n83316 );
and ( n83318 , n42188 , n56996 );
or ( n83319 , n83317 , n83318 );
and ( n83320 , n83311 , n83319 );
not ( n83321 , n57016 );
not ( n83322 , n57018 );
and ( n83323 , n83322 , n83319 );
and ( n83324 , n42216 , n57018 );
or ( n83325 , n83323 , n83324 );
and ( n83326 , n83321 , n83325 );
and ( n83327 , n42224 , n57016 );
or ( n83328 , n83326 , n83327 );
and ( n83329 , n83328 , n32475 );
or ( n83330 , n83320 , n83329 );
and ( n83331 , n83330 , n32486 );
and ( n83332 , n31826 , n41278 );
or ( n83333 , C0 , n83301 , n83310 , n83331 , n83332 );
buf ( n83334 , n83333 );
buf ( n83335 , n83334 );
buf ( n83336 , n31655 );
buf ( n83337 , n30987 );
buf ( n83338 , n30987 );
buf ( n83339 , n30987 );
buf ( n83340 , n31655 );
buf ( n83341 , n31655 );
not ( n83342 , n34150 );
and ( n83343 , n83342 , n32765 );
not ( n83344 , n59105 );
and ( n83345 , n83344 , n32765 );
and ( n83346 , n32789 , n59105 );
or ( n83347 , n83345 , n83346 );
and ( n83348 , n83347 , n34150 );
or ( n83349 , n83343 , n83348 );
and ( n83350 , n83349 , n33381 );
not ( n83351 , n59113 );
not ( n83352 , n59105 );
and ( n83353 , n83352 , n32765 );
and ( n83354 , n34301 , n59105 );
or ( n83355 , n83353 , n83354 );
and ( n83356 , n83351 , n83355 );
and ( n83357 , n34301 , n59113 );
or ( n83358 , n83356 , n83357 );
and ( n83359 , n83358 , n33375 );
not ( n83360 , n32968 );
not ( n83361 , n59113 );
not ( n83362 , n59105 );
and ( n83363 , n83362 , n32765 );
and ( n83364 , n34301 , n59105 );
or ( n83365 , n83363 , n83364 );
and ( n83366 , n83361 , n83365 );
and ( n83367 , n34301 , n59113 );
or ( n83368 , n83366 , n83367 );
and ( n83369 , n83360 , n83368 );
not ( n83370 , n59133 );
not ( n83371 , n59135 );
and ( n83372 , n83371 , n83368 );
and ( n83373 , n34761 , n59135 );
or ( n83374 , n83372 , n83373 );
and ( n83375 , n83370 , n83374 );
and ( n83376 , n35050 , n59133 );
or ( n83377 , n83375 , n83376 );
and ( n83378 , n83377 , n32968 );
or ( n83379 , n83369 , n83378 );
and ( n83380 , n83379 , n33370 );
and ( n83381 , n32765 , n35062 );
or ( n83382 , C0 , n83350 , n83359 , n83380 , n83381 );
buf ( n83383 , n83382 );
buf ( n83384 , n83383 );
buf ( n83385 , n31655 );
buf ( n83386 , n31655 );
not ( n83387 , n43755 );
and ( n83388 , n83387 , n43445 );
xor ( n83389 , n50498 , n50507 );
and ( n83390 , n83389 , n43755 );
or ( n83391 , n83388 , n83390 );
and ( n83392 , n83391 , n43774 );
not ( n83393 , n44663 );
and ( n83394 , n83393 , n44357 );
xor ( n83395 , n50516 , n50525 );
and ( n83396 , n83395 , n44663 );
or ( n83397 , n83394 , n83396 );
and ( n83398 , n83397 , n44682 );
and ( n83399 , n75085 , n44695 );
or ( n83400 , n83392 , n83398 , n83399 );
buf ( n83401 , n83400 );
buf ( n83402 , n83401 );
buf ( n83403 , n30987 );
buf ( n83404 , n30987 );
buf ( n83405 , n30987 );
buf ( n83406 , n30987 );
buf ( n83407 , n31655 );
not ( n83408 , n34150 );
and ( n83409 , n83408 , n32832 );
not ( n83410 , n59105 );
and ( n83411 , n83410 , n32832 );
and ( n83412 , n32856 , n59105 );
or ( n83413 , n83411 , n83412 );
and ( n83414 , n83413 , n34150 );
or ( n83415 , n83409 , n83414 );
and ( n83416 , n83415 , n33381 );
not ( n83417 , n59113 );
not ( n83418 , n59105 );
and ( n83419 , n83418 , n32832 );
and ( n83420 , n48160 , n59105 );
or ( n83421 , n83419 , n83420 );
and ( n83422 , n83417 , n83421 );
and ( n83423 , n48160 , n59113 );
or ( n83424 , n83422 , n83423 );
and ( n83425 , n83424 , n33375 );
not ( n83426 , n32968 );
not ( n83427 , n59113 );
not ( n83428 , n59105 );
and ( n83429 , n83428 , n32832 );
and ( n83430 , n48160 , n59105 );
or ( n83431 , n83429 , n83430 );
and ( n83432 , n83427 , n83431 );
and ( n83433 , n48160 , n59113 );
or ( n83434 , n83432 , n83433 );
and ( n83435 , n83426 , n83434 );
not ( n83436 , n59133 );
not ( n83437 , n59135 );
and ( n83438 , n83437 , n83434 );
and ( n83439 , n48186 , n59135 );
or ( n83440 , n83438 , n83439 );
and ( n83441 , n83436 , n83440 );
and ( n83442 , n48196 , n59133 );
or ( n83443 , n83441 , n83442 );
and ( n83444 , n83443 , n32968 );
or ( n83445 , n83435 , n83444 );
and ( n83446 , n83445 , n33370 );
and ( n83447 , n32832 , n35062 );
or ( n83448 , C0 , n83416 , n83425 , n83446 , n83447 );
buf ( n83449 , n83448 );
buf ( n83450 , n83449 );
buf ( n83451 , n31655 );
buf ( n83452 , n31655 );
buf ( n83453 , n30987 );
and ( n83454 , n49089 , n48639 );
not ( n83455 , n48642 );
and ( n83456 , n83455 , n48609 );
and ( n83457 , n49089 , n48642 );
or ( n83458 , n83456 , n83457 );
and ( n83459 , n83458 , n32890 );
not ( n83460 , n48648 );
and ( n83461 , n83460 , n48609 );
and ( n83462 , n49089 , n48648 );
or ( n83463 , n83461 , n83462 );
and ( n83464 , n83463 , n32924 );
not ( n83465 , n48654 );
and ( n83466 , n83465 , n48609 );
and ( n83467 , n49089 , n48654 );
or ( n83468 , n83466 , n83467 );
and ( n83469 , n83468 , n33038 );
not ( n83470 , n48660 );
and ( n83471 , n83470 , n48609 );
and ( n83472 , n49089 , n48660 );
or ( n83473 , n83471 , n83472 );
and ( n83474 , n83473 , n33172 );
not ( n83475 , n41576 );
and ( n83476 , n83475 , n48609 );
and ( n83477 , n48923 , n41576 );
or ( n83478 , n83476 , n83477 );
and ( n83479 , n83478 , n33189 );
not ( n83480 , n48730 );
and ( n83481 , n83480 , n48609 );
and ( n83482 , n48923 , n48730 );
or ( n83483 , n83481 , n83482 );
and ( n83484 , n83483 , n33187 );
not ( n83485 , n48765 );
and ( n83486 , n83485 , n48609 );
and ( n83487 , n50780 , n48765 );
or ( n83488 , n83486 , n83487 );
and ( n83489 , n83488 , n33180 );
not ( n83490 , n49054 );
and ( n83491 , n83490 , n48609 );
and ( n83492 , n50793 , n49054 );
or ( n83493 , n83491 , n83492 );
and ( n83494 , n83493 , n33178 );
and ( n83495 , n49208 , n49275 );
or ( n83496 , n83454 , n83459 , n83464 , n83469 , n83474 , n83479 , n83484 , n83489 , n83494 , n83495 );
and ( n83497 , n83496 , n33208 );
and ( n83498 , n33002 , n35056 );
and ( n83499 , n48609 , n49286 );
or ( n83500 , C0 , n83497 , n83498 , n83499 );
buf ( n83501 , n83500 );
buf ( n83502 , n83501 );
buf ( n83503 , n30987 );
buf ( n83504 , n31655 );
not ( n83505 , n41532 );
and ( n83506 , n83505 , n34369 );
buf ( n83507 , RI15b53970_717);
and ( n83508 , n83507 , n41532 );
or ( n83509 , n83506 , n83508 );
buf ( n83510 , n83509 );
buf ( n83511 , n83510 );
buf ( n83512 , n31655 );
buf ( n83513 , n30987 );
xor ( n83514 , n54142 , n78382 );
and ( n83515 , n83514 , n33199 );
not ( n83516 , n48648 );
and ( n83517 , n83516 , n54142 );
and ( n83518 , n34427 , n48648 );
or ( n83519 , n83517 , n83518 );
and ( n83520 , n83519 , n32924 );
not ( n83521 , n48660 );
and ( n83522 , n83521 , n54142 );
and ( n83523 , n65095 , n48660 );
or ( n83524 , n83522 , n83523 );
and ( n83525 , n83524 , n33172 );
not ( n83526 , n48730 );
and ( n83527 , n83526 , n54142 );
xor ( n83528 , n58540 , n78401 );
and ( n83529 , n83528 , n48730 );
or ( n83530 , n83527 , n83529 );
and ( n83531 , n83530 , n33187 );
and ( n83532 , n54142 , n54713 );
or ( n83533 , n83515 , n83520 , n83525 , n83531 , n83532 );
and ( n83534 , n83533 , n33208 );
and ( n83535 , n54142 , n39805 );
or ( n83536 , C0 , n83534 , n83535 );
buf ( n83537 , n83536 );
buf ( n83538 , n83537 );
buf ( n83539 , n30987 );
buf ( n83540 , n31655 );
buf ( n83541 , n31655 );
not ( n83542 , n46356 );
and ( n83543 , n83542 , n31323 );
not ( n83544 , n55263 );
and ( n83545 , n83544 , n31323 );
and ( n83546 , n31339 , n55263 );
or ( n83547 , n83545 , n83546 );
and ( n83548 , n83547 , n46356 );
or ( n83549 , n83543 , n83548 );
and ( n83550 , n83549 , n31649 );
not ( n83551 , n55271 );
not ( n83552 , n55263 );
and ( n83553 , n83552 , n31323 );
and ( n83554 , n47449 , n55263 );
or ( n83555 , n83553 , n83554 );
and ( n83556 , n83551 , n83555 );
and ( n83557 , n47449 , n55271 );
or ( n83558 , n83556 , n83557 );
and ( n83559 , n83558 , n31643 );
not ( n83560 , n31452 );
not ( n83561 , n55271 );
not ( n83562 , n55263 );
and ( n83563 , n83562 , n31323 );
and ( n83564 , n47449 , n55263 );
or ( n83565 , n83563 , n83564 );
and ( n83566 , n83561 , n83565 );
and ( n83567 , n47449 , n55271 );
or ( n83568 , n83566 , n83567 );
and ( n83569 , n83560 , n83568 );
not ( n83570 , n55291 );
not ( n83571 , n55293 );
and ( n83572 , n83571 , n83568 );
and ( n83573 , n47485 , n55293 );
or ( n83574 , n83572 , n83573 );
and ( n83575 , n83570 , n83574 );
and ( n83576 , n47503 , n55291 );
or ( n83577 , n83575 , n83576 );
and ( n83578 , n83577 , n31452 );
or ( n83579 , n83569 , n83578 );
and ( n83580 , n83579 , n31638 );
and ( n83581 , n31323 , n47277 );
or ( n83582 , C0 , n83550 , n83559 , n83580 , n83581 );
buf ( n83583 , n83582 );
buf ( n83584 , n83583 );
xor ( n83585 , n46107 , n49987 );
and ( n83586 , n83585 , n32431 );
not ( n83587 , n50002 );
and ( n83588 , n83587 , n46107 );
and ( n83589 , n40269 , n50002 );
or ( n83590 , n83588 , n83589 );
and ( n83591 , n83590 , n32419 );
not ( n83592 , n50008 );
and ( n83593 , n83592 , n46107 );
not ( n83594 , n47910 );
and ( n83595 , n83594 , n63070 );
and ( n83596 , n63086 , n47910 );
or ( n83597 , n83595 , n83596 );
and ( n83598 , n83597 , n50008 );
or ( n83599 , n83593 , n83598 );
and ( n83600 , n83599 , n32415 );
not ( n83601 , n50067 );
and ( n83602 , n83601 , n46107 );
and ( n83603 , n31998 , n50067 );
or ( n83604 , n83602 , n83603 );
and ( n83605 , n83604 , n32411 );
and ( n83606 , n46107 , n50098 );
or ( n83607 , n83586 , n83591 , n83600 , n83605 , n83606 );
and ( n83608 , n83607 , n32456 );
and ( n83609 , n46107 , n47409 );
or ( n83610 , C0 , n83608 , n83609 );
buf ( n83611 , n83610 );
buf ( n83612 , n83611 );
buf ( n83613 , n30987 );
buf ( n83614 , n31655 );
buf ( n83615 , n55526 );
buf ( n83616 , n31655 );
not ( n83617 , n40163 );
and ( n83618 , n83617 , n31994 );
not ( n83619 , n75905 );
and ( n83620 , n83619 , n31994 );
and ( n83621 , n32165 , n75905 );
or ( n83622 , n83620 , n83621 );
and ( n83623 , n83622 , n40163 );
or ( n83624 , n83618 , n83623 );
and ( n83625 , n83624 , n32498 );
not ( n83626 , n75913 );
not ( n83627 , n75905 );
and ( n83628 , n83627 , n31994 );
and ( n83629 , n59005 , n75905 );
or ( n83630 , n83628 , n83629 );
and ( n83631 , n83626 , n83630 );
and ( n83632 , n59005 , n75913 );
or ( n83633 , n83631 , n83632 );
and ( n83634 , n83633 , n32473 );
not ( n83635 , n32475 );
not ( n83636 , n75913 );
not ( n83637 , n75905 );
and ( n83638 , n83637 , n31994 );
and ( n83639 , n59005 , n75905 );
or ( n83640 , n83638 , n83639 );
and ( n83641 , n83636 , n83640 );
and ( n83642 , n59005 , n75913 );
or ( n83643 , n83641 , n83642 );
and ( n83644 , n83635 , n83643 );
not ( n83645 , n75933 );
not ( n83646 , n75935 );
and ( n83647 , n83646 , n83643 );
and ( n83648 , n59029 , n75935 );
or ( n83649 , n83647 , n83648 );
and ( n83650 , n83645 , n83649 );
and ( n83651 , n59037 , n75933 );
or ( n83652 , n83650 , n83651 );
and ( n83653 , n83652 , n32475 );
or ( n83654 , n83644 , n83653 );
and ( n83655 , n83654 , n32486 );
and ( n83656 , n31994 , n41278 );
or ( n83657 , C0 , n83625 , n83634 , n83655 , n83656 );
buf ( n83658 , n83657 );
buf ( n83659 , n83658 );
buf ( n83660 , n30987 );
buf ( n83661 , n30987 );
xor ( n83662 , n35439 , n39944 );
and ( n83663 , n83662 , n31550 );
not ( n83664 , n39979 );
and ( n83665 , n83664 , n35439 );
and ( n83666 , n77283 , n39979 );
or ( n83667 , n83665 , n83666 );
and ( n83668 , n83667 , n31538 );
and ( n83669 , n35439 , n40143 );
or ( n83670 , n83663 , n83668 , n83669 );
and ( n83671 , n83670 , n31557 );
and ( n83672 , n35439 , n40154 );
or ( n83673 , C0 , n83671 , n83672 );
buf ( n83674 , n83673 );
buf ( n83675 , n83674 );
buf ( n83676 , n30987 );
and ( n83677 , n52176 , n31645 );
not ( n83678 , n45274 );
and ( n83679 , n83678 , n66889 );
and ( n83680 , n83277 , n45274 );
or ( n83681 , n83679 , n83680 );
and ( n83682 , n83681 , n31373 );
not ( n83683 , n45280 );
and ( n83684 , n83683 , n66889 );
and ( n83685 , n83277 , n45280 );
or ( n83686 , n83684 , n83685 );
and ( n83687 , n83686 , n31468 );
and ( n83688 , n66889 , n45802 );
or ( n83689 , n83682 , n83687 , n83688 );
and ( n83690 , n83689 , n31557 );
and ( n83691 , n66889 , n45808 );
or ( n83692 , C0 , n83677 , n83690 , n83691 );
buf ( n83693 , n83692 );
buf ( n83694 , n83693 );
buf ( n83695 , n31655 );
not ( n83696 , n40163 );
and ( n83697 , n83696 , n31830 );
not ( n83698 , n56287 );
and ( n83699 , n83698 , n31830 );
and ( n83700 , n32235 , n56287 );
or ( n83701 , n83699 , n83700 );
and ( n83702 , n83701 , n40163 );
or ( n83703 , n83697 , n83702 );
and ( n83704 , n83703 , n32498 );
not ( n83705 , n56295 );
not ( n83706 , n56287 );
and ( n83707 , n83706 , n31830 );
and ( n83708 , n42188 , n56287 );
or ( n83709 , n83707 , n83708 );
and ( n83710 , n83705 , n83709 );
and ( n83711 , n42188 , n56295 );
or ( n83712 , n83710 , n83711 );
and ( n83713 , n83712 , n32473 );
not ( n83714 , n32475 );
not ( n83715 , n56295 );
not ( n83716 , n56287 );
and ( n83717 , n83716 , n31830 );
and ( n83718 , n42188 , n56287 );
or ( n83719 , n83717 , n83718 );
and ( n83720 , n83715 , n83719 );
and ( n83721 , n42188 , n56295 );
or ( n83722 , n83720 , n83721 );
and ( n83723 , n83714 , n83722 );
not ( n83724 , n56315 );
not ( n83725 , n56317 );
and ( n83726 , n83725 , n83722 );
and ( n83727 , n42216 , n56317 );
or ( n83728 , n83726 , n83727 );
and ( n83729 , n83724 , n83728 );
and ( n83730 , n42224 , n56315 );
or ( n83731 , n83729 , n83730 );
and ( n83732 , n83731 , n32475 );
or ( n83733 , n83723 , n83732 );
and ( n83734 , n83733 , n32486 );
and ( n83735 , n31830 , n41278 );
or ( n83736 , C0 , n83704 , n83713 , n83734 , n83735 );
buf ( n83737 , n83736 );
buf ( n83738 , n83737 );
not ( n83739 , n31437 );
and ( n83740 , n83739 , n58634 );
not ( n83741 , n41809 );
and ( n83742 , n83741 , n41662 );
xor ( n83743 , n41816 , n41824 );
and ( n83744 , n83743 , n41809 );
or ( n83745 , n83742 , n83744 );
and ( n83746 , n83745 , n31437 );
or ( n83747 , n83740 , n83746 );
and ( n83748 , n83747 , n31468 );
not ( n83749 , n41837 );
and ( n83750 , n83749 , n58634 );
and ( n83751 , n58640 , n41837 );
or ( n83752 , n83750 , n83751 );
and ( n83753 , n83752 , n31521 );
and ( n83754 , n58634 , n42158 );
or ( n83755 , n83748 , n83753 , n83754 );
and ( n83756 , n83755 , n31557 );
and ( n83757 , n58634 , n40154 );
or ( n83758 , C0 , n83756 , n83757 );
buf ( n83759 , n83758 );
buf ( n83760 , n83759 );
not ( n83761 , n40163 );
and ( n83762 , n83761 , n31966 );
not ( n83763 , n56988 );
and ( n83764 , n83763 , n31966 );
and ( n83765 , n32165 , n56988 );
or ( n83766 , n83764 , n83765 );
and ( n83767 , n83766 , n40163 );
or ( n83768 , n83762 , n83767 );
and ( n83769 , n83768 , n32498 );
not ( n83770 , n56996 );
not ( n83771 , n56988 );
and ( n83772 , n83771 , n31966 );
and ( n83773 , n59005 , n56988 );
or ( n83774 , n83772 , n83773 );
and ( n83775 , n83770 , n83774 );
and ( n83776 , n59005 , n56996 );
or ( n83777 , n83775 , n83776 );
and ( n83778 , n83777 , n32473 );
not ( n83779 , n32475 );
not ( n83780 , n56996 );
not ( n83781 , n56988 );
and ( n83782 , n83781 , n31966 );
and ( n83783 , n59005 , n56988 );
or ( n83784 , n83782 , n83783 );
and ( n83785 , n83780 , n83784 );
and ( n83786 , n59005 , n56996 );
or ( n83787 , n83785 , n83786 );
and ( n83788 , n83779 , n83787 );
not ( n83789 , n57016 );
not ( n83790 , n57018 );
and ( n83791 , n83790 , n83787 );
and ( n83792 , n59029 , n57018 );
or ( n83793 , n83791 , n83792 );
and ( n83794 , n83789 , n83793 );
and ( n83795 , n59037 , n57016 );
or ( n83796 , n83794 , n83795 );
and ( n83797 , n83796 , n32475 );
or ( n83798 , n83788 , n83797 );
and ( n83799 , n83798 , n32486 );
and ( n83800 , n31966 , n41278 );
or ( n83801 , C0 , n83769 , n83778 , n83799 , n83800 );
buf ( n83802 , n83801 );
buf ( n83803 , n83802 );
buf ( n83804 , n31655 );
buf ( n83805 , n30987 );
buf ( n83806 , n31655 );
xor ( n83807 , n34042 , n39936 );
and ( n83808 , n83807 , n31550 );
not ( n83809 , n39979 );
and ( n83810 , n83809 , n34042 );
and ( n83811 , n31307 , n42330 );
and ( n83812 , n31309 , n42332 );
and ( n83813 , n31311 , n42334 );
and ( n83814 , n31313 , n42336 );
and ( n83815 , n31315 , n42338 );
and ( n83816 , n31317 , n42340 );
and ( n83817 , n31319 , n42342 );
and ( n83818 , n31321 , n42344 );
and ( n83819 , n31323 , n42346 );
and ( n83820 , n31325 , n42348 );
and ( n83821 , n31327 , n42350 );
and ( n83822 , n31329 , n42352 );
and ( n83823 , n31331 , n42354 );
and ( n83824 , n31333 , n42356 );
and ( n83825 , n31335 , n42358 );
and ( n83826 , n31337 , n42360 );
or ( n83827 , n83811 , n83812 , n83813 , n83814 , n83815 , n83816 , n83817 , n83818 , n83819 , n83820 , n83821 , n83822 , n83823 , n83824 , n83825 , n83826 );
and ( n83828 , n83827 , n39979 );
or ( n83829 , n83810 , n83828 );
and ( n83830 , n83829 , n31538 );
and ( n83831 , n34042 , n40143 );
or ( n83832 , n83808 , n83830 , n83831 );
and ( n83833 , n83832 , n31557 );
and ( n83834 , n34042 , n40154 );
or ( n83835 , C0 , n83833 , n83834 );
buf ( n83836 , n83835 );
buf ( n83837 , n83836 );
buf ( n83838 , n30987 );
buf ( n83839 , n30987 );
not ( n83840 , n40163 );
and ( n83841 , n83840 , n31992 );
not ( n83842 , n42238 );
and ( n83843 , n83842 , n31992 );
and ( n83844 , n32165 , n42238 );
or ( n83845 , n83843 , n83844 );
and ( n83846 , n83845 , n40163 );
or ( n83847 , n83841 , n83846 );
and ( n83848 , n83847 , n32498 );
not ( n83849 , n42247 );
not ( n83850 , n42238 );
and ( n83851 , n83850 , n31992 );
and ( n83852 , n59005 , n42238 );
or ( n83853 , n83851 , n83852 );
and ( n83854 , n83849 , n83853 );
and ( n83855 , n59005 , n42247 );
or ( n83856 , n83854 , n83855 );
and ( n83857 , n83856 , n32473 );
not ( n83858 , n32475 );
not ( n83859 , n42247 );
not ( n83860 , n42238 );
and ( n83861 , n83860 , n31992 );
and ( n83862 , n59005 , n42238 );
or ( n83863 , n83861 , n83862 );
and ( n83864 , n83859 , n83863 );
and ( n83865 , n59005 , n42247 );
or ( n83866 , n83864 , n83865 );
and ( n83867 , n83858 , n83866 );
not ( n83868 , n42273 );
not ( n83869 , n42276 );
and ( n83870 , n83869 , n83866 );
and ( n83871 , n59029 , n42276 );
or ( n83872 , n83870 , n83871 );
and ( n83873 , n83868 , n83872 );
and ( n83874 , n59037 , n42273 );
or ( n83875 , n83873 , n83874 );
and ( n83876 , n83875 , n32475 );
or ( n83877 , n83867 , n83876 );
and ( n83878 , n83877 , n32486 );
and ( n83879 , n31992 , n41278 );
or ( n83880 , C0 , n83848 , n83857 , n83878 , n83879 );
buf ( n83881 , n83880 );
buf ( n83882 , n83881 );
buf ( n83883 , n31655 );
and ( n83884 , n69808 , n33377 );
not ( n83885 , n48545 );
and ( n83886 , n83885 , n65367 );
buf ( n83887 , n83886 );
and ( n83888 , n83887 , n32890 );
not ( n83889 , n48557 );
and ( n83890 , n83889 , n65367 );
and ( n83891 , n69814 , n48557 );
or ( n83892 , n83890 , n83891 );
and ( n83893 , n83892 , n33038 );
and ( n83894 , n65367 , n48571 );
or ( n83895 , n83888 , n83893 , n83894 );
and ( n83896 , n83895 , n33208 );
and ( n83897 , n65367 , n48577 );
or ( n83898 , C0 , n83884 , n83896 , n83897 );
buf ( n83899 , n83898 );
buf ( n83900 , n83899 );
buf ( n83901 , n31655 );
buf ( n83902 , n30987 );
buf ( n83903 , n30987 );
xor ( n83904 , n46224 , n49996 );
and ( n83905 , n83904 , n32431 );
not ( n83906 , n50002 );
and ( n83907 , n83906 , n46224 );
and ( n83908 , n40493 , n50002 );
or ( n83909 , n83907 , n83908 );
and ( n83910 , n83909 , n32419 );
not ( n83911 , n50008 );
and ( n83912 , n83911 , n46224 );
not ( n83913 , n47910 );
and ( n83914 , n83913 , n69391 );
not ( n83915 , n48101 );
and ( n83916 , n83915 , n48049 );
xor ( n83917 , n50019 , n50026 );
and ( n83918 , n83917 , n48101 );
or ( n83919 , n83916 , n83918 );
and ( n83920 , n83919 , n47910 );
or ( n83921 , n83914 , n83920 );
and ( n83922 , n83921 , n50008 );
or ( n83923 , n83912 , n83922 );
and ( n83924 , n83923 , n32415 );
not ( n83925 , n50067 );
and ( n83926 , n83925 , n46224 );
and ( n83927 , n72653 , n50067 );
or ( n83928 , n83926 , n83927 );
and ( n83929 , n83928 , n32411 );
and ( n83930 , n46224 , n50098 );
or ( n83931 , n83905 , n83910 , n83924 , n83929 , n83930 );
and ( n83932 , n83931 , n32456 );
and ( n83933 , n46224 , n47409 );
or ( n83934 , C0 , n83932 , n83933 );
buf ( n83935 , n83934 );
buf ( n83936 , n83935 );
buf ( n83937 , n31655 );
not ( n83938 , n46356 );
and ( n83939 , n83938 , n31292 );
not ( n83940 , n50109 );
and ( n83941 , n83940 , n31292 );
and ( n83942 , n31306 , n50109 );
or ( n83943 , n83941 , n83942 );
and ( n83944 , n83943 , n46356 );
or ( n83945 , n83939 , n83944 );
and ( n83946 , n83945 , n31649 );
not ( n83947 , n50117 );
not ( n83948 , n50109 );
and ( n83949 , n83948 , n31292 );
and ( n83950 , n58061 , n50109 );
or ( n83951 , n83949 , n83950 );
and ( n83952 , n83947 , n83951 );
and ( n83953 , n58061 , n50117 );
or ( n83954 , n83952 , n83953 );
and ( n83955 , n83954 , n31643 );
not ( n83956 , n31452 );
not ( n83957 , n50117 );
not ( n83958 , n50109 );
and ( n83959 , n83958 , n31292 );
and ( n83960 , n58061 , n50109 );
or ( n83961 , n83959 , n83960 );
and ( n83962 , n83957 , n83961 );
and ( n83963 , n58061 , n50117 );
or ( n83964 , n83962 , n83963 );
and ( n83965 , n83956 , n83964 );
not ( n83966 , n50142 );
not ( n83967 , n50144 );
and ( n83968 , n83967 , n83964 );
and ( n83969 , n58085 , n50144 );
or ( n83970 , n83968 , n83969 );
and ( n83971 , n83966 , n83970 );
and ( n83972 , n58093 , n50142 );
or ( n83973 , n83971 , n83972 );
and ( n83974 , n83973 , n31452 );
or ( n83975 , n83965 , n83974 );
and ( n83976 , n83975 , n31638 );
and ( n83977 , n31292 , n47277 );
or ( n83978 , C0 , n83946 , n83955 , n83976 , n83977 );
buf ( n83979 , n83978 );
buf ( n83980 , n83979 );
buf ( n83981 , n30987 );
buf ( n83982 , n31655 );
buf ( n83983 , n30987 );
not ( n83984 , n40163 );
and ( n83985 , n83984 , n31968 );
not ( n83986 , n42171 );
and ( n83987 , n83986 , n31968 );
and ( n83988 , n32165 , n42171 );
or ( n83989 , n83987 , n83988 );
and ( n83990 , n83989 , n40163 );
or ( n83991 , n83985 , n83990 );
and ( n83992 , n83991 , n32498 );
not ( n83993 , n42180 );
not ( n83994 , n42171 );
and ( n83995 , n83994 , n31968 );
and ( n83996 , n59005 , n42171 );
or ( n83997 , n83995 , n83996 );
and ( n83998 , n83993 , n83997 );
and ( n83999 , n59005 , n42180 );
or ( n84000 , n83998 , n83999 );
and ( n84001 , n84000 , n32473 );
not ( n84002 , n32475 );
not ( n84003 , n42180 );
not ( n84004 , n42171 );
and ( n84005 , n84004 , n31968 );
and ( n84006 , n59005 , n42171 );
or ( n84007 , n84005 , n84006 );
and ( n84008 , n84003 , n84007 );
and ( n84009 , n59005 , n42180 );
or ( n84010 , n84008 , n84009 );
and ( n84011 , n84002 , n84010 );
not ( n84012 , n42206 );
not ( n84013 , n42209 );
and ( n84014 , n84013 , n84010 );
and ( n84015 , n59029 , n42209 );
or ( n84016 , n84014 , n84015 );
and ( n84017 , n84012 , n84016 );
and ( n84018 , n59037 , n42206 );
or ( n84019 , n84017 , n84018 );
and ( n84020 , n84019 , n32475 );
or ( n84021 , n84011 , n84020 );
and ( n84022 , n84021 , n32486 );
and ( n84023 , n31968 , n41278 );
or ( n84024 , C0 , n83992 , n84001 , n84022 , n84023 );
buf ( n84025 , n84024 );
buf ( n84026 , n84025 );
buf ( n84027 , n31655 );
not ( n84028 , n31437 );
and ( n84029 , n84028 , n65626 );
and ( n84030 , n81122 , n31437 );
or ( n84031 , n84029 , n84030 );
and ( n84032 , n84031 , n31468 );
not ( n84033 , n41837 );
and ( n84034 , n84033 , n65626 );
and ( n84035 , n65632 , n41837 );
or ( n84036 , n84034 , n84035 );
and ( n84037 , n84036 , n31521 );
and ( n84038 , n65626 , n42158 );
or ( n84039 , n84032 , n84037 , n84038 );
and ( n84040 , n84039 , n31557 );
and ( n84041 , n65626 , n40154 );
or ( n84042 , C0 , n84040 , n84041 );
buf ( n84043 , n84042 );
buf ( n84044 , n84043 );
and ( n84045 , n31569 , n31007 );
not ( n84046 , n31077 );
and ( n84047 , n84046 , n35395 );
buf ( n84048 , n84047 );
and ( n84049 , n84048 , n31373 );
not ( n84050 , n31402 );
and ( n84051 , n84050 , n35395 );
buf ( n84052 , n84051 );
and ( n84053 , n84052 , n31408 );
not ( n84054 , n31437 );
and ( n84055 , n84054 , n35395 );
not ( n84056 , n31455 );
and ( n84057 , n84056 , n35439 );
xor ( n84058 , n35395 , n35403 );
and ( n84059 , n84058 , n31455 );
or ( n84060 , n84057 , n84059 );
and ( n84061 , n84060 , n31437 );
or ( n84062 , n84055 , n84061 );
and ( n84063 , n84062 , n31468 );
not ( n84064 , n31497 );
and ( n84065 , n84064 , n35395 );
not ( n84066 , n31454 );
not ( n84067 , n31501 );
and ( n84068 , n84067 , n35439 );
xor ( n84069 , n35440 , n35453 );
and ( n84070 , n84069 , n31501 );
or ( n84071 , n84068 , n84070 );
and ( n84072 , n84066 , n84071 );
and ( n84073 , n84058 , n31454 );
or ( n84074 , n84072 , n84073 );
and ( n84075 , n84074 , n31497 );
or ( n84076 , n84065 , n84075 );
and ( n84077 , n84076 , n31521 );
and ( n84078 , n35395 , n31553 );
or ( n84079 , n84049 , n84053 , n84063 , n84077 , n84078 );
and ( n84080 , n84079 , n31557 );
not ( n84081 , n31452 );
not ( n84082 , n31619 );
and ( n84083 , n84082 , n35494 );
xor ( n84084 , n35495 , n35507 );
and ( n84085 , n84084 , n31619 );
or ( n84086 , n84083 , n84085 );
and ( n84087 , n84081 , n84086 );
and ( n84088 , n35395 , n31452 );
or ( n84089 , n84087 , n84088 );
and ( n84090 , n84089 , n31638 );
and ( n84091 , n35395 , n31650 );
or ( n84092 , C0 , n84045 , n84080 , n84090 , C0 , n84091 );
buf ( n84093 , n84092 );
buf ( n84094 , n84093 );
not ( n84095 , n33419 );
and ( n84096 , n84095 , n31575 );
and ( n84097 , n56788 , n33419 );
or ( n84098 , n84096 , n84097 );
and ( n84099 , n84098 , n31529 );
not ( n84100 , n33734 );
and ( n84101 , n84100 , n31575 );
and ( n84102 , n56799 , n33734 );
or ( n84103 , n84101 , n84102 );
and ( n84104 , n84103 , n31527 );
and ( n84105 , n31575 , n33942 );
or ( n84106 , n84099 , n84104 , n84105 );
and ( n84107 , n84106 , n31557 );
and ( n84108 , n34095 , n31643 );
not ( n84109 , n31452 );
and ( n84110 , n84109 , n34095 );
xor ( n84111 , n31575 , n33962 );
and ( n84112 , n84111 , n31452 );
or ( n84113 , n84110 , n84112 );
and ( n84114 , n84113 , n31638 );
and ( n84115 , n33999 , n33973 );
and ( n84116 , n31575 , n33978 );
or ( n84117 , C0 , n84107 , n84108 , n84114 , n84115 , n84116 );
buf ( n84118 , n84117 );
buf ( n84119 , n84118 );
buf ( n84120 , n30987 );
buf ( n84121 , n31655 );
buf ( n84122 , n31655 );
buf ( n84123 , n30987 );
buf ( n84124 , n31655 );
and ( n84125 , n57090 , n31645 );
not ( n84126 , n45274 );
and ( n84127 , n84126 , n64906 );
buf ( n84128 , n84127 );
and ( n84129 , n84128 , n31373 );
not ( n84130 , n45280 );
and ( n84131 , n84130 , n64906 );
and ( n84132 , n57096 , n45280 );
or ( n84133 , n84131 , n84132 );
and ( n84134 , n84133 , n31468 );
and ( n84135 , n64906 , n45802 );
or ( n84136 , n84129 , n84134 , n84135 );
and ( n84137 , n84136 , n31557 );
and ( n84138 , n64906 , n45808 );
or ( n84139 , C0 , n84125 , n84137 , n84138 );
buf ( n84140 , n84139 );
buf ( n84141 , n84140 );
not ( n84142 , n40163 );
and ( n84143 , n84142 , n31904 );
not ( n84144 , n54629 );
and ( n84145 , n84144 , n31904 );
and ( n84146 , n32200 , n54629 );
or ( n84147 , n84145 , n84146 );
and ( n84148 , n84147 , n40163 );
or ( n84149 , n84143 , n84148 );
and ( n84150 , n84149 , n32498 );
not ( n84151 , n54637 );
not ( n84152 , n54629 );
and ( n84153 , n84152 , n31904 );
and ( n84154 , n53243 , n54629 );
or ( n84155 , n84153 , n84154 );
and ( n84156 , n84151 , n84155 );
and ( n84157 , n53243 , n54637 );
or ( n84158 , n84156 , n84157 );
and ( n84159 , n84158 , n32473 );
not ( n84160 , n32475 );
not ( n84161 , n54637 );
not ( n84162 , n54629 );
and ( n84163 , n84162 , n31904 );
and ( n84164 , n53243 , n54629 );
or ( n84165 , n84163 , n84164 );
and ( n84166 , n84161 , n84165 );
and ( n84167 , n53243 , n54637 );
or ( n84168 , n84166 , n84167 );
and ( n84169 , n84160 , n84168 );
not ( n84170 , n54657 );
not ( n84171 , n54659 );
and ( n84172 , n84171 , n84168 );
and ( n84173 , n53269 , n54659 );
or ( n84174 , n84172 , n84173 );
and ( n84175 , n84170 , n84174 );
and ( n84176 , n53277 , n54657 );
or ( n84177 , n84175 , n84176 );
and ( n84178 , n84177 , n32475 );
or ( n84179 , n84169 , n84178 );
and ( n84180 , n84179 , n32486 );
and ( n84181 , n31904 , n41278 );
or ( n84182 , C0 , n84150 , n84159 , n84180 , n84181 );
buf ( n84183 , n84182 );
buf ( n84184 , n84183 );
buf ( n84185 , n30987 );
buf ( n84186 , n31655 );
and ( n84187 , n46036 , n32500 );
not ( n84188 , n35211 );
and ( n84189 , n84188 , n37569 );
buf ( n84190 , n84189 );
and ( n84191 , n84190 , n32421 );
not ( n84192 , n35245 );
and ( n84193 , n84192 , n37569 );
buf ( n84194 , n84193 );
and ( n84195 , n84194 , n32419 );
not ( n84196 , n35278 );
and ( n84197 , n84196 , n37569 );
not ( n84198 , n35295 );
and ( n84199 , n84198 , n49599 );
xor ( n84200 , n37569 , n49531 );
and ( n84201 , n84200 , n35295 );
or ( n84202 , n84199 , n84201 );
and ( n84203 , n84202 , n35278 );
or ( n84204 , n84197 , n84203 );
and ( n84205 , n84204 , n32417 );
not ( n84206 , n35331 );
and ( n84207 , n84206 , n37569 );
not ( n84208 , n35294 );
not ( n84209 , n45995 );
and ( n84210 , n84209 , n49599 );
xor ( n84211 , n49600 , n49617 );
and ( n84212 , n84211 , n45995 );
or ( n84213 , n84210 , n84212 );
and ( n84214 , n84208 , n84213 );
and ( n84215 , n84200 , n35294 );
or ( n84216 , n84214 , n84215 );
and ( n84217 , n84216 , n35331 );
or ( n84218 , n84207 , n84217 );
and ( n84219 , n84218 , n32415 );
and ( n84220 , n37569 , n35354 );
or ( n84221 , n84191 , n84195 , n84205 , n84219 , n84220 );
and ( n84222 , n84221 , n32456 );
not ( n84223 , n32475 );
not ( n84224 , n46060 );
and ( n84225 , n84224 , n49689 );
xor ( n84226 , n49690 , n49711 );
and ( n84227 , n84226 , n46060 );
or ( n84228 , n84225 , n84227 );
and ( n84229 , n84223 , n84228 );
and ( n84230 , n37569 , n32475 );
or ( n84231 , n84229 , n84230 );
and ( n84232 , n84231 , n32486 );
buf ( n84233 , n32489 );
and ( n84234 , n37569 , n35367 );
or ( n84235 , C0 , n84187 , n84222 , n84232 , n84233 , n84234 );
buf ( n84236 , n84235 );
buf ( n84237 , n84236 );
buf ( n84238 , n30987 );
not ( n84239 , n48765 );
and ( n84240 , n84239 , n33214 );
and ( n84241 , n73988 , n48765 );
or ( n84242 , n84240 , n84241 );
and ( n84243 , n84242 , n33180 );
not ( n84244 , n49054 );
and ( n84245 , n84244 , n33214 );
and ( n84246 , n73999 , n49054 );
or ( n84247 , n84245 , n84246 );
and ( n84248 , n84247 , n33178 );
and ( n84249 , n33214 , n49774 );
or ( n84250 , n84243 , n84248 , n84249 );
and ( n84251 , n84250 , n33208 );
and ( n84252 , n33279 , n33375 );
not ( n84253 , n32968 );
and ( n84254 , n84253 , n33279 );
xor ( n84255 , n33214 , n66021 );
and ( n84256 , n84255 , n32968 );
or ( n84257 , n84254 , n84256 );
and ( n84258 , n84257 , n33370 );
and ( n84259 , n32977 , n35056 );
and ( n84260 , n33214 , n49794 );
or ( n84261 , C0 , n84251 , n84252 , n84258 , n84259 , n84260 );
buf ( n84262 , n84261 );
buf ( n84263 , n84262 );
buf ( n84264 , n30987 );
buf ( n84265 , n31655 );
buf ( n84266 , n39348 );
and ( n84267 , n33758 , n48455 );
not ( n84268 , n48457 );
and ( n84269 , n84268 , n33423 );
and ( n84270 , n33758 , n48457 );
or ( n84271 , n84269 , n84270 );
and ( n84272 , n84271 , n31373 );
not ( n84273 , n44807 );
and ( n84274 , n84273 , n33423 );
and ( n84275 , n33758 , n44807 );
or ( n84276 , n84274 , n84275 );
and ( n84277 , n84276 , n31408 );
not ( n84278 , n48468 );
and ( n84279 , n84278 , n33423 );
and ( n84280 , n33758 , n48468 );
or ( n84281 , n84279 , n84280 );
and ( n84282 , n84281 , n31468 );
not ( n84283 , n44817 );
and ( n84284 , n84283 , n33423 );
and ( n84285 , n33758 , n44817 );
or ( n84286 , n84284 , n84285 );
and ( n84287 , n84286 , n31521 );
not ( n84288 , n39979 );
and ( n84289 , n84288 , n33423 );
and ( n84290 , n33465 , n39979 );
or ( n84291 , n84289 , n84290 );
and ( n84292 , n84291 , n31538 );
not ( n84293 , n45059 );
and ( n84294 , n84293 , n33423 );
and ( n84295 , n33465 , n45059 );
or ( n84296 , n84294 , n84295 );
and ( n84297 , n84296 , n31536 );
not ( n84298 , n33419 );
and ( n84299 , n84298 , n33423 );
and ( n84300 , n66534 , n33419 );
or ( n84301 , n84299 , n84300 );
and ( n84302 , n84301 , n31529 );
not ( n84303 , n33734 );
and ( n84304 , n84303 , n33423 );
and ( n84305 , n66545 , n33734 );
or ( n84306 , n84304 , n84305 );
and ( n84307 , n84306 , n31527 );
and ( n84308 , n33843 , n48513 );
or ( n84309 , n84267 , n84272 , n84277 , n84282 , n84287 , n84292 , n84297 , n84302 , n84307 , n84308 );
and ( n84310 , n84309 , n31557 );
and ( n84311 , n35396 , n33973 );
and ( n84312 , n33423 , n48524 );
or ( n84313 , C0 , n84310 , n84311 , n84312 );
buf ( n84314 , n84313 );
buf ( n84315 , n84314 );
buf ( n84316 , n31655 );
buf ( n84317 , n30987 );
not ( n84318 , n38443 );
and ( n84319 , n84318 , n38405 );
xor ( n84320 , n69917 , n69920 );
and ( n84321 , n84320 , n38443 );
or ( n84322 , n84319 , n84321 );
and ( n84323 , n84322 , n38450 );
not ( n84324 , n39339 );
and ( n84325 , n84324 , n39305 );
xor ( n84326 , n69931 , n69934 );
and ( n84327 , n84326 , n39339 );
or ( n84328 , n84325 , n84327 );
and ( n84329 , n84328 , n39346 );
and ( n84330 , n40159 , n39359 );
or ( n84331 , n84323 , n84329 , n84330 );
buf ( n84332 , n84331 );
buf ( n84333 , n84332 );
buf ( n84334 , n31655 );
and ( n84335 , n47658 , n50275 );
not ( n84336 , n50278 );
and ( n84337 , n84336 , n47571 );
and ( n84338 , n47658 , n50278 );
or ( n84339 , n84337 , n84338 );
and ( n84340 , n84339 , n32421 );
not ( n84341 , n50002 );
and ( n84342 , n84341 , n47571 );
and ( n84343 , n47658 , n50002 );
or ( n84344 , n84342 , n84343 );
and ( n84345 , n84344 , n32419 );
not ( n84346 , n50289 );
and ( n84347 , n84346 , n47571 );
and ( n84348 , n47658 , n50289 );
or ( n84349 , n84347 , n84348 );
and ( n84350 , n84349 , n32417 );
not ( n84351 , n50008 );
and ( n84352 , n84351 , n47571 );
and ( n84353 , n47658 , n50008 );
or ( n84354 , n84352 , n84353 );
and ( n84355 , n84354 , n32415 );
not ( n84356 , n47331 );
and ( n84357 , n84356 , n47571 );
and ( n84358 , n47603 , n47331 );
or ( n84359 , n84357 , n84358 );
and ( n84360 , n84359 , n32413 );
not ( n84361 , n50067 );
and ( n84362 , n84361 , n47571 );
and ( n84363 , n47603 , n50067 );
or ( n84364 , n84362 , n84363 );
and ( n84365 , n84364 , n32411 );
not ( n84366 , n31728 );
and ( n84367 , n84366 , n47571 );
xor ( n84368 , n47603 , n47626 );
and ( n84369 , n84368 , n31728 );
or ( n84370 , n84367 , n84369 );
and ( n84371 , n84370 , n32253 );
not ( n84372 , n32283 );
and ( n84373 , n84372 , n47571 );
not ( n84374 , n31823 );
xor ( n84375 , n47658 , n47681 );
and ( n84376 , n84374 , n84375 );
xnor ( n84377 , n47708 , n47731 );
and ( n84378 , n84377 , n31823 );
or ( n84379 , n84376 , n84378 );
and ( n84380 , n84379 , n32283 );
or ( n84381 , n84373 , n84380 );
and ( n84382 , n84381 , n32398 );
and ( n84383 , n47708 , n50334 );
or ( n84384 , n84335 , n84340 , n84345 , n84350 , n84355 , n84360 , n84365 , n84371 , n84382 , n84383 );
and ( n84385 , n84384 , n32456 );
and ( n84386 , n37549 , n32489 );
and ( n84387 , n47571 , n50345 );
or ( n84388 , C0 , n84385 , n84386 , n84387 );
buf ( n84389 , n84388 );
buf ( n84390 , n84389 );
buf ( n84391 , n30987 );
not ( n84392 , n36587 );
and ( n84393 , n84392 , n36532 );
xor ( n84394 , n61940 , n61945 );
and ( n84395 , n84394 , n36587 );
or ( n84396 , n84393 , n84395 );
and ( n84397 , n84396 , n36596 );
not ( n84398 , n37485 );
and ( n84399 , n84398 , n37434 );
xor ( n84400 , n61956 , n61961 );
and ( n84401 , n84400 , n37485 );
or ( n84402 , n84399 , n84401 );
and ( n84403 , n84402 , n37494 );
and ( n84404 , n41865 , n37506 );
or ( n84405 , n84397 , n84403 , n84404 );
buf ( n84406 , n84405 );
buf ( n84407 , n84406 );
not ( n84408 , n31728 );
and ( n84409 , n84408 , n46031 );
and ( n84410 , n58965 , n31728 );
or ( n84411 , n84409 , n84410 );
and ( n84412 , n84411 , n32253 );
not ( n84413 , n32283 );
and ( n84414 , n84413 , n46031 );
and ( n84415 , n58976 , n32283 );
or ( n84416 , n84414 , n84415 );
and ( n84417 , n84416 , n32398 );
and ( n84418 , n46031 , n32436 );
or ( n84419 , n84412 , n84417 , n84418 );
and ( n84420 , n84419 , n32456 );
and ( n84421 , n49679 , n32473 );
not ( n84422 , n32475 );
and ( n84423 , n84422 , n49679 );
xor ( n84424 , n46031 , n47755 );
and ( n84425 , n84424 , n32475 );
or ( n84426 , n84423 , n84425 );
and ( n84427 , n84426 , n32486 );
and ( n84428 , n37559 , n32489 );
and ( n84429 , n46031 , n32501 );
or ( n84430 , C0 , n84420 , n84421 , n84427 , n84428 , n84429 );
buf ( n84431 , n84430 );
buf ( n84432 , n84431 );
buf ( n84433 , n31655 );
buf ( n84434 , n30987 );
and ( n84435 , n33219 , n32528 );
not ( n84436 , n32598 );
and ( n84437 , n84436 , n32982 );
buf ( n84438 , n84437 );
and ( n84439 , n84438 , n32890 );
not ( n84440 , n32919 );
and ( n84441 , n84440 , n32982 );
buf ( n84442 , n84441 );
and ( n84443 , n84442 , n32924 );
not ( n84444 , n32953 );
and ( n84445 , n84444 , n32982 );
not ( n84446 , n32971 );
and ( n84447 , n84446 , n33089 );
xor ( n84448 , n32982 , n33023 );
and ( n84449 , n84448 , n32971 );
or ( n84450 , n84447 , n84449 );
and ( n84451 , n84450 , n32953 );
or ( n84452 , n84445 , n84451 );
and ( n84453 , n84452 , n33038 );
not ( n84454 , n33067 );
and ( n84455 , n84454 , n32982 );
not ( n84456 , n32970 );
not ( n84457 , n33071 );
and ( n84458 , n84457 , n33089 );
xor ( n84459 , n33090 , n33155 );
and ( n84460 , n84459 , n33071 );
or ( n84461 , n84458 , n84460 );
and ( n84462 , n84456 , n84461 );
and ( n84463 , n84448 , n32970 );
or ( n84464 , n84462 , n84463 );
and ( n84465 , n84464 , n33067 );
or ( n84466 , n84455 , n84465 );
and ( n84467 , n84466 , n33172 );
and ( n84468 , n32982 , n33204 );
or ( n84469 , n84439 , n84443 , n84453 , n84467 , n84468 );
and ( n84470 , n84469 , n33208 );
not ( n84471 , n32968 );
not ( n84472 , n33270 );
and ( n84473 , n84472 , n33289 );
xor ( n84474 , n33290 , n33355 );
and ( n84475 , n84474 , n33270 );
or ( n84476 , n84473 , n84475 );
and ( n84477 , n84471 , n84476 );
and ( n84478 , n32982 , n32968 );
or ( n84479 , n84477 , n84478 );
and ( n84480 , n84479 , n33370 );
and ( n84481 , n32982 , n33382 );
or ( n84482 , C0 , n84435 , n84470 , n84480 , C0 , n84481 );
buf ( n84483 , n84482 );
buf ( n84484 , n84483 );
buf ( n84485 , n30987 );
buf ( n84486 , n31655 );
not ( n84487 , n38443 );
and ( n84488 , n84487 , n38150 );
xor ( n84489 , n53473 , n53496 );
and ( n84490 , n84489 , n38443 );
or ( n84491 , n84488 , n84490 );
and ( n84492 , n84491 , n38450 );
not ( n84493 , n39339 );
and ( n84494 , n84493 , n39050 );
xor ( n84495 , n53529 , n53552 );
and ( n84496 , n84495 , n39339 );
or ( n84497 , n84494 , n84496 );
and ( n84498 , n84497 , n39346 );
and ( n84499 , n40211 , n39359 );
or ( n84500 , n84492 , n84498 , n84499 );
buf ( n84501 , n84500 );
buf ( n84502 , n84501 );
buf ( n84503 , n31655 );
and ( n84504 , n33499 , n46356 );
buf ( n84505 , n84504 );
and ( n84506 , n84505 , n31649 );
and ( n84507 , n52552 , n31647 );
and ( n84508 , n63691 , n31557 );
and ( n84509 , n31014 , n61220 );
or ( n84510 , C0 , n84506 , n84507 , n84508 , n84509 );
buf ( n84511 , n84510 );
buf ( n84512 , n84511 );
buf ( n84513 , n30987 );
buf ( n84514 , n30987 );
buf ( n84515 , n31655 );
buf ( n84516 , n31655 );
buf ( n84517 , n30987 );
not ( n84518 , n31728 );
and ( n84519 , n84518 , n46023 );
and ( n84520 , n50312 , n31728 );
or ( n84521 , n84519 , n84520 );
and ( n84522 , n84521 , n32253 );
not ( n84523 , n32283 );
and ( n84524 , n84523 , n46023 );
and ( n84525 , n50323 , n32283 );
or ( n84526 , n84524 , n84525 );
and ( n84527 , n84526 , n32398 );
and ( n84528 , n46023 , n32436 );
or ( n84529 , n84522 , n84527 , n84528 );
and ( n84530 , n84529 , n32456 );
and ( n84531 , n49663 , n32473 );
not ( n84532 , n32475 );
and ( n84533 , n84532 , n49663 );
xor ( n84534 , n46023 , n47763 );
and ( n84535 , n84534 , n32475 );
or ( n84536 , n84533 , n84535 );
and ( n84537 , n84536 , n32486 );
and ( n84538 , n37543 , n32489 );
and ( n84539 , n46023 , n32501 );
or ( n84540 , C0 , n84530 , n84531 , n84537 , n84538 , n84539 );
buf ( n84541 , n84540 );
buf ( n84542 , n84541 );
and ( n84543 , n33227 , n32528 );
not ( n84544 , n32598 );
and ( n84545 , n84544 , n32990 );
buf ( n84546 , n84545 );
and ( n84547 , n84546 , n32890 );
not ( n84548 , n32919 );
and ( n84549 , n84548 , n32990 );
buf ( n84550 , n84549 );
and ( n84551 , n84550 , n32924 );
not ( n84552 , n32953 );
and ( n84553 , n84552 , n32990 );
not ( n84554 , n32971 );
and ( n84555 , n84554 , n33105 );
xor ( n84556 , n32990 , n33015 );
and ( n84557 , n84556 , n32971 );
or ( n84558 , n84555 , n84557 );
and ( n84559 , n84558 , n32953 );
or ( n84560 , n84553 , n84559 );
and ( n84561 , n84560 , n33038 );
not ( n84562 , n33067 );
and ( n84563 , n84562 , n32990 );
not ( n84564 , n32970 );
not ( n84565 , n33071 );
and ( n84566 , n84565 , n33105 );
xor ( n84567 , n33106 , n33147 );
and ( n84568 , n84567 , n33071 );
or ( n84569 , n84566 , n84568 );
and ( n84570 , n84564 , n84569 );
and ( n84571 , n84556 , n32970 );
or ( n84572 , n84570 , n84571 );
and ( n84573 , n84572 , n33067 );
or ( n84574 , n84563 , n84573 );
and ( n84575 , n84574 , n33172 );
and ( n84576 , n32990 , n33204 );
or ( n84577 , n84547 , n84551 , n84561 , n84575 , n84576 );
and ( n84578 , n84577 , n33208 );
not ( n84579 , n32968 );
not ( n84580 , n33270 );
and ( n84581 , n84580 , n33305 );
xor ( n84582 , n33306 , n33347 );
and ( n84583 , n84582 , n33270 );
or ( n84584 , n84581 , n84583 );
and ( n84585 , n84579 , n84584 );
and ( n84586 , n32990 , n32968 );
or ( n84587 , n84585 , n84586 );
and ( n84588 , n84587 , n33370 );
buf ( n84589 , n35056 );
and ( n84590 , n32990 , n33382 );
or ( n84591 , C0 , n84543 , n84578 , n84588 , n84589 , n84590 );
buf ( n84592 , n84591 );
buf ( n84593 , n84592 );
buf ( n84594 , n30987 );
buf ( n84595 , n31655 );
buf ( n84596 , n30987 );
not ( n84597 , n45274 );
and ( n84598 , n84597 , n35534 );
buf ( n84599 , n84598 );
and ( n84600 , n84599 , n31373 );
not ( n84601 , n45280 );
and ( n84602 , n84601 , n35534 );
buf ( n84603 , n84602 );
and ( n84604 , n84603 , n31468 );
and ( n84605 , n35534 , n45802 );
or ( n84606 , n84600 , n84604 , n84605 );
and ( n84607 , n84606 , n31557 );
and ( n84608 , n35534 , n45808 );
or ( n84609 , C0 , C0 , n84607 , n84608 );
buf ( n84610 , n84609 );
buf ( n84611 , n84610 );
not ( n84612 , n40163 );
and ( n84613 , n84612 , n31793 );
not ( n84614 , n52903 );
and ( n84615 , n84614 , n31793 );
and ( n84616 , n32252 , n52903 );
or ( n84617 , n84615 , n84616 );
and ( n84618 , n84617 , n40163 );
or ( n84619 , n84613 , n84618 );
and ( n84620 , n84619 , n32498 );
not ( n84621 , n52911 );
not ( n84622 , n52903 );
and ( n84623 , n84622 , n31793 );
and ( n84624 , n40393 , n52903 );
or ( n84625 , n84623 , n84624 );
and ( n84626 , n84621 , n84625 );
and ( n84627 , n40393 , n52911 );
or ( n84628 , n84626 , n84627 );
and ( n84629 , n84628 , n32473 );
not ( n84630 , n32475 );
not ( n84631 , n52911 );
not ( n84632 , n52903 );
and ( n84633 , n84632 , n31793 );
and ( n84634 , n40393 , n52903 );
or ( n84635 , n84633 , n84634 );
and ( n84636 , n84631 , n84635 );
and ( n84637 , n40393 , n52911 );
or ( n84638 , n84636 , n84637 );
and ( n84639 , n84630 , n84638 );
not ( n84640 , n52931 );
not ( n84641 , n52933 );
and ( n84642 , n84641 , n84638 );
and ( n84643 , n40972 , n52933 );
or ( n84644 , n84642 , n84643 );
and ( n84645 , n84640 , n84644 );
and ( n84646 , n41267 , n52931 );
or ( n84647 , n84645 , n84646 );
and ( n84648 , n84647 , n32475 );
or ( n84649 , n84639 , n84648 );
and ( n84650 , n84649 , n32486 );
and ( n84651 , n31793 , n41278 );
or ( n84652 , C0 , n84620 , n84629 , n84650 , n84651 );
buf ( n84653 , n84652 );
buf ( n84654 , n84653 );
not ( n84655 , n43755 );
and ( n84656 , n84655 , n43649 );
xor ( n84657 , n52304 , n52325 );
and ( n84658 , n84657 , n43755 );
or ( n84659 , n84656 , n84658 );
and ( n84660 , n84659 , n43774 );
not ( n84661 , n44663 );
and ( n84662 , n84661 , n44561 );
xor ( n84663 , n52342 , n52363 );
and ( n84664 , n84663 , n44663 );
or ( n84665 , n84662 , n84664 );
and ( n84666 , n84665 , n44682 );
and ( n84667 , n73635 , n44695 );
or ( n84668 , n84660 , n84666 , n84667 );
buf ( n84669 , n84668 );
buf ( n84670 , n84669 );
buf ( n84671 , n30987 );
buf ( n84672 , n31655 );
buf ( n84673 , n31655 );
buf ( n84674 , n30987 );
buf ( n84675 , n30987 );
buf ( n84676 , n31655 );
buf ( n84677 , n31655 );
buf ( n84678 , n30987 );
not ( n84679 , n32953 );
and ( n84680 , n84679 , n80800 );
and ( n84681 , n80814 , n32953 );
or ( n84682 , n84680 , n84681 );
and ( n84683 , n84682 , n33038 );
not ( n84684 , n48660 );
and ( n84685 , n84684 , n80800 );
and ( n84686 , n79824 , n48660 );
or ( n84687 , n84685 , n84686 );
and ( n84688 , n84687 , n33172 );
and ( n84689 , n80800 , n39795 );
or ( n84690 , n84683 , n84688 , n84689 );
and ( n84691 , n84690 , n33208 );
and ( n84692 , n80800 , n39805 );
or ( n84693 , C0 , n84691 , n84692 );
buf ( n84694 , n84693 );
buf ( n84695 , n84694 );
buf ( n84696 , n30987 );
buf ( n84697 , n31655 );
not ( n84698 , n31437 );
and ( n84699 , n84698 , n66042 );
and ( n84700 , n66054 , n31437 );
or ( n84701 , n84699 , n84700 );
and ( n84702 , n84701 , n31468 );
not ( n84703 , n44817 );
and ( n84704 , n84703 , n66042 );
and ( n84705 , n82943 , n44817 );
or ( n84706 , n84704 , n84705 );
and ( n84707 , n84706 , n31521 );
and ( n84708 , n66042 , n42158 );
or ( n84709 , n84702 , n84707 , n84708 );
and ( n84710 , n84709 , n31557 );
and ( n84711 , n66042 , n40154 );
or ( n84712 , C0 , n84710 , n84711 );
buf ( n84713 , n84712 );
buf ( n84714 , n84713 );
and ( n84715 , n47667 , n50275 );
not ( n84716 , n50278 );
and ( n84717 , n84716 , n47580 );
and ( n84718 , n47667 , n50278 );
or ( n84719 , n84717 , n84718 );
and ( n84720 , n84719 , n32421 );
not ( n84721 , n50002 );
and ( n84722 , n84721 , n47580 );
and ( n84723 , n47667 , n50002 );
or ( n84724 , n84722 , n84723 );
and ( n84725 , n84724 , n32419 );
not ( n84726 , n50289 );
and ( n84727 , n84726 , n47580 );
and ( n84728 , n47667 , n50289 );
or ( n84729 , n84727 , n84728 );
and ( n84730 , n84729 , n32417 );
not ( n84731 , n50008 );
and ( n84732 , n84731 , n47580 );
and ( n84733 , n47667 , n50008 );
or ( n84734 , n84732 , n84733 );
and ( n84735 , n84734 , n32415 );
not ( n84736 , n47331 );
and ( n84737 , n84736 , n47580 );
and ( n84738 , n47612 , n47331 );
or ( n84739 , n84737 , n84738 );
and ( n84740 , n84739 , n32413 );
not ( n84741 , n50067 );
and ( n84742 , n84741 , n47580 );
and ( n84743 , n47612 , n50067 );
or ( n84744 , n84742 , n84743 );
and ( n84745 , n84744 , n32411 );
not ( n84746 , n31728 );
and ( n84747 , n84746 , n47580 );
and ( n84748 , n60771 , n31728 );
or ( n84749 , n84747 , n84748 );
and ( n84750 , n84749 , n32253 );
not ( n84751 , n32283 );
and ( n84752 , n84751 , n47580 );
and ( n84753 , n60782 , n32283 );
or ( n84754 , n84752 , n84753 );
and ( n84755 , n84754 , n32398 );
and ( n84756 , n47717 , n50334 );
or ( n84757 , n84715 , n84720 , n84725 , n84730 , n84735 , n84740 , n84745 , n84750 , n84755 , n84756 );
and ( n84758 , n84757 , n32456 );
and ( n84759 , n37567 , n32489 );
and ( n84760 , n47580 , n50345 );
or ( n84761 , C0 , n84758 , n84759 , n84760 );
buf ( n84762 , n84761 );
buf ( n84763 , n84762 );
buf ( n84764 , n31655 );
buf ( n84765 , n30987 );
buf ( n84766 , n30987 );
buf ( n84767 , n31655 );
and ( n84768 , n56473 , n81346 );
xor ( n84769 , n56471 , n84768 );
and ( n84770 , n84769 , n48639 );
not ( n84771 , n48642 );
and ( n84772 , n84771 , n56471 );
and ( n84773 , n84769 , n48642 );
or ( n84774 , n84772 , n84773 );
and ( n84775 , n84774 , n32890 );
not ( n84776 , n48648 );
and ( n84777 , n84776 , n56471 );
and ( n84778 , n84769 , n48648 );
or ( n84779 , n84777 , n84778 );
and ( n84780 , n84779 , n32924 );
not ( n84781 , n48654 );
and ( n84782 , n84781 , n56471 );
and ( n84783 , n84769 , n48654 );
or ( n84784 , n84782 , n84783 );
and ( n84785 , n84784 , n33038 );
not ( n84786 , n48660 );
and ( n84787 , n84786 , n56471 );
and ( n84788 , n84769 , n48660 );
or ( n84789 , n84787 , n84788 );
and ( n84790 , n84789 , n33172 );
not ( n84791 , n41576 );
and ( n84792 , n84791 , n56471 );
and ( n84793 , n56473 , n81336 );
xor ( n84794 , n56471 , n84793 );
and ( n84795 , n84794 , n41576 );
or ( n84796 , n84792 , n84795 );
and ( n84797 , n84796 , n33189 );
not ( n84798 , n48730 );
and ( n84799 , n84798 , n56471 );
and ( n84800 , n84794 , n48730 );
or ( n84801 , n84799 , n84800 );
and ( n84802 , n84801 , n33187 );
not ( n84803 , n48765 );
and ( n84804 , n84803 , n56471 );
and ( n84805 , n81337 , n81338 );
xor ( n84806 , n84794 , n84805 );
and ( n84807 , n84806 , n48765 );
or ( n84808 , n84804 , n84807 );
and ( n84809 , n84808 , n33180 );
not ( n84810 , n49054 );
and ( n84811 , n84810 , n56471 );
not ( n84812 , n48845 );
and ( n84813 , n81347 , n81348 );
xor ( n84814 , n84769 , n84813 );
and ( n84815 , n84812 , n84814 );
and ( n84816 , n56473 , n81351 );
xor ( n84817 , n56471 , n84816 );
or ( n84818 , n81352 , n81353 );
xnor ( n84819 , n84817 , n84818 );
and ( n84820 , n84819 , n48845 );
or ( n84821 , n84815 , n84820 );
and ( n84822 , n84821 , n49054 );
or ( n84823 , n84811 , n84822 );
and ( n84824 , n84823 , n33178 );
and ( n84825 , n84817 , n49275 );
or ( n84826 , n84770 , n84775 , n84780 , n84785 , n84790 , n84797 , n84802 , n84809 , n84824 , n84825 );
and ( n84827 , n84826 , n33208 );
and ( n84828 , n35592 , n35056 );
and ( n84829 , n56471 , n49286 );
or ( n84830 , C0 , n84827 , n84828 , n84829 );
buf ( n84831 , n84830 );
buf ( n84832 , n84831 );
buf ( n84833 , n31655 );
buf ( n84834 , n30987 );
not ( n84835 , n33133 );
and ( n84836 , n84835 , n33201 );
not ( n84837 , n41576 );
and ( n84838 , n84837 , n33133 );
buf ( n84839 , n32652 );
and ( n84840 , n84839 , n41576 );
or ( n84841 , n84838 , n84840 );
and ( n84842 , n84841 , n33189 );
and ( n84843 , n33133 , n41592 );
or ( n84844 , n84836 , n84842 , n84843 );
and ( n84845 , n84844 , n33208 );
and ( n84846 , n33133 , n39805 );
or ( n84847 , C0 , n84845 , n84846 );
buf ( n84848 , n84847 );
buf ( n84849 , n84848 );
buf ( n84850 , n30987 );
buf ( n84851 , n31655 );
not ( n84852 , n41532 );
and ( n84853 , n84852 , n34260 );
and ( n84854 , n65190 , n41532 );
or ( n84855 , n84853 , n84854 );
buf ( n84856 , n84855 );
buf ( n84857 , n84856 );
buf ( n84858 , n31655 );
buf ( n84859 , n30987 );
and ( n84860 , n42610 , n33377 );
not ( n84861 , n48545 );
buf ( n84862 , RI15b47580_299);
and ( n84863 , n84861 , n84862 );
and ( n84864 , n42642 , n48545 );
or ( n84865 , n84863 , n84864 );
and ( n84866 , n84865 , n32890 );
not ( n84867 , n48557 );
and ( n84868 , n84867 , n84862 );
and ( n84869 , n42642 , n48557 );
or ( n84870 , n84868 , n84869 );
and ( n84871 , n84870 , n33038 );
and ( n84872 , n84862 , n48571 );
or ( n84873 , n84866 , n84871 , n84872 );
and ( n84874 , n84873 , n33208 );
and ( n84875 , n84862 , n48577 );
or ( n84876 , C0 , n84860 , n84874 , n84875 );
buf ( n84877 , n84876 );
buf ( n84878 , n84877 );
buf ( n84879 , n30987 );
buf ( n84880 , n31655 );
buf ( n84881 , n30987 );
xor ( n84882 , n41717 , n44784 );
and ( n84883 , n84882 , n31548 );
not ( n84884 , n44807 );
and ( n84885 , n84884 , n41717 );
and ( n84886 , n42014 , n44807 );
or ( n84887 , n84885 , n84886 );
and ( n84888 , n84887 , n31408 );
not ( n84889 , n44817 );
and ( n84890 , n84889 , n41717 );
not ( n84891 , n41835 );
buf ( n84892 , RI15b53010_697);
and ( n84893 , n84891 , n84892 );
not ( n84894 , n42124 );
and ( n84895 , n84894 , n42024 );
xor ( n84896 , n49379 , n49380 );
and ( n84897 , n84896 , n42124 );
or ( n84898 , n84895 , n84897 );
and ( n84899 , n84898 , n41835 );
or ( n84900 , n84893 , n84899 );
and ( n84901 , n84900 , n44817 );
or ( n84902 , n84890 , n84901 );
and ( n84903 , n84902 , n31521 );
not ( n84904 , n45059 );
and ( n84905 , n84904 , n41717 );
and ( n84906 , n69086 , n45059 );
or ( n84907 , n84905 , n84906 );
and ( n84908 , n84907 , n31536 );
and ( n84909 , n41717 , n45148 );
or ( n84910 , n84883 , n84888 , n84903 , n84908 , n84909 );
and ( n84911 , n84910 , n31557 );
and ( n84912 , n41717 , n40154 );
or ( n84913 , C0 , n84911 , n84912 );
buf ( n84914 , n84913 );
buf ( n84915 , n84914 );
buf ( n84916 , n31655 );
not ( n84917 , n40163 );
and ( n84918 , n84917 , n31802 );
not ( n84919 , n49298 );
and ( n84920 , n84919 , n31802 );
and ( n84921 , n32252 , n49298 );
or ( n84922 , n84920 , n84921 );
and ( n84923 , n84922 , n40163 );
or ( n84924 , n84918 , n84923 );
and ( n84925 , n84924 , n32498 );
not ( n84926 , n49306 );
not ( n84927 , n49298 );
and ( n84928 , n84927 , n31802 );
and ( n84929 , n40393 , n49298 );
or ( n84930 , n84928 , n84929 );
and ( n84931 , n84926 , n84930 );
and ( n84932 , n40393 , n49306 );
or ( n84933 , n84931 , n84932 );
and ( n84934 , n84933 , n32473 );
not ( n84935 , n32475 );
not ( n84936 , n49306 );
not ( n84937 , n49298 );
and ( n84938 , n84937 , n31802 );
and ( n84939 , n40393 , n49298 );
or ( n84940 , n84938 , n84939 );
and ( n84941 , n84936 , n84940 );
and ( n84942 , n40393 , n49306 );
or ( n84943 , n84941 , n84942 );
and ( n84944 , n84935 , n84943 );
not ( n84945 , n49331 );
not ( n84946 , n49333 );
and ( n84947 , n84946 , n84943 );
and ( n84948 , n40972 , n49333 );
or ( n84949 , n84947 , n84948 );
and ( n84950 , n84945 , n84949 );
and ( n84951 , n41267 , n49331 );
or ( n84952 , n84950 , n84951 );
and ( n84953 , n84952 , n32475 );
or ( n84954 , n84944 , n84953 );
and ( n84955 , n84954 , n32486 );
and ( n84956 , n31802 , n41278 );
or ( n84957 , C0 , n84925 , n84934 , n84955 , n84956 );
buf ( n84958 , n84957 );
buf ( n84959 , n84958 );
buf ( n84960 , n30987 );
buf ( n84961 , n31655 );
and ( n84962 , n63843 , n31557 );
and ( n84963 , n63812 , n40154 );
or ( n84964 , C0 , n84962 , n84963 );
buf ( n84965 , n84964 );
buf ( n84966 , n84965 );
buf ( n84967 , n30987 );
not ( n84968 , n38443 );
and ( n84969 , n84968 , n38116 );
xor ( n84970 , n53475 , n53494 );
and ( n84971 , n84970 , n38443 );
or ( n84972 , n84969 , n84971 );
and ( n84973 , n84972 , n38450 );
not ( n84974 , n39339 );
and ( n84975 , n84974 , n39016 );
xor ( n84976 , n53531 , n53550 );
and ( n84977 , n84976 , n39339 );
or ( n84978 , n84975 , n84977 );
and ( n84979 , n84978 , n39346 );
and ( n84980 , n40209 , n39359 );
or ( n84981 , n84973 , n84979 , n84980 );
buf ( n84982 , n84981 );
buf ( n84983 , n84982 );
buf ( n84984 , n31655 );
not ( n84985 , n46356 );
and ( n84986 , n84985 , n31315 );
not ( n84987 , n78324 );
and ( n84988 , n84987 , n31315 );
and ( n84989 , n31339 , n78324 );
or ( n84990 , n84988 , n84989 );
and ( n84991 , n84990 , n46356 );
or ( n84992 , n84986 , n84991 );
and ( n84993 , n84992 , n31649 );
not ( n84994 , n78332 );
not ( n84995 , n78324 );
and ( n84996 , n84995 , n31315 );
and ( n84997 , n47449 , n78324 );
or ( n84998 , n84996 , n84997 );
and ( n84999 , n84994 , n84998 );
and ( n85000 , n47449 , n78332 );
or ( n85001 , n84999 , n85000 );
and ( n85002 , n85001 , n31643 );
not ( n85003 , n31452 );
not ( n85004 , n78332 );
not ( n85005 , n78324 );
and ( n85006 , n85005 , n31315 );
and ( n85007 , n47449 , n78324 );
or ( n85008 , n85006 , n85007 );
and ( n85009 , n85004 , n85008 );
and ( n85010 , n47449 , n78332 );
or ( n85011 , n85009 , n85010 );
and ( n85012 , n85003 , n85011 );
not ( n85013 , n78352 );
not ( n85014 , n78354 );
and ( n85015 , n85014 , n85011 );
and ( n85016 , n47485 , n78354 );
or ( n85017 , n85015 , n85016 );
and ( n85018 , n85013 , n85017 );
and ( n85019 , n47503 , n78352 );
or ( n85020 , n85018 , n85019 );
and ( n85021 , n85020 , n31452 );
or ( n85022 , n85012 , n85021 );
and ( n85023 , n85022 , n31638 );
and ( n85024 , n31315 , n47277 );
or ( n85025 , C0 , n84993 , n85002 , n85023 , n85024 );
buf ( n85026 , n85025 );
buf ( n85027 , n85026 );
buf ( n85028 , n30987 );
buf ( n85029 , RI15b5e938_1092);
and ( n85030 , n85029 , n32494 );
not ( n85031 , n46083 );
and ( n85032 , n85031 , n66716 );
xor ( n85033 , n46286 , n46092 );
and ( n85034 , n72078 , n72079 );
and ( n85035 , n85033 , n85034 );
buf ( n85036 , n85035 );
and ( n85037 , n85036 , n46290 );
buf ( n85038 , n85037 );
and ( n85039 , n85038 , n46083 );
or ( n85040 , n85032 , n85039 );
and ( n85041 , n85040 , n32421 );
not ( n85042 , n46326 );
and ( n85043 , n85042 , n66716 );
not ( n85044 , n51396 );
and ( n85045 , n85044 , n50945 );
xor ( n85046 , n51405 , n51155 );
and ( n85047 , n85046 , n51396 );
or ( n85048 , n85045 , n85047 );
and ( n85049 , n85048 , n46326 );
or ( n85050 , n85043 , n85049 );
and ( n85051 , n85050 , n32417 );
and ( n85052 , n66716 , n46340 );
or ( n85053 , n85041 , n85051 , n85052 );
and ( n85054 , n85053 , n32456 );
and ( n85055 , n66716 , n46349 );
or ( n85056 , C0 , n85030 , n85054 , n85055 );
buf ( n85057 , n85056 );
buf ( n85058 , n85057 );
buf ( n85059 , n31655 );
and ( n85060 , n49060 , n48639 );
not ( n85061 , n48642 );
and ( n85062 , n85061 , n48585 );
and ( n85063 , n49060 , n48642 );
or ( n85064 , n85062 , n85063 );
and ( n85065 , n85064 , n32890 );
not ( n85066 , n48648 );
and ( n85067 , n85066 , n48585 );
and ( n85068 , n49060 , n48648 );
or ( n85069 , n85067 , n85068 );
and ( n85070 , n85069 , n32924 );
not ( n85071 , n48654 );
and ( n85072 , n85071 , n48585 );
and ( n85073 , n49060 , n48654 );
or ( n85074 , n85072 , n85073 );
and ( n85075 , n85074 , n33038 );
not ( n85076 , n48660 );
and ( n85077 , n85076 , n48585 );
and ( n85078 , n49060 , n48660 );
or ( n85079 , n85077 , n85078 );
and ( n85080 , n85079 , n33172 );
not ( n85081 , n41576 );
and ( n85082 , n85081 , n48585 );
and ( n85083 , n48770 , n41576 );
or ( n85084 , n85082 , n85083 );
and ( n85085 , n85084 , n33189 );
not ( n85086 , n48730 );
and ( n85087 , n85086 , n48585 );
and ( n85088 , n48770 , n48730 );
or ( n85089 , n85087 , n85088 );
and ( n85090 , n85089 , n33187 );
not ( n85091 , n48765 );
and ( n85092 , n85091 , n48585 );
and ( n85093 , n71977 , n48765 );
or ( n85094 , n85092 , n85093 );
and ( n85095 , n85094 , n33180 );
not ( n85096 , n49054 );
and ( n85097 , n85096 , n48585 );
and ( n85098 , n71988 , n49054 );
or ( n85099 , n85097 , n85098 );
and ( n85100 , n85099 , n33178 );
and ( n85101 , n49169 , n49275 );
or ( n85102 , n85060 , n85065 , n85070 , n85075 , n85080 , n85085 , n85090 , n85095 , n85100 , n85101 );
and ( n85103 , n85102 , n33208 );
and ( n85104 , n32978 , n35056 );
and ( n85105 , n48585 , n49286 );
or ( n85106 , C0 , n85103 , n85104 , n85105 );
buf ( n85107 , n85106 );
buf ( n85108 , n85107 );
buf ( n85109 , n30987 );
buf ( n85110 , n30987 );
buf ( n85111 , n31655 );
buf ( n85112 , n31655 );
buf ( n85113 , n30987 );
buf ( n85114 , n31655 );
not ( n85115 , n48545 );
and ( n85116 , n85115 , n35539 );
buf ( n85117 , n85116 );
and ( n85118 , n85117 , n32890 );
not ( n85119 , n48557 );
and ( n85120 , n85119 , n35539 );
buf ( n85121 , n85120 );
and ( n85122 , n85121 , n33038 );
and ( n85123 , n35539 , n48571 );
or ( n85124 , n85118 , n85122 , n85123 );
and ( n85125 , n85124 , n33208 );
and ( n85126 , n35539 , n48577 );
or ( n85127 , C0 , C0 , n85125 , n85126 );
buf ( n85128 , n85127 );
buf ( n85129 , n85128 );
buf ( n85130 , n30987 );
buf ( n85131 , n31655 );
buf ( n85132 , n30987 );
not ( n85133 , n34150 );
and ( n85134 , n85133 , n32534 );
and ( n85135 , n34183 , n34150 );
or ( n85136 , n85134 , n85135 );
and ( n85137 , n85136 , n33381 );
not ( n85138 , n56687 );
not ( n85139 , n56464 );
and ( n85140 , n85139 , n32534 );
buf ( n85141 , n85140 );
and ( n85142 , n85138 , n85141 );
buf ( n85143 , n85142 );
and ( n85144 , n85143 , n33379 );
and ( n85145 , n34349 , n33375 );
not ( n85146 , n32968 );
and ( n85147 , n85146 , n34349 );
and ( n85148 , n34344 , n59867 );
xor ( n85149 , n34354 , n85148 );
not ( n85150 , n85149 );
buf ( n85151 , n85150 );
not ( n85152 , n85151 );
and ( n85153 , n85152 , n32968 );
or ( n85154 , n85147 , n85153 );
and ( n85155 , n85154 , n33370 );
and ( n85156 , n32534 , n56699 );
or ( n85157 , C0 , n85137 , n85144 , n85145 , n85155 , n85156 );
buf ( n85158 , n85157 );
buf ( n85159 , n85158 );
not ( n85160 , n34150 );
and ( n85161 , n85160 , n32677 );
not ( n85162 , n56413 );
and ( n85163 , n85162 , n32677 );
and ( n85164 , n32689 , n56413 );
or ( n85165 , n85163 , n85164 );
and ( n85166 , n85165 , n34150 );
or ( n85167 , n85161 , n85166 );
and ( n85168 , n85167 , n33381 );
not ( n85169 , n56421 );
not ( n85170 , n56413 );
and ( n85171 , n85170 , n32677 );
and ( n85172 , n50682 , n56413 );
or ( n85173 , n85171 , n85172 );
and ( n85174 , n85169 , n85173 );
and ( n85175 , n50682 , n56421 );
or ( n85176 , n85174 , n85175 );
and ( n85177 , n85176 , n33375 );
not ( n85178 , n32968 );
not ( n85179 , n56421 );
not ( n85180 , n56413 );
and ( n85181 , n85180 , n32677 );
and ( n85182 , n50682 , n56413 );
or ( n85183 , n85181 , n85182 );
and ( n85184 , n85179 , n85183 );
and ( n85185 , n50682 , n56421 );
or ( n85186 , n85184 , n85185 );
and ( n85187 , n85178 , n85186 );
not ( n85188 , n56441 );
not ( n85189 , n56443 );
and ( n85190 , n85189 , n85186 );
and ( n85191 , n50706 , n56443 );
or ( n85192 , n85190 , n85191 );
and ( n85193 , n85188 , n85192 );
and ( n85194 , n50714 , n56441 );
or ( n85195 , n85193 , n85194 );
and ( n85196 , n85195 , n32968 );
or ( n85197 , n85187 , n85196 );
and ( n85198 , n85197 , n33370 );
and ( n85199 , n32677 , n35062 );
or ( n85200 , C0 , n85168 , n85177 , n85198 , n85199 );
buf ( n85201 , n85200 );
buf ( n85202 , n85201 );
buf ( n85203 , n30987 );
buf ( n85204 , n31655 );
buf ( n85205 , n31655 );
buf ( n85206 , n30987 );
buf ( n85207 , n54731 );
not ( n85208 , n34150 );
and ( n85209 , n85208 , n32877 );
not ( n85210 , n56413 );
and ( n85211 , n85210 , n32877 );
and ( n85212 , n32889 , n56413 );
or ( n85213 , n85211 , n85212 );
and ( n85214 , n85213 , n34150 );
or ( n85215 , n85209 , n85214 );
and ( n85216 , n85215 , n33381 );
not ( n85217 , n56421 );
not ( n85218 , n56413 );
and ( n85219 , n85218 , n32877 );
and ( n85220 , n52819 , n56413 );
or ( n85221 , n85219 , n85220 );
and ( n85222 , n85217 , n85221 );
and ( n85223 , n52819 , n56421 );
or ( n85224 , n85222 , n85223 );
and ( n85225 , n85224 , n33375 );
not ( n85226 , n32968 );
not ( n85227 , n56421 );
not ( n85228 , n56413 );
and ( n85229 , n85228 , n32877 );
and ( n85230 , n52819 , n56413 );
or ( n85231 , n85229 , n85230 );
and ( n85232 , n85227 , n85231 );
and ( n85233 , n52819 , n56421 );
or ( n85234 , n85232 , n85233 );
and ( n85235 , n85226 , n85234 );
not ( n85236 , n56441 );
not ( n85237 , n56443 );
and ( n85238 , n85237 , n85234 );
and ( n85239 , n52845 , n56443 );
or ( n85240 , n85238 , n85239 );
and ( n85241 , n85236 , n85240 );
and ( n85242 , n52855 , n56441 );
or ( n85243 , n85241 , n85242 );
and ( n85244 , n85243 , n32968 );
or ( n85245 , n85235 , n85244 );
and ( n85246 , n85245 , n33370 );
and ( n85247 , n32877 , n35062 );
or ( n85248 , C0 , n85216 , n85225 , n85246 , n85247 );
buf ( n85249 , n85248 );
buf ( n85250 , n85249 );
buf ( n85251 , n30987 );
buf ( n85252 , n31655 );
buf ( n85253 , n31655 );
not ( n85254 , n46356 );
and ( n85255 , n85254 , n31321 );
not ( n85256 , n48214 );
and ( n85257 , n85256 , n31321 );
and ( n85258 , n31339 , n48214 );
or ( n85259 , n85257 , n85258 );
and ( n85260 , n85259 , n46356 );
or ( n85261 , n85255 , n85260 );
and ( n85262 , n85261 , n31649 );
not ( n85263 , n48223 );
not ( n85264 , n48214 );
and ( n85265 , n85264 , n31321 );
and ( n85266 , n47449 , n48214 );
or ( n85267 , n85265 , n85266 );
and ( n85268 , n85263 , n85267 );
and ( n85269 , n47449 , n48223 );
or ( n85270 , n85268 , n85269 );
and ( n85271 , n85270 , n31643 );
not ( n85272 , n31452 );
not ( n85273 , n48223 );
not ( n85274 , n48214 );
and ( n85275 , n85274 , n31321 );
and ( n85276 , n47449 , n48214 );
or ( n85277 , n85275 , n85276 );
and ( n85278 , n85273 , n85277 );
and ( n85279 , n47449 , n48223 );
or ( n85280 , n85278 , n85279 );
and ( n85281 , n85272 , n85280 );
not ( n85282 , n48244 );
not ( n85283 , n48247 );
and ( n85284 , n85283 , n85280 );
and ( n85285 , n47485 , n48247 );
or ( n85286 , n85284 , n85285 );
and ( n85287 , n85282 , n85286 );
and ( n85288 , n47503 , n48244 );
or ( n85289 , n85287 , n85288 );
and ( n85290 , n85289 , n31452 );
or ( n85291 , n85281 , n85290 );
and ( n85292 , n85291 , n31638 );
and ( n85293 , n31321 , n47277 );
or ( n85294 , C0 , n85262 , n85271 , n85292 , n85293 );
buf ( n85295 , n85294 );
buf ( n85296 , n85295 );
buf ( n85297 , n31655 );
buf ( n85298 , n30987 );
buf ( n85299 , n67704 );
buf ( n85300 , n67668 );
or ( n85301 , C0 , C0 , C0 , n85299 , n85300 );
and ( n85302 , n85301 , n67701 );
buf ( n85303 , n79276 );
buf ( n85304 , n67704 );
buf ( n85305 , n67668 );
or ( n85306 , C0 , C0 , n85303 , n85304 , n85305 );
and ( n85307 , n85306 , n67737 );
or ( n85308 , C0 , C0 , n85302 , n85307 );
buf ( n85309 , n85308 );
buf ( n85310 , n85309 );
buf ( n85311 , n31655 );
buf ( n85312 , n31655 );
xor ( n85313 , n44772 , n44795 );
and ( n85314 , n85313 , n31548 );
not ( n85315 , n44807 );
and ( n85316 , n85315 , n44772 );
and ( n85317 , n46657 , n44807 );
or ( n85318 , n85316 , n85317 );
and ( n85319 , n85318 , n31408 );
not ( n85320 , n44817 );
and ( n85321 , n85320 , n44772 );
and ( n85322 , n51741 , n44817 );
or ( n85323 , n85321 , n85322 );
and ( n85324 , n85323 , n31521 );
not ( n85325 , n45059 );
and ( n85326 , n85325 , n44772 );
and ( n85327 , n78002 , n45059 );
or ( n85328 , n85326 , n85327 );
and ( n85329 , n85328 , n31536 );
and ( n85330 , n44772 , n45148 );
or ( n85331 , n85314 , n85319 , n85324 , n85329 , n85330 );
and ( n85332 , n85331 , n31557 );
and ( n85333 , n44772 , n40154 );
or ( n85334 , C0 , n85332 , n85333 );
buf ( n85335 , n85334 );
buf ( n85336 , n85335 );
not ( n85337 , n40163 );
and ( n85338 , n85337 , n31916 );
not ( n85339 , n55888 );
and ( n85340 , n85339 , n31916 );
and ( n85341 , n32200 , n55888 );
or ( n85342 , n85340 , n85341 );
and ( n85343 , n85342 , n40163 );
or ( n85344 , n85338 , n85343 );
and ( n85345 , n85344 , n32498 );
not ( n85346 , n55896 );
not ( n85347 , n55888 );
and ( n85348 , n85347 , n31916 );
and ( n85349 , n53243 , n55888 );
or ( n85350 , n85348 , n85349 );
and ( n85351 , n85346 , n85350 );
and ( n85352 , n53243 , n55896 );
or ( n85353 , n85351 , n85352 );
and ( n85354 , n85353 , n32473 );
not ( n85355 , n32475 );
not ( n85356 , n55896 );
not ( n85357 , n55888 );
and ( n85358 , n85357 , n31916 );
and ( n85359 , n53243 , n55888 );
or ( n85360 , n85358 , n85359 );
and ( n85361 , n85356 , n85360 );
and ( n85362 , n53243 , n55896 );
or ( n85363 , n85361 , n85362 );
and ( n85364 , n85355 , n85363 );
not ( n85365 , n55916 );
not ( n85366 , n55918 );
and ( n85367 , n85366 , n85363 );
and ( n85368 , n53269 , n55918 );
or ( n85369 , n85367 , n85368 );
and ( n85370 , n85365 , n85369 );
and ( n85371 , n53277 , n55916 );
or ( n85372 , n85370 , n85371 );
and ( n85373 , n85372 , n32475 );
or ( n85374 , n85364 , n85373 );
and ( n85375 , n85374 , n32486 );
and ( n85376 , n31916 , n41278 );
or ( n85377 , C0 , n85345 , n85354 , n85375 , n85376 );
buf ( n85378 , n85377 );
buf ( n85379 , n85378 );
buf ( n85380 , n30987 );
buf ( n85381 , n30987 );
buf ( n85382 , n31655 );
buf ( n85383 , n31655 );
not ( n85384 , n33419 );
and ( n85385 , n85384 , n31569 );
and ( n85386 , n53433 , n33419 );
or ( n85387 , n85385 , n85386 );
and ( n85388 , n85387 , n31529 );
not ( n85389 , n33734 );
and ( n85390 , n85389 , n31569 );
and ( n85391 , n53444 , n33734 );
or ( n85392 , n85390 , n85391 );
and ( n85393 , n85392 , n31527 );
and ( n85394 , n31569 , n33942 );
or ( n85395 , n85388 , n85393 , n85394 );
and ( n85396 , n85395 , n31557 );
and ( n85397 , n35494 , n31643 );
not ( n85398 , n31452 );
and ( n85399 , n85398 , n35494 );
xor ( n85400 , n31569 , n42437 );
and ( n85401 , n85400 , n31452 );
or ( n85402 , n85399 , n85401 );
and ( n85403 , n85402 , n31638 );
and ( n85404 , n35395 , n33973 );
and ( n85405 , n31569 , n33978 );
or ( n85406 , C0 , n85396 , n85397 , n85403 , n85404 , n85405 );
buf ( n85407 , n85406 );
buf ( n85408 , n85407 );
and ( n85409 , n31575 , n31007 );
not ( n85410 , n31077 );
and ( n85411 , n85410 , n33999 );
buf ( n85412 , n85411 );
and ( n85413 , n85412 , n31373 );
not ( n85414 , n31402 );
and ( n85415 , n85414 , n33999 );
buf ( n85416 , n85415 );
and ( n85417 , n85416 , n31408 );
not ( n85418 , n31437 );
and ( n85419 , n85418 , n33999 );
not ( n85420 , n31455 );
and ( n85421 , n85420 , n34038 );
xor ( n85422 , n33999 , n34024 );
and ( n85423 , n85422 , n31455 );
or ( n85424 , n85421 , n85423 );
and ( n85425 , n85424 , n31437 );
or ( n85426 , n85419 , n85425 );
and ( n85427 , n85426 , n31468 );
not ( n85428 , n31497 );
and ( n85429 , n85428 , n33999 );
not ( n85430 , n31454 );
not ( n85431 , n31501 );
and ( n85432 , n85431 , n34038 );
xor ( n85433 , n34039 , n34076 );
and ( n85434 , n85433 , n31501 );
or ( n85435 , n85432 , n85434 );
and ( n85436 , n85430 , n85435 );
and ( n85437 , n85422 , n31454 );
or ( n85438 , n85436 , n85437 );
and ( n85439 , n85438 , n31497 );
or ( n85440 , n85429 , n85439 );
and ( n85441 , n85440 , n31521 );
and ( n85442 , n33999 , n31553 );
or ( n85443 , n85413 , n85417 , n85427 , n85441 , n85442 );
and ( n85444 , n85443 , n31557 );
not ( n85445 , n31452 );
not ( n85446 , n31619 );
and ( n85447 , n85446 , n34095 );
xor ( n85448 , n34096 , n34133 );
and ( n85449 , n85448 , n31619 );
or ( n85450 , n85447 , n85449 );
and ( n85451 , n85445 , n85450 );
and ( n85452 , n33999 , n31452 );
or ( n85453 , n85451 , n85452 );
and ( n85454 , n85453 , n31638 );
buf ( n85455 , n33973 );
and ( n85456 , n33999 , n31650 );
or ( n85457 , C0 , n85409 , n85444 , n85454 , n85455 , n85456 );
buf ( n85458 , n85457 );
buf ( n85459 , n85458 );
buf ( n85460 , n30987 );
buf ( n85461 , n30987 );
buf ( n85462 , n31655 );
buf ( n85463 , n67277 );
buf ( n85464 , n53832 );
or ( n85465 , C0 , C0 , C0 , n85463 , n85464 );
and ( n85466 , n85465 , n53828 );
buf ( n85467 , n53758 );
buf ( n85468 , n67277 );
buf ( n85469 , n53832 );
or ( n85470 , C0 , C0 , n85467 , n85468 , n85469 );
and ( n85471 , n85470 , n53864 );
or ( n85472 , C0 , C0 , n85466 , n85471 );
buf ( n85473 , n85472 );
buf ( n85474 , n85473 );
not ( n85475 , n40163 );
and ( n85476 , n85475 , n31796 );
not ( n85477 , n52120 );
and ( n85478 , n85477 , n31796 );
and ( n85479 , n32252 , n52120 );
or ( n85480 , n85478 , n85479 );
and ( n85481 , n85480 , n40163 );
or ( n85482 , n85476 , n85481 );
and ( n85483 , n85482 , n32498 );
not ( n85484 , n52128 );
not ( n85485 , n52120 );
and ( n85486 , n85485 , n31796 );
and ( n85487 , n40393 , n52120 );
or ( n85488 , n85486 , n85487 );
and ( n85489 , n85484 , n85488 );
and ( n85490 , n40393 , n52128 );
or ( n85491 , n85489 , n85490 );
and ( n85492 , n85491 , n32473 );
not ( n85493 , n32475 );
not ( n85494 , n52128 );
not ( n85495 , n52120 );
and ( n85496 , n85495 , n31796 );
and ( n85497 , n40393 , n52120 );
or ( n85498 , n85496 , n85497 );
and ( n85499 , n85494 , n85498 );
and ( n85500 , n40393 , n52128 );
or ( n85501 , n85499 , n85500 );
and ( n85502 , n85493 , n85501 );
not ( n85503 , n52148 );
not ( n85504 , n52150 );
and ( n85505 , n85504 , n85501 );
and ( n85506 , n40972 , n52150 );
or ( n85507 , n85505 , n85506 );
and ( n85508 , n85503 , n85507 );
and ( n85509 , n41267 , n52148 );
or ( n85510 , n85508 , n85509 );
and ( n85511 , n85510 , n32475 );
or ( n85512 , n85502 , n85511 );
and ( n85513 , n85512 , n32486 );
and ( n85514 , n31796 , n41278 );
or ( n85515 , C0 , n85483 , n85492 , n85513 , n85514 );
buf ( n85516 , n85515 );
buf ( n85517 , n85516 );
buf ( n85518 , n30987 );
buf ( n85519 , n30987 );
buf ( n85520 , n31655 );
and ( n85521 , n50596 , n31645 );
not ( n85522 , n45274 );
and ( n85523 , n85522 , n68204 );
and ( n85524 , n70773 , n45274 );
or ( n85525 , n85523 , n85524 );
and ( n85526 , n85525 , n31373 );
not ( n85527 , n45280 );
and ( n85528 , n85527 , n68204 );
and ( n85529 , n70773 , n45280 );
or ( n85530 , n85528 , n85529 );
and ( n85531 , n85530 , n31468 );
and ( n85532 , n68204 , n45802 );
or ( n85533 , n85526 , n85531 , n85532 );
and ( n85534 , n85533 , n31557 );
and ( n85535 , n68204 , n45808 );
or ( n85536 , C0 , n85521 , n85534 , n85535 );
buf ( n85537 , n85536 );
buf ( n85538 , n85537 );
not ( n85539 , n40163 );
and ( n85540 , n85539 , n31865 );
not ( n85541 , n56287 );
and ( n85542 , n85541 , n31865 );
and ( n85543 , n32218 , n56287 );
or ( n85544 , n85542 , n85543 );
and ( n85545 , n85544 , n40163 );
or ( n85546 , n85540 , n85545 );
and ( n85547 , n85546 , n32498 );
not ( n85548 , n56295 );
not ( n85549 , n56287 );
and ( n85550 , n85549 , n31865 );
and ( n85551 , n42255 , n56287 );
or ( n85552 , n85550 , n85551 );
and ( n85553 , n85548 , n85552 );
and ( n85554 , n42255 , n56295 );
or ( n85555 , n85553 , n85554 );
and ( n85556 , n85555 , n32473 );
not ( n85557 , n32475 );
not ( n85558 , n56295 );
not ( n85559 , n56287 );
and ( n85560 , n85559 , n31865 );
and ( n85561 , n42255 , n56287 );
or ( n85562 , n85560 , n85561 );
and ( n85563 , n85558 , n85562 );
and ( n85564 , n42255 , n56295 );
or ( n85565 , n85563 , n85564 );
and ( n85566 , n85557 , n85565 );
not ( n85567 , n56315 );
not ( n85568 , n56317 );
and ( n85569 , n85568 , n85565 );
and ( n85570 , n42283 , n56317 );
or ( n85571 , n85569 , n85570 );
and ( n85572 , n85567 , n85571 );
and ( n85573 , n42291 , n56315 );
or ( n85574 , n85572 , n85573 );
and ( n85575 , n85574 , n32475 );
or ( n85576 , n85566 , n85575 );
and ( n85577 , n85576 , n32486 );
and ( n85578 , n31865 , n41278 );
or ( n85579 , C0 , n85547 , n85556 , n85577 , n85578 );
buf ( n85580 , n85579 );
buf ( n85581 , n85580 );
buf ( n85582 , n30987 );
buf ( n85583 , n31655 );
buf ( n85584 , n30987 );
xor ( n85585 , n33119 , n52219 );
and ( n85586 , n85585 , n33201 );
not ( n85587 , n41576 );
and ( n85588 , n85587 , n33119 );
buf ( n85589 , n32887 );
and ( n85590 , n85589 , n41576 );
or ( n85591 , n85588 , n85590 );
and ( n85592 , n85591 , n33189 );
and ( n85593 , n33119 , n41592 );
or ( n85594 , n85586 , n85592 , n85593 );
and ( n85595 , n85594 , n33208 );
and ( n85596 , n33119 , n39805 );
or ( n85597 , C0 , n85595 , n85596 );
buf ( n85598 , n85597 );
buf ( n85599 , n85598 );
buf ( n85600 , n30987 );
buf ( n85601 , n31655 );
not ( n85602 , n50828 );
not ( n85603 , n50834 );
and ( n85604 , n85603 , n40242 );
and ( n85605 , n35534 , n50834 );
or ( n85606 , n85604 , n85605 );
and ( n85607 , n85602 , n85606 );
and ( n85608 , n35530 , n50828 );
or ( n85609 , n85607 , n85608 );
buf ( n85610 , n85609 );
buf ( n85611 , n85610 );
not ( n85612 , n43755 );
and ( n85613 , n85612 , n42868 );
xor ( n85614 , n43764 , n43259 );
and ( n85615 , n85614 , n43755 );
or ( n85616 , n85613 , n85615 );
and ( n85617 , n85616 , n43774 );
not ( n85618 , n44663 );
and ( n85619 , n85618 , n43793 );
xor ( n85620 , n44672 , n44171 );
and ( n85621 , n85620 , n44663 );
or ( n85622 , n85619 , n85621 );
and ( n85623 , n85622 , n44682 );
buf ( n85624 , RI15b45078_220);
and ( n85625 , n85624 , n44695 );
or ( n85626 , n85617 , n85623 , n85625 );
buf ( n85627 , n85626 );
buf ( n85628 , n85627 );
buf ( n85629 , n30987 );
buf ( n85630 , n30987 );
buf ( n85631 , n31655 );
buf ( n85632 , n31655 );
buf ( n85633 , n40215 );
buf ( n85634 , n31655 );
not ( n85635 , n48765 );
and ( n85636 , n85635 , n33218 );
and ( n85637 , n78449 , n48765 );
or ( n85638 , n85636 , n85637 );
and ( n85639 , n85638 , n33180 );
not ( n85640 , n49054 );
and ( n85641 , n85640 , n33218 );
and ( n85642 , n78460 , n49054 );
or ( n85643 , n85641 , n85642 );
and ( n85644 , n85643 , n33178 );
and ( n85645 , n33218 , n49774 );
or ( n85646 , n85639 , n85644 , n85645 );
and ( n85647 , n85646 , n33208 );
and ( n85648 , n33287 , n33375 );
not ( n85649 , n32968 );
and ( n85650 , n85649 , n33287 );
xor ( n85651 , n33218 , n59700 );
and ( n85652 , n85651 , n32968 );
or ( n85653 , n85650 , n85652 );
and ( n85654 , n85653 , n33370 );
and ( n85655 , n32981 , n35056 );
and ( n85656 , n33218 , n49794 );
or ( n85657 , C0 , n85647 , n85648 , n85654 , n85655 , n85656 );
buf ( n85658 , n85657 );
buf ( n85659 , n85658 );
buf ( n85660 , n30987 );
buf ( n85661 , n30987 );
buf ( n85662 , n31655 );
and ( n85663 , n46032 , n32500 );
not ( n85664 , n35211 );
and ( n85665 , n85664 , n37561 );
buf ( n85666 , n85665 );
and ( n85667 , n85666 , n32421 );
not ( n85668 , n35245 );
and ( n85669 , n85668 , n37561 );
buf ( n85670 , n85669 );
and ( n85671 , n85670 , n32419 );
not ( n85672 , n35278 );
and ( n85673 , n85672 , n37561 );
not ( n85674 , n35295 );
and ( n85675 , n85674 , n49591 );
xor ( n85676 , n37561 , n49535 );
and ( n85677 , n85676 , n35295 );
or ( n85678 , n85675 , n85677 );
and ( n85679 , n85678 , n35278 );
or ( n85680 , n85673 , n85679 );
and ( n85681 , n85680 , n32417 );
not ( n85682 , n35331 );
and ( n85683 , n85682 , n37561 );
not ( n85684 , n35294 );
not ( n85685 , n45995 );
and ( n85686 , n85685 , n49591 );
xor ( n85687 , n49592 , n49621 );
and ( n85688 , n85687 , n45995 );
or ( n85689 , n85686 , n85688 );
and ( n85690 , n85684 , n85689 );
and ( n85691 , n85676 , n35294 );
or ( n85692 , n85690 , n85691 );
and ( n85693 , n85692 , n35331 );
or ( n85694 , n85683 , n85693 );
and ( n85695 , n85694 , n32415 );
and ( n85696 , n37561 , n35354 );
or ( n85697 , n85667 , n85671 , n85681 , n85695 , n85696 );
and ( n85698 , n85697 , n32456 );
not ( n85699 , n32475 );
not ( n85700 , n46060 );
and ( n85701 , n85700 , n49681 );
xor ( n85702 , n49682 , n49715 );
and ( n85703 , n85702 , n46060 );
or ( n85704 , n85701 , n85703 );
and ( n85705 , n85699 , n85704 );
and ( n85706 , n37561 , n32475 );
or ( n85707 , n85705 , n85706 );
and ( n85708 , n85707 , n32486 );
buf ( n85709 , n32489 );
and ( n85710 , n37561 , n35367 );
or ( n85711 , C0 , n85663 , n85698 , n85708 , n85709 , n85710 );
buf ( n85712 , n85711 );
buf ( n85713 , n85712 );
buf ( n85714 , n30987 );
buf ( n85715 , n30987 );
and ( n85716 , n49073 , n48639 );
not ( n85717 , n48642 );
and ( n85718 , n85717 , n48598 );
and ( n85719 , n49073 , n48642 );
or ( n85720 , n85718 , n85719 );
and ( n85721 , n85720 , n32890 );
not ( n85722 , n48648 );
and ( n85723 , n85722 , n48598 );
and ( n85724 , n49073 , n48648 );
or ( n85725 , n85723 , n85724 );
and ( n85726 , n85725 , n32924 );
not ( n85727 , n48654 );
and ( n85728 , n85727 , n48598 );
and ( n85729 , n49073 , n48654 );
or ( n85730 , n85728 , n85729 );
and ( n85731 , n85730 , n33038 );
not ( n85732 , n48660 );
and ( n85733 , n85732 , n48598 );
and ( n85734 , n49073 , n48660 );
or ( n85735 , n85733 , n85734 );
and ( n85736 , n85735 , n33172 );
not ( n85737 , n41576 );
and ( n85738 , n85737 , n48598 );
and ( n85739 , n48783 , n41576 );
or ( n85740 , n85738 , n85739 );
and ( n85741 , n85740 , n33189 );
not ( n85742 , n48730 );
and ( n85743 , n85742 , n48598 );
and ( n85744 , n48783 , n48730 );
or ( n85745 , n85743 , n85744 );
and ( n85746 , n85745 , n33187 );
not ( n85747 , n48765 );
and ( n85748 , n85747 , n48598 );
xor ( n85749 , n48783 , n49005 );
and ( n85750 , n85749 , n48765 );
or ( n85751 , n85748 , n85750 );
and ( n85752 , n85751 , n33180 );
not ( n85753 , n49054 );
and ( n85754 , n85753 , n48598 );
not ( n85755 , n48845 );
xor ( n85756 , n49073 , n49119 );
and ( n85757 , n85755 , n85756 );
xnor ( n85758 , n49182 , n49245 );
and ( n85759 , n85758 , n48845 );
or ( n85760 , n85757 , n85759 );
and ( n85761 , n85760 , n49054 );
or ( n85762 , n85754 , n85761 );
and ( n85763 , n85762 , n33178 );
and ( n85764 , n49182 , n49275 );
or ( n85765 , n85716 , n85721 , n85726 , n85731 , n85736 , n85741 , n85746 , n85752 , n85763 , n85764 );
and ( n85766 , n85765 , n33208 );
and ( n85767 , n32991 , n35056 );
and ( n85768 , n48598 , n49286 );
or ( n85769 , C0 , n85766 , n85767 , n85768 );
buf ( n85770 , n85769 );
buf ( n85771 , n85770 );
buf ( n85772 , n31655 );
buf ( n85773 , n31655 );
buf ( n85774 , n31655 );
not ( n85775 , n36587 );
and ( n85776 , n85775 , n36447 );
xor ( n85777 , n50174 , n50213 );
and ( n85778 , n85777 , n36587 );
or ( n85779 , n85776 , n85778 );
and ( n85780 , n85779 , n36596 );
not ( n85781 , n37485 );
and ( n85782 , n85781 , n37349 );
xor ( n85783 , n50224 , n50263 );
and ( n85784 , n85783 , n37485 );
or ( n85785 , n85782 , n85784 );
and ( n85786 , n85785 , n37494 );
and ( n85787 , n41860 , n37506 );
or ( n85788 , n85780 , n85786 , n85787 );
buf ( n85789 , n85788 );
buf ( n85790 , n85789 );
and ( n85791 , n50443 , n50275 );
not ( n85792 , n50278 );
and ( n85793 , n85792 , n50411 );
and ( n85794 , n50443 , n50278 );
or ( n85795 , n85793 , n85794 );
and ( n85796 , n85795 , n32421 );
not ( n85797 , n50002 );
and ( n85798 , n85797 , n50411 );
and ( n85799 , n50443 , n50002 );
or ( n85800 , n85798 , n85799 );
and ( n85801 , n85800 , n32419 );
not ( n85802 , n50289 );
and ( n85803 , n85802 , n50411 );
and ( n85804 , n50443 , n50289 );
or ( n85805 , n85803 , n85804 );
and ( n85806 , n85805 , n32417 );
not ( n85807 , n50008 );
and ( n85808 , n85807 , n50411 );
and ( n85809 , n50443 , n50008 );
or ( n85810 , n85808 , n85809 );
and ( n85811 , n85810 , n32415 );
not ( n85812 , n47331 );
and ( n85813 , n85812 , n50411 );
and ( n85814 , n50421 , n47331 );
or ( n85815 , n85813 , n85814 );
and ( n85816 , n85815 , n32413 );
not ( n85817 , n50067 );
and ( n85818 , n85817 , n50411 );
and ( n85819 , n50421 , n50067 );
or ( n85820 , n85818 , n85819 );
and ( n85821 , n85820 , n32411 );
not ( n85822 , n31728 );
and ( n85823 , n85822 , n50411 );
and ( n85824 , n71290 , n31728 );
or ( n85825 , n85823 , n85824 );
and ( n85826 , n85825 , n32253 );
not ( n85827 , n32283 );
and ( n85828 , n85827 , n50411 );
and ( n85829 , n71301 , n32283 );
or ( n85830 , n85828 , n85829 );
and ( n85831 , n85830 , n32398 );
and ( n85832 , n50460 , n50334 );
or ( n85833 , n85791 , n85796 , n85801 , n85806 , n85811 , n85816 , n85821 , n85826 , n85831 , n85832 );
and ( n85834 , n85833 , n32456 );
and ( n85835 , n37539 , n32489 );
and ( n85836 , n50411 , n50345 );
or ( n85837 , C0 , n85834 , n85835 , n85836 );
buf ( n85838 , n85837 );
buf ( n85839 , n85838 );
buf ( n85840 , n30987 );
buf ( n85841 , n30987 );
buf ( n85842 , n30987 );
and ( n85843 , n49071 , n48639 );
not ( n85844 , n48642 );
and ( n85845 , n85844 , n48596 );
and ( n85846 , n49071 , n48642 );
or ( n85847 , n85845 , n85846 );
and ( n85848 , n85847 , n32890 );
not ( n85849 , n48648 );
and ( n85850 , n85849 , n48596 );
and ( n85851 , n49071 , n48648 );
or ( n85852 , n85850 , n85851 );
and ( n85853 , n85852 , n32924 );
not ( n85854 , n48654 );
and ( n85855 , n85854 , n48596 );
and ( n85856 , n49071 , n48654 );
or ( n85857 , n85855 , n85856 );
and ( n85858 , n85857 , n33038 );
not ( n85859 , n48660 );
and ( n85860 , n85859 , n48596 );
and ( n85861 , n49071 , n48660 );
or ( n85862 , n85860 , n85861 );
and ( n85863 , n85862 , n33172 );
not ( n85864 , n41576 );
and ( n85865 , n85864 , n48596 );
and ( n85866 , n48781 , n41576 );
or ( n85867 , n85865 , n85866 );
and ( n85868 , n85867 , n33189 );
not ( n85869 , n48730 );
and ( n85870 , n85869 , n48596 );
and ( n85871 , n48781 , n48730 );
or ( n85872 , n85870 , n85871 );
and ( n85873 , n85872 , n33187 );
not ( n85874 , n48765 );
and ( n85875 , n85874 , n48596 );
xor ( n85876 , n48781 , n49007 );
and ( n85877 , n85876 , n48765 );
or ( n85878 , n85875 , n85877 );
and ( n85879 , n85878 , n33180 );
not ( n85880 , n49054 );
and ( n85881 , n85880 , n48596 );
not ( n85882 , n48845 );
xor ( n85883 , n49071 , n49121 );
and ( n85884 , n85882 , n85883 );
xnor ( n85885 , n49180 , n49247 );
and ( n85886 , n85885 , n48845 );
or ( n85887 , n85884 , n85886 );
and ( n85888 , n85887 , n49054 );
or ( n85889 , n85881 , n85888 );
and ( n85890 , n85889 , n33178 );
and ( n85891 , n49180 , n49275 );
or ( n85892 , n85843 , n85848 , n85853 , n85858 , n85863 , n85868 , n85873 , n85879 , n85890 , n85891 );
and ( n85893 , n85892 , n33208 );
and ( n85894 , n32989 , n35056 );
and ( n85895 , n48596 , n49286 );
or ( n85896 , C0 , n85893 , n85894 , n85895 );
buf ( n85897 , n85896 );
buf ( n85898 , n85897 );
buf ( n85899 , n31655 );
buf ( n85900 , n31655 );
buf ( n85901 , n31655 );
not ( n85902 , n46356 );
and ( n85903 , n85902 , n31117 );
not ( n85904 , n50109 );
and ( n85905 , n85904 , n31117 );
and ( n85906 , n31138 , n50109 );
or ( n85907 , n85905 , n85906 );
and ( n85908 , n85907 , n46356 );
or ( n85909 , n85903 , n85908 );
and ( n85910 , n85909 , n31649 );
not ( n85911 , n50117 );
not ( n85912 , n50109 );
and ( n85913 , n85912 , n31117 );
and ( n85914 , n56920 , n50109 );
or ( n85915 , n85913 , n85914 );
and ( n85916 , n85911 , n85915 );
and ( n85917 , n56920 , n50117 );
or ( n85918 , n85916 , n85917 );
and ( n85919 , n85918 , n31643 );
not ( n85920 , n31452 );
not ( n85921 , n50117 );
not ( n85922 , n50109 );
and ( n85923 , n85922 , n31117 );
and ( n85924 , n56920 , n50109 );
or ( n85925 , n85923 , n85924 );
and ( n85926 , n85921 , n85925 );
and ( n85927 , n56920 , n50117 );
or ( n85928 , n85926 , n85927 );
and ( n85929 , n85920 , n85928 );
not ( n85930 , n50142 );
not ( n85931 , n50144 );
and ( n85932 , n85931 , n85928 );
and ( n85933 , n56946 , n50144 );
or ( n85934 , n85932 , n85933 );
and ( n85935 , n85930 , n85934 );
and ( n85936 , n56954 , n50142 );
or ( n85937 , n85935 , n85936 );
and ( n85938 , n85937 , n31452 );
or ( n85939 , n85929 , n85938 );
and ( n85940 , n85939 , n31638 );
and ( n85941 , n31117 , n47277 );
or ( n85942 , C0 , n85910 , n85919 , n85940 , n85941 );
buf ( n85943 , n85942 );
buf ( n85944 , n85943 );
buf ( n85945 , n30987 );
xor ( n85946 , n50900 , n64709 );
and ( n85947 , n85946 , n32431 );
not ( n85948 , n50002 );
and ( n85949 , n85948 , n50900 );
and ( n85950 , n40457 , n50002 );
or ( n85951 , n85949 , n85950 );
and ( n85952 , n85951 , n32419 );
not ( n85953 , n50008 );
and ( n85954 , n85953 , n50900 );
not ( n85955 , n51594 );
and ( n85956 , n85955 , n51423 );
xor ( n85957 , n51603 , n40244 );
and ( n85958 , n85957 , n51594 );
or ( n85959 , n85956 , n85958 );
and ( n85960 , n85959 , n50008 );
or ( n85961 , n85954 , n85960 );
and ( n85962 , n85961 , n32415 );
not ( n85963 , n50067 );
and ( n85964 , n85963 , n50900 );
and ( n85965 , n32036 , n60510 );
and ( n85966 , n32038 , n60512 );
and ( n85967 , n32040 , n60514 );
and ( n85968 , n32042 , n60516 );
and ( n85969 , n32044 , n60518 );
and ( n85970 , n32046 , n60520 );
and ( n85971 , n32048 , n60522 );
and ( n85972 , n32050 , n60524 );
and ( n85973 , n32052 , n60526 );
and ( n85974 , n32054 , n60528 );
and ( n85975 , n32056 , n60530 );
and ( n85976 , n32058 , n60532 );
and ( n85977 , n32060 , n60534 );
and ( n85978 , n32062 , n60536 );
and ( n85979 , n32064 , n60538 );
and ( n85980 , n32066 , n60540 );
or ( n85981 , n85965 , n85966 , n85967 , n85968 , n85969 , n85970 , n85971 , n85972 , n85973 , n85974 , n85975 , n85976 , n85977 , n85978 , n85979 , n85980 );
and ( n85982 , n85981 , n50067 );
or ( n85983 , n85964 , n85982 );
and ( n85984 , n85983 , n32411 );
and ( n85985 , n50900 , n50098 );
or ( n85986 , n85947 , n85952 , n85962 , n85984 , n85985 );
and ( n85987 , n85986 , n32456 );
and ( n85988 , n50900 , n47409 );
or ( n85989 , C0 , n85987 , n85988 );
buf ( n85990 , n85989 );
buf ( n85991 , n85990 );
buf ( n85992 , n31655 );
buf ( n85993 , n31655 );
not ( n85994 , n35542 );
and ( n85995 , n85994 , n41845 );
and ( n85996 , n44684 , n35542 );
or ( n85997 , n85995 , n85996 );
buf ( n85998 , n85997 );
buf ( n85999 , n85998 );
buf ( n86000 , n30987 );
and ( n86001 , n33240 , n32528 );
not ( n86002 , n32598 );
and ( n86003 , n86002 , n33003 );
and ( n86004 , n48795 , n32598 );
or ( n86005 , n86003 , n86004 );
and ( n86006 , n86005 , n32890 );
not ( n86007 , n32919 );
and ( n86008 , n86007 , n33003 );
and ( n86009 , n48795 , n32919 );
or ( n86010 , n86008 , n86009 );
and ( n86011 , n86010 , n32924 );
not ( n86012 , n32953 );
and ( n86013 , n86012 , n33003 );
not ( n86014 , n32971 );
and ( n86015 , n86014 , n33131 );
not ( n86016 , n33003 );
and ( n86017 , n86016 , n32971 );
or ( n86018 , n86015 , n86017 );
and ( n86019 , n86018 , n32953 );
or ( n86020 , n86013 , n86019 );
and ( n86021 , n86020 , n33038 );
not ( n86022 , n33067 );
and ( n86023 , n86022 , n33003 );
not ( n86024 , n32970 );
not ( n86025 , n33071 );
and ( n86026 , n86025 , n33131 );
xor ( n86027 , n33132 , n33134 );
and ( n86028 , n86027 , n33071 );
or ( n86029 , n86026 , n86028 );
and ( n86030 , n86024 , n86029 );
and ( n86031 , n86016 , n32970 );
or ( n86032 , n86030 , n86031 );
and ( n86033 , n86032 , n33067 );
or ( n86034 , n86023 , n86033 );
and ( n86035 , n86034 , n33172 );
and ( n86036 , n33003 , n33204 );
or ( n86037 , n86006 , n86011 , n86021 , n86035 , n86036 );
and ( n86038 , n86037 , n33208 );
not ( n86039 , n32968 );
not ( n86040 , n33270 );
and ( n86041 , n86040 , n33331 );
xor ( n86042 , n33332 , n33334 );
and ( n86043 , n86042 , n33270 );
or ( n86044 , n86041 , n86043 );
and ( n86045 , n86039 , n86044 );
and ( n86046 , n33003 , n32968 );
or ( n86047 , n86045 , n86046 );
and ( n86048 , n86047 , n33370 );
and ( n86049 , n33003 , n33382 );
or ( n86050 , C0 , n86001 , n86038 , n86048 , C0 , n86049 );
buf ( n86051 , n86050 );
buf ( n86052 , n86051 );
buf ( n86053 , n30987 );
buf ( n86054 , n31655 );
and ( n86055 , n32460 , n32500 );
not ( n86056 , n35211 );
and ( n86057 , n86056 , n37579 );
and ( n86058 , n31658 , n58320 );
and ( n86059 , n86058 , n35211 );
or ( n86060 , n86057 , n86059 );
and ( n86061 , n86060 , n32421 );
not ( n86062 , n35245 );
and ( n86063 , n86062 , n37579 );
and ( n86064 , n86058 , n35245 );
or ( n86065 , n86063 , n86064 );
and ( n86066 , n86065 , n32419 );
not ( n86067 , n35278 );
and ( n86068 , n86067 , n37579 );
not ( n86069 , n35295 );
and ( n86070 , n86069 , n47288 );
xor ( n86071 , n37579 , n49525 );
and ( n86072 , n86071 , n35295 );
or ( n86073 , n86070 , n86072 );
and ( n86074 , n86073 , n35278 );
or ( n86075 , n86068 , n86074 );
and ( n86076 , n86075 , n32417 );
not ( n86077 , n35331 );
and ( n86078 , n86077 , n37579 );
not ( n86079 , n35294 );
not ( n86080 , n45995 );
and ( n86081 , n86080 , n47288 );
xor ( n86082 , n49606 , n49611 );
and ( n86083 , n86082 , n45995 );
or ( n86084 , n86081 , n86083 );
and ( n86085 , n86079 , n86084 );
and ( n86086 , n86071 , n35294 );
or ( n86087 , n86085 , n86086 );
and ( n86088 , n86087 , n35331 );
or ( n86089 , n86078 , n86088 );
and ( n86090 , n86089 , n32415 );
and ( n86091 , n37579 , n35354 );
or ( n86092 , n86061 , n86066 , n86076 , n86090 , n86091 );
and ( n86093 , n86092 , n32456 );
not ( n86094 , n32475 );
not ( n86095 , n46060 );
and ( n86096 , n86095 , n49697 );
xor ( n86097 , n49698 , n49705 );
and ( n86098 , n86097 , n46060 );
or ( n86099 , n86096 , n86098 );
and ( n86100 , n86094 , n86099 );
and ( n86101 , n37579 , n32475 );
or ( n86102 , n86100 , n86101 );
and ( n86103 , n86102 , n32486 );
buf ( n86104 , n32489 );
and ( n86105 , n37579 , n35367 );
or ( n86106 , C0 , n86055 , n86093 , n86103 , n86104 , n86105 );
buf ( n86107 , n86106 );
buf ( n86108 , n86107 );
buf ( n86109 , n30987 );
not ( n86110 , n34150 );
and ( n86111 , n86110 , n32751 );
not ( n86112 , n56140 );
and ( n86113 , n86112 , n32751 );
and ( n86114 , n32755 , n56140 );
or ( n86115 , n86113 , n86114 );
and ( n86116 , n86115 , n34150 );
or ( n86117 , n86111 , n86116 );
and ( n86118 , n86117 , n33381 );
not ( n86119 , n56148 );
not ( n86120 , n56140 );
and ( n86121 , n86120 , n32751 );
and ( n86122 , n35083 , n56140 );
or ( n86123 , n86121 , n86122 );
and ( n86124 , n86119 , n86123 );
and ( n86125 , n35083 , n56148 );
or ( n86126 , n86124 , n86125 );
and ( n86127 , n86126 , n33375 );
not ( n86128 , n32968 );
not ( n86129 , n56148 );
not ( n86130 , n56140 );
and ( n86131 , n86130 , n32751 );
and ( n86132 , n35083 , n56140 );
or ( n86133 , n86131 , n86132 );
and ( n86134 , n86129 , n86133 );
and ( n86135 , n35083 , n56148 );
or ( n86136 , n86134 , n86135 );
and ( n86137 , n86128 , n86136 );
not ( n86138 , n56168 );
not ( n86139 , n56170 );
and ( n86140 , n86139 , n86136 );
and ( n86141 , n35107 , n56170 );
or ( n86142 , n86140 , n86141 );
and ( n86143 , n86138 , n86142 );
and ( n86144 , n35115 , n56168 );
or ( n86145 , n86143 , n86144 );
and ( n86146 , n86145 , n32968 );
or ( n86147 , n86137 , n86146 );
and ( n86148 , n86147 , n33370 );
and ( n86149 , n32751 , n35062 );
or ( n86150 , C0 , n86118 , n86127 , n86148 , n86149 );
buf ( n86151 , n86150 );
buf ( n86152 , n86151 );
not ( n86153 , n34150 );
and ( n86154 , n86153 , n32781 );
not ( n86155 , n56093 );
and ( n86156 , n86155 , n32781 );
and ( n86157 , n32789 , n56093 );
or ( n86158 , n86156 , n86157 );
and ( n86159 , n86158 , n34150 );
or ( n86160 , n86154 , n86159 );
and ( n86161 , n86160 , n33381 );
not ( n86162 , n56101 );
not ( n86163 , n56093 );
and ( n86164 , n86163 , n32781 );
and ( n86165 , n34301 , n56093 );
or ( n86166 , n86164 , n86165 );
and ( n86167 , n86162 , n86166 );
and ( n86168 , n34301 , n56101 );
or ( n86169 , n86167 , n86168 );
and ( n86170 , n86169 , n33375 );
not ( n86171 , n32968 );
not ( n86172 , n56101 );
not ( n86173 , n56093 );
and ( n86174 , n86173 , n32781 );
and ( n86175 , n34301 , n56093 );
or ( n86176 , n86174 , n86175 );
and ( n86177 , n86172 , n86176 );
and ( n86178 , n34301 , n56101 );
or ( n86179 , n86177 , n86178 );
and ( n86180 , n86171 , n86179 );
not ( n86181 , n56121 );
not ( n86182 , n56123 );
and ( n86183 , n86182 , n86179 );
and ( n86184 , n34761 , n56123 );
or ( n86185 , n86183 , n86184 );
and ( n86186 , n86181 , n86185 );
and ( n86187 , n35050 , n56121 );
or ( n86188 , n86186 , n86187 );
and ( n86189 , n86188 , n32968 );
or ( n86190 , n86180 , n86189 );
and ( n86191 , n86190 , n33370 );
and ( n86192 , n32781 , n35062 );
or ( n86193 , C0 , n86161 , n86170 , n86191 , n86192 );
buf ( n86194 , n86193 );
buf ( n86195 , n86194 );
buf ( n86196 , n30987 );
buf ( n86197 , n31655 );
buf ( n86198 , n31655 );
buf ( n86199 , n31655 );
not ( n86200 , n31437 );
and ( n86201 , n86200 , n51807 );
and ( n86202 , n68689 , n31437 );
or ( n86203 , n86201 , n86202 );
and ( n86204 , n86203 , n31468 );
not ( n86205 , n41837 );
and ( n86206 , n86205 , n51807 );
and ( n86207 , n51813 , n41837 );
or ( n86208 , n86206 , n86207 );
and ( n86209 , n86208 , n31521 );
and ( n86210 , n51807 , n42158 );
or ( n86211 , n86204 , n86209 , n86210 );
and ( n86212 , n86211 , n31557 );
and ( n86213 , n51807 , n40154 );
or ( n86214 , C0 , n86212 , n86213 );
buf ( n86215 , n86214 );
buf ( n86216 , n86215 );
not ( n86217 , n40163 );
and ( n86218 , n86217 , n31933 );
not ( n86219 , n42171 );
and ( n86220 , n86219 , n31933 );
and ( n86221 , n32183 , n42171 );
or ( n86222 , n86220 , n86221 );
and ( n86223 , n86222 , n40163 );
or ( n86224 , n86218 , n86223 );
and ( n86225 , n86224 , n32498 );
not ( n86226 , n42180 );
not ( n86227 , n42171 );
and ( n86228 , n86227 , n31933 );
and ( n86229 , n45178 , n42171 );
or ( n86230 , n86228 , n86229 );
and ( n86231 , n86226 , n86230 );
and ( n86232 , n45178 , n42180 );
or ( n86233 , n86231 , n86232 );
and ( n86234 , n86233 , n32473 );
not ( n86235 , n32475 );
not ( n86236 , n42180 );
not ( n86237 , n42171 );
and ( n86238 , n86237 , n31933 );
and ( n86239 , n45178 , n42171 );
or ( n86240 , n86238 , n86239 );
and ( n86241 , n86236 , n86240 );
and ( n86242 , n45178 , n42180 );
or ( n86243 , n86241 , n86242 );
and ( n86244 , n86235 , n86243 );
not ( n86245 , n42206 );
not ( n86246 , n42209 );
and ( n86247 , n86246 , n86243 );
and ( n86248 , n45206 , n42209 );
or ( n86249 , n86247 , n86248 );
and ( n86250 , n86245 , n86249 );
and ( n86251 , n45214 , n42206 );
or ( n86252 , n86250 , n86251 );
and ( n86253 , n86252 , n32475 );
or ( n86254 , n86244 , n86253 );
and ( n86255 , n86254 , n32486 );
and ( n86256 , n31933 , n41278 );
or ( n86257 , C0 , n86225 , n86234 , n86255 , n86256 );
buf ( n86258 , n86257 );
buf ( n86259 , n86258 );
buf ( n86260 , n30987 );
not ( n86261 , n46356 );
and ( n86262 , n86261 , n31317 );
not ( n86263 , n53353 );
and ( n86264 , n86263 , n31317 );
and ( n86265 , n31339 , n53353 );
or ( n86266 , n86264 , n86265 );
and ( n86267 , n86266 , n46356 );
or ( n86268 , n86262 , n86267 );
and ( n86269 , n86268 , n31649 );
not ( n86270 , n53361 );
not ( n86271 , n53353 );
and ( n86272 , n86271 , n31317 );
and ( n86273 , n47449 , n53353 );
or ( n86274 , n86272 , n86273 );
and ( n86275 , n86270 , n86274 );
and ( n86276 , n47449 , n53361 );
or ( n86277 , n86275 , n86276 );
and ( n86278 , n86277 , n31643 );
not ( n86279 , n31452 );
not ( n86280 , n53361 );
not ( n86281 , n53353 );
and ( n86282 , n86281 , n31317 );
and ( n86283 , n47449 , n53353 );
or ( n86284 , n86282 , n86283 );
and ( n86285 , n86280 , n86284 );
and ( n86286 , n47449 , n53361 );
or ( n86287 , n86285 , n86286 );
and ( n86288 , n86279 , n86287 );
not ( n86289 , n53381 );
not ( n86290 , n53383 );
and ( n86291 , n86290 , n86287 );
and ( n86292 , n47485 , n53383 );
or ( n86293 , n86291 , n86292 );
and ( n86294 , n86289 , n86293 );
and ( n86295 , n47503 , n53381 );
or ( n86296 , n86294 , n86295 );
and ( n86297 , n86296 , n31452 );
or ( n86298 , n86288 , n86297 );
and ( n86299 , n86298 , n31638 );
and ( n86300 , n31317 , n47277 );
or ( n86301 , C0 , n86269 , n86278 , n86299 , n86300 );
buf ( n86302 , n86301 );
buf ( n86303 , n86302 );
buf ( n86304 , n31655 );
buf ( n86305 , n30987 );
and ( n86306 , n65160 , n32494 );
not ( n86307 , n46083 );
buf ( n86308 , RI15b60300_1147);
and ( n86309 , n86307 , n86308 );
buf ( n86310 , n86309 );
and ( n86311 , n86310 , n32421 );
not ( n86312 , n46326 );
and ( n86313 , n86312 , n86308 );
and ( n86314 , n65166 , n46326 );
or ( n86315 , n86313 , n86314 );
and ( n86316 , n86315 , n32417 );
and ( n86317 , n86308 , n46340 );
or ( n86318 , n86311 , n86316 , n86317 );
and ( n86319 , n86318 , n32456 );
and ( n86320 , n86308 , n46349 );
or ( n86321 , C0 , n86306 , n86319 , n86320 );
buf ( n86322 , n86321 );
buf ( n86323 , n86322 );
buf ( n86324 , n31655 );
not ( n86325 , n32953 );
and ( n86326 , n86325 , n73768 );
and ( n86327 , n73776 , n32953 );
or ( n86328 , n86326 , n86327 );
and ( n86329 , n86328 , n33038 );
not ( n86330 , n39586 );
and ( n86331 , n86330 , n73768 );
not ( n86332 , n39775 );
and ( n86333 , n86332 , n39687 );
xor ( n86334 , n42656 , n42669 );
and ( n86335 , n86334 , n39775 );
or ( n86336 , n86333 , n86335 );
and ( n86337 , n86336 , n39586 );
or ( n86338 , n86331 , n86337 );
and ( n86339 , n86338 , n33172 );
and ( n86340 , n73768 , n39795 );
or ( n86341 , n86329 , n86339 , n86340 );
and ( n86342 , n86341 , n33208 );
and ( n86343 , n73768 , n39805 );
or ( n86344 , C0 , n86342 , n86343 );
buf ( n86345 , n86344 );
buf ( n86346 , n86345 );
buf ( n86347 , n31655 );
buf ( n86348 , n30987 );
buf ( n86349 , n30987 );
buf ( n86350 , n31655 );
buf ( n86351 , n40210 );
buf ( n86352 , n31655 );
xor ( n86353 , n35425 , n62856 );
and ( n86354 , n86353 , n31550 );
not ( n86355 , n39979 );
and ( n86356 , n86355 , n35425 );
and ( n86357 , n45095 , n76770 );
xor ( n86358 , n45078 , n86357 );
and ( n86359 , n86358 , n39979 );
or ( n86360 , n86356 , n86359 );
and ( n86361 , n86360 , n31538 );
and ( n86362 , n35425 , n40143 );
or ( n86363 , n86354 , n86361 , n86362 );
and ( n86364 , n86363 , n31557 );
and ( n86365 , n35425 , n40154 );
or ( n86366 , C0 , n86364 , n86365 );
buf ( n86367 , n86366 );
buf ( n86368 , n86367 );
not ( n86369 , n40163 );
and ( n86370 , n86369 , n31961 );
not ( n86371 , n40166 );
and ( n86372 , n86371 , n31961 );
and ( n86373 , n32183 , n40166 );
or ( n86374 , n86372 , n86373 );
and ( n86375 , n86374 , n40163 );
or ( n86376 , n86370 , n86375 );
and ( n86377 , n86376 , n32498 );
not ( n86378 , n40195 );
not ( n86379 , n40166 );
and ( n86380 , n86379 , n31961 );
and ( n86381 , n45178 , n40166 );
or ( n86382 , n86380 , n86381 );
and ( n86383 , n86378 , n86382 );
and ( n86384 , n45178 , n40195 );
or ( n86385 , n86383 , n86384 );
and ( n86386 , n86385 , n32473 );
not ( n86387 , n32475 );
not ( n86388 , n40195 );
not ( n86389 , n40166 );
and ( n86390 , n86389 , n31961 );
and ( n86391 , n45178 , n40166 );
or ( n86392 , n86390 , n86391 );
and ( n86393 , n86388 , n86392 );
and ( n86394 , n45178 , n40195 );
or ( n86395 , n86393 , n86394 );
and ( n86396 , n86387 , n86395 );
not ( n86397 , n40446 );
not ( n86398 , n40448 );
and ( n86399 , n86398 , n86395 );
and ( n86400 , n45206 , n40448 );
or ( n86401 , n86399 , n86400 );
and ( n86402 , n86397 , n86401 );
and ( n86403 , n45214 , n40446 );
or ( n86404 , n86402 , n86403 );
and ( n86405 , n86404 , n32475 );
or ( n86406 , n86396 , n86405 );
and ( n86407 , n86406 , n32486 );
and ( n86408 , n31961 , n41278 );
or ( n86409 , C0 , n86377 , n86386 , n86407 , n86408 );
buf ( n86410 , n86409 );
buf ( n86411 , n86410 );
buf ( n86412 , n30987 );
buf ( n86413 , n30987 );
and ( n86414 , n33781 , n48455 );
not ( n86415 , n48457 );
and ( n86416 , n86415 , n33441 );
and ( n86417 , n33781 , n48457 );
or ( n86418 , n86416 , n86417 );
and ( n86419 , n86418 , n31373 );
not ( n86420 , n44807 );
and ( n86421 , n86420 , n33441 );
and ( n86422 , n33781 , n44807 );
or ( n86423 , n86421 , n86422 );
and ( n86424 , n86423 , n31408 );
not ( n86425 , n48468 );
and ( n86426 , n86425 , n33441 );
and ( n86427 , n33781 , n48468 );
or ( n86428 , n86426 , n86427 );
and ( n86429 , n86428 , n31468 );
not ( n86430 , n44817 );
and ( n86431 , n86430 , n33441 );
and ( n86432 , n33781 , n44817 );
or ( n86433 , n86431 , n86432 );
and ( n86434 , n86433 , n31521 );
not ( n86435 , n39979 );
and ( n86436 , n86435 , n33441 );
and ( n86437 , n33611 , n39979 );
or ( n86438 , n86436 , n86437 );
and ( n86439 , n86438 , n31538 );
not ( n86440 , n45059 );
and ( n86441 , n86440 , n33441 );
and ( n86442 , n33611 , n45059 );
or ( n86443 , n86441 , n86442 );
and ( n86444 , n86443 , n31536 );
not ( n86445 , n33419 );
and ( n86446 , n86445 , n33441 );
and ( n86447 , n55808 , n33419 );
or ( n86448 , n86446 , n86447 );
and ( n86449 , n86448 , n31529 );
not ( n86450 , n33734 );
and ( n86451 , n86450 , n33441 );
and ( n86452 , n55821 , n33734 );
or ( n86453 , n86451 , n86452 );
and ( n86454 , n86453 , n31527 );
and ( n86455 , n33876 , n48513 );
or ( n86456 , n86414 , n86419 , n86424 , n86429 , n86434 , n86439 , n86444 , n86449 , n86454 , n86455 );
and ( n86457 , n86456 , n31557 );
and ( n86458 , n31459 , n33973 );
and ( n86459 , n33441 , n48524 );
or ( n86460 , C0 , n86457 , n86458 , n86459 );
buf ( n86461 , n86460 );
buf ( n86462 , n86461 );
buf ( n86463 , n31655 );
buf ( n86464 , n30987 );
not ( n86465 , n35278 );
and ( n86466 , n86465 , n53316 );
and ( n86467 , n53339 , n35278 );
or ( n86468 , n86466 , n86467 );
and ( n86469 , n86468 , n32417 );
not ( n86470 , n50008 );
and ( n86471 , n86470 , n53316 );
and ( n86472 , n72987 , n50008 );
or ( n86473 , n86471 , n86472 );
and ( n86474 , n86473 , n32415 );
and ( n86475 , n53316 , n48133 );
or ( n86476 , n86469 , n86474 , n86475 );
and ( n86477 , n86476 , n32456 );
and ( n86478 , n53316 , n47409 );
or ( n86479 , C0 , n86477 , n86478 );
buf ( n86480 , n86479 );
buf ( n86481 , n86480 );
not ( n86482 , n39369 );
and ( n86483 , n86482 , n33199 );
not ( n86484 , n48648 );
and ( n86485 , n86484 , n39369 );
and ( n86486 , n34188 , n48648 );
or ( n86487 , n86485 , n86486 );
and ( n86488 , n86487 , n32924 );
not ( n86489 , n48660 );
and ( n86490 , n86489 , n39369 );
not ( n86491 , n39584 );
buf ( n86492 , RI15b46770_269);
and ( n86493 , n86491 , n86492 );
not ( n86494 , n39775 );
and ( n86495 , n86494 , n39592 );
xor ( n86496 , n39779 , n34193 );
and ( n86497 , n86496 , n39775 );
or ( n86498 , n86495 , n86497 );
and ( n86499 , n86498 , n39584 );
or ( n86500 , n86493 , n86499 );
and ( n86501 , n86500 , n48660 );
or ( n86502 , n86490 , n86501 );
and ( n86503 , n86502 , n33172 );
not ( n86504 , n48730 );
and ( n86505 , n86504 , n39369 );
and ( n86506 , n48978 , n48730 );
or ( n86507 , n86505 , n86506 );
and ( n86508 , n86507 , n33187 );
and ( n86509 , n39369 , n54713 );
or ( n86510 , n86483 , n86488 , n86503 , n86508 , n86509 );
and ( n86511 , n86510 , n33208 );
and ( n86512 , n39369 , n39805 );
or ( n86513 , C0 , n86511 , n86512 );
buf ( n86514 , n86513 );
buf ( n86515 , n86514 );
buf ( n86516 , n31655 );
buf ( n86517 , n30987 );
buf ( n86518 , n30987 );
buf ( n86519 , n31655 );
buf ( n86520 , n40220 );
buf ( n86521 , n30987 );
buf ( n86522 , n30987 );
not ( n86523 , n34150 );
and ( n86524 , n86523 , n32773 );
not ( n86525 , n57038 );
and ( n86526 , n86525 , n32773 );
and ( n86527 , n32789 , n57038 );
or ( n86528 , n86526 , n86527 );
and ( n86529 , n86528 , n34150 );
or ( n86530 , n86524 , n86529 );
and ( n86531 , n86530 , n33381 );
not ( n86532 , n57046 );
not ( n86533 , n57038 );
and ( n86534 , n86533 , n32773 );
and ( n86535 , n34301 , n57038 );
or ( n86536 , n86534 , n86535 );
and ( n86537 , n86532 , n86536 );
and ( n86538 , n34301 , n57046 );
or ( n86539 , n86537 , n86538 );
and ( n86540 , n86539 , n33375 );
not ( n86541 , n32968 );
not ( n86542 , n57046 );
not ( n86543 , n57038 );
and ( n86544 , n86543 , n32773 );
and ( n86545 , n34301 , n57038 );
or ( n86546 , n86544 , n86545 );
and ( n86547 , n86542 , n86546 );
and ( n86548 , n34301 , n57046 );
or ( n86549 , n86547 , n86548 );
and ( n86550 , n86541 , n86549 );
not ( n86551 , n57066 );
not ( n86552 , n57068 );
and ( n86553 , n86552 , n86549 );
and ( n86554 , n34761 , n57068 );
or ( n86555 , n86553 , n86554 );
and ( n86556 , n86551 , n86555 );
and ( n86557 , n35050 , n57066 );
or ( n86558 , n86556 , n86557 );
and ( n86559 , n86558 , n32968 );
or ( n86560 , n86550 , n86559 );
and ( n86561 , n86560 , n33370 );
and ( n86562 , n32773 , n35062 );
or ( n86563 , C0 , n86531 , n86540 , n86561 , n86562 );
buf ( n86564 , n86563 );
buf ( n86565 , n86564 );
buf ( n86566 , n31655 );
buf ( n86567 , n31655 );
buf ( n86568 , n30987 );
buf ( n86569 , n30987 );
not ( n86570 , n34150 );
and ( n86571 , n86570 , n32698 );
not ( n86572 , n59105 );
and ( n86573 , n86572 , n32698 );
and ( n86574 , n32722 , n59105 );
or ( n86575 , n86573 , n86574 );
and ( n86576 , n86575 , n34150 );
or ( n86577 , n86571 , n86576 );
and ( n86578 , n86577 , n33381 );
not ( n86579 , n59113 );
not ( n86580 , n59105 );
and ( n86581 , n86580 , n32698 );
and ( n86582 , n42565 , n59105 );
or ( n86583 , n86581 , n86582 );
and ( n86584 , n86579 , n86583 );
and ( n86585 , n42565 , n59113 );
or ( n86586 , n86584 , n86585 );
and ( n86587 , n86586 , n33375 );
not ( n86588 , n32968 );
not ( n86589 , n59113 );
not ( n86590 , n59105 );
and ( n86591 , n86590 , n32698 );
and ( n86592 , n42565 , n59105 );
or ( n86593 , n86591 , n86592 );
and ( n86594 , n86589 , n86593 );
and ( n86595 , n42565 , n59113 );
or ( n86596 , n86594 , n86595 );
and ( n86597 , n86588 , n86596 );
not ( n86598 , n59133 );
not ( n86599 , n59135 );
and ( n86600 , n86599 , n86596 );
and ( n86601 , n42589 , n59135 );
or ( n86602 , n86600 , n86601 );
and ( n86603 , n86598 , n86602 );
and ( n86604 , n42597 , n59133 );
or ( n86605 , n86603 , n86604 );
and ( n86606 , n86605 , n32968 );
or ( n86607 , n86597 , n86606 );
and ( n86608 , n86607 , n33370 );
and ( n86609 , n32698 , n35062 );
or ( n86610 , C0 , n86578 , n86587 , n86608 , n86609 );
buf ( n86611 , n86610 );
buf ( n86612 , n86611 );
buf ( n86613 , n31655 );
buf ( n86614 , n31655 );
buf ( n86615 , n31655 );
not ( n86616 , n36587 );
and ( n86617 , n86616 , n36124 );
xor ( n86618 , n50193 , n50194 );
and ( n86619 , n86618 , n36587 );
or ( n86620 , n86617 , n86619 );
and ( n86621 , n86620 , n36596 );
not ( n86622 , n37485 );
and ( n86623 , n86622 , n37026 );
xor ( n86624 , n50243 , n50244 );
and ( n86625 , n86624 , n37485 );
or ( n86626 , n86623 , n86625 );
and ( n86627 , n86626 , n37494 );
and ( n86628 , n41841 , n37506 );
or ( n86629 , n86621 , n86627 , n86628 );
buf ( n86630 , n86629 );
buf ( n86631 , n86630 );
buf ( n86632 , n30987 );
buf ( n86633 , RI15b60a80_1163);
and ( n86634 , n86633 , n48531 );
and ( n86635 , n50826 , n39359 );
or ( n86636 , n86634 , n86635 );
buf ( n86637 , n86636 );
buf ( n86638 , n86637 );
xor ( n86639 , n54144 , n78381 );
and ( n86640 , n86639 , n33199 );
not ( n86641 , n48648 );
and ( n86642 , n86641 , n54144 );
and ( n86643 , n34429 , n48648 );
or ( n86644 , n86642 , n86643 );
and ( n86645 , n86644 , n32924 );
not ( n86646 , n48660 );
and ( n86647 , n86646 , n54144 );
and ( n86648 , n64077 , n48660 );
or ( n86649 , n86647 , n86648 );
and ( n86650 , n86649 , n33172 );
not ( n86651 , n48730 );
and ( n86652 , n86651 , n54144 );
xor ( n86653 , n58557 , n78400 );
and ( n86654 , n86653 , n48730 );
or ( n86655 , n86652 , n86654 );
and ( n86656 , n86655 , n33187 );
and ( n86657 , n54144 , n54713 );
or ( n86658 , n86640 , n86645 , n86650 , n86656 , n86657 );
and ( n86659 , n86658 , n33208 );
and ( n86660 , n54144 , n39805 );
or ( n86661 , C0 , n86659 , n86660 );
buf ( n86662 , n86661 );
buf ( n86663 , n86662 );
buf ( n86664 , n30987 );
buf ( n86665 , n31655 );
buf ( n86666 , n30987 );
buf ( n86667 , n31655 );
not ( n86668 , n41532 );
and ( n86669 , n86668 , n34367 );
and ( n86670 , n62428 , n41532 );
or ( n86671 , n86669 , n86670 );
buf ( n86672 , n86671 );
buf ( n86673 , n86672 );
buf ( n86674 , n30987 );
buf ( n86675 , n30987 );
not ( n86676 , n34150 );
and ( n86677 , n86676 , n32615 );
not ( n86678 , n59574 );
and ( n86679 , n86678 , n32615 );
and ( n86680 , n32655 , n59574 );
or ( n86681 , n86679 , n86680 );
and ( n86682 , n86681 , n34150 );
or ( n86683 , n86677 , n86682 );
and ( n86684 , n86683 , n33381 );
not ( n86685 , n59582 );
not ( n86686 , n59574 );
and ( n86687 , n86686 , n32615 );
and ( n86688 , n56044 , n59574 );
or ( n86689 , n86687 , n86688 );
and ( n86690 , n86685 , n86689 );
and ( n86691 , n56044 , n59582 );
or ( n86692 , n86690 , n86691 );
and ( n86693 , n86692 , n33375 );
not ( n86694 , n32968 );
not ( n86695 , n59582 );
not ( n86696 , n59574 );
and ( n86697 , n86696 , n32615 );
and ( n86698 , n56044 , n59574 );
or ( n86699 , n86697 , n86698 );
and ( n86700 , n86695 , n86699 );
and ( n86701 , n56044 , n59582 );
or ( n86702 , n86700 , n86701 );
and ( n86703 , n86694 , n86702 );
not ( n86704 , n59602 );
not ( n86705 , n59604 );
and ( n86706 , n86705 , n86702 );
and ( n86707 , n56068 , n59604 );
or ( n86708 , n86706 , n86707 );
and ( n86709 , n86704 , n86708 );
and ( n86710 , n56076 , n59602 );
or ( n86711 , n86709 , n86710 );
and ( n86712 , n86711 , n32968 );
or ( n86713 , n86703 , n86712 );
and ( n86714 , n86713 , n33370 );
and ( n86715 , n32615 , n35062 );
or ( n86716 , C0 , n86684 , n86693 , n86714 , n86715 );
buf ( n86717 , n86716 );
buf ( n86718 , n86717 );
buf ( n86719 , n31655 );
buf ( n86720 , n31655 );
buf ( n86721 , n31655 );
not ( n86722 , n46356 );
and ( n86723 , n86722 , n31280 );
not ( n86724 , n46362 );
and ( n86725 , n86724 , n31280 );
and ( n86726 , n31306 , n46362 );
or ( n86727 , n86725 , n86726 );
and ( n86728 , n86727 , n46356 );
or ( n86729 , n86723 , n86728 );
and ( n86730 , n86729 , n31649 );
not ( n86731 , n46393 );
not ( n86732 , n46362 );
and ( n86733 , n86732 , n31280 );
and ( n86734 , n58061 , n46362 );
or ( n86735 , n86733 , n86734 );
and ( n86736 , n86731 , n86735 );
and ( n86737 , n58061 , n46393 );
or ( n86738 , n86736 , n86737 );
and ( n86739 , n86738 , n31643 );
not ( n86740 , n31452 );
not ( n86741 , n46393 );
not ( n86742 , n46362 );
and ( n86743 , n86742 , n31280 );
and ( n86744 , n58061 , n46362 );
or ( n86745 , n86743 , n86744 );
and ( n86746 , n86741 , n86745 );
and ( n86747 , n58061 , n46393 );
or ( n86748 , n86746 , n86747 );
and ( n86749 , n86740 , n86748 );
not ( n86750 , n46550 );
not ( n86751 , n46554 );
and ( n86752 , n86751 , n86748 );
and ( n86753 , n58085 , n46554 );
or ( n86754 , n86752 , n86753 );
and ( n86755 , n86750 , n86754 );
and ( n86756 , n58093 , n46550 );
or ( n86757 , n86755 , n86756 );
and ( n86758 , n86757 , n31452 );
or ( n86759 , n86749 , n86758 );
and ( n86760 , n86759 , n31638 );
and ( n86761 , n31280 , n47277 );
or ( n86762 , C0 , n86730 , n86739 , n86760 , n86761 );
buf ( n86763 , n86762 );
buf ( n86764 , n86763 );
buf ( n86765 , n30987 );
and ( n86766 , n61466 , n32494 );
not ( n86767 , n46083 );
and ( n86768 , n86767 , n74198 );
not ( n86769 , n46290 );
and ( n86770 , n86769 , n46208 );
xor ( n86771 , n46297 , n46315 );
and ( n86772 , n86771 , n46290 );
or ( n86773 , n86770 , n86772 );
and ( n86774 , n86773 , n46083 );
or ( n86775 , n86768 , n86774 );
and ( n86776 , n86775 , n32421 );
not ( n86777 , n46326 );
and ( n86778 , n86777 , n74198 );
and ( n86779 , n86773 , n46326 );
or ( n86780 , n86778 , n86779 );
and ( n86781 , n86780 , n32417 );
and ( n86782 , n74198 , n46340 );
or ( n86783 , n86776 , n86781 , n86782 );
and ( n86784 , n86783 , n32456 );
and ( n86785 , n74198 , n46349 );
or ( n86786 , C0 , n86766 , n86784 , n86785 );
buf ( n86787 , n86786 );
buf ( n86788 , n86787 );
buf ( n86789 , n31655 );
buf ( n86790 , n31655 );
buf ( n86791 , n30987 );
xor ( n86792 , n33105 , n56361 );
and ( n86793 , n86792 , n33201 );
not ( n86794 , n41576 );
and ( n86795 , n86794 , n33105 );
and ( n86796 , n82803 , n41576 );
or ( n86797 , n86795 , n86796 );
and ( n86798 , n86797 , n33189 );
and ( n86799 , n33105 , n41592 );
or ( n86800 , n86793 , n86798 , n86799 );
and ( n86801 , n86800 , n33208 );
and ( n86802 , n33105 , n39805 );
or ( n86803 , C0 , n86801 , n86802 );
buf ( n86804 , n86803 );
buf ( n86805 , n86804 );
buf ( n86806 , n30987 );
buf ( n86807 , n31655 );
not ( n86808 , n50828 );
not ( n86809 , n50834 );
and ( n86810 , n86809 , n40597 );
and ( n86811 , n74778 , n50834 );
or ( n86812 , n86810 , n86811 );
and ( n86813 , n86808 , n86812 );
and ( n86814 , n86308 , n50828 );
or ( n86815 , n86813 , n86814 );
buf ( n86816 , n86815 );
buf ( n86817 , n86816 );
buf ( n86818 , n31655 );
xor ( n86819 , n34056 , n39929 );
and ( n86820 , n86819 , n31550 );
not ( n86821 , n39979 );
and ( n86822 , n86821 , n34056 );
buf ( n86823 , n31370 );
and ( n86824 , n86823 , n39979 );
or ( n86825 , n86822 , n86824 );
and ( n86826 , n86825 , n31538 );
and ( n86827 , n34056 , n40143 );
or ( n86828 , n86820 , n86826 , n86827 );
and ( n86829 , n86828 , n31557 );
and ( n86830 , n34056 , n40154 );
or ( n86831 , C0 , n86829 , n86830 );
buf ( n86832 , n86831 );
buf ( n86833 , n86832 );
not ( n86834 , n40163 );
and ( n86835 , n86834 , n32025 );
not ( n86836 , n57233 );
and ( n86837 , n86836 , n32025 );
and ( n86838 , n32147 , n57233 );
or ( n86839 , n86837 , n86838 );
and ( n86840 , n86839 , n40163 );
or ( n86841 , n86835 , n86840 );
and ( n86842 , n86841 , n32498 );
not ( n86843 , n57241 );
not ( n86844 , n57233 );
and ( n86845 , n86844 , n32025 );
and ( n86846 , n49314 , n57233 );
or ( n86847 , n86845 , n86846 );
and ( n86848 , n86843 , n86847 );
and ( n86849 , n49314 , n57241 );
or ( n86850 , n86848 , n86849 );
and ( n86851 , n86850 , n32473 );
not ( n86852 , n32475 );
not ( n86853 , n57241 );
not ( n86854 , n57233 );
and ( n86855 , n86854 , n32025 );
and ( n86856 , n49314 , n57233 );
or ( n86857 , n86855 , n86856 );
and ( n86858 , n86853 , n86857 );
and ( n86859 , n49314 , n57241 );
or ( n86860 , n86858 , n86859 );
and ( n86861 , n86852 , n86860 );
not ( n86862 , n57261 );
not ( n86863 , n57263 );
and ( n86864 , n86863 , n86860 );
and ( n86865 , n49340 , n57263 );
or ( n86866 , n86864 , n86865 );
and ( n86867 , n86862 , n86866 );
and ( n86868 , n49348 , n57261 );
or ( n86869 , n86867 , n86868 );
and ( n86870 , n86869 , n32475 );
or ( n86871 , n86861 , n86870 );
and ( n86872 , n86871 , n32486 );
and ( n86873 , n32025 , n41278 );
or ( n86874 , C0 , n86842 , n86851 , n86872 , n86873 );
buf ( n86875 , n86874 );
buf ( n86876 , n86875 );
buf ( n86877 , n30987 );
buf ( n86878 , n30987 );
not ( n86879 , n34150 );
and ( n86880 , n86879 , n32803 );
not ( n86881 , n57872 );
and ( n86882 , n86881 , n32803 );
and ( n86883 , n32823 , n57872 );
or ( n86884 , n86882 , n86883 );
and ( n86885 , n86884 , n34150 );
or ( n86886 , n86880 , n86885 );
and ( n86887 , n86886 , n33381 );
not ( n86888 , n57880 );
not ( n86889 , n57872 );
and ( n86890 , n86889 , n32803 );
and ( n86891 , n41464 , n57872 );
or ( n86892 , n86890 , n86891 );
and ( n86893 , n86888 , n86892 );
and ( n86894 , n41464 , n57880 );
or ( n86895 , n86893 , n86894 );
and ( n86896 , n86895 , n33375 );
not ( n86897 , n32968 );
not ( n86898 , n57880 );
not ( n86899 , n57872 );
and ( n86900 , n86899 , n32803 );
and ( n86901 , n41464 , n57872 );
or ( n86902 , n86900 , n86901 );
and ( n86903 , n86898 , n86902 );
and ( n86904 , n41464 , n57880 );
or ( n86905 , n86903 , n86904 );
and ( n86906 , n86897 , n86905 );
not ( n86907 , n57900 );
not ( n86908 , n57902 );
and ( n86909 , n86908 , n86905 );
and ( n86910 , n41490 , n57902 );
or ( n86911 , n86909 , n86910 );
and ( n86912 , n86907 , n86911 );
and ( n86913 , n41500 , n57900 );
or ( n86914 , n86912 , n86913 );
and ( n86915 , n86914 , n32968 );
or ( n86916 , n86906 , n86915 );
and ( n86917 , n86916 , n33370 );
and ( n86918 , n32803 , n35062 );
or ( n86919 , C0 , n86887 , n86896 , n86917 , n86918 );
buf ( n86920 , n86919 );
buf ( n86921 , n86920 );
buf ( n86922 , n30987 );
buf ( n86923 , n30987 );
buf ( n86924 , n31655 );
buf ( n86925 , n31655 );
not ( n86926 , n46356 );
and ( n86927 , n86926 , n31129 );
not ( n86928 , n47423 );
and ( n86929 , n86928 , n31129 );
and ( n86930 , n31138 , n47423 );
or ( n86931 , n86929 , n86930 );
and ( n86932 , n86931 , n46356 );
or ( n86933 , n86927 , n86932 );
and ( n86934 , n86933 , n31649 );
not ( n86935 , n47431 );
not ( n86936 , n47423 );
and ( n86937 , n86936 , n31129 );
and ( n86938 , n56920 , n47423 );
or ( n86939 , n86937 , n86938 );
and ( n86940 , n86935 , n86939 );
and ( n86941 , n56920 , n47431 );
or ( n86942 , n86940 , n86941 );
and ( n86943 , n86942 , n31643 );
not ( n86944 , n31452 );
not ( n86945 , n47431 );
not ( n86946 , n47423 );
and ( n86947 , n86946 , n31129 );
and ( n86948 , n56920 , n47423 );
or ( n86949 , n86947 , n86948 );
and ( n86950 , n86945 , n86949 );
and ( n86951 , n56920 , n47431 );
or ( n86952 , n86950 , n86951 );
and ( n86953 , n86944 , n86952 );
not ( n86954 , n47466 );
not ( n86955 , n47468 );
and ( n86956 , n86955 , n86952 );
and ( n86957 , n56946 , n47468 );
or ( n86958 , n86956 , n86957 );
and ( n86959 , n86954 , n86958 );
and ( n86960 , n56954 , n47466 );
or ( n86961 , n86959 , n86960 );
and ( n86962 , n86961 , n31452 );
or ( n86963 , n86953 , n86962 );
and ( n86964 , n86963 , n31638 );
and ( n86965 , n31129 , n47277 );
or ( n86966 , C0 , n86934 , n86943 , n86964 , n86965 );
buf ( n86967 , n86966 );
buf ( n86968 , n86967 );
buf ( n86969 , n31655 );
buf ( n86970 , n30987 );
buf ( n86971 , n30987 );
xor ( n86972 , n49589 , n60311 );
and ( n86973 , n86972 , n32433 );
not ( n86974 , n47331 );
and ( n86975 , n86974 , n49589 );
and ( n86976 , n85981 , n47331 );
or ( n86977 , n86975 , n86976 );
and ( n86978 , n86977 , n32413 );
and ( n86979 , n49589 , n47402 );
or ( n86980 , n86973 , n86978 , n86979 );
and ( n86981 , n86980 , n32456 );
and ( n86982 , n49589 , n47409 );
or ( n86983 , C0 , n86981 , n86982 );
buf ( n86984 , n86983 );
buf ( n86985 , n86984 );
buf ( n86986 , n31655 );
buf ( n86987 , n30987 );
not ( n86988 , n43755 );
and ( n86989 , n86988 , n43343 );
xor ( n86990 , n43759 , n43769 );
and ( n86991 , n86990 , n43755 );
or ( n86992 , n86989 , n86991 );
and ( n86993 , n86992 , n43774 );
not ( n86994 , n44663 );
and ( n86995 , n86994 , n44255 );
xor ( n86996 , n44667 , n44677 );
and ( n86997 , n86996 , n44663 );
or ( n86998 , n86995 , n86997 );
and ( n86999 , n86998 , n44682 );
and ( n87000 , n79658 , n44695 );
or ( n87001 , n86993 , n86999 , n87000 );
buf ( n87002 , n87001 );
buf ( n87003 , n87002 );
buf ( n87004 , n30987 );
buf ( n87005 , n31655 );
buf ( n87006 , n31655 );
and ( n87007 , n33488 , n46356 );
buf ( n87008 , n87007 );
and ( n87009 , n87008 , n31649 );
and ( n87010 , n52610 , n31647 );
and ( n87011 , n63734 , n31557 );
and ( n87012 , n31022 , n61220 );
or ( n87013 , C0 , n87009 , n87010 , n87011 , n87012 );
buf ( n87014 , n87013 );
buf ( n87015 , n87014 );
buf ( n87016 , n31655 );
buf ( n87017 , n30987 );
not ( n87018 , n38443 );
and ( n87019 , n87018 , n38184 );
xor ( n87020 , n53471 , n53498 );
and ( n87021 , n87020 , n38443 );
or ( n87022 , n87019 , n87021 );
and ( n87023 , n87022 , n38450 );
not ( n87024 , n39339 );
and ( n87025 , n87024 , n39084 );
xor ( n87026 , n53527 , n53554 );
and ( n87027 , n87026 , n39339 );
or ( n87028 , n87025 , n87027 );
and ( n87029 , n87028 , n39346 );
and ( n87030 , n40213 , n39359 );
or ( n87031 , n87023 , n87029 , n87030 );
buf ( n87032 , n87031 );
buf ( n87033 , n87032 );
buf ( n87034 , n31655 );
not ( n87035 , n31437 );
and ( n87036 , n87035 , n45272 );
and ( n87037 , n45790 , n31437 );
or ( n87038 , n87036 , n87037 );
and ( n87039 , n87038 , n31468 );
not ( n87040 , n44817 );
and ( n87041 , n87040 , n45272 );
not ( n87042 , n44994 );
and ( n87043 , n87042 , n44930 );
xor ( n87044 , n45001 , n45019 );
and ( n87045 , n87044 , n44994 );
or ( n87046 , n87043 , n87045 );
and ( n87047 , n87046 , n44817 );
or ( n87048 , n87041 , n87047 );
and ( n87049 , n87048 , n31521 );
and ( n87050 , n45272 , n42158 );
or ( n87051 , n87039 , n87049 , n87050 );
and ( n87052 , n87051 , n31557 );
and ( n87053 , n45272 , n40154 );
or ( n87054 , C0 , n87052 , n87053 );
buf ( n87055 , n87054 );
buf ( n87056 , n87055 );
and ( n87057 , n32300 , n50275 );
not ( n87058 , n50278 );
and ( n87059 , n87058 , n31736 );
and ( n87060 , n32300 , n50278 );
or ( n87061 , n87059 , n87060 );
and ( n87062 , n87061 , n32421 );
not ( n87063 , n50002 );
and ( n87064 , n87063 , n31736 );
and ( n87065 , n32300 , n50002 );
or ( n87066 , n87064 , n87065 );
and ( n87067 , n87066 , n32419 );
not ( n87068 , n50289 );
and ( n87069 , n87068 , n31736 );
and ( n87070 , n32300 , n50289 );
or ( n87071 , n87069 , n87070 );
and ( n87072 , n87071 , n32417 );
not ( n87073 , n50008 );
and ( n87074 , n87073 , n31736 );
and ( n87075 , n32300 , n50008 );
or ( n87076 , n87074 , n87075 );
and ( n87077 , n87076 , n32415 );
not ( n87078 , n47331 );
and ( n87079 , n87078 , n31736 );
and ( n87080 , n31895 , n47331 );
or ( n87081 , n87079 , n87080 );
and ( n87082 , n87081 , n32413 );
not ( n87083 , n50067 );
and ( n87084 , n87083 , n31736 );
and ( n87085 , n31895 , n50067 );
or ( n87086 , n87084 , n87085 );
and ( n87087 , n87086 , n32411 );
not ( n87088 , n31728 );
and ( n87089 , n87088 , n31736 );
and ( n87090 , n57953 , n31728 );
or ( n87091 , n87089 , n87090 );
and ( n87092 , n87091 , n32253 );
not ( n87093 , n32283 );
and ( n87094 , n87093 , n31736 );
and ( n87095 , n57966 , n32283 );
or ( n87096 , n87094 , n87095 );
and ( n87097 , n87096 , n32398 );
and ( n87098 , n32352 , n50334 );
or ( n87099 , n87057 , n87062 , n87067 , n87072 , n87077 , n87082 , n87087 , n87092 , n87097 , n87098 );
and ( n87100 , n87099 , n32456 );
and ( n87101 , n37581 , n32489 );
and ( n87102 , n31736 , n50345 );
or ( n87103 , C0 , n87100 , n87101 , n87102 );
buf ( n87104 , n87103 );
buf ( n87105 , n87104 );
buf ( n87106 , n30987 );
buf ( n87107 , n31655 );
buf ( n87108 , n30987 );
xor ( n87109 , n33111 , n52223 );
and ( n87110 , n87109 , n33201 );
not ( n87111 , n41576 );
and ( n87112 , n87111 , n33111 );
and ( n87113 , n81541 , n41576 );
or ( n87114 , n87112 , n87113 );
and ( n87115 , n87114 , n33189 );
and ( n87116 , n33111 , n41592 );
or ( n87117 , n87110 , n87115 , n87116 );
and ( n87118 , n87117 , n33208 );
and ( n87119 , n33111 , n39805 );
or ( n87120 , C0 , n87118 , n87119 );
buf ( n87121 , n87120 );
buf ( n87122 , n87121 );
buf ( n87123 , n30987 );
buf ( n87124 , n31655 );
not ( n87125 , n50828 );
not ( n87126 , n50834 );
and ( n87127 , n87126 , n40576 );
and ( n87128 , n59978 , n50834 );
or ( n87129 , n87127 , n87128 );
and ( n87130 , n87125 , n87129 );
and ( n87131 , n53319 , n50828 );
or ( n87132 , n87130 , n87131 );
buf ( n87133 , n87132 );
buf ( n87134 , n87133 );
buf ( n87135 , n70982 );
buf ( n87136 , n30987 );
not ( n87137 , n48765 );
and ( n87138 , n87137 , n33228 );
and ( n87139 , n85749 , n48765 );
or ( n87140 , n87138 , n87139 );
and ( n87141 , n87140 , n33180 );
not ( n87142 , n49054 );
and ( n87143 , n87142 , n33228 );
and ( n87144 , n85760 , n49054 );
or ( n87145 , n87143 , n87144 );
and ( n87146 , n87145 , n33178 );
and ( n87147 , n33228 , n49774 );
or ( n87148 , n87141 , n87146 , n87147 );
and ( n87149 , n87148 , n33208 );
and ( n87150 , n33307 , n33375 );
not ( n87151 , n32968 );
and ( n87152 , n87151 , n33307 );
xor ( n87153 , n33228 , n53901 );
and ( n87154 , n87153 , n32968 );
or ( n87155 , n87152 , n87154 );
and ( n87156 , n87155 , n33370 );
and ( n87157 , n32991 , n35056 );
and ( n87158 , n33228 , n49794 );
or ( n87159 , C0 , n87149 , n87150 , n87156 , n87157 , n87158 );
buf ( n87160 , n87159 );
buf ( n87161 , n87160 );
buf ( n87162 , n31655 );
buf ( n87163 , n30987 );
buf ( n87164 , n31655 );
and ( n87165 , n46022 , n32500 );
not ( n87166 , n35211 );
and ( n87167 , n87166 , n37541 );
buf ( n87168 , n87167 );
and ( n87169 , n87168 , n32421 );
not ( n87170 , n35245 );
and ( n87171 , n87170 , n37541 );
buf ( n87172 , n87171 );
and ( n87173 , n87172 , n32419 );
not ( n87174 , n35278 );
and ( n87175 , n87174 , n37541 );
not ( n87176 , n35295 );
and ( n87177 , n87176 , n49571 );
xor ( n87178 , n37541 , n49545 );
and ( n87179 , n87178 , n35295 );
or ( n87180 , n87177 , n87179 );
and ( n87181 , n87180 , n35278 );
or ( n87182 , n87175 , n87181 );
and ( n87183 , n87182 , n32417 );
not ( n87184 , n35331 );
and ( n87185 , n87184 , n37541 );
not ( n87186 , n35294 );
not ( n87187 , n45995 );
and ( n87188 , n87187 , n49571 );
xor ( n87189 , n49572 , n49631 );
and ( n87190 , n87189 , n45995 );
or ( n87191 , n87188 , n87190 );
and ( n87192 , n87186 , n87191 );
and ( n87193 , n87178 , n35294 );
or ( n87194 , n87192 , n87193 );
and ( n87195 , n87194 , n35331 );
or ( n87196 , n87185 , n87195 );
and ( n87197 , n87196 , n32415 );
and ( n87198 , n37541 , n35354 );
or ( n87199 , n87169 , n87173 , n87183 , n87197 , n87198 );
and ( n87200 , n87199 , n32456 );
not ( n87201 , n32475 );
not ( n87202 , n46060 );
and ( n87203 , n87202 , n47745 );
xor ( n87204 , n49662 , n49725 );
and ( n87205 , n87204 , n46060 );
or ( n87206 , n87203 , n87205 );
and ( n87207 , n87201 , n87206 );
and ( n87208 , n37541 , n32475 );
or ( n87209 , n87207 , n87208 );
and ( n87210 , n87209 , n32486 );
and ( n87211 , n37541 , n35367 );
or ( n87212 , C0 , n87165 , n87200 , n87210 , C0 , n87211 );
buf ( n87213 , n87212 );
buf ( n87214 , n87213 );
buf ( n87215 , n31655 );
buf ( n87216 , n81144 );
xor ( n87217 , n35437 , n39945 );
and ( n87218 , n87217 , n31550 );
not ( n87219 , n39979 );
and ( n87220 , n87219 , n35437 );
xor ( n87221 , n40069 , n40127 );
and ( n87222 , n87221 , n39979 );
or ( n87223 , n87220 , n87222 );
and ( n87224 , n87223 , n31538 );
and ( n87225 , n35437 , n40143 );
or ( n87226 , n87218 , n87224 , n87225 );
and ( n87227 , n87226 , n31557 );
and ( n87228 , n35437 , n40154 );
or ( n87229 , C0 , n87227 , n87228 );
buf ( n87230 , n87229 );
buf ( n87231 , n87230 );
not ( n87232 , n40163 );
and ( n87233 , n87232 , n32029 );
not ( n87234 , n75905 );
and ( n87235 , n87234 , n32029 );
and ( n87236 , n32147 , n75905 );
or ( n87237 , n87235 , n87236 );
and ( n87238 , n87237 , n40163 );
or ( n87239 , n87233 , n87238 );
and ( n87240 , n87239 , n32498 );
not ( n87241 , n75913 );
not ( n87242 , n75905 );
and ( n87243 , n87242 , n32029 );
and ( n87244 , n49314 , n75905 );
or ( n87245 , n87243 , n87244 );
and ( n87246 , n87241 , n87245 );
and ( n87247 , n49314 , n75913 );
or ( n87248 , n87246 , n87247 );
and ( n87249 , n87248 , n32473 );
not ( n87250 , n32475 );
not ( n87251 , n75913 );
not ( n87252 , n75905 );
and ( n87253 , n87252 , n32029 );
and ( n87254 , n49314 , n75905 );
or ( n87255 , n87253 , n87254 );
and ( n87256 , n87251 , n87255 );
and ( n87257 , n49314 , n75913 );
or ( n87258 , n87256 , n87257 );
and ( n87259 , n87250 , n87258 );
not ( n87260 , n75933 );
not ( n87261 , n75935 );
and ( n87262 , n87261 , n87258 );
and ( n87263 , n49340 , n75935 );
or ( n87264 , n87262 , n87263 );
and ( n87265 , n87260 , n87264 );
and ( n87266 , n49348 , n75933 );
or ( n87267 , n87265 , n87266 );
and ( n87268 , n87267 , n32475 );
or ( n87269 , n87259 , n87268 );
and ( n87270 , n87269 , n32486 );
and ( n87271 , n32029 , n41278 );
or ( n87272 , C0 , n87240 , n87249 , n87270 , n87271 );
buf ( n87273 , n87272 );
buf ( n87274 , n87273 );
buf ( n87275 , n30987 );
buf ( n87276 , n30987 );
buf ( n87277 , n31655 );
not ( n87278 , n36587 );
and ( n87279 , n87278 , n36209 );
xor ( n87280 , n50188 , n50199 );
and ( n87281 , n87280 , n36587 );
or ( n87282 , n87279 , n87281 );
and ( n87283 , n87282 , n36596 );
not ( n87284 , n37485 );
and ( n87285 , n87284 , n37111 );
xor ( n87286 , n50238 , n50249 );
and ( n87287 , n87286 , n37485 );
or ( n87288 , n87285 , n87287 );
and ( n87289 , n87288 , n37494 );
and ( n87290 , n41846 , n37506 );
or ( n87291 , n87283 , n87289 , n87290 );
buf ( n87292 , n87291 );
buf ( n87293 , n87292 );
buf ( n87294 , n30987 );
not ( n87295 , n35292 );
and ( n87296 , n87295 , n32442 );
buf ( n87297 , n35292 );
or ( n87298 , n87296 , n87297 );
and ( n87299 , n87298 , n32494 );
not ( n87300 , n76230 );
not ( n87301 , n76232 );
and ( n87302 , n87301 , n32442 );
buf ( n87303 , n76232 );
or ( n87304 , n87302 , n87303 );
and ( n87305 , n87304 , n32417 );
and ( n87306 , n32442 , n76244 );
or ( n87307 , n87305 , n87306 );
and ( n87308 , n87300 , n87307 );
buf ( n87309 , n76230 );
or ( n87310 , n87308 , n87309 );
and ( n87311 , n87310 , n32456 );
buf ( n87312 , n32473 );
not ( n87313 , n76252 );
and ( n87314 , n87313 , n32492 );
and ( n87315 , n32475 , n32486 );
or ( n87316 , C0 , C0 , C0 , n87299 , n87311 , n87312 , n87314 , n87315 , C0 , C0 );
buf ( n87317 , n87316 );
buf ( n87318 , n87317 );
buf ( n87319 , n31655 );
not ( n87320 , n46356 );
and ( n87321 , n87320 , n31199 );
not ( n87322 , n47423 );
and ( n87323 , n87322 , n31199 );
and ( n87324 , n31205 , n47423 );
or ( n87325 , n87323 , n87324 );
and ( n87326 , n87325 , n46356 );
or ( n87327 , n87321 , n87326 );
and ( n87328 , n87327 , n31649 );
not ( n87329 , n47431 );
not ( n87330 , n47423 );
and ( n87331 , n87330 , n31199 );
and ( n87332 , n50125 , n47423 );
or ( n87333 , n87331 , n87332 );
and ( n87334 , n87329 , n87333 );
and ( n87335 , n50125 , n47431 );
or ( n87336 , n87334 , n87335 );
and ( n87337 , n87336 , n31643 );
not ( n87338 , n31452 );
not ( n87339 , n47431 );
not ( n87340 , n47423 );
and ( n87341 , n87340 , n31199 );
and ( n87342 , n50125 , n47423 );
or ( n87343 , n87341 , n87342 );
and ( n87344 , n87339 , n87343 );
and ( n87345 , n50125 , n47431 );
or ( n87346 , n87344 , n87345 );
and ( n87347 , n87338 , n87346 );
not ( n87348 , n47466 );
not ( n87349 , n47468 );
and ( n87350 , n87349 , n87346 );
and ( n87351 , n50151 , n47468 );
or ( n87352 , n87350 , n87351 );
and ( n87353 , n87348 , n87352 );
and ( n87354 , n50159 , n47466 );
or ( n87355 , n87353 , n87354 );
and ( n87356 , n87355 , n31452 );
or ( n87357 , n87347 , n87356 );
and ( n87358 , n87357 , n31638 );
and ( n87359 , n31199 , n47277 );
or ( n87360 , C0 , n87328 , n87337 , n87358 , n87359 );
buf ( n87361 , n87360 );
buf ( n87362 , n87361 );
buf ( n87363 , n30987 );
buf ( n87364 , n30987 );
xor ( n87365 , n49593 , n60309 );
and ( n87366 , n87365 , n32433 );
not ( n87367 , n47331 );
and ( n87368 , n87367 , n49593 );
and ( n87369 , n50086 , n47331 );
or ( n87370 , n87368 , n87369 );
and ( n87371 , n87370 , n32413 );
and ( n87372 , n49593 , n47402 );
or ( n87373 , n87366 , n87371 , n87372 );
and ( n87374 , n87373 , n32456 );
and ( n87375 , n49593 , n47409 );
or ( n87376 , C0 , n87374 , n87375 );
buf ( n87377 , n87376 );
buf ( n87378 , n87377 );
buf ( n87379 , n31655 );
buf ( n87380 , n30987 );
buf ( n87381 , n75453 );
buf ( n87382 , n31655 );
not ( n87383 , n48765 );
and ( n87384 , n87383 , n33227 );
and ( n87385 , n62345 , n48765 );
or ( n87386 , n87384 , n87385 );
and ( n87387 , n87386 , n33180 );
not ( n87388 , n49054 );
and ( n87389 , n87388 , n33227 );
and ( n87390 , n62356 , n49054 );
or ( n87391 , n87389 , n87390 );
and ( n87392 , n87391 , n33178 );
and ( n87393 , n33227 , n49774 );
or ( n87394 , n87387 , n87392 , n87393 );
and ( n87395 , n87394 , n33208 );
and ( n87396 , n33305 , n33375 );
not ( n87397 , n32968 );
and ( n87398 , n87397 , n33305 );
xor ( n87399 , n33227 , n53902 );
and ( n87400 , n87399 , n32968 );
or ( n87401 , n87398 , n87400 );
and ( n87402 , n87401 , n33370 );
and ( n87403 , n32990 , n35056 );
and ( n87404 , n33227 , n49794 );
or ( n87405 , C0 , n87395 , n87396 , n87402 , n87403 , n87404 );
buf ( n87406 , n87405 );
buf ( n87407 , n87406 );
buf ( n87408 , n30987 );
buf ( n87409 , n31655 );
and ( n87410 , n46023 , n32500 );
not ( n87411 , n35211 );
and ( n87412 , n87411 , n37543 );
buf ( n87413 , n87412 );
and ( n87414 , n87413 , n32421 );
not ( n87415 , n35245 );
and ( n87416 , n87415 , n37543 );
buf ( n87417 , n87416 );
and ( n87418 , n87417 , n32419 );
not ( n87419 , n35278 );
and ( n87420 , n87419 , n37543 );
not ( n87421 , n35295 );
and ( n87422 , n87421 , n49573 );
xor ( n87423 , n37543 , n49544 );
and ( n87424 , n87423 , n35295 );
or ( n87425 , n87422 , n87424 );
and ( n87426 , n87425 , n35278 );
or ( n87427 , n87420 , n87426 );
and ( n87428 , n87427 , n32417 );
not ( n87429 , n35331 );
and ( n87430 , n87429 , n37543 );
not ( n87431 , n35294 );
not ( n87432 , n45995 );
and ( n87433 , n87432 , n49573 );
xor ( n87434 , n49574 , n49630 );
and ( n87435 , n87434 , n45995 );
or ( n87436 , n87433 , n87435 );
and ( n87437 , n87431 , n87436 );
and ( n87438 , n87423 , n35294 );
or ( n87439 , n87437 , n87438 );
and ( n87440 , n87439 , n35331 );
or ( n87441 , n87430 , n87440 );
and ( n87442 , n87441 , n32415 );
and ( n87443 , n37543 , n35354 );
or ( n87444 , n87414 , n87418 , n87428 , n87442 , n87443 );
and ( n87445 , n87444 , n32456 );
not ( n87446 , n32475 );
not ( n87447 , n46060 );
and ( n87448 , n87447 , n49663 );
xor ( n87449 , n49664 , n49724 );
and ( n87450 , n87449 , n46060 );
or ( n87451 , n87448 , n87450 );
and ( n87452 , n87446 , n87451 );
and ( n87453 , n37543 , n32475 );
or ( n87454 , n87452 , n87453 );
and ( n87455 , n87454 , n32486 );
and ( n87456 , n37543 , n35367 );
or ( n87457 , C0 , n87410 , n87445 , n87455 , C0 , n87456 );
buf ( n87458 , n87457 );
buf ( n87459 , n87458 );
buf ( n87460 , n31655 );
xor ( n87461 , n41782 , n44789 );
and ( n87462 , n87461 , n31548 );
not ( n87463 , n44807 );
and ( n87464 , n87463 , n41782 );
and ( n87465 , n42094 , n44807 );
or ( n87466 , n87464 , n87465 );
and ( n87467 , n87466 , n31408 );
not ( n87468 , n44817 );
and ( n87469 , n87468 , n41782 );
not ( n87470 , n41835 );
and ( n87471 , n87470 , n62425 );
and ( n87472 , n82209 , n41835 );
or ( n87473 , n87471 , n87472 );
and ( n87474 , n87473 , n44817 );
or ( n87475 , n87469 , n87474 );
and ( n87476 , n87475 , n31521 );
not ( n87477 , n45059 );
and ( n87478 , n87477 , n41782 );
and ( n87479 , n83827 , n45059 );
or ( n87480 , n87478 , n87479 );
and ( n87481 , n87480 , n31536 );
and ( n87482 , n41782 , n45148 );
or ( n87483 , n87462 , n87467 , n87476 , n87481 , n87482 );
and ( n87484 , n87483 , n31557 );
and ( n87485 , n41782 , n40154 );
or ( n87486 , C0 , n87484 , n87485 );
buf ( n87487 , n87486 );
buf ( n87488 , n87487 );
not ( n87489 , n40163 );
and ( n87490 , n87489 , n31984 );
not ( n87491 , n49298 );
and ( n87492 , n87491 , n31984 );
and ( n87493 , n32165 , n49298 );
or ( n87494 , n87492 , n87493 );
and ( n87495 , n87494 , n40163 );
or ( n87496 , n87490 , n87495 );
and ( n87497 , n87496 , n32498 );
not ( n87498 , n49306 );
not ( n87499 , n49298 );
and ( n87500 , n87499 , n31984 );
and ( n87501 , n59005 , n49298 );
or ( n87502 , n87500 , n87501 );
and ( n87503 , n87498 , n87502 );
and ( n87504 , n59005 , n49306 );
or ( n87505 , n87503 , n87504 );
and ( n87506 , n87505 , n32473 );
not ( n87507 , n32475 );
not ( n87508 , n49306 );
not ( n87509 , n49298 );
and ( n87510 , n87509 , n31984 );
and ( n87511 , n59005 , n49298 );
or ( n87512 , n87510 , n87511 );
and ( n87513 , n87508 , n87512 );
and ( n87514 , n59005 , n49306 );
or ( n87515 , n87513 , n87514 );
and ( n87516 , n87507 , n87515 );
not ( n87517 , n49331 );
not ( n87518 , n49333 );
and ( n87519 , n87518 , n87515 );
and ( n87520 , n59029 , n49333 );
or ( n87521 , n87519 , n87520 );
and ( n87522 , n87517 , n87521 );
and ( n87523 , n59037 , n49331 );
or ( n87524 , n87522 , n87523 );
and ( n87525 , n87524 , n32475 );
or ( n87526 , n87516 , n87525 );
and ( n87527 , n87526 , n32486 );
and ( n87528 , n31984 , n41278 );
or ( n87529 , C0 , n87497 , n87506 , n87527 , n87528 );
buf ( n87530 , n87529 );
buf ( n87531 , n87530 );
buf ( n87532 , n30987 );
buf ( n87533 , n30987 );
buf ( n87534 , n31655 );
and ( n87535 , n81623 , n31645 );
not ( n87536 , n45274 );
and ( n87537 , n87536 , n74228 );
buf ( n87538 , n87537 );
and ( n87539 , n87538 , n31373 );
not ( n87540 , n45280 );
and ( n87541 , n87540 , n74228 );
and ( n87542 , n81629 , n45280 );
or ( n87543 , n87541 , n87542 );
and ( n87544 , n87543 , n31468 );
and ( n87545 , n74228 , n45802 );
or ( n87546 , n87539 , n87544 , n87545 );
and ( n87547 , n87546 , n31557 );
and ( n87548 , n74228 , n45808 );
or ( n87549 , C0 , n87535 , n87547 , n87548 );
buf ( n87550 , n87549 );
buf ( n87551 , n87550 );
not ( n87552 , n40163 );
and ( n87553 , n87552 , n31976 );
not ( n87554 , n45227 );
and ( n87555 , n87554 , n31976 );
and ( n87556 , n32165 , n45227 );
or ( n87557 , n87555 , n87556 );
and ( n87558 , n87557 , n40163 );
or ( n87559 , n87553 , n87558 );
and ( n87560 , n87559 , n32498 );
not ( n87561 , n45235 );
not ( n87562 , n45227 );
and ( n87563 , n87562 , n31976 );
and ( n87564 , n59005 , n45227 );
or ( n87565 , n87563 , n87564 );
and ( n87566 , n87561 , n87565 );
and ( n87567 , n59005 , n45235 );
or ( n87568 , n87566 , n87567 );
and ( n87569 , n87568 , n32473 );
not ( n87570 , n32475 );
not ( n87571 , n45235 );
not ( n87572 , n45227 );
and ( n87573 , n87572 , n31976 );
and ( n87574 , n59005 , n45227 );
or ( n87575 , n87573 , n87574 );
and ( n87576 , n87571 , n87575 );
and ( n87577 , n59005 , n45235 );
or ( n87578 , n87576 , n87577 );
and ( n87579 , n87570 , n87578 );
not ( n87580 , n45255 );
not ( n87581 , n45257 );
and ( n87582 , n87581 , n87578 );
and ( n87583 , n59029 , n45257 );
or ( n87584 , n87582 , n87583 );
and ( n87585 , n87580 , n87584 );
and ( n87586 , n59037 , n45255 );
or ( n87587 , n87585 , n87586 );
and ( n87588 , n87587 , n32475 );
or ( n87589 , n87579 , n87588 );
and ( n87590 , n87589 , n32486 );
and ( n87591 , n31976 , n41278 );
or ( n87592 , C0 , n87560 , n87569 , n87590 , n87591 );
buf ( n87593 , n87592 );
buf ( n87594 , n87593 );
buf ( n87595 , n30987 );
buf ( n87596 , n30987 );
buf ( n87597 , n31655 );
xor ( n87598 , n34044 , n39935 );
and ( n87599 , n87598 , n31550 );
not ( n87600 , n39979 );
and ( n87601 , n87600 , n34044 );
and ( n87602 , n76137 , n39979 );
or ( n87603 , n87601 , n87602 );
and ( n87604 , n87603 , n31538 );
and ( n87605 , n34044 , n40143 );
or ( n87606 , n87599 , n87604 , n87605 );
and ( n87607 , n87606 , n31557 );
and ( n87608 , n34044 , n40154 );
or ( n87609 , C0 , n87607 , n87608 );
buf ( n87610 , n87609 );
buf ( n87611 , n87610 );
not ( n87612 , n40163 );
and ( n87613 , n87612 , n31957 );
not ( n87614 , n42238 );
and ( n87615 , n87614 , n31957 );
and ( n87616 , n32183 , n42238 );
or ( n87617 , n87615 , n87616 );
and ( n87618 , n87617 , n40163 );
or ( n87619 , n87613 , n87618 );
and ( n87620 , n87619 , n32498 );
not ( n87621 , n42247 );
not ( n87622 , n42238 );
and ( n87623 , n87622 , n31957 );
and ( n87624 , n45178 , n42238 );
or ( n87625 , n87623 , n87624 );
and ( n87626 , n87621 , n87625 );
and ( n87627 , n45178 , n42247 );
or ( n87628 , n87626 , n87627 );
and ( n87629 , n87628 , n32473 );
not ( n87630 , n32475 );
not ( n87631 , n42247 );
not ( n87632 , n42238 );
and ( n87633 , n87632 , n31957 );
and ( n87634 , n45178 , n42238 );
or ( n87635 , n87633 , n87634 );
and ( n87636 , n87631 , n87635 );
and ( n87637 , n45178 , n42247 );
or ( n87638 , n87636 , n87637 );
and ( n87639 , n87630 , n87638 );
not ( n87640 , n42273 );
not ( n87641 , n42276 );
and ( n87642 , n87641 , n87638 );
and ( n87643 , n45206 , n42276 );
or ( n87644 , n87642 , n87643 );
and ( n87645 , n87640 , n87644 );
and ( n87646 , n45214 , n42273 );
or ( n87647 , n87645 , n87646 );
and ( n87648 , n87647 , n32475 );
or ( n87649 , n87639 , n87648 );
and ( n87650 , n87649 , n32486 );
and ( n87651 , n31957 , n41278 );
or ( n87652 , C0 , n87620 , n87629 , n87650 , n87651 );
buf ( n87653 , n87652 );
buf ( n87654 , n87653 );
buf ( n87655 , n30987 );
buf ( n87656 , n30987 );
buf ( n87657 , n31655 );
xor ( n87658 , n39467 , n54971 );
and ( n87659 , n87658 , n33199 );
not ( n87660 , n48648 );
and ( n87661 , n87660 , n39467 );
and ( n87662 , n34379 , n48648 );
or ( n87663 , n87661 , n87662 );
and ( n87664 , n87663 , n32924 );
not ( n87665 , n48660 );
and ( n87666 , n87665 , n39467 );
not ( n87667 , n39584 );
and ( n87668 , n87667 , n73768 );
and ( n87669 , n86336 , n39584 );
or ( n87670 , n87668 , n87669 );
and ( n87671 , n87670 , n48660 );
or ( n87672 , n87666 , n87671 );
and ( n87673 , n87672 , n33172 );
not ( n87674 , n48730 );
and ( n87675 , n87674 , n39467 );
and ( n87676 , n32603 , n52252 );
and ( n87677 , n32607 , n52254 );
and ( n87678 , n32611 , n52256 );
and ( n87679 , n32615 , n52258 );
and ( n87680 , n32618 , n52260 );
and ( n87681 , n32622 , n52262 );
and ( n87682 , n32625 , n52264 );
and ( n87683 , n32628 , n52266 );
and ( n87684 , n32631 , n52268 );
and ( n87685 , n32634 , n52270 );
and ( n87686 , n32637 , n52272 );
and ( n87687 , n32640 , n52274 );
and ( n87688 , n32643 , n52276 );
and ( n87689 , n32646 , n52278 );
and ( n87690 , n32649 , n52280 );
and ( n87691 , n32652 , n52282 );
or ( n87692 , n87676 , n87677 , n87678 , n87679 , n87680 , n87681 , n87682 , n87683 , n87684 , n87685 , n87686 , n87687 , n87688 , n87689 , n87690 , n87691 );
and ( n87693 , n87692 , n48730 );
or ( n87694 , n87675 , n87693 );
and ( n87695 , n87694 , n33187 );
and ( n87696 , n39467 , n54713 );
or ( n87697 , n87659 , n87664 , n87673 , n87695 , n87696 );
and ( n87698 , n87697 , n33208 );
and ( n87699 , n39467 , n39805 );
or ( n87700 , C0 , n87698 , n87699 );
buf ( n87701 , n87700 );
buf ( n87702 , n87701 );
buf ( n87703 , n30987 );
buf ( n87704 , n30987 );
buf ( n87705 , n31655 );
not ( n87706 , n41532 );
and ( n87707 , n87706 , n34417 );
and ( n87708 , n35533 , n41532 );
or ( n87709 , n87707 , n87708 );
buf ( n87710 , n87709 );
buf ( n87711 , n87710 );
buf ( n87712 , n42734 );
buf ( n87713 , n42736 );
buf ( n87714 , n66430 );
or ( n87715 , n87712 , n87713 , n87714 , C0 );
and ( n87716 , n87715 , n42771 );
buf ( n87717 , n42734 );
buf ( n87718 , n42736 );
buf ( n87719 , n66430 );
or ( n87720 , C0 , n87717 , n87718 , n87719 , C0 );
and ( n87721 , n87720 , n42806 );
buf ( n87722 , n42734 );
buf ( n87723 , n42736 );
buf ( n87724 , n66430 );
or ( n87725 , C0 , n87722 , n87723 , n87724 , C0 );
and ( n87726 , n87725 , n42842 );
or ( n87727 , C0 , n87716 , n87721 , n87726 );
buf ( n87728 , n87727 );
buf ( n87729 , n87728 );
buf ( n87730 , n30987 );
buf ( n87731 , n31655 );
buf ( n87732 , n30987 );
buf ( n87733 , n31655 );
buf ( n87734 , n30987 );
not ( n87735 , n34150 );
and ( n87736 , n87735 , n32753 );
not ( n87737 , n56239 );
and ( n87738 , n87737 , n32753 );
and ( n87739 , n32755 , n56239 );
or ( n87740 , n87738 , n87739 );
and ( n87741 , n87740 , n34150 );
or ( n87742 , n87736 , n87741 );
and ( n87743 , n87742 , n33381 );
not ( n87744 , n56247 );
not ( n87745 , n56239 );
and ( n87746 , n87745 , n32753 );
and ( n87747 , n35083 , n56239 );
or ( n87748 , n87746 , n87747 );
and ( n87749 , n87744 , n87748 );
and ( n87750 , n35083 , n56247 );
or ( n87751 , n87749 , n87750 );
and ( n87752 , n87751 , n33375 );
not ( n87753 , n32968 );
not ( n87754 , n56247 );
not ( n87755 , n56239 );
and ( n87756 , n87755 , n32753 );
and ( n87757 , n35083 , n56239 );
or ( n87758 , n87756 , n87757 );
and ( n87759 , n87754 , n87758 );
and ( n87760 , n35083 , n56247 );
or ( n87761 , n87759 , n87760 );
and ( n87762 , n87753 , n87761 );
not ( n87763 , n56267 );
not ( n87764 , n56269 );
and ( n87765 , n87764 , n87761 );
and ( n87766 , n35107 , n56269 );
or ( n87767 , n87765 , n87766 );
and ( n87768 , n87763 , n87767 );
and ( n87769 , n35115 , n56267 );
or ( n87770 , n87768 , n87769 );
and ( n87771 , n87770 , n32968 );
or ( n87772 , n87762 , n87771 );
and ( n87773 , n87772 , n33370 );
and ( n87774 , n32753 , n35062 );
or ( n87775 , C0 , n87743 , n87752 , n87773 , n87774 );
buf ( n87776 , n87775 );
buf ( n87777 , n87776 );
not ( n87778 , n34150 );
and ( n87779 , n87778 , n32779 );
not ( n87780 , n56192 );
and ( n87781 , n87780 , n32779 );
and ( n87782 , n32789 , n56192 );
or ( n87783 , n87781 , n87782 );
and ( n87784 , n87783 , n34150 );
or ( n87785 , n87779 , n87784 );
and ( n87786 , n87785 , n33381 );
not ( n87787 , n56200 );
not ( n87788 , n56192 );
and ( n87789 , n87788 , n32779 );
and ( n87790 , n34301 , n56192 );
or ( n87791 , n87789 , n87790 );
and ( n87792 , n87787 , n87791 );
and ( n87793 , n34301 , n56200 );
or ( n87794 , n87792 , n87793 );
and ( n87795 , n87794 , n33375 );
not ( n87796 , n32968 );
not ( n87797 , n56200 );
not ( n87798 , n56192 );
and ( n87799 , n87798 , n32779 );
and ( n87800 , n34301 , n56192 );
or ( n87801 , n87799 , n87800 );
and ( n87802 , n87797 , n87801 );
and ( n87803 , n34301 , n56200 );
or ( n87804 , n87802 , n87803 );
and ( n87805 , n87796 , n87804 );
not ( n87806 , n56220 );
not ( n87807 , n56222 );
and ( n87808 , n87807 , n87804 );
and ( n87809 , n34761 , n56222 );
or ( n87810 , n87808 , n87809 );
and ( n87811 , n87806 , n87810 );
and ( n87812 , n35050 , n56220 );
or ( n87813 , n87811 , n87812 );
and ( n87814 , n87813 , n32968 );
or ( n87815 , n87805 , n87814 );
and ( n87816 , n87815 , n33370 );
and ( n87817 , n32779 , n35062 );
or ( n87818 , C0 , n87786 , n87795 , n87816 , n87817 );
buf ( n87819 , n87818 );
buf ( n87820 , n87819 );
buf ( n87821 , n30987 );
buf ( n87822 , n31655 );
buf ( n87823 , n31655 );
buf ( n87824 , n31655 );
buf ( n87825 , n30987 );
not ( n87826 , n46356 );
and ( n87827 , n87826 , n31170 );
not ( n87828 , n60564 );
and ( n87829 , n87828 , n31170 );
and ( n87830 , n31172 , n60564 );
or ( n87831 , n87829 , n87830 );
and ( n87832 , n87831 , n46356 );
or ( n87833 , n87827 , n87832 );
and ( n87834 , n87833 , n31649 );
not ( n87835 , n60572 );
not ( n87836 , n60564 );
and ( n87837 , n87836 , n31170 );
and ( n87838 , n46495 , n60564 );
or ( n87839 , n87837 , n87838 );
and ( n87840 , n87835 , n87839 );
and ( n87841 , n46495 , n60572 );
or ( n87842 , n87840 , n87841 );
and ( n87843 , n87842 , n31643 );
not ( n87844 , n31452 );
not ( n87845 , n60572 );
not ( n87846 , n60564 );
and ( n87847 , n87846 , n31170 );
and ( n87848 , n46495 , n60564 );
or ( n87849 , n87847 , n87848 );
and ( n87850 , n87845 , n87849 );
and ( n87851 , n46495 , n60572 );
or ( n87852 , n87850 , n87851 );
and ( n87853 , n87844 , n87852 );
not ( n87854 , n60592 );
not ( n87855 , n60594 );
and ( n87856 , n87855 , n87852 );
and ( n87857 , n46984 , n60594 );
or ( n87858 , n87856 , n87857 );
and ( n87859 , n87854 , n87858 );
and ( n87860 , n47267 , n60592 );
or ( n87861 , n87859 , n87860 );
and ( n87862 , n87861 , n31452 );
or ( n87863 , n87853 , n87862 );
and ( n87864 , n87863 , n31638 );
and ( n87865 , n31170 , n47277 );
or ( n87866 , C0 , n87834 , n87843 , n87864 , n87865 );
buf ( n87867 , n87866 );
buf ( n87868 , n87867 );
buf ( n87869 , n30987 );
and ( n87870 , n49563 , n60324 );
and ( n87871 , n49521 , n87870 );
xor ( n87872 , n45995 , n87871 );
and ( n87873 , n87872 , n32433 );
not ( n87874 , n47331 );
and ( n87875 , n87874 , n45995 );
buf ( n87876 , n87875 );
and ( n87877 , n87876 , n32413 );
and ( n87878 , n45995 , n47402 );
or ( n87879 , n87873 , n87877 , n87878 );
and ( n87880 , n87879 , n32456 );
and ( n87881 , n45995 , n47409 );
or ( n87882 , C0 , n87880 , n87881 );
buf ( n87883 , n87882 );
buf ( n87884 , n87883 );
buf ( n87885 , n31655 );
buf ( n87886 , n35538 );
buf ( n87887 , n30987 );
not ( n87888 , n48765 );
and ( n87889 , n87888 , n33229 );
and ( n87890 , n64487 , n48765 );
or ( n87891 , n87889 , n87890 );
and ( n87892 , n87891 , n33180 );
not ( n87893 , n49054 );
and ( n87894 , n87893 , n33229 );
and ( n87895 , n64498 , n49054 );
or ( n87896 , n87894 , n87895 );
and ( n87897 , n87896 , n33178 );
and ( n87898 , n33229 , n49774 );
or ( n87899 , n87892 , n87897 , n87898 );
and ( n87900 , n87899 , n33208 );
and ( n87901 , n33309 , n33375 );
not ( n87902 , n32968 );
and ( n87903 , n87902 , n33309 );
xor ( n87904 , n33229 , n53900 );
and ( n87905 , n87904 , n32968 );
or ( n87906 , n87903 , n87905 );
and ( n87907 , n87906 , n33370 );
and ( n87908 , n32992 , n35056 );
and ( n87909 , n33229 , n49794 );
or ( n87910 , C0 , n87900 , n87901 , n87907 , n87908 , n87909 );
buf ( n87911 , n87910 );
buf ( n87912 , n87911 );
buf ( n87913 , n31655 );
buf ( n87914 , n30987 );
buf ( n87915 , n31655 );
and ( n87916 , n46021 , n32500 );
not ( n87917 , n35211 );
and ( n87918 , n87917 , n37539 );
buf ( n87919 , n87918 );
and ( n87920 , n87919 , n32421 );
not ( n87921 , n35245 );
and ( n87922 , n87921 , n37539 );
buf ( n87923 , n87922 );
and ( n87924 , n87923 , n32419 );
not ( n87925 , n35278 );
and ( n87926 , n87925 , n37539 );
not ( n87927 , n35295 );
and ( n87928 , n87927 , n49569 );
xor ( n87929 , n37539 , n49546 );
and ( n87930 , n87929 , n35295 );
or ( n87931 , n87928 , n87930 );
and ( n87932 , n87931 , n35278 );
or ( n87933 , n87926 , n87932 );
and ( n87934 , n87933 , n32417 );
not ( n87935 , n35331 );
and ( n87936 , n87935 , n37539 );
not ( n87937 , n35294 );
not ( n87938 , n45995 );
and ( n87939 , n87938 , n49569 );
xor ( n87940 , n49570 , n49632 );
and ( n87941 , n87940 , n45995 );
or ( n87942 , n87939 , n87941 );
and ( n87943 , n87937 , n87942 );
and ( n87944 , n87929 , n35294 );
or ( n87945 , n87943 , n87944 );
and ( n87946 , n87945 , n35331 );
or ( n87947 , n87936 , n87946 );
and ( n87948 , n87947 , n32415 );
and ( n87949 , n37539 , n35354 );
or ( n87950 , n87920 , n87924 , n87934 , n87948 , n87949 );
and ( n87951 , n87950 , n32456 );
not ( n87952 , n32475 );
not ( n87953 , n46060 );
and ( n87954 , n87953 , n49660 );
xor ( n87955 , n49661 , n49726 );
and ( n87956 , n87955 , n46060 );
or ( n87957 , n87954 , n87956 );
and ( n87958 , n87952 , n87957 );
and ( n87959 , n37539 , n32475 );
or ( n87960 , n87958 , n87959 );
and ( n87961 , n87960 , n32486 );
and ( n87962 , n37539 , n35367 );
or ( n87963 , C0 , n87916 , n87951 , n87961 , C0 , n87962 );
buf ( n87964 , n87963 );
buf ( n87965 , n87964 );
and ( n87966 , n33230 , n32528 );
not ( n87967 , n32598 );
and ( n87968 , n87967 , n32993 );
buf ( n87969 , n87968 );
and ( n87970 , n87969 , n32890 );
not ( n87971 , n32919 );
and ( n87972 , n87971 , n32993 );
buf ( n87973 , n87972 );
and ( n87974 , n87973 , n32924 );
not ( n87975 , n32953 );
and ( n87976 , n87975 , n32993 );
not ( n87977 , n32971 );
and ( n87978 , n87977 , n33111 );
xor ( n87979 , n32993 , n33012 );
and ( n87980 , n87979 , n32971 );
or ( n87981 , n87978 , n87980 );
and ( n87982 , n87981 , n32953 );
or ( n87983 , n87976 , n87982 );
and ( n87984 , n87983 , n33038 );
not ( n87985 , n33067 );
and ( n87986 , n87985 , n32993 );
not ( n87987 , n32970 );
not ( n87988 , n33071 );
and ( n87989 , n87988 , n33111 );
xor ( n87990 , n33112 , n33144 );
and ( n87991 , n87990 , n33071 );
or ( n87992 , n87989 , n87991 );
and ( n87993 , n87987 , n87992 );
and ( n87994 , n87979 , n32970 );
or ( n87995 , n87993 , n87994 );
and ( n87996 , n87995 , n33067 );
or ( n87997 , n87986 , n87996 );
and ( n87998 , n87997 , n33172 );
and ( n87999 , n32993 , n33204 );
or ( n88000 , n87970 , n87974 , n87984 , n87998 , n87999 );
and ( n88001 , n88000 , n33208 );
not ( n88002 , n32968 );
not ( n88003 , n33270 );
and ( n88004 , n88003 , n33311 );
xor ( n88005 , n33312 , n33344 );
and ( n88006 , n88005 , n33270 );
or ( n88007 , n88004 , n88006 );
and ( n88008 , n88002 , n88007 );
and ( n88009 , n32993 , n32968 );
or ( n88010 , n88008 , n88009 );
and ( n88011 , n88010 , n33370 );
buf ( n88012 , n35056 );
and ( n88013 , n32993 , n33382 );
or ( n88014 , C0 , n87966 , n88001 , n88011 , n88012 , n88013 );
buf ( n88015 , n88014 );
buf ( n88016 , n88015 );
buf ( n88017 , n30987 );
buf ( n88018 , n31655 );
buf ( n88019 , n30987 );
buf ( n88020 , n31655 );
not ( n88021 , n31728 );
and ( n88022 , n88021 , n46020 );
and ( n88023 , n80363 , n31728 );
or ( n88024 , n88022 , n88023 );
and ( n88025 , n88024 , n32253 );
not ( n88026 , n32283 );
and ( n88027 , n88026 , n46020 );
and ( n88028 , n80374 , n32283 );
or ( n88029 , n88027 , n88028 );
and ( n88030 , n88029 , n32398 );
and ( n88031 , n46020 , n32436 );
or ( n88032 , n88025 , n88030 , n88031 );
and ( n88033 , n88032 , n32456 );
and ( n88034 , n49658 , n32473 );
not ( n88035 , n32475 );
and ( n88036 , n88035 , n49658 );
xor ( n88037 , n46020 , n50479 );
and ( n88038 , n88037 , n32475 );
or ( n88039 , n88036 , n88038 );
and ( n88040 , n88039 , n32486 );
and ( n88041 , n37537 , n32489 );
and ( n88042 , n46020 , n32501 );
or ( n88043 , C0 , n88033 , n88034 , n88040 , n88041 , n88042 );
buf ( n88044 , n88043 );
buf ( n88045 , n88044 );
buf ( n88046 , n30987 );
not ( n88047 , n35542 );
and ( n88048 , n88047 , n41858 );
and ( n88049 , n69550 , n35542 );
or ( n88050 , n88048 , n88049 );
buf ( n88051 , n88050 );
buf ( n88052 , n88051 );
not ( n88053 , n34150 );
and ( n88054 , n88053 , n32775 );
not ( n88055 , n56836 );
and ( n88056 , n88055 , n32775 );
and ( n88057 , n32789 , n56836 );
or ( n88058 , n88056 , n88057 );
and ( n88059 , n88058 , n34150 );
or ( n88060 , n88054 , n88059 );
and ( n88061 , n88060 , n33381 );
not ( n88062 , n56844 );
not ( n88063 , n56836 );
and ( n88064 , n88063 , n32775 );
and ( n88065 , n34301 , n56836 );
or ( n88066 , n88064 , n88065 );
and ( n88067 , n88062 , n88066 );
and ( n88068 , n34301 , n56844 );
or ( n88069 , n88067 , n88068 );
and ( n88070 , n88069 , n33375 );
not ( n88071 , n32968 );
not ( n88072 , n56844 );
not ( n88073 , n56836 );
and ( n88074 , n88073 , n32775 );
and ( n88075 , n34301 , n56836 );
or ( n88076 , n88074 , n88075 );
and ( n88077 , n88072 , n88076 );
and ( n88078 , n34301 , n56844 );
or ( n88079 , n88077 , n88078 );
and ( n88080 , n88071 , n88079 );
not ( n88081 , n56864 );
not ( n88082 , n56866 );
and ( n88083 , n88082 , n88079 );
and ( n88084 , n34761 , n56866 );
or ( n88085 , n88083 , n88084 );
and ( n88086 , n88081 , n88085 );
and ( n88087 , n35050 , n56864 );
or ( n88088 , n88086 , n88087 );
and ( n88089 , n88088 , n32968 );
or ( n88090 , n88080 , n88089 );
and ( n88091 , n88090 , n33370 );
and ( n88092 , n32775 , n35062 );
or ( n88093 , C0 , n88061 , n88070 , n88091 , n88092 );
buf ( n88094 , n88093 );
buf ( n88095 , n88094 );
buf ( n88096 , n30987 );
buf ( n88097 , n31655 );
buf ( n88098 , n31655 );
buf ( n88099 , n31655 );
xor ( n88100 , n33091 , n58388 );
and ( n88101 , n88100 , n33201 );
not ( n88102 , n41576 );
and ( n88103 , n88102 , n33091 );
and ( n88104 , n55247 , n41576 );
or ( n88105 , n88103 , n88104 );
and ( n88106 , n88105 , n33189 );
and ( n88107 , n33091 , n41592 );
or ( n88108 , n88101 , n88106 , n88107 );
and ( n88109 , n88108 , n33208 );
and ( n88110 , n33091 , n39805 );
or ( n88111 , C0 , n88109 , n88110 );
buf ( n88112 , n88111 );
buf ( n88113 , n88112 );
buf ( n88114 , n30987 );
buf ( n88115 , n30987 );
buf ( n88116 , n31655 );
not ( n88117 , n50828 );
not ( n88118 , n50834 );
and ( n88119 , n88118 , n40646 );
and ( n88120 , n54960 , n50834 );
or ( n88121 , n88119 , n88120 );
and ( n88122 , n88117 , n88121 );
and ( n88123 , n82380 , n50828 );
or ( n88124 , n88122 , n88123 );
buf ( n88125 , n88124 );
buf ( n88126 , n88125 );
buf ( n88127 , n31655 );
buf ( n88128 , n30987 );
xor ( n88129 , n33131 , n33133 );
and ( n88130 , n88129 , n33201 );
not ( n88131 , n41576 );
and ( n88132 , n88131 , n33131 );
buf ( n88133 , n32687 );
and ( n88134 , n88133 , n41576 );
or ( n88135 , n88132 , n88134 );
and ( n88136 , n88135 , n33189 );
and ( n88137 , n33131 , n41592 );
or ( n88138 , n88130 , n88136 , n88137 );
and ( n88139 , n88138 , n33208 );
and ( n88140 , n33131 , n39805 );
or ( n88141 , C0 , n88139 , n88140 );
buf ( n88142 , n88141 );
buf ( n88143 , n88142 );
buf ( n88144 , n30987 );
buf ( n88145 , n31655 );
not ( n88146 , n41532 );
and ( n88147 , n88146 , n34247 );
and ( n88148 , n56336 , n41532 );
or ( n88149 , n88147 , n88148 );
buf ( n88150 , n88149 );
buf ( n88151 , n88150 );
and ( n88152 , n57514 , n48455 );
not ( n88153 , n48457 );
and ( n88154 , n88153 , n52400 );
and ( n88155 , n57514 , n48457 );
or ( n88156 , n88154 , n88155 );
and ( n88157 , n88156 , n31373 );
not ( n88158 , n44807 );
and ( n88159 , n88158 , n52400 );
and ( n88160 , n57514 , n44807 );
or ( n88161 , n88159 , n88160 );
and ( n88162 , n88161 , n31408 );
not ( n88163 , n48468 );
and ( n88164 , n88163 , n52400 );
and ( n88165 , n57514 , n48468 );
or ( n88166 , n88164 , n88165 );
and ( n88167 , n88166 , n31468 );
not ( n88168 , n44817 );
and ( n88169 , n88168 , n52400 );
and ( n88170 , n57514 , n44817 );
or ( n88171 , n88169 , n88170 );
and ( n88172 , n88171 , n31521 );
not ( n88173 , n39979 );
and ( n88174 , n88173 , n52400 );
and ( n88175 , n57502 , n39979 );
or ( n88176 , n88174 , n88175 );
and ( n88177 , n88176 , n31538 );
not ( n88178 , n45059 );
and ( n88179 , n88178 , n52400 );
and ( n88180 , n57502 , n45059 );
or ( n88181 , n88179 , n88180 );
and ( n88182 , n88181 , n31536 );
not ( n88183 , n33419 );
and ( n88184 , n88183 , n52400 );
and ( n88185 , n75231 , n33419 );
or ( n88186 , n88184 , n88185 );
and ( n88187 , n88186 , n31529 );
not ( n88188 , n33734 );
and ( n88189 , n88188 , n52400 );
and ( n88190 , n75242 , n33734 );
or ( n88191 , n88189 , n88190 );
and ( n88192 , n88191 , n31527 );
and ( n88193 , n57525 , n48513 );
or ( n88194 , n88152 , n88157 , n88162 , n88167 , n88172 , n88177 , n88182 , n88187 , n88192 , n88193 );
and ( n88195 , n88194 , n31557 );
and ( n88196 , n35389 , n33973 );
and ( n88197 , n52400 , n48524 );
or ( n88198 , C0 , n88195 , n88196 , n88197 );
buf ( n88199 , n88198 );
buf ( n88200 , n88199 );
buf ( n88201 , n31655 );
buf ( n88202 , n30987 );
not ( n88203 , n38443 );
and ( n88204 , n88203 , n38269 );
xor ( n88205 , n53466 , n53503 );
and ( n88206 , n88205 , n38443 );
or ( n88207 , n88204 , n88206 );
and ( n88208 , n88207 , n38450 );
not ( n88209 , n39339 );
and ( n88210 , n88209 , n39169 );
xor ( n88211 , n53522 , n53559 );
and ( n88212 , n88211 , n39339 );
or ( n88213 , n88210 , n88212 );
and ( n88214 , n88213 , n39346 );
and ( n88215 , n40218 , n39359 );
or ( n88216 , n88208 , n88214 , n88215 );
buf ( n88217 , n88216 );
buf ( n88218 , n88217 );
buf ( n88219 , n30987 );
not ( n88220 , n34150 );
and ( n88221 , n88220 , n32795 );
not ( n88222 , n60126 );
and ( n88223 , n88222 , n32795 );
and ( n88224 , n32823 , n60126 );
or ( n88225 , n88223 , n88224 );
and ( n88226 , n88225 , n34150 );
or ( n88227 , n88221 , n88226 );
and ( n88228 , n88227 , n33381 );
not ( n88229 , n60134 );
not ( n88230 , n60126 );
and ( n88231 , n88230 , n32795 );
and ( n88232 , n41464 , n60126 );
or ( n88233 , n88231 , n88232 );
and ( n88234 , n88229 , n88233 );
and ( n88235 , n41464 , n60134 );
or ( n88236 , n88234 , n88235 );
and ( n88237 , n88236 , n33375 );
not ( n88238 , n32968 );
not ( n88239 , n60134 );
not ( n88240 , n60126 );
and ( n88241 , n88240 , n32795 );
and ( n88242 , n41464 , n60126 );
or ( n88243 , n88241 , n88242 );
and ( n88244 , n88239 , n88243 );
and ( n88245 , n41464 , n60134 );
or ( n88246 , n88244 , n88245 );
and ( n88247 , n88238 , n88246 );
not ( n88248 , n60154 );
not ( n88249 , n60156 );
and ( n88250 , n88249 , n88246 );
and ( n88251 , n41490 , n60156 );
or ( n88252 , n88250 , n88251 );
and ( n88253 , n88248 , n88252 );
and ( n88254 , n41500 , n60154 );
or ( n88255 , n88253 , n88254 );
and ( n88256 , n88255 , n32968 );
or ( n88257 , n88247 , n88256 );
and ( n88258 , n88257 , n33370 );
and ( n88259 , n32795 , n35062 );
or ( n88260 , C0 , n88228 , n88237 , n88258 , n88259 );
buf ( n88261 , n88260 );
buf ( n88262 , n88261 );
buf ( n88263 , n30987 );
buf ( n88264 , n31655 );
buf ( n88265 , n31655 );
buf ( n88266 , n40205 );
not ( n88267 , n46356 );
and ( n88268 , n88267 , n31298 );
not ( n88269 , n49427 );
and ( n88270 , n88269 , n31298 );
and ( n88271 , n31306 , n49427 );
or ( n88272 , n88270 , n88271 );
and ( n88273 , n88272 , n46356 );
or ( n88274 , n88268 , n88273 );
and ( n88275 , n88274 , n31649 );
not ( n88276 , n49435 );
not ( n88277 , n49427 );
and ( n88278 , n88277 , n31298 );
and ( n88279 , n58061 , n49427 );
or ( n88280 , n88278 , n88279 );
and ( n88281 , n88276 , n88280 );
and ( n88282 , n58061 , n49435 );
or ( n88283 , n88281 , n88282 );
and ( n88284 , n88283 , n31643 );
not ( n88285 , n31452 );
not ( n88286 , n49435 );
not ( n88287 , n49427 );
and ( n88288 , n88287 , n31298 );
and ( n88289 , n58061 , n49427 );
or ( n88290 , n88288 , n88289 );
and ( n88291 , n88286 , n88290 );
and ( n88292 , n58061 , n49435 );
or ( n88293 , n88291 , n88292 );
and ( n88294 , n88285 , n88293 );
not ( n88295 , n49460 );
not ( n88296 , n49462 );
and ( n88297 , n88296 , n88293 );
and ( n88298 , n58085 , n49462 );
or ( n88299 , n88297 , n88298 );
and ( n88300 , n88295 , n88299 );
and ( n88301 , n58093 , n49460 );
or ( n88302 , n88300 , n88301 );
and ( n88303 , n88302 , n31452 );
or ( n88304 , n88294 , n88303 );
and ( n88305 , n88304 , n31638 );
and ( n88306 , n31298 , n47277 );
or ( n88307 , C0 , n88275 , n88284 , n88305 , n88306 );
buf ( n88308 , n88307 );
buf ( n88309 , n88308 );
buf ( n88310 , n31655 );
buf ( n88311 , n30987 );
xor ( n88312 , n47290 , n47292 );
and ( n88313 , n88312 , n32433 );
not ( n88314 , n47331 );
and ( n88315 , n88314 , n47290 );
buf ( n88316 , n31961 );
and ( n88317 , n88316 , n47331 );
or ( n88318 , n88315 , n88317 );
and ( n88319 , n88318 , n32413 );
and ( n88320 , n47290 , n47402 );
or ( n88321 , n88313 , n88319 , n88320 );
and ( n88322 , n88321 , n32456 );
and ( n88323 , n47290 , n47409 );
or ( n88324 , C0 , n88322 , n88323 );
buf ( n88325 , n88324 );
buf ( n88326 , n88325 );
buf ( n88327 , n31655 );
not ( n88328 , n32953 );
and ( n88329 , n88328 , n74642 );
and ( n88330 , n74650 , n32953 );
or ( n88331 , n88329 , n88330 );
and ( n88332 , n88331 , n33038 );
not ( n88333 , n39586 );
and ( n88334 , n88333 , n74642 );
and ( n88335 , n81517 , n39586 );
or ( n88336 , n88334 , n88335 );
and ( n88337 , n88336 , n33172 );
and ( n88338 , n74642 , n39795 );
or ( n88339 , n88332 , n88337 , n88338 );
and ( n88340 , n88339 , n33208 );
and ( n88341 , n74642 , n39805 );
or ( n88342 , C0 , n88340 , n88341 );
buf ( n88343 , n88342 );
buf ( n88344 , n88343 );
buf ( n88345 , n31655 );
buf ( n88346 , n30987 );
buf ( n88347 , n30987 );
buf ( n88348 , n31655 );
and ( n88349 , n33224 , n32528 );
not ( n88350 , n32598 );
and ( n88351 , n88350 , n32987 );
buf ( n88352 , n88351 );
and ( n88353 , n88352 , n32890 );
not ( n88354 , n32919 );
and ( n88355 , n88354 , n32987 );
buf ( n88356 , n88355 );
and ( n88357 , n88356 , n32924 );
not ( n88358 , n32953 );
and ( n88359 , n88358 , n32987 );
not ( n88360 , n32971 );
and ( n88361 , n88360 , n33099 );
xor ( n88362 , n32987 , n33018 );
and ( n88363 , n88362 , n32971 );
or ( n88364 , n88361 , n88363 );
and ( n88365 , n88364 , n32953 );
or ( n88366 , n88359 , n88365 );
and ( n88367 , n88366 , n33038 );
not ( n88368 , n33067 );
and ( n88369 , n88368 , n32987 );
not ( n88370 , n32970 );
not ( n88371 , n33071 );
and ( n88372 , n88371 , n33099 );
xor ( n88373 , n33100 , n33150 );
and ( n88374 , n88373 , n33071 );
or ( n88375 , n88372 , n88374 );
and ( n88376 , n88370 , n88375 );
and ( n88377 , n88362 , n32970 );
or ( n88378 , n88376 , n88377 );
and ( n88379 , n88378 , n33067 );
or ( n88380 , n88369 , n88379 );
and ( n88381 , n88380 , n33172 );
and ( n88382 , n32987 , n33204 );
or ( n88383 , n88353 , n88357 , n88367 , n88381 , n88382 );
and ( n88384 , n88383 , n33208 );
not ( n88385 , n32968 );
not ( n88386 , n33270 );
and ( n88387 , n88386 , n33299 );
xor ( n88388 , n33300 , n33350 );
and ( n88389 , n88388 , n33270 );
or ( n88390 , n88387 , n88389 );
and ( n88391 , n88385 , n88390 );
and ( n88392 , n32987 , n32968 );
or ( n88393 , n88391 , n88392 );
and ( n88394 , n88393 , n33370 );
buf ( n88395 , n35056 );
and ( n88396 , n32987 , n33382 );
or ( n88397 , C0 , n88349 , n88384 , n88394 , n88395 , n88396 );
buf ( n88398 , n88397 );
buf ( n88399 , n88398 );
buf ( n88400 , n30987 );
buf ( n88401 , n31655 );
buf ( n88402 , n30987 );
buf ( n88403 , n31655 );
not ( n88404 , n31728 );
and ( n88405 , n88404 , n46026 );
and ( n88406 , n84368 , n31728 );
or ( n88407 , n88405 , n88406 );
and ( n88408 , n88407 , n32253 );
not ( n88409 , n32283 );
and ( n88410 , n88409 , n46026 );
and ( n88411 , n84379 , n32283 );
or ( n88412 , n88410 , n88411 );
and ( n88413 , n88412 , n32398 );
and ( n88414 , n46026 , n32436 );
or ( n88415 , n88408 , n88413 , n88414 );
and ( n88416 , n88415 , n32456 );
and ( n88417 , n49669 , n32473 );
not ( n88418 , n32475 );
and ( n88419 , n88418 , n49669 );
xor ( n88420 , n46026 , n47760 );
and ( n88421 , n88420 , n32475 );
or ( n88422 , n88419 , n88421 );
and ( n88423 , n88422 , n32486 );
and ( n88424 , n37549 , n32489 );
and ( n88425 , n46026 , n32501 );
or ( n88426 , C0 , n88416 , n88417 , n88423 , n88424 , n88425 );
buf ( n88427 , n88426 );
buf ( n88428 , n88427 );
buf ( n88429 , n31655 );
buf ( n88430 , n30987 );
and ( n88431 , n72102 , n33377 );
not ( n88432 , n48545 );
buf ( n88433 , RI15b473a0_295);
and ( n88434 , n88432 , n88433 );
and ( n88435 , n72108 , n48545 );
or ( n88436 , n88434 , n88435 );
and ( n88437 , n88436 , n32890 );
not ( n88438 , n48557 );
and ( n88439 , n88438 , n88433 );
and ( n88440 , n72108 , n48557 );
or ( n88441 , n88439 , n88440 );
and ( n88442 , n88441 , n33038 );
and ( n88443 , n88433 , n48571 );
or ( n88444 , n88437 , n88442 , n88443 );
and ( n88445 , n88444 , n33208 );
and ( n88446 , n88433 , n48577 );
or ( n88447 , C0 , n88431 , n88445 , n88446 );
buf ( n88448 , n88447 );
buf ( n88449 , n88448 );
buf ( n88450 , n30987 );
buf ( n88451 , n31655 );
buf ( n88452 , n30987 );
buf ( n88453 , RI15b47760_303);
buf ( n88454 , n88453 );
buf ( n88455 , n31655 );
not ( n88456 , n48765 );
and ( n88457 , n88456 , n33226 );
and ( n88458 , n85876 , n48765 );
or ( n88459 , n88457 , n88458 );
and ( n88460 , n88459 , n33180 );
not ( n88461 , n49054 );
and ( n88462 , n88461 , n33226 );
and ( n88463 , n85887 , n49054 );
or ( n88464 , n88462 , n88463 );
and ( n88465 , n88464 , n33178 );
and ( n88466 , n33226 , n49774 );
or ( n88467 , n88460 , n88465 , n88466 );
and ( n88468 , n88467 , n33208 );
and ( n88469 , n33303 , n33375 );
not ( n88470 , n32968 );
and ( n88471 , n88470 , n33303 );
xor ( n88472 , n33226 , n53903 );
and ( n88473 , n88472 , n32968 );
or ( n88474 , n88471 , n88473 );
and ( n88475 , n88474 , n33370 );
and ( n88476 , n32989 , n35056 );
and ( n88477 , n33226 , n49794 );
or ( n88478 , C0 , n88468 , n88469 , n88475 , n88476 , n88477 );
buf ( n88479 , n88478 );
buf ( n88480 , n88479 );
buf ( n88481 , n30987 );
buf ( n88482 , n31655 );
and ( n88483 , n46024 , n32500 );
not ( n88484 , n35211 );
and ( n88485 , n88484 , n37545 );
buf ( n88486 , n88485 );
and ( n88487 , n88486 , n32421 );
not ( n88488 , n35245 );
and ( n88489 , n88488 , n37545 );
buf ( n88490 , n88489 );
and ( n88491 , n88490 , n32419 );
not ( n88492 , n35278 );
and ( n88493 , n88492 , n37545 );
not ( n88494 , n35295 );
and ( n88495 , n88494 , n49575 );
xor ( n88496 , n37545 , n49543 );
and ( n88497 , n88496 , n35295 );
or ( n88498 , n88495 , n88497 );
and ( n88499 , n88498 , n35278 );
or ( n88500 , n88493 , n88499 );
and ( n88501 , n88500 , n32417 );
not ( n88502 , n35331 );
and ( n88503 , n88502 , n37545 );
not ( n88504 , n35294 );
not ( n88505 , n45995 );
and ( n88506 , n88505 , n49575 );
xor ( n88507 , n49576 , n49629 );
and ( n88508 , n88507 , n45995 );
or ( n88509 , n88506 , n88508 );
and ( n88510 , n88504 , n88509 );
and ( n88511 , n88496 , n35294 );
or ( n88512 , n88510 , n88511 );
and ( n88513 , n88512 , n35331 );
or ( n88514 , n88503 , n88513 );
and ( n88515 , n88514 , n32415 );
and ( n88516 , n37545 , n35354 );
or ( n88517 , n88487 , n88491 , n88501 , n88515 , n88516 );
and ( n88518 , n88517 , n32456 );
not ( n88519 , n32475 );
not ( n88520 , n46060 );
and ( n88521 , n88520 , n49665 );
xor ( n88522 , n49666 , n49723 );
and ( n88523 , n88522 , n46060 );
or ( n88524 , n88521 , n88523 );
and ( n88525 , n88519 , n88524 );
and ( n88526 , n37545 , n32475 );
or ( n88527 , n88525 , n88526 );
and ( n88528 , n88527 , n32486 );
and ( n88529 , n37545 , n35367 );
or ( n88530 , C0 , n88483 , n88518 , n88528 , C0 , n88529 );
buf ( n88531 , n88530 );
buf ( n88532 , n88531 );
buf ( n88533 , n31655 );
and ( n88534 , n51843 , n31645 );
not ( n88535 , n45274 );
and ( n88536 , n88535 , n59536 );
and ( n88537 , n56970 , n45274 );
or ( n88538 , n88536 , n88537 );
and ( n88539 , n88538 , n31373 );
not ( n88540 , n45280 );
and ( n88541 , n88540 , n59536 );
and ( n88542 , n56970 , n45280 );
or ( n88543 , n88541 , n88542 );
and ( n88544 , n88543 , n31468 );
and ( n88545 , n59536 , n45802 );
or ( n88546 , n88539 , n88544 , n88545 );
and ( n88547 , n88546 , n31557 );
and ( n88548 , n59536 , n45808 );
or ( n88549 , C0 , n88534 , n88547 , n88548 );
buf ( n88550 , n88549 );
buf ( n88551 , n88550 );
not ( n88552 , n40163 );
and ( n88553 , n88552 , n31900 );
not ( n88554 , n56287 );
and ( n88555 , n88554 , n31900 );
and ( n88556 , n32200 , n56287 );
or ( n88557 , n88555 , n88556 );
and ( n88558 , n88557 , n40163 );
or ( n88559 , n88553 , n88558 );
and ( n88560 , n88559 , n32498 );
not ( n88561 , n56295 );
not ( n88562 , n56287 );
and ( n88563 , n88562 , n31900 );
and ( n88564 , n53243 , n56287 );
or ( n88565 , n88563 , n88564 );
and ( n88566 , n88561 , n88565 );
and ( n88567 , n53243 , n56295 );
or ( n88568 , n88566 , n88567 );
and ( n88569 , n88568 , n32473 );
not ( n88570 , n32475 );
not ( n88571 , n56295 );
not ( n88572 , n56287 );
and ( n88573 , n88572 , n31900 );
and ( n88574 , n53243 , n56287 );
or ( n88575 , n88573 , n88574 );
and ( n88576 , n88571 , n88575 );
and ( n88577 , n53243 , n56295 );
or ( n88578 , n88576 , n88577 );
and ( n88579 , n88570 , n88578 );
not ( n88580 , n56315 );
not ( n88581 , n56317 );
and ( n88582 , n88581 , n88578 );
and ( n88583 , n53269 , n56317 );
or ( n88584 , n88582 , n88583 );
and ( n88585 , n88580 , n88584 );
and ( n88586 , n53277 , n56315 );
or ( n88587 , n88585 , n88586 );
and ( n88588 , n88587 , n32475 );
or ( n88589 , n88579 , n88588 );
and ( n88590 , n88589 , n32486 );
and ( n88591 , n31900 , n41278 );
or ( n88592 , C0 , n88560 , n88569 , n88590 , n88591 );
buf ( n88593 , n88592 );
buf ( n88594 , n88593 );
buf ( n88595 , n30987 );
buf ( n88596 , n40225 );
not ( n88597 , n46356 );
and ( n88598 , n88597 , n31195 );
not ( n88599 , n56904 );
and ( n88600 , n88599 , n31195 );
and ( n88601 , n31205 , n56904 );
or ( n88602 , n88600 , n88601 );
and ( n88603 , n88602 , n46356 );
or ( n88604 , n88598 , n88603 );
and ( n88605 , n88604 , n31649 );
not ( n88606 , n56912 );
not ( n88607 , n56904 );
and ( n88608 , n88607 , n31195 );
and ( n88609 , n50125 , n56904 );
or ( n88610 , n88608 , n88609 );
and ( n88611 , n88606 , n88610 );
and ( n88612 , n50125 , n56912 );
or ( n88613 , n88611 , n88612 );
and ( n88614 , n88613 , n31643 );
not ( n88615 , n31452 );
not ( n88616 , n56912 );
not ( n88617 , n56904 );
and ( n88618 , n88617 , n31195 );
and ( n88619 , n50125 , n56904 );
or ( n88620 , n88618 , n88619 );
and ( n88621 , n88616 , n88620 );
and ( n88622 , n50125 , n56912 );
or ( n88623 , n88621 , n88622 );
and ( n88624 , n88615 , n88623 );
not ( n88625 , n56937 );
not ( n88626 , n56939 );
and ( n88627 , n88626 , n88623 );
and ( n88628 , n50151 , n56939 );
or ( n88629 , n88627 , n88628 );
and ( n88630 , n88625 , n88629 );
and ( n88631 , n50159 , n56937 );
or ( n88632 , n88630 , n88631 );
and ( n88633 , n88632 , n31452 );
or ( n88634 , n88624 , n88633 );
and ( n88635 , n88634 , n31638 );
and ( n88636 , n31195 , n47277 );
or ( n88637 , C0 , n88605 , n88614 , n88635 , n88636 );
buf ( n88638 , n88637 );
buf ( n88639 , n88638 );
buf ( n88640 , n31655 );
buf ( n88641 , n30987 );
and ( n88642 , n50949 , n83089 );
xor ( n88643 , n50947 , n88642 );
and ( n88644 , n88643 , n32431 );
not ( n88645 , n50002 );
and ( n88646 , n88645 , n50947 );
and ( n88647 , n40557 , n50002 );
or ( n88648 , n88646 , n88647 );
and ( n88649 , n88648 , n32419 );
not ( n88650 , n50008 );
and ( n88651 , n88650 , n50947 );
and ( n88652 , n71274 , n50008 );
or ( n88653 , n88651 , n88652 );
and ( n88654 , n88653 , n32415 );
not ( n88655 , n50067 );
and ( n88656 , n88655 , n50947 );
and ( n88657 , n31750 , n60350 );
and ( n88658 , n31778 , n60352 );
and ( n88659 , n31781 , n60354 );
and ( n88660 , n31784 , n60356 );
and ( n88661 , n31787 , n60358 );
and ( n88662 , n31790 , n60360 );
and ( n88663 , n31793 , n60362 );
and ( n88664 , n31796 , n60364 );
and ( n88665 , n31799 , n60366 );
and ( n88666 , n31802 , n60368 );
and ( n88667 , n31805 , n60370 );
and ( n88668 , n31808 , n60372 );
and ( n88669 , n31811 , n60374 );
and ( n88670 , n31814 , n60376 );
and ( n88671 , n31817 , n60378 );
and ( n88672 , n31820 , n60380 );
or ( n88673 , n88657 , n88658 , n88659 , n88660 , n88661 , n88662 , n88663 , n88664 , n88665 , n88666 , n88667 , n88668 , n88669 , n88670 , n88671 , n88672 );
and ( n88674 , n60382 , n83104 );
xor ( n88675 , n88673 , n88674 );
and ( n88676 , n88675 , n50067 );
or ( n88677 , n88656 , n88676 );
and ( n88678 , n88677 , n32411 );
and ( n88679 , n50947 , n50098 );
or ( n88680 , n88644 , n88649 , n88654 , n88678 , n88679 );
and ( n88681 , n88680 , n32456 );
and ( n88682 , n50947 , n47409 );
or ( n88683 , C0 , n88681 , n88682 );
buf ( n88684 , n88683 );
buf ( n88685 , n88684 );
buf ( n88686 , n31655 );
buf ( n88687 , n31655 );
not ( n88688 , n46356 );
and ( n88689 , n88688 , n31348 );
not ( n88690 , n78324 );
and ( n88691 , n88690 , n31348 );
and ( n88692 , n31372 , n78324 );
or ( n88693 , n88691 , n88692 );
and ( n88694 , n88693 , n46356 );
or ( n88695 , n88689 , n88694 );
and ( n88696 , n88695 , n31649 );
not ( n88697 , n78332 );
not ( n88698 , n78324 );
and ( n88699 , n88698 , n31348 );
and ( n88700 , n47849 , n78324 );
or ( n88701 , n88699 , n88700 );
and ( n88702 , n88697 , n88701 );
and ( n88703 , n47849 , n78332 );
or ( n88704 , n88702 , n88703 );
and ( n88705 , n88704 , n31643 );
not ( n88706 , n31452 );
not ( n88707 , n78332 );
not ( n88708 , n78324 );
and ( n88709 , n88708 , n31348 );
and ( n88710 , n47849 , n78324 );
or ( n88711 , n88709 , n88710 );
and ( n88712 , n88707 , n88711 );
and ( n88713 , n47849 , n78332 );
or ( n88714 , n88712 , n88713 );
and ( n88715 , n88706 , n88714 );
not ( n88716 , n78352 );
not ( n88717 , n78354 );
and ( n88718 , n88717 , n88714 );
and ( n88719 , n47877 , n78354 );
or ( n88720 , n88718 , n88719 );
and ( n88721 , n88716 , n88720 );
and ( n88722 , n47887 , n78352 );
or ( n88723 , n88721 , n88722 );
and ( n88724 , n88723 , n31452 );
or ( n88725 , n88715 , n88724 );
and ( n88726 , n88725 , n31638 );
and ( n88727 , n31348 , n47277 );
or ( n88728 , C0 , n88696 , n88705 , n88726 , n88727 );
buf ( n88729 , n88728 );
buf ( n88730 , n88729 );
buf ( n88731 , n30987 );
buf ( n88732 , RI15b5f748_1122);
and ( n88733 , n88732 , n32494 );
not ( n88734 , n46083 );
buf ( n88735 , RI15b5fec8_1138);
and ( n88736 , n88734 , n88735 );
not ( n88737 , n46290 );
and ( n88738 , n88737 , n46286 );
xor ( n88739 , n85033 , n85034 );
and ( n88740 , n88739 , n46290 );
or ( n88741 , n88738 , n88740 );
and ( n88742 , n88741 , n46083 );
or ( n88743 , n88736 , n88742 );
and ( n88744 , n88743 , n32421 );
not ( n88745 , n46326 );
and ( n88746 , n88745 , n88735 );
and ( n88747 , n88741 , n46326 );
or ( n88748 , n88746 , n88747 );
and ( n88749 , n88748 , n32417 );
and ( n88750 , n88735 , n46340 );
or ( n88751 , n88744 , n88749 , n88750 );
and ( n88752 , n88751 , n32456 );
and ( n88753 , n88735 , n46349 );
or ( n88754 , C0 , n88733 , n88752 , n88753 );
buf ( n88755 , n88754 );
buf ( n88756 , n88755 );
buf ( n88757 , n31655 );
buf ( n88758 , n31655 );
buf ( n88759 , n30987 );
and ( n88760 , n72876 , n33377 );
not ( n88761 , n48545 );
and ( n88762 , n88761 , n47517 );
buf ( n88763 , n88762 );
and ( n88764 , n88763 , n32890 );
not ( n88765 , n48557 );
and ( n88766 , n88765 , n47517 );
and ( n88767 , n72882 , n48557 );
or ( n88768 , n88766 , n88767 );
and ( n88769 , n88768 , n33038 );
and ( n88770 , n47517 , n48571 );
or ( n88771 , n88764 , n88769 , n88770 );
and ( n88772 , n88771 , n33208 );
and ( n88773 , n47517 , n48577 );
or ( n88774 , C0 , n88760 , n88772 , n88773 );
buf ( n88775 , n88774 );
buf ( n88776 , n88775 );
buf ( n88777 , n30987 );
buf ( n88778 , n31655 );
not ( n88779 , n46356 );
and ( n88780 , n88779 , n31244 );
not ( n88781 , n55473 );
and ( n88782 , n88781 , n31244 );
and ( n88783 , n31272 , n55473 );
or ( n88784 , n88782 , n88783 );
and ( n88785 , n88784 , n46356 );
or ( n88786 , n88780 , n88785 );
and ( n88787 , n88786 , n31649 );
not ( n88788 , n55481 );
not ( n88789 , n55473 );
and ( n88790 , n88789 , n31244 );
and ( n88791 , n49443 , n55473 );
or ( n88792 , n88790 , n88791 );
and ( n88793 , n88788 , n88792 );
and ( n88794 , n49443 , n55481 );
or ( n88795 , n88793 , n88794 );
and ( n88796 , n88795 , n31643 );
not ( n88797 , n31452 );
not ( n88798 , n55481 );
not ( n88799 , n55473 );
and ( n88800 , n88799 , n31244 );
and ( n88801 , n49443 , n55473 );
or ( n88802 , n88800 , n88801 );
and ( n88803 , n88798 , n88802 );
and ( n88804 , n49443 , n55481 );
or ( n88805 , n88803 , n88804 );
and ( n88806 , n88797 , n88805 );
not ( n88807 , n55501 );
not ( n88808 , n55503 );
and ( n88809 , n88808 , n88805 );
and ( n88810 , n49469 , n55503 );
or ( n88811 , n88809 , n88810 );
and ( n88812 , n88807 , n88811 );
and ( n88813 , n49477 , n55501 );
or ( n88814 , n88812 , n88813 );
and ( n88815 , n88814 , n31452 );
or ( n88816 , n88806 , n88815 );
and ( n88817 , n88816 , n31638 );
and ( n88818 , n31244 , n47277 );
or ( n88819 , C0 , n88787 , n88796 , n88817 , n88818 );
buf ( n88820 , n88819 );
buf ( n88821 , n88820 );
buf ( n88822 , n31655 );
buf ( n88823 , n30987 );
and ( n88824 , n63070 , n32494 );
not ( n88825 , n46083 );
and ( n88826 , n88825 , n82409 );
and ( n88827 , n63076 , n46083 );
or ( n88828 , n88826 , n88827 );
and ( n88829 , n88828 , n32421 );
not ( n88830 , n46326 );
and ( n88831 , n88830 , n82409 );
and ( n88832 , n63076 , n46326 );
or ( n88833 , n88831 , n88832 );
and ( n88834 , n88833 , n32417 );
and ( n88835 , n82409 , n46340 );
or ( n88836 , n88829 , n88834 , n88835 );
and ( n88837 , n88836 , n32456 );
and ( n88838 , n82409 , n46349 );
or ( n88839 , C0 , n88824 , n88837 , n88838 );
buf ( n88840 , n88839 );
buf ( n88841 , n88840 );
buf ( n88842 , n31655 );
not ( n88843 , n46356 );
and ( n88844 , n88843 , n31144 );
not ( n88845 , n55473 );
and ( n88846 , n88845 , n31144 );
and ( n88847 , n31172 , n55473 );
or ( n88848 , n88846 , n88847 );
and ( n88849 , n88848 , n46356 );
or ( n88850 , n88844 , n88849 );
and ( n88851 , n88850 , n31649 );
not ( n88852 , n55481 );
not ( n88853 , n55473 );
and ( n88854 , n88853 , n31144 );
and ( n88855 , n46495 , n55473 );
or ( n88856 , n88854 , n88855 );
and ( n88857 , n88852 , n88856 );
and ( n88858 , n46495 , n55481 );
or ( n88859 , n88857 , n88858 );
and ( n88860 , n88859 , n31643 );
not ( n88861 , n31452 );
not ( n88862 , n55481 );
not ( n88863 , n55473 );
and ( n88864 , n88863 , n31144 );
and ( n88865 , n46495 , n55473 );
or ( n88866 , n88864 , n88865 );
and ( n88867 , n88862 , n88866 );
and ( n88868 , n46495 , n55481 );
or ( n88869 , n88867 , n88868 );
and ( n88870 , n88861 , n88869 );
not ( n88871 , n55501 );
not ( n88872 , n55503 );
and ( n88873 , n88872 , n88869 );
and ( n88874 , n46984 , n55503 );
or ( n88875 , n88873 , n88874 );
and ( n88876 , n88871 , n88875 );
and ( n88877 , n47267 , n55501 );
or ( n88878 , n88876 , n88877 );
and ( n88879 , n88878 , n31452 );
or ( n88880 , n88870 , n88879 );
and ( n88881 , n88880 , n31638 );
and ( n88882 , n31144 , n47277 );
or ( n88883 , C0 , n88851 , n88860 , n88881 , n88882 );
buf ( n88884 , n88883 );
buf ( n88885 , n88884 );
buf ( n88886 , n31655 );
buf ( n88887 , n30987 );
and ( n88888 , n64257 , n32494 );
not ( n88889 , n46083 );
and ( n88890 , n88889 , n66819 );
and ( n88891 , n64263 , n46083 );
or ( n88892 , n88890 , n88891 );
and ( n88893 , n88892 , n32421 );
not ( n88894 , n46326 );
and ( n88895 , n88894 , n66819 );
and ( n88896 , n64263 , n46326 );
or ( n88897 , n88895 , n88896 );
and ( n88898 , n88897 , n32417 );
and ( n88899 , n66819 , n46340 );
or ( n88900 , n88893 , n88898 , n88899 );
and ( n88901 , n88900 , n32456 );
and ( n88902 , n66819 , n46349 );
or ( n88903 , C0 , n88888 , n88901 , n88902 );
buf ( n88904 , n88903 );
buf ( n88905 , n88904 );
buf ( n88906 , n31655 );
not ( n88907 , n35542 );
and ( n88908 , n88907 , n41864 );
buf ( n88909 , RI15b45c30_245);
and ( n88910 , n88909 , n35542 );
or ( n88911 , n88908 , n88910 );
buf ( n88912 , n88911 );
buf ( n88913 , n88912 );
buf ( n88914 , n31655 );
not ( n88915 , n33419 );
and ( n88916 , n88915 , n31589 );
xor ( n88917 , n33630 , n33647 );
xor ( n88918 , n88917 , n33667 );
and ( n88919 , n88918 , n33419 );
or ( n88920 , n88916 , n88919 );
and ( n88921 , n88920 , n31529 );
not ( n88922 , n33734 );
and ( n88923 , n88922 , n31589 );
not ( n88924 , n33533 );
xor ( n88925 , n33783 , n33647 );
xor ( n88926 , n88925 , n33785 );
and ( n88927 , n88924 , n88926 );
xor ( n88928 , n33880 , n33882 );
xor ( n88929 , n88928 , n33887 );
and ( n88930 , n88929 , n33533 );
or ( n88931 , n88927 , n88930 );
and ( n88932 , n88931 , n33734 );
or ( n88933 , n88923 , n88932 );
and ( n88934 , n88933 , n31527 );
and ( n88935 , n31589 , n33942 );
or ( n88936 , n88921 , n88934 , n88935 );
and ( n88937 , n88936 , n31557 );
and ( n88938 , n31626 , n31643 );
not ( n88939 , n31452 );
and ( n88940 , n88939 , n31626 );
and ( n88941 , n31589 , n31452 );
or ( n88942 , n88940 , n88941 );
and ( n88943 , n88942 , n31638 );
and ( n88944 , n31460 , n33973 );
and ( n88945 , n31589 , n33978 );
or ( n88946 , C0 , n88937 , n88938 , n88943 , n88944 , n88945 );
buf ( n88947 , n88946 );
buf ( n88948 , n88947 );
not ( n88949 , n40163 );
and ( n88950 , n88949 , n31657 );
buf ( n88951 , n88950 );
and ( n88952 , n88951 , n32498 );
not ( n88953 , n55780 );
not ( n88954 , n55558 );
and ( n88955 , n88954 , n31657 );
buf ( n88956 , n88955 );
and ( n88957 , n88953 , n88956 );
buf ( n88958 , n88957 );
and ( n88959 , n88958 , n32496 );
and ( n88960 , n31657 , n55800 );
or ( n88961 , C0 , n88952 , n88959 , C0 , C0 , n88960 );
buf ( n88962 , n88961 );
buf ( n88963 , n88962 );
buf ( n88964 , n30987 );
buf ( n88965 , n30987 );
buf ( n88966 , n31655 );
not ( n88967 , n31077 );
and ( n88968 , n75795 , n88967 );
and ( n88969 , n88968 , n31373 );
not ( n88970 , n31402 );
and ( n88971 , n75795 , n88970 );
and ( n88972 , n88971 , n31408 );
not ( n88973 , n31437 );
and ( n88974 , n88973 , n75795 );
buf ( n88975 , n31437 );
or ( n88976 , n88974 , n88975 );
and ( n88977 , n88976 , n31468 );
not ( n88978 , n31497 );
and ( n88979 , n88978 , n75795 );
buf ( n88980 , n31497 );
or ( n88981 , n88979 , n88980 );
and ( n88982 , n88981 , n31521 );
and ( n88983 , n75795 , n31553 );
or ( n88984 , n88969 , n88972 , n88977 , n88982 , n88983 );
and ( n88985 , n88984 , n31557 );
and ( n88986 , n75795 , n52894 );
buf ( n88987 , n52896 );
or ( n88988 , C0 , n88985 , n88986 , n88987 );
buf ( n88989 , n88988 );
buf ( n88990 , n88989 );
not ( n88991 , n40163 );
and ( n88992 , n88991 , n31908 );
not ( n88993 , n52903 );
and ( n88994 , n88993 , n31908 );
and ( n88995 , n32200 , n52903 );
or ( n88996 , n88994 , n88995 );
and ( n88997 , n88996 , n40163 );
or ( n88998 , n88992 , n88997 );
and ( n88999 , n88998 , n32498 );
not ( n89000 , n52911 );
not ( n89001 , n52903 );
and ( n89002 , n89001 , n31908 );
and ( n89003 , n53243 , n52903 );
or ( n89004 , n89002 , n89003 );
and ( n89005 , n89000 , n89004 );
and ( n89006 , n53243 , n52911 );
or ( n89007 , n89005 , n89006 );
and ( n89008 , n89007 , n32473 );
not ( n89009 , n32475 );
not ( n89010 , n52911 );
not ( n89011 , n52903 );
and ( n89012 , n89011 , n31908 );
and ( n89013 , n53243 , n52903 );
or ( n89014 , n89012 , n89013 );
and ( n89015 , n89010 , n89014 );
and ( n89016 , n53243 , n52911 );
or ( n89017 , n89015 , n89016 );
and ( n89018 , n89009 , n89017 );
not ( n89019 , n52931 );
not ( n89020 , n52933 );
and ( n89021 , n89020 , n89017 );
and ( n89022 , n53269 , n52933 );
or ( n89023 , n89021 , n89022 );
and ( n89024 , n89019 , n89023 );
and ( n89025 , n53277 , n52931 );
or ( n89026 , n89024 , n89025 );
and ( n89027 , n89026 , n32475 );
or ( n89028 , n89018 , n89027 );
and ( n89029 , n89028 , n32486 );
and ( n89030 , n31908 , n41278 );
or ( n89031 , C0 , n88999 , n89008 , n89029 , n89030 );
buf ( n89032 , n89031 );
buf ( n89033 , n89032 );
buf ( n89034 , n30987 );
buf ( n89035 , n30987 );
not ( n89036 , n32953 );
and ( n89037 , n89036 , n65456 );
and ( n89038 , n65476 , n32953 );
or ( n89039 , n89037 , n89038 );
and ( n89040 , n89039 , n33038 );
not ( n89041 , n48660 );
and ( n89042 , n89041 , n65456 );
and ( n89043 , n55367 , n48660 );
or ( n89044 , n89042 , n89043 );
and ( n89045 , n89044 , n33172 );
and ( n89046 , n65456 , n39795 );
or ( n89047 , n89040 , n89045 , n89046 );
and ( n89048 , n89047 , n33208 );
and ( n89049 , n65456 , n39805 );
or ( n89050 , C0 , n89048 , n89049 );
buf ( n89051 , n89050 );
buf ( n89052 , n89051 );
buf ( n89053 , n30987 );
buf ( n89054 , n30987 );
buf ( n89055 , n31655 );
buf ( n89056 , n31655 );
buf ( n89057 , n30987 );
buf ( n89058 , n30987 );
not ( n89059 , n34150 );
and ( n89060 , n89059 , n32801 );
not ( n89061 , n58762 );
and ( n89062 , n89061 , n32801 );
and ( n89063 , n32823 , n58762 );
or ( n89064 , n89062 , n89063 );
and ( n89065 , n89064 , n34150 );
or ( n89066 , n89060 , n89065 );
and ( n89067 , n89066 , n33381 );
not ( n89068 , n58770 );
not ( n89069 , n58762 );
and ( n89070 , n89069 , n32801 );
and ( n89071 , n41464 , n58762 );
or ( n89072 , n89070 , n89071 );
and ( n89073 , n89068 , n89072 );
and ( n89074 , n41464 , n58770 );
or ( n89075 , n89073 , n89074 );
and ( n89076 , n89075 , n33375 );
not ( n89077 , n32968 );
not ( n89078 , n58770 );
not ( n89079 , n58762 );
and ( n89080 , n89079 , n32801 );
and ( n89081 , n41464 , n58762 );
or ( n89082 , n89080 , n89081 );
and ( n89083 , n89078 , n89082 );
and ( n89084 , n41464 , n58770 );
or ( n89085 , n89083 , n89084 );
and ( n89086 , n89077 , n89085 );
not ( n89087 , n58790 );
not ( n89088 , n58792 );
and ( n89089 , n89088 , n89085 );
and ( n89090 , n41490 , n58792 );
or ( n89091 , n89089 , n89090 );
and ( n89092 , n89087 , n89091 );
and ( n89093 , n41500 , n58790 );
or ( n89094 , n89092 , n89093 );
and ( n89095 , n89094 , n32968 );
or ( n89096 , n89086 , n89095 );
and ( n89097 , n89096 , n33370 );
and ( n89098 , n32801 , n35062 );
or ( n89099 , C0 , n89067 , n89076 , n89097 , n89098 );
buf ( n89100 , n89099 );
buf ( n89101 , n89100 );
buf ( n89102 , n31655 );
buf ( n89103 , n31655 );
buf ( n89104 , n31655 );
not ( n89105 , n31451 );
and ( n89106 , n89105 , n30993 );
buf ( n89107 , n89106 );
and ( n89108 , n89107 , n31645 );
not ( n89109 , n63845 );
not ( n89110 , n63847 );
and ( n89111 , n89110 , n30993 );
buf ( n89112 , n63847 );
or ( n89113 , n89111 , n89112 );
and ( n89114 , n89113 , n31468 );
and ( n89115 , n30993 , n63859 );
or ( n89116 , n89114 , n89115 );
and ( n89117 , n89109 , n89116 );
buf ( n89118 , n63845 );
or ( n89119 , n89117 , n89118 );
and ( n89120 , n89119 , n31557 );
and ( n89121 , n59060 , n31641 );
not ( n89122 , n31452 );
and ( n89123 , n89122 , n31638 );
not ( n89124 , n59060 );
and ( n89125 , n89124 , n31640 );
or ( n89126 , C0 , C0 , C0 , n89108 , n89120 , C0 , n89121 , n89123 , n89125 , C0 );
buf ( n89127 , n89126 );
buf ( n89128 , n89127 );
buf ( n89129 , n30987 );
not ( n89130 , n38443 );
and ( n89131 , n89130 , n38082 );
xor ( n89132 , n53477 , n53492 );
and ( n89133 , n89132 , n38443 );
or ( n89134 , n89131 , n89133 );
and ( n89135 , n89134 , n38450 );
not ( n89136 , n39339 );
and ( n89137 , n89136 , n38982 );
xor ( n89138 , n53533 , n53548 );
and ( n89139 , n89138 , n39339 );
or ( n89140 , n89137 , n89139 );
and ( n89141 , n89140 , n39346 );
and ( n89142 , n40207 , n39359 );
or ( n89143 , n89135 , n89141 , n89142 );
buf ( n89144 , n89143 );
buf ( n89145 , n89144 );
not ( n89146 , n46356 );
and ( n89147 , n89146 , n31156 );
not ( n89148 , n55263 );
and ( n89149 , n89148 , n31156 );
and ( n89150 , n31172 , n55263 );
or ( n89151 , n89149 , n89150 );
and ( n89152 , n89151 , n46356 );
or ( n89153 , n89147 , n89152 );
and ( n89154 , n89153 , n31649 );
not ( n89155 , n55271 );
not ( n89156 , n55263 );
and ( n89157 , n89156 , n31156 );
and ( n89158 , n46495 , n55263 );
or ( n89159 , n89157 , n89158 );
and ( n89160 , n89155 , n89159 );
and ( n89161 , n46495 , n55271 );
or ( n89162 , n89160 , n89161 );
and ( n89163 , n89162 , n31643 );
not ( n89164 , n31452 );
not ( n89165 , n55271 );
not ( n89166 , n55263 );
and ( n89167 , n89166 , n31156 );
and ( n89168 , n46495 , n55263 );
or ( n89169 , n89167 , n89168 );
and ( n89170 , n89165 , n89169 );
and ( n89171 , n46495 , n55271 );
or ( n89172 , n89170 , n89171 );
and ( n89173 , n89164 , n89172 );
not ( n89174 , n55291 );
not ( n89175 , n55293 );
and ( n89176 , n89175 , n89172 );
and ( n89177 , n46984 , n55293 );
or ( n89178 , n89176 , n89177 );
and ( n89179 , n89174 , n89178 );
and ( n89180 , n47267 , n55291 );
or ( n89181 , n89179 , n89180 );
and ( n89182 , n89181 , n31452 );
or ( n89183 , n89173 , n89182 );
and ( n89184 , n89183 , n31638 );
and ( n89185 , n31156 , n47277 );
or ( n89186 , C0 , n89154 , n89163 , n89184 , n89185 );
buf ( n89187 , n89186 );
buf ( n89188 , n89187 );
buf ( n89189 , n31655 );
buf ( n89190 , n30987 );
xor ( n89191 , n46172 , n49992 );
and ( n89192 , n89191 , n32431 );
not ( n89193 , n50002 );
and ( n89194 , n89193 , n46172 );
and ( n89195 , n40359 , n50002 );
or ( n89196 , n89194 , n89195 );
and ( n89197 , n89196 , n32419 );
not ( n89198 , n50008 );
and ( n89199 , n89198 , n46172 );
not ( n89200 , n47910 );
and ( n89201 , n89200 , n47900 );
and ( n89202 , n48121 , n47910 );
or ( n89203 , n89201 , n89202 );
and ( n89204 , n89203 , n50008 );
or ( n89205 , n89199 , n89204 );
and ( n89206 , n89205 , n32415 );
not ( n89207 , n50067 );
and ( n89208 , n89207 , n46172 );
and ( n89209 , n31823 , n50067 );
or ( n89210 , n89208 , n89209 );
and ( n89211 , n89210 , n32411 );
and ( n89212 , n46172 , n50098 );
or ( n89213 , n89192 , n89197 , n89206 , n89211 , n89212 );
and ( n89214 , n89213 , n32456 );
and ( n89215 , n46172 , n47409 );
or ( n89216 , C0 , n89214 , n89215 );
buf ( n89217 , n89216 );
buf ( n89218 , n89217 );
buf ( n89219 , n31655 );
and ( n89220 , n49075 , n48639 );
not ( n89221 , n48642 );
and ( n89222 , n89221 , n48600 );
and ( n89223 , n49075 , n48642 );
or ( n89224 , n89222 , n89223 );
and ( n89225 , n89224 , n32890 );
not ( n89226 , n48648 );
and ( n89227 , n89226 , n48600 );
and ( n89228 , n49075 , n48648 );
or ( n89229 , n89227 , n89228 );
and ( n89230 , n89229 , n32924 );
not ( n89231 , n48654 );
and ( n89232 , n89231 , n48600 );
and ( n89233 , n49075 , n48654 );
or ( n89234 , n89232 , n89233 );
and ( n89235 , n89234 , n33038 );
not ( n89236 , n48660 );
and ( n89237 , n89236 , n48600 );
and ( n89238 , n49075 , n48660 );
or ( n89239 , n89237 , n89238 );
and ( n89240 , n89239 , n33172 );
not ( n89241 , n41576 );
and ( n89242 , n89241 , n48600 );
and ( n89243 , n48785 , n41576 );
or ( n89244 , n89242 , n89243 );
and ( n89245 , n89244 , n33189 );
not ( n89246 , n48730 );
and ( n89247 , n89246 , n48600 );
and ( n89248 , n48785 , n48730 );
or ( n89249 , n89247 , n89248 );
and ( n89250 , n89249 , n33187 );
not ( n89251 , n48765 );
and ( n89252 , n89251 , n48600 );
xor ( n89253 , n48785 , n49003 );
and ( n89254 , n89253 , n48765 );
or ( n89255 , n89252 , n89254 );
and ( n89256 , n89255 , n33180 );
not ( n89257 , n49054 );
and ( n89258 , n89257 , n48600 );
not ( n89259 , n48845 );
xor ( n89260 , n49075 , n49117 );
and ( n89261 , n89259 , n89260 );
xnor ( n89262 , n49184 , n49243 );
and ( n89263 , n89262 , n48845 );
or ( n89264 , n89261 , n89263 );
and ( n89265 , n89264 , n49054 );
or ( n89266 , n89258 , n89265 );
and ( n89267 , n89266 , n33178 );
and ( n89268 , n49184 , n49275 );
or ( n89269 , n89220 , n89225 , n89230 , n89235 , n89240 , n89245 , n89250 , n89256 , n89267 , n89268 );
and ( n89270 , n89269 , n33208 );
and ( n89271 , n32993 , n35056 );
and ( n89272 , n48600 , n49286 );
or ( n89273 , C0 , n89270 , n89271 , n89272 );
buf ( n89274 , n89273 );
buf ( n89275 , n89274 );
buf ( n89276 , n30987 );
buf ( n89277 , n30987 );
buf ( n89278 , n31655 );
buf ( n89279 , n31655 );
buf ( n89280 , n30987 );
not ( n89281 , n34150 );
and ( n89282 , n89281 , n32824 );
not ( n89283 , n56708 );
and ( n89284 , n89283 , n32824 );
and ( n89285 , n32856 , n56708 );
or ( n89286 , n89284 , n89285 );
and ( n89287 , n89286 , n34150 );
or ( n89288 , n89282 , n89287 );
and ( n89289 , n89288 , n33381 );
not ( n89290 , n56716 );
not ( n89291 , n56708 );
and ( n89292 , n89291 , n32824 );
and ( n89293 , n48160 , n56708 );
or ( n89294 , n89292 , n89293 );
and ( n89295 , n89290 , n89294 );
and ( n89296 , n48160 , n56716 );
or ( n89297 , n89295 , n89296 );
and ( n89298 , n89297 , n33375 );
not ( n89299 , n32968 );
not ( n89300 , n56716 );
not ( n89301 , n56708 );
and ( n89302 , n89301 , n32824 );
and ( n89303 , n48160 , n56708 );
or ( n89304 , n89302 , n89303 );
and ( n89305 , n89300 , n89304 );
and ( n89306 , n48160 , n56716 );
or ( n89307 , n89305 , n89306 );
and ( n89308 , n89299 , n89307 );
not ( n89309 , n56736 );
not ( n89310 , n56738 );
and ( n89311 , n89310 , n89307 );
and ( n89312 , n48186 , n56738 );
or ( n89313 , n89311 , n89312 );
and ( n89314 , n89309 , n89313 );
and ( n89315 , n48196 , n56736 );
or ( n89316 , n89314 , n89315 );
and ( n89317 , n89316 , n32968 );
or ( n89318 , n89308 , n89317 );
and ( n89319 , n89318 , n33370 );
and ( n89320 , n32824 , n35062 );
or ( n89321 , C0 , n89289 , n89298 , n89319 , n89320 );
buf ( n89322 , n89321 );
buf ( n89323 , n89322 );
buf ( n89324 , n30987 );
buf ( n89325 , n31655 );
buf ( n89326 , n31655 );
buf ( n89327 , n31655 );
not ( n89328 , n31437 );
and ( n89329 , n89328 , n53287 );
and ( n89330 , n53300 , n31437 );
or ( n89331 , n89329 , n89330 );
and ( n89332 , n89331 , n31468 );
not ( n89333 , n41837 );
and ( n89334 , n89333 , n53287 );
not ( n89335 , n42124 );
and ( n89336 , n89335 , n42040 );
xor ( n89337 , n49378 , n49381 );
and ( n89338 , n89337 , n42124 );
or ( n89339 , n89336 , n89338 );
and ( n89340 , n89339 , n41837 );
or ( n89341 , n89334 , n89340 );
and ( n89342 , n89341 , n31521 );
and ( n89343 , n53287 , n42158 );
or ( n89344 , n89332 , n89342 , n89343 );
and ( n89345 , n89344 , n31557 );
and ( n89346 , n53287 , n40154 );
or ( n89347 , C0 , n89345 , n89346 );
buf ( n89348 , n89347 );
buf ( n89349 , n89348 );
not ( n89350 , n40163 );
and ( n89351 , n89350 , n31898 );
not ( n89352 , n42171 );
and ( n89353 , n89352 , n31898 );
and ( n89354 , n32200 , n42171 );
or ( n89355 , n89353 , n89354 );
and ( n89356 , n89355 , n40163 );
or ( n89357 , n89351 , n89356 );
and ( n89358 , n89357 , n32498 );
not ( n89359 , n42180 );
not ( n89360 , n42171 );
and ( n89361 , n89360 , n31898 );
and ( n89362 , n53243 , n42171 );
or ( n89363 , n89361 , n89362 );
and ( n89364 , n89359 , n89363 );
and ( n89365 , n53243 , n42180 );
or ( n89366 , n89364 , n89365 );
and ( n89367 , n89366 , n32473 );
not ( n89368 , n32475 );
not ( n89369 , n42180 );
not ( n89370 , n42171 );
and ( n89371 , n89370 , n31898 );
and ( n89372 , n53243 , n42171 );
or ( n89373 , n89371 , n89372 );
and ( n89374 , n89369 , n89373 );
and ( n89375 , n53243 , n42180 );
or ( n89376 , n89374 , n89375 );
and ( n89377 , n89368 , n89376 );
not ( n89378 , n42206 );
not ( n89379 , n42209 );
and ( n89380 , n89379 , n89376 );
and ( n89381 , n53269 , n42209 );
or ( n89382 , n89380 , n89381 );
and ( n89383 , n89378 , n89382 );
and ( n89384 , n53277 , n42206 );
or ( n89385 , n89383 , n89384 );
and ( n89386 , n89385 , n32475 );
or ( n89387 , n89377 , n89386 );
and ( n89388 , n89387 , n32486 );
and ( n89389 , n31898 , n41278 );
or ( n89390 , C0 , n89358 , n89367 , n89388 , n89389 );
buf ( n89391 , n89390 );
buf ( n89392 , n89391 );
buf ( n89393 , n30987 );
not ( n89394 , n35542 );
and ( n89395 , n89394 , n41852 );
and ( n89396 , n74110 , n35542 );
or ( n89397 , n89395 , n89396 );
buf ( n89398 , n89397 );
buf ( n89399 , n89398 );
buf ( n89400 , n31655 );
not ( n89401 , n33419 );
and ( n89402 , n89401 , n31587 );
and ( n89403 , n71869 , n33419 );
or ( n89404 , n89402 , n89403 );
and ( n89405 , n89404 , n31529 );
not ( n89406 , n33734 );
and ( n89407 , n89406 , n31587 );
and ( n89408 , n71882 , n33734 );
or ( n89409 , n89407 , n89408 );
and ( n89410 , n89409 , n31527 );
and ( n89411 , n31587 , n33942 );
or ( n89412 , n89405 , n89410 , n89411 );
and ( n89413 , n89412 , n31557 );
and ( n89414 , n34119 , n31643 );
not ( n89415 , n31452 );
and ( n89416 , n89415 , n34119 );
xor ( n89417 , n31587 , n33950 );
and ( n89418 , n89417 , n31452 );
or ( n89419 , n89416 , n89418 );
and ( n89420 , n89419 , n31638 );
and ( n89421 , n34011 , n33973 );
and ( n89422 , n31587 , n33978 );
or ( n89423 , C0 , n89413 , n89414 , n89420 , n89421 , n89422 );
buf ( n89424 , n89423 );
buf ( n89425 , n89424 );
not ( n89426 , n40163 );
and ( n89427 , n89426 , n31669 );
and ( n89428 , n40182 , n40163 );
or ( n89429 , n89427 , n89428 );
and ( n89430 , n89429 , n32498 );
not ( n89431 , n55780 );
not ( n89432 , n55558 );
and ( n89433 , n89432 , n31669 );
buf ( n89434 , n89433 );
and ( n89435 , n89431 , n89434 );
buf ( n89436 , n89435 );
and ( n89437 , n89436 , n32496 );
and ( n89438 , n40421 , n32473 );
not ( n89439 , n32475 );
and ( n89440 , n89439 , n40421 );
xor ( n89441 , n40425 , n40417 );
not ( n89442 , n89441 );
buf ( n89443 , n89442 );
not ( n89444 , n89443 );
and ( n89445 , n89444 , n32475 );
or ( n89446 , n89440 , n89445 );
and ( n89447 , n89446 , n32486 );
and ( n89448 , n31669 , n55800 );
or ( n89449 , C0 , n89430 , n89437 , n89438 , n89447 , n89448 );
buf ( n89450 , n89449 );
buf ( n89451 , n89450 );
buf ( n89452 , n30987 );
buf ( n89453 , n30987 );
buf ( n89454 , n30987 );
buf ( n89455 , n30987 );
not ( n89456 , n43755 );
and ( n89457 , n89456 , n43751 );
xor ( n89458 , n43751 , n43259 );
and ( n89459 , n52299 , n52330 );
xor ( n89460 , n89458 , n89459 );
and ( n89461 , n89460 , n43755 );
or ( n89462 , n89457 , n89461 );
and ( n89463 , n89462 , n43774 );
not ( n89464 , n44663 );
and ( n89465 , n89464 , n44659 );
xor ( n89466 , n44659 , n44171 );
and ( n89467 , n52337 , n52368 );
xor ( n89468 , n89466 , n89467 );
and ( n89469 , n89468 , n44663 );
or ( n89470 , n89465 , n89469 );
and ( n89471 , n89470 , n44682 );
and ( n89472 , n75493 , n44695 );
or ( n89473 , n89463 , n89471 , n89472 );
buf ( n89474 , n89473 );
buf ( n89475 , n89474 );
buf ( n89476 , n31655 );
buf ( n89477 , n31655 );
buf ( n89478 , n31655 );
xor ( n89479 , n33077 , n58395 );
and ( n89480 , n89479 , n33201 );
not ( n89481 , n41576 );
and ( n89482 , n89481 , n33077 );
xor ( n89483 , n58489 , n58596 );
and ( n89484 , n89483 , n41576 );
or ( n89485 , n89482 , n89484 );
and ( n89486 , n89485 , n33189 );
and ( n89487 , n33077 , n41592 );
or ( n89488 , n89480 , n89486 , n89487 );
and ( n89489 , n89488 , n33208 );
and ( n89490 , n33077 , n39805 );
or ( n89491 , C0 , n89489 , n89490 );
buf ( n89492 , n89491 );
buf ( n89493 , n89492 );
buf ( n89494 , n30987 );
buf ( n89495 , n30987 );
buf ( n89496 , n31655 );
not ( n89497 , n50828 );
not ( n89498 , n50834 );
and ( n89499 , n89498 , n40498 );
and ( n89500 , n53290 , n50834 );
or ( n89501 , n89499 , n89500 );
and ( n89502 , n89497 , n89501 );
and ( n89503 , n77679 , n50828 );
or ( n89504 , n89502 , n89503 );
buf ( n89505 , n89504 );
buf ( n89506 , n89505 );
xor ( n89507 , n33095 , n58386 );
and ( n89508 , n89507 , n33201 );
not ( n89509 , n41576 );
and ( n89510 , n89509 , n33095 );
and ( n89511 , n73036 , n41576 );
or ( n89512 , n89510 , n89511 );
and ( n89513 , n89512 , n33189 );
and ( n89514 , n33095 , n41592 );
or ( n89515 , n89508 , n89513 , n89514 );
and ( n89516 , n89515 , n33208 );
and ( n89517 , n33095 , n39805 );
or ( n89518 , C0 , n89516 , n89517 );
buf ( n89519 , n89518 );
buf ( n89520 , n89519 );
buf ( n89521 , n31655 );
buf ( n89522 , n30987 );
buf ( n89523 , n30987 );
buf ( n89524 , n31655 );
not ( n89525 , n50828 );
not ( n89526 , n50834 );
and ( n89527 , n89526 , n40632 );
and ( n89528 , n54606 , n50834 );
or ( n89529 , n89527 , n89528 );
and ( n89530 , n89525 , n89529 );
and ( n89531 , n78758 , n50828 );
or ( n89532 , n89530 , n89531 );
buf ( n89533 , n89532 );
buf ( n89534 , n89533 );
buf ( n89535 , n30987 );
not ( n89536 , n48765 );
and ( n89537 , n89536 , n33230 );
and ( n89538 , n89253 , n48765 );
or ( n89539 , n89537 , n89538 );
and ( n89540 , n89539 , n33180 );
not ( n89541 , n49054 );
and ( n89542 , n89541 , n33230 );
and ( n89543 , n89264 , n49054 );
or ( n89544 , n89542 , n89543 );
and ( n89545 , n89544 , n33178 );
and ( n89546 , n33230 , n49774 );
or ( n89547 , n89540 , n89545 , n89546 );
and ( n89548 , n89547 , n33208 );
and ( n89549 , n33311 , n33375 );
not ( n89550 , n32968 );
and ( n89551 , n89550 , n33311 );
xor ( n89552 , n33230 , n53899 );
and ( n89553 , n89552 , n32968 );
or ( n89554 , n89551 , n89553 );
and ( n89555 , n89554 , n33370 );
and ( n89556 , n32993 , n35056 );
and ( n89557 , n33230 , n49794 );
or ( n89558 , C0 , n89548 , n89549 , n89555 , n89556 , n89557 );
buf ( n89559 , n89558 );
buf ( n89560 , n89559 );
buf ( n89561 , n31655 );
buf ( n89562 , n30987 );
buf ( n89563 , n31655 );
and ( n89564 , n46020 , n32500 );
not ( n89565 , n35211 );
and ( n89566 , n89565 , n37537 );
buf ( n89567 , n89566 );
and ( n89568 , n89567 , n32421 );
not ( n89569 , n35245 );
and ( n89570 , n89569 , n37537 );
buf ( n89571 , n89570 );
and ( n89572 , n89571 , n32419 );
not ( n89573 , n35278 );
and ( n89574 , n89573 , n37537 );
not ( n89575 , n35295 );
and ( n89576 , n89575 , n49567 );
xor ( n89577 , n37537 , n49547 );
and ( n89578 , n89577 , n35295 );
or ( n89579 , n89576 , n89578 );
and ( n89580 , n89579 , n35278 );
or ( n89581 , n89574 , n89580 );
and ( n89582 , n89581 , n32417 );
not ( n89583 , n35331 );
and ( n89584 , n89583 , n37537 );
not ( n89585 , n35294 );
not ( n89586 , n45995 );
and ( n89587 , n89586 , n49567 );
xor ( n89588 , n49568 , n49633 );
and ( n89589 , n89588 , n45995 );
or ( n89590 , n89587 , n89589 );
and ( n89591 , n89585 , n89590 );
and ( n89592 , n89577 , n35294 );
or ( n89593 , n89591 , n89592 );
and ( n89594 , n89593 , n35331 );
or ( n89595 , n89584 , n89594 );
and ( n89596 , n89595 , n32415 );
and ( n89597 , n37537 , n35354 );
or ( n89598 , n89568 , n89572 , n89582 , n89596 , n89597 );
and ( n89599 , n89598 , n32456 );
not ( n89600 , n32475 );
not ( n89601 , n46060 );
and ( n89602 , n89601 , n49658 );
xor ( n89603 , n49659 , n49727 );
and ( n89604 , n89603 , n46060 );
or ( n89605 , n89602 , n89604 );
and ( n89606 , n89600 , n89605 );
and ( n89607 , n37537 , n32475 );
or ( n89608 , n89606 , n89607 );
and ( n89609 , n89608 , n32486 );
and ( n89610 , n37537 , n35367 );
or ( n89611 , C0 , n89564 , n89599 , n89609 , C0 , n89610 );
buf ( n89612 , n89611 );
buf ( n89613 , n89612 );
and ( n89614 , n49069 , n48639 );
not ( n89615 , n48642 );
and ( n89616 , n89615 , n48594 );
and ( n89617 , n49069 , n48642 );
or ( n89618 , n89616 , n89617 );
and ( n89619 , n89618 , n32890 );
not ( n89620 , n48648 );
and ( n89621 , n89620 , n48594 );
and ( n89622 , n49069 , n48648 );
or ( n89623 , n89621 , n89622 );
and ( n89624 , n89623 , n32924 );
not ( n89625 , n48654 );
and ( n89626 , n89625 , n48594 );
and ( n89627 , n49069 , n48654 );
or ( n89628 , n89626 , n89627 );
and ( n89629 , n89628 , n33038 );
not ( n89630 , n48660 );
and ( n89631 , n89630 , n48594 );
and ( n89632 , n49069 , n48660 );
or ( n89633 , n89631 , n89632 );
and ( n89634 , n89633 , n33172 );
not ( n89635 , n41576 );
and ( n89636 , n89635 , n48594 );
and ( n89637 , n48779 , n41576 );
or ( n89638 , n89636 , n89637 );
and ( n89639 , n89638 , n33189 );
not ( n89640 , n48730 );
and ( n89641 , n89640 , n48594 );
and ( n89642 , n48779 , n48730 );
or ( n89643 , n89641 , n89642 );
and ( n89644 , n89643 , n33187 );
not ( n89645 , n48765 );
and ( n89646 , n89645 , n48594 );
xor ( n89647 , n48779 , n49009 );
and ( n89648 , n89647 , n48765 );
or ( n89649 , n89646 , n89648 );
and ( n89650 , n89649 , n33180 );
not ( n89651 , n49054 );
and ( n89652 , n89651 , n48594 );
not ( n89653 , n48845 );
xor ( n89654 , n49069 , n49123 );
and ( n89655 , n89653 , n89654 );
xnor ( n89656 , n49178 , n49249 );
and ( n89657 , n89656 , n48845 );
or ( n89658 , n89655 , n89657 );
and ( n89659 , n89658 , n49054 );
or ( n89660 , n89652 , n89659 );
and ( n89661 , n89660 , n33178 );
and ( n89662 , n49178 , n49275 );
or ( n89663 , n89614 , n89619 , n89624 , n89629 , n89634 , n89639 , n89644 , n89650 , n89661 , n89662 );
and ( n89664 , n89663 , n33208 );
and ( n89665 , n32987 , n35056 );
and ( n89666 , n48594 , n49286 );
or ( n89667 , C0 , n89664 , n89665 , n89666 );
buf ( n89668 , n89667 );
buf ( n89669 , n89668 );
buf ( n89670 , n30987 );
buf ( n89671 , n30987 );
buf ( n89672 , n31655 );
buf ( n89673 , n31655 );
buf ( n89674 , n30987 );
buf ( n89675 , n30987 );
not ( n89676 , n34150 );
and ( n89677 , n89676 , n32797 );
not ( n89678 , n59574 );
and ( n89679 , n89678 , n32797 );
and ( n89680 , n32823 , n59574 );
or ( n89681 , n89679 , n89680 );
and ( n89682 , n89681 , n34150 );
or ( n89683 , n89677 , n89682 );
and ( n89684 , n89683 , n33381 );
not ( n89685 , n59582 );
not ( n89686 , n59574 );
and ( n89687 , n89686 , n32797 );
and ( n89688 , n41464 , n59574 );
or ( n89689 , n89687 , n89688 );
and ( n89690 , n89685 , n89689 );
and ( n89691 , n41464 , n59582 );
or ( n89692 , n89690 , n89691 );
and ( n89693 , n89692 , n33375 );
not ( n89694 , n32968 );
not ( n89695 , n59582 );
not ( n89696 , n59574 );
and ( n89697 , n89696 , n32797 );
and ( n89698 , n41464 , n59574 );
or ( n89699 , n89697 , n89698 );
and ( n89700 , n89695 , n89699 );
and ( n89701 , n41464 , n59582 );
or ( n89702 , n89700 , n89701 );
and ( n89703 , n89694 , n89702 );
not ( n89704 , n59602 );
not ( n89705 , n59604 );
and ( n89706 , n89705 , n89702 );
and ( n89707 , n41490 , n59604 );
or ( n89708 , n89706 , n89707 );
and ( n89709 , n89704 , n89708 );
and ( n89710 , n41500 , n59602 );
or ( n89711 , n89709 , n89710 );
and ( n89712 , n89711 , n32968 );
or ( n89713 , n89703 , n89712 );
and ( n89714 , n89713 , n33370 );
and ( n89715 , n32797 , n35062 );
or ( n89716 , C0 , n89684 , n89693 , n89714 , n89715 );
buf ( n89717 , n89716 );
buf ( n89718 , n89717 );
buf ( n89719 , n31655 );
buf ( n89720 , n31655 );
buf ( n89721 , n31655 );
xor ( n89722 , n31457 , n39925 );
and ( n89723 , n89722 , n31550 );
not ( n89724 , n39979 );
and ( n89725 , n89724 , n31457 );
buf ( n89726 , n31236 );
and ( n89727 , n89726 , n39979 );
or ( n89728 , n89725 , n89727 );
and ( n89729 , n89728 , n31538 );
and ( n89730 , n31457 , n40143 );
or ( n89731 , n89723 , n89729 , n89730 );
and ( n89732 , n89731 , n31557 );
and ( n89733 , n31457 , n40154 );
or ( n89734 , C0 , n89732 , n89733 );
buf ( n89735 , n89734 );
buf ( n89736 , n89735 );
not ( n89737 , n40163 );
and ( n89738 , n89737 , n31885 );
not ( n89739 , n57233 );
and ( n89740 , n89739 , n31885 );
and ( n89741 , n32218 , n57233 );
or ( n89742 , n89740 , n89741 );
and ( n89743 , n89742 , n40163 );
or ( n89744 , n89738 , n89743 );
and ( n89745 , n89744 , n32498 );
not ( n89746 , n57241 );
not ( n89747 , n57233 );
and ( n89748 , n89747 , n31885 );
and ( n89749 , n42255 , n57233 );
or ( n89750 , n89748 , n89749 );
and ( n89751 , n89746 , n89750 );
and ( n89752 , n42255 , n57241 );
or ( n89753 , n89751 , n89752 );
and ( n89754 , n89753 , n32473 );
not ( n89755 , n32475 );
not ( n89756 , n57241 );
not ( n89757 , n57233 );
and ( n89758 , n89757 , n31885 );
and ( n89759 , n42255 , n57233 );
or ( n89760 , n89758 , n89759 );
and ( n89761 , n89756 , n89760 );
and ( n89762 , n42255 , n57241 );
or ( n89763 , n89761 , n89762 );
and ( n89764 , n89755 , n89763 );
not ( n89765 , n57261 );
not ( n89766 , n57263 );
and ( n89767 , n89766 , n89763 );
and ( n89768 , n42283 , n57263 );
or ( n89769 , n89767 , n89768 );
and ( n89770 , n89765 , n89769 );
and ( n89771 , n42291 , n57261 );
or ( n89772 , n89770 , n89771 );
and ( n89773 , n89772 , n32475 );
or ( n89774 , n89764 , n89773 );
and ( n89775 , n89774 , n32486 );
and ( n89776 , n31885 , n41278 );
or ( n89777 , C0 , n89745 , n89754 , n89775 , n89776 );
buf ( n89778 , n89777 );
buf ( n89779 , n89778 );
buf ( n89780 , n30987 );
buf ( n89781 , n30987 );
buf ( n89782 , n31655 );
not ( n89783 , n52869 );
and ( n89784 , n89783 , n58921 );
and ( n89785 , n41525 , n37506 );
or ( n89786 , n89784 , n89785 );
buf ( n89787 , n89786 );
buf ( n89788 , n89787 );
and ( n89789 , n47662 , n50275 );
not ( n89790 , n50278 );
and ( n89791 , n89790 , n47575 );
and ( n89792 , n47662 , n50278 );
or ( n89793 , n89791 , n89792 );
and ( n89794 , n89793 , n32421 );
not ( n89795 , n50002 );
and ( n89796 , n89795 , n47575 );
and ( n89797 , n47662 , n50002 );
or ( n89798 , n89796 , n89797 );
and ( n89799 , n89798 , n32419 );
not ( n89800 , n50289 );
and ( n89801 , n89800 , n47575 );
and ( n89802 , n47662 , n50289 );
or ( n89803 , n89801 , n89802 );
and ( n89804 , n89803 , n32417 );
not ( n89805 , n50008 );
and ( n89806 , n89805 , n47575 );
and ( n89807 , n47662 , n50008 );
or ( n89808 , n89806 , n89807 );
and ( n89809 , n89808 , n32415 );
not ( n89810 , n47331 );
and ( n89811 , n89810 , n47575 );
and ( n89812 , n47607 , n47331 );
or ( n89813 , n89811 , n89812 );
and ( n89814 , n89813 , n32413 );
not ( n89815 , n50067 );
and ( n89816 , n89815 , n47575 );
and ( n89817 , n47607 , n50067 );
or ( n89818 , n89816 , n89817 );
and ( n89819 , n89818 , n32411 );
not ( n89820 , n31728 );
and ( n89821 , n89820 , n47575 );
xor ( n89822 , n47607 , n47622 );
and ( n89823 , n89822 , n31728 );
or ( n89824 , n89821 , n89823 );
and ( n89825 , n89824 , n32253 );
not ( n89826 , n32283 );
and ( n89827 , n89826 , n47575 );
not ( n89828 , n31823 );
xor ( n89829 , n47662 , n47677 );
and ( n89830 , n89828 , n89829 );
xnor ( n89831 , n47712 , n47727 );
and ( n89832 , n89831 , n31823 );
or ( n89833 , n89830 , n89832 );
and ( n89834 , n89833 , n32283 );
or ( n89835 , n89827 , n89834 );
and ( n89836 , n89835 , n32398 );
and ( n89837 , n47712 , n50334 );
or ( n89838 , n89789 , n89794 , n89799 , n89804 , n89809 , n89814 , n89819 , n89825 , n89836 , n89837 );
and ( n89839 , n89838 , n32456 );
and ( n89840 , n37557 , n32489 );
and ( n89841 , n47575 , n50345 );
or ( n89842 , C0 , n89839 , n89840 , n89841 );
buf ( n89843 , n89842 );
buf ( n89844 , n89843 );
buf ( n89845 , n30987 );
buf ( n89846 , n30987 );
buf ( n89847 , n30987 );
not ( n89848 , n43755 );
and ( n89849 , n89848 , n43530 );
xor ( n89850 , n52311 , n52318 );
and ( n89851 , n89850 , n43755 );
or ( n89852 , n89849 , n89851 );
and ( n89853 , n89852 , n43774 );
not ( n89854 , n44663 );
and ( n89855 , n89854 , n44442 );
xor ( n89856 , n52349 , n52356 );
and ( n89857 , n89856 , n44663 );
or ( n89858 , n89855 , n89857 );
and ( n89859 , n89858 , n44682 );
and ( n89860 , n66317 , n44695 );
or ( n89861 , n89853 , n89859 , n89860 );
buf ( n89862 , n89861 );
buf ( n89863 , n89862 );
buf ( n89864 , n31655 );
buf ( n89865 , n31655 );
buf ( n89866 , n31655 );
and ( n89867 , n61336 , n33377 );
not ( n89868 , n48545 );
and ( n89869 , n89868 , n62168 );
and ( n89870 , n72475 , n48545 );
or ( n89871 , n89869 , n89870 );
and ( n89872 , n89871 , n32890 );
not ( n89873 , n48557 );
and ( n89874 , n89873 , n62168 );
and ( n89875 , n72475 , n48557 );
or ( n89876 , n89874 , n89875 );
and ( n89877 , n89876 , n33038 );
and ( n89878 , n62168 , n48571 );
or ( n89879 , n89872 , n89877 , n89878 );
and ( n89880 , n89879 , n33208 );
and ( n89881 , n62168 , n48577 );
or ( n89882 , C0 , n89867 , n89880 , n89881 );
buf ( n89883 , n89882 );
buf ( n89884 , n89883 );
buf ( n89885 , n30987 );
buf ( n89886 , n30987 );
buf ( n89887 , n31655 );
buf ( n89888 , n31655 );
buf ( n89889 , n31655 );
not ( n89890 , n33419 );
and ( n89891 , n89890 , n31565 );
and ( n89892 , n57318 , n33419 );
or ( n89893 , n89891 , n89892 );
and ( n89894 , n89893 , n31529 );
not ( n89895 , n33734 );
and ( n89896 , n89895 , n31565 );
and ( n89897 , n57333 , n33734 );
or ( n89898 , n89896 , n89897 );
and ( n89899 , n89898 , n31527 );
and ( n89900 , n31565 , n33942 );
or ( n89901 , n89894 , n89899 , n89900 );
and ( n89902 , n89901 , n31557 );
and ( n89903 , n35486 , n31643 );
not ( n89904 , n31452 );
and ( n89905 , n89904 , n35486 );
xor ( n89906 , n31565 , n59435 );
and ( n89907 , n89906 , n31452 );
or ( n89908 , n89905 , n89907 );
and ( n89909 , n89908 , n31638 );
and ( n89910 , n35391 , n33973 );
and ( n89911 , n31565 , n33978 );
or ( n89912 , C0 , n89902 , n89903 , n89909 , n89910 , n89911 );
buf ( n89913 , n89912 );
buf ( n89914 , n89913 );
and ( n89915 , n31579 , n31007 );
not ( n89916 , n31077 );
and ( n89917 , n89916 , n34003 );
buf ( n89918 , n89917 );
and ( n89919 , n89918 , n31373 );
not ( n89920 , n31402 );
and ( n89921 , n89920 , n34003 );
buf ( n89922 , n89921 );
and ( n89923 , n89922 , n31408 );
not ( n89924 , n31437 );
and ( n89925 , n89924 , n34003 );
not ( n89926 , n31455 );
and ( n89927 , n89926 , n34046 );
xor ( n89928 , n34003 , n34020 );
and ( n89929 , n89928 , n31455 );
or ( n89930 , n89927 , n89929 );
and ( n89931 , n89930 , n31437 );
or ( n89932 , n89925 , n89931 );
and ( n89933 , n89932 , n31468 );
not ( n89934 , n31497 );
and ( n89935 , n89934 , n34003 );
not ( n89936 , n31454 );
not ( n89937 , n31501 );
and ( n89938 , n89937 , n34046 );
xor ( n89939 , n34047 , n34072 );
and ( n89940 , n89939 , n31501 );
or ( n89941 , n89938 , n89940 );
and ( n89942 , n89936 , n89941 );
and ( n89943 , n89928 , n31454 );
or ( n89944 , n89942 , n89943 );
and ( n89945 , n89944 , n31497 );
or ( n89946 , n89935 , n89945 );
and ( n89947 , n89946 , n31521 );
and ( n89948 , n34003 , n31553 );
or ( n89949 , n89919 , n89923 , n89933 , n89947 , n89948 );
and ( n89950 , n89949 , n31557 );
not ( n89951 , n31452 );
not ( n89952 , n31619 );
and ( n89953 , n89952 , n34103 );
xor ( n89954 , n34104 , n34129 );
and ( n89955 , n89954 , n31619 );
or ( n89956 , n89953 , n89955 );
and ( n89957 , n89951 , n89956 );
and ( n89958 , n34003 , n31452 );
or ( n89959 , n89957 , n89958 );
and ( n89960 , n89959 , n31638 );
buf ( n89961 , n33973 );
and ( n89962 , n34003 , n31650 );
or ( n89963 , C0 , n89915 , n89950 , n89960 , n89961 , n89962 );
buf ( n89964 , n89963 );
buf ( n89965 , n89964 );
buf ( n89966 , n30987 );
buf ( n89967 , n30987 );
buf ( n89968 , n30987 );
buf ( n89969 , n30987 );
not ( n89970 , n43755 );
and ( n89971 , n89970 , n43564 );
xor ( n89972 , n52309 , n52320 );
and ( n89973 , n89972 , n43755 );
or ( n89974 , n89971 , n89973 );
and ( n89975 , n89974 , n43774 );
not ( n89976 , n44663 );
and ( n89977 , n89976 , n44476 );
xor ( n89978 , n52347 , n52358 );
and ( n89979 , n89978 , n44663 );
or ( n89980 , n89977 , n89979 );
and ( n89981 , n89980 , n44682 );
and ( n89982 , n81328 , n44695 );
or ( n89983 , n89975 , n89981 , n89982 );
buf ( n89984 , n89983 );
buf ( n89985 , n89984 );
buf ( n89986 , n31655 );
buf ( n89987 , n31655 );
not ( n89988 , n46356 );
and ( n89989 , n89988 , n31335 );
not ( n89990 , n61975 );
and ( n89991 , n89990 , n31335 );
and ( n89992 , n31339 , n61975 );
or ( n89993 , n89991 , n89992 );
and ( n89994 , n89993 , n46356 );
or ( n89995 , n89989 , n89994 );
and ( n89996 , n89995 , n31649 );
not ( n89997 , n61983 );
not ( n89998 , n61975 );
and ( n89999 , n89998 , n31335 );
and ( n90000 , n47449 , n61975 );
or ( n90001 , n89999 , n90000 );
and ( n90002 , n89997 , n90001 );
and ( n90003 , n47449 , n61983 );
or ( n90004 , n90002 , n90003 );
and ( n90005 , n90004 , n31643 );
not ( n90006 , n31452 );
not ( n90007 , n61983 );
not ( n90008 , n61975 );
and ( n90009 , n90008 , n31335 );
and ( n90010 , n47449 , n61975 );
or ( n90011 , n90009 , n90010 );
and ( n90012 , n90007 , n90011 );
and ( n90013 , n47449 , n61983 );
or ( n90014 , n90012 , n90013 );
and ( n90015 , n90006 , n90014 );
not ( n90016 , n62003 );
not ( n90017 , n62005 );
and ( n90018 , n90017 , n90014 );
and ( n90019 , n47485 , n62005 );
or ( n90020 , n90018 , n90019 );
and ( n90021 , n90016 , n90020 );
and ( n90022 , n47503 , n62003 );
or ( n90023 , n90021 , n90022 );
and ( n90024 , n90023 , n31452 );
or ( n90025 , n90015 , n90024 );
and ( n90026 , n90025 , n31638 );
and ( n90027 , n31335 , n47277 );
or ( n90028 , C0 , n89996 , n90005 , n90026 , n90027 );
buf ( n90029 , n90028 );
buf ( n90030 , n90029 );
buf ( n90031 , n31655 );
buf ( n90032 , n30987 );
buf ( n90033 , n30987 );
xor ( n90034 , n49585 , n60313 );
and ( n90035 , n90034 , n32433 );
not ( n90036 , n47331 );
and ( n90037 , n90036 , n49585 );
and ( n90038 , n75172 , n47331 );
or ( n90039 , n90037 , n90038 );
and ( n90040 , n90039 , n32413 );
and ( n90041 , n49585 , n47402 );
or ( n90042 , n90035 , n90040 , n90041 );
and ( n90043 , n90042 , n32456 );
and ( n90044 , n49585 , n47409 );
or ( n90045 , C0 , n90043 , n90044 );
buf ( n90046 , n90045 );
buf ( n90047 , n90046 );
buf ( n90048 , n31655 );
buf ( n90049 , n31655 );
xor ( n90050 , n33087 , n58390 );
and ( n90051 , n90050 , n33201 );
not ( n90052 , n41576 );
and ( n90053 , n90052 , n33087 );
xor ( n90054 , n58574 , n58591 );
and ( n90055 , n90054 , n41576 );
or ( n90056 , n90053 , n90055 );
and ( n90057 , n90056 , n33189 );
and ( n90058 , n33087 , n41592 );
or ( n90059 , n90051 , n90057 , n90058 );
and ( n90060 , n90059 , n33208 );
and ( n90061 , n33087 , n39805 );
or ( n90062 , C0 , n90060 , n90061 );
buf ( n90063 , n90062 );
buf ( n90064 , n90063 );
buf ( n90065 , n30987 );
buf ( n90066 , n30987 );
buf ( n90067 , n31655 );
not ( n90068 , n50828 );
not ( n90069 , n50834 );
and ( n90070 , n90069 , n40463 );
and ( n90071 , n78185 , n50834 );
or ( n90072 , n90070 , n90071 );
and ( n90073 , n90068 , n90072 );
and ( n90074 , n88735 , n50828 );
or ( n90075 , n90073 , n90074 );
buf ( n90076 , n90075 );
buf ( n90077 , n90076 );
buf ( n90078 , n31655 );
not ( n90079 , n31509 );
and ( n90080 , n90079 , n31550 );
not ( n90081 , n39979 );
and ( n90082 , n90081 , n31509 );
buf ( n90083 , n31135 );
and ( n90084 , n90083 , n39979 );
or ( n90085 , n90082 , n90084 );
and ( n90086 , n90085 , n31538 );
and ( n90087 , n31509 , n40143 );
or ( n90088 , n90080 , n90086 , n90087 );
and ( n90089 , n90088 , n31557 );
and ( n90090 , n31509 , n40154 );
or ( n90091 , C0 , n90089 , n90090 );
buf ( n90092 , n90091 );
buf ( n90093 , n90092 );
not ( n90094 , n40163 );
and ( n90095 , n90094 , n32058 );
not ( n90096 , n45161 );
and ( n90097 , n90096 , n32058 );
and ( n90098 , n32130 , n45161 );
or ( n90099 , n90097 , n90098 );
and ( n90100 , n90099 , n40163 );
or ( n90101 , n90095 , n90100 );
and ( n90102 , n90101 , n32498 );
not ( n90103 , n45170 );
not ( n90104 , n45161 );
and ( n90105 , n90104 , n32058 );
and ( n90106 , n45833 , n45161 );
or ( n90107 , n90105 , n90106 );
and ( n90108 , n90103 , n90107 );
and ( n90109 , n45833 , n45170 );
or ( n90110 , n90108 , n90109 );
and ( n90111 , n90110 , n32473 );
not ( n90112 , n32475 );
not ( n90113 , n45170 );
not ( n90114 , n45161 );
and ( n90115 , n90114 , n32058 );
and ( n90116 , n45833 , n45161 );
or ( n90117 , n90115 , n90116 );
and ( n90118 , n90113 , n90117 );
and ( n90119 , n45833 , n45170 );
or ( n90120 , n90118 , n90119 );
and ( n90121 , n90112 , n90120 );
not ( n90122 , n45196 );
not ( n90123 , n45199 );
and ( n90124 , n90123 , n90120 );
and ( n90125 , n45857 , n45199 );
or ( n90126 , n90124 , n90125 );
and ( n90127 , n90122 , n90126 );
and ( n90128 , n45865 , n45196 );
or ( n90129 , n90127 , n90128 );
and ( n90130 , n90129 , n32475 );
or ( n90131 , n90121 , n90130 );
and ( n90132 , n90131 , n32486 );
and ( n90133 , n32058 , n41278 );
or ( n90134 , C0 , n90102 , n90111 , n90132 , n90133 );
buf ( n90135 , n90134 );
buf ( n90136 , n90135 );
buf ( n90137 , n30987 );
buf ( n90138 , n30987 );
not ( n90139 , n46356 );
and ( n90140 , n90139 , n31284 );
not ( n90141 , n53353 );
and ( n90142 , n90141 , n31284 );
and ( n90143 , n31306 , n53353 );
or ( n90144 , n90142 , n90143 );
and ( n90145 , n90144 , n46356 );
or ( n90146 , n90140 , n90145 );
and ( n90147 , n90146 , n31649 );
not ( n90148 , n53361 );
not ( n90149 , n53353 );
and ( n90150 , n90149 , n31284 );
and ( n90151 , n58061 , n53353 );
or ( n90152 , n90150 , n90151 );
and ( n90153 , n90148 , n90152 );
and ( n90154 , n58061 , n53361 );
or ( n90155 , n90153 , n90154 );
and ( n90156 , n90155 , n31643 );
not ( n90157 , n31452 );
not ( n90158 , n53361 );
not ( n90159 , n53353 );
and ( n90160 , n90159 , n31284 );
and ( n90161 , n58061 , n53353 );
or ( n90162 , n90160 , n90161 );
and ( n90163 , n90158 , n90162 );
and ( n90164 , n58061 , n53361 );
or ( n90165 , n90163 , n90164 );
and ( n90166 , n90157 , n90165 );
not ( n90167 , n53381 );
not ( n90168 , n53383 );
and ( n90169 , n90168 , n90165 );
and ( n90170 , n58085 , n53383 );
or ( n90171 , n90169 , n90170 );
and ( n90172 , n90167 , n90171 );
and ( n90173 , n58093 , n53381 );
or ( n90174 , n90172 , n90173 );
and ( n90175 , n90174 , n31452 );
or ( n90176 , n90166 , n90175 );
and ( n90177 , n90176 , n31638 );
and ( n90178 , n31284 , n47277 );
or ( n90179 , C0 , n90147 , n90156 , n90177 , n90178 );
buf ( n90180 , n90179 );
buf ( n90181 , n90180 );
buf ( n90182 , n31655 );
buf ( n90183 , n30987 );
and ( n90184 , n71895 , n32494 );
not ( n90185 , n46083 );
and ( n90186 , n90185 , n71601 );
buf ( n90187 , n90186 );
and ( n90188 , n90187 , n32421 );
not ( n90189 , n46326 );
and ( n90190 , n90189 , n71601 );
and ( n90191 , n71901 , n46326 );
or ( n90192 , n90190 , n90191 );
and ( n90193 , n90192 , n32417 );
and ( n90194 , n71601 , n46340 );
or ( n90195 , n90188 , n90193 , n90194 );
and ( n90196 , n90195 , n32456 );
and ( n90197 , n71601 , n46349 );
or ( n90198 , C0 , n90184 , n90196 , n90197 );
buf ( n90199 , n90198 );
buf ( n90200 , n90199 );
buf ( n90201 , n31655 );
buf ( n90202 , n31655 );
not ( n90203 , n46356 );
and ( n90204 , n90203 , n31352 );
not ( n90205 , n52734 );
and ( n90206 , n90205 , n31352 );
and ( n90207 , n31372 , n52734 );
or ( n90208 , n90206 , n90207 );
and ( n90209 , n90208 , n46356 );
or ( n90210 , n90204 , n90209 );
and ( n90211 , n90210 , n31649 );
not ( n90212 , n52742 );
not ( n90213 , n52734 );
and ( n90214 , n90213 , n31352 );
and ( n90215 , n47849 , n52734 );
or ( n90216 , n90214 , n90215 );
and ( n90217 , n90212 , n90216 );
and ( n90218 , n47849 , n52742 );
or ( n90219 , n90217 , n90218 );
and ( n90220 , n90219 , n31643 );
not ( n90221 , n31452 );
not ( n90222 , n52742 );
not ( n90223 , n52734 );
and ( n90224 , n90223 , n31352 );
and ( n90225 , n47849 , n52734 );
or ( n90226 , n90224 , n90225 );
and ( n90227 , n90222 , n90226 );
and ( n90228 , n47849 , n52742 );
or ( n90229 , n90227 , n90228 );
and ( n90230 , n90221 , n90229 );
not ( n90231 , n52762 );
not ( n90232 , n52764 );
and ( n90233 , n90232 , n90229 );
and ( n90234 , n47877 , n52764 );
or ( n90235 , n90233 , n90234 );
and ( n90236 , n90231 , n90235 );
and ( n90237 , n47887 , n52762 );
or ( n90238 , n90236 , n90237 );
and ( n90239 , n90238 , n31452 );
or ( n90240 , n90230 , n90239 );
and ( n90241 , n90240 , n31638 );
and ( n90242 , n31352 , n47277 );
or ( n90243 , C0 , n90211 , n90220 , n90241 , n90242 );
buf ( n90244 , n90243 );
buf ( n90245 , n90244 );
buf ( n90246 , n30987 );
not ( n90247 , n46083 );
and ( n90248 , n90247 , n35530 );
buf ( n90249 , n90248 );
and ( n90250 , n90249 , n32421 );
not ( n90251 , n46326 );
and ( n90252 , n90251 , n35530 );
buf ( n90253 , n90252 );
and ( n90254 , n90253 , n32417 );
and ( n90255 , n35530 , n46340 );
or ( n90256 , n90250 , n90254 , n90255 );
and ( n90257 , n90256 , n32456 );
and ( n90258 , n35530 , n46349 );
or ( n90259 , C0 , C0 , n90257 , n90258 );
buf ( n90260 , n90259 );
buf ( n90261 , n90260 );
buf ( n90262 , n31655 );
buf ( n90263 , n30987 );
buf ( n90264 , n84862 );
buf ( n90265 , n31655 );
not ( n90266 , n48765 );
and ( n90267 , n90266 , n33225 );
and ( n90268 , n64831 , n48765 );
or ( n90269 , n90267 , n90268 );
and ( n90270 , n90269 , n33180 );
not ( n90271 , n49054 );
and ( n90272 , n90271 , n33225 );
and ( n90273 , n64842 , n49054 );
or ( n90274 , n90272 , n90273 );
and ( n90275 , n90274 , n33178 );
and ( n90276 , n33225 , n49774 );
or ( n90277 , n90270 , n90275 , n90276 );
and ( n90278 , n90277 , n33208 );
and ( n90279 , n33301 , n33375 );
not ( n90280 , n32968 );
and ( n90281 , n90280 , n33301 );
xor ( n90282 , n33225 , n53904 );
and ( n90283 , n90282 , n32968 );
or ( n90284 , n90281 , n90283 );
and ( n90285 , n90284 , n33370 );
and ( n90286 , n32988 , n35056 );
and ( n90287 , n33225 , n49794 );
or ( n90288 , C0 , n90278 , n90279 , n90285 , n90286 , n90287 );
buf ( n90289 , n90288 );
buf ( n90290 , n90289 );
buf ( n90291 , n30987 );
buf ( n90292 , n31655 );
and ( n90293 , n46025 , n32500 );
not ( n90294 , n35211 );
and ( n90295 , n90294 , n37547 );
buf ( n90296 , n90295 );
and ( n90297 , n90296 , n32421 );
not ( n90298 , n35245 );
and ( n90299 , n90298 , n37547 );
buf ( n90300 , n90299 );
and ( n90301 , n90300 , n32419 );
not ( n90302 , n35278 );
and ( n90303 , n90302 , n37547 );
not ( n90304 , n35295 );
and ( n90305 , n90304 , n49577 );
xor ( n90306 , n37547 , n49542 );
and ( n90307 , n90306 , n35295 );
or ( n90308 , n90305 , n90307 );
and ( n90309 , n90308 , n35278 );
or ( n90310 , n90303 , n90309 );
and ( n90311 , n90310 , n32417 );
not ( n90312 , n35331 );
and ( n90313 , n90312 , n37547 );
not ( n90314 , n35294 );
not ( n90315 , n45995 );
and ( n90316 , n90315 , n49577 );
xor ( n90317 , n49578 , n49628 );
and ( n90318 , n90317 , n45995 );
or ( n90319 , n90316 , n90318 );
and ( n90320 , n90314 , n90319 );
and ( n90321 , n90306 , n35294 );
or ( n90322 , n90320 , n90321 );
and ( n90323 , n90322 , n35331 );
or ( n90324 , n90313 , n90323 );
and ( n90325 , n90324 , n32415 );
and ( n90326 , n37547 , n35354 );
or ( n90327 , n90297 , n90301 , n90311 , n90325 , n90326 );
and ( n90328 , n90327 , n32456 );
not ( n90329 , n32475 );
not ( n90330 , n46060 );
and ( n90331 , n90330 , n49667 );
xor ( n90332 , n49668 , n49722 );
and ( n90333 , n90332 , n46060 );
or ( n90334 , n90331 , n90333 );
and ( n90335 , n90329 , n90334 );
and ( n90336 , n37547 , n32475 );
or ( n90337 , n90335 , n90336 );
and ( n90338 , n90337 , n32486 );
and ( n90339 , n37547 , n35367 );
or ( n90340 , C0 , n90293 , n90328 , n90338 , C0 , n90339 );
buf ( n90341 , n90340 );
buf ( n90342 , n90341 );
or ( n90343 , n44688 , n44690 );
and ( n90344 , n52719 , n90343 );
buf ( n90345 , n44686 );
and ( n90346 , n32968 , n62377 );
or ( n90347 , n90344 , n90345 , n90346 );
buf ( n90348 , n90347 );
buf ( n90349 , n90348 );
buf ( n90350 , n30987 );
buf ( n90351 , n31655 );
buf ( n90352 , n30987 );
buf ( n90353 , n31655 );
buf ( n90354 , n31655 );
buf ( n90355 , n30987 );
not ( n90356 , n32953 );
and ( n90357 , n90356 , n86492 );
not ( n90358 , n39572 );
and ( n90359 , n90358 , n39373 );
xor ( n90360 , n39576 , n39374 );
and ( n90361 , n90360 , n39572 );
or ( n90362 , n90359 , n90361 );
and ( n90363 , n90362 , n32953 );
or ( n90364 , n90357 , n90363 );
and ( n90365 , n90364 , n33038 );
not ( n90366 , n39586 );
and ( n90367 , n90366 , n86492 );
and ( n90368 , n86498 , n39586 );
or ( n90369 , n90367 , n90368 );
and ( n90370 , n90369 , n33172 );
and ( n90371 , n86492 , n39795 );
or ( n90372 , n90365 , n90370 , n90371 );
and ( n90373 , n90372 , n33208 );
and ( n90374 , n86492 , n39805 );
or ( n90375 , C0 , n90373 , n90374 );
buf ( n90376 , n90375 );
buf ( n90377 , n90376 );
buf ( n90378 , n30987 );
buf ( n90379 , n31655 );
buf ( n90380 , n30987 );
not ( n90381 , n48765 );
and ( n90382 , n90381 , n33238 );
xor ( n90383 , n48904 , n48921 );
xor ( n90384 , n90383 , n48985 );
and ( n90385 , n90384 , n48765 );
or ( n90386 , n90382 , n90385 );
and ( n90387 , n90386 , n33180 );
not ( n90388 , n49054 );
and ( n90389 , n90388 , n33238 );
not ( n90390 , n48845 );
xor ( n90391 , n49087 , n48921 );
xor ( n90392 , n90391 , n49099 );
and ( n90393 , n90390 , n90392 );
xor ( n90394 , n49204 , n49206 );
xor ( n90395 , n90394 , n49225 );
and ( n90396 , n90395 , n48845 );
or ( n90397 , n90393 , n90396 );
and ( n90398 , n90397 , n49054 );
or ( n90399 , n90389 , n90398 );
and ( n90400 , n90399 , n33178 );
and ( n90401 , n33238 , n49774 );
or ( n90402 , n90387 , n90400 , n90401 );
and ( n90403 , n90402 , n33208 );
and ( n90404 , n33327 , n33375 );
not ( n90405 , n32968 );
and ( n90406 , n90405 , n33327 );
xor ( n90407 , n33238 , n33239 );
and ( n90408 , n90407 , n32968 );
or ( n90409 , n90406 , n90408 );
and ( n90410 , n90409 , n33370 );
and ( n90411 , n33001 , n35056 );
and ( n90412 , n33238 , n49794 );
or ( n90413 , C0 , n90403 , n90404 , n90410 , n90411 , n90412 );
buf ( n90414 , n90413 );
buf ( n90415 , n90414 );
buf ( n90416 , n31655 );
buf ( n90417 , n30987 );
buf ( n90418 , n31655 );
not ( n90419 , n50828 );
not ( n90420 , n50834 );
and ( n90421 , n90420 , n40285 );
and ( n90422 , n41535 , n50834 );
or ( n90423 , n90421 , n90422 );
and ( n90424 , n90419 , n90423 );
and ( n90425 , n73105 , n50828 );
or ( n90426 , n90424 , n90425 );
buf ( n90427 , n90426 );
buf ( n90428 , n90427 );
and ( n90429 , n42403 , n48455 );
not ( n90430 , n48457 );
and ( n90431 , n90430 , n42376 );
and ( n90432 , n42403 , n48457 );
or ( n90433 , n90431 , n90432 );
and ( n90434 , n90433 , n31373 );
not ( n90435 , n44807 );
and ( n90436 , n90435 , n42376 );
and ( n90437 , n42403 , n44807 );
or ( n90438 , n90436 , n90437 );
and ( n90439 , n90438 , n31408 );
not ( n90440 , n48468 );
and ( n90441 , n90440 , n42376 );
and ( n90442 , n42403 , n48468 );
or ( n90443 , n90441 , n90442 );
and ( n90444 , n90443 , n31468 );
not ( n90445 , n44817 );
and ( n90446 , n90445 , n42376 );
and ( n90447 , n42403 , n44817 );
or ( n90448 , n90446 , n90447 );
and ( n90449 , n90448 , n31521 );
not ( n90450 , n39979 );
and ( n90451 , n90450 , n42376 );
and ( n90452 , n42384 , n39979 );
or ( n90453 , n90451 , n90452 );
and ( n90454 , n90453 , n31538 );
not ( n90455 , n45059 );
and ( n90456 , n90455 , n42376 );
and ( n90457 , n42384 , n45059 );
or ( n90458 , n90456 , n90457 );
and ( n90459 , n90458 , n31536 );
not ( n90460 , n33419 );
and ( n90461 , n90460 , n42376 );
and ( n90462 , n42392 , n33419 );
or ( n90463 , n90461 , n90462 );
and ( n90464 , n90463 , n31529 );
not ( n90465 , n33734 );
and ( n90466 , n90465 , n42376 );
and ( n90467 , n42427 , n33734 );
or ( n90468 , n90466 , n90467 );
and ( n90469 , n90468 , n31527 );
and ( n90470 , n42417 , n48513 );
or ( n90471 , n90429 , n90434 , n90439 , n90444 , n90449 , n90454 , n90459 , n90464 , n90469 , n90470 );
and ( n90472 , n90471 , n31557 );
and ( n90473 , n35392 , n33973 );
and ( n90474 , n42376 , n48524 );
or ( n90475 , C0 , n90472 , n90473 , n90474 );
buf ( n90476 , n90475 );
buf ( n90477 , n90476 );
buf ( n90478 , n31655 );
buf ( n90479 , n30987 );
not ( n90480 , n38443 );
and ( n90481 , n90480 , n38320 );
xor ( n90482 , n53463 , n53506 );
and ( n90483 , n90482 , n38443 );
or ( n90484 , n90481 , n90483 );
and ( n90485 , n90484 , n38450 );
not ( n90486 , n39339 );
and ( n90487 , n90486 , n39220 );
xor ( n90488 , n53519 , n53562 );
and ( n90489 , n90488 , n39339 );
or ( n90490 , n90487 , n90489 );
and ( n90491 , n90490 , n39346 );
and ( n90492 , n40221 , n39359 );
or ( n90493 , n90485 , n90491 , n90492 );
buf ( n90494 , n90493 );
buf ( n90495 , n90494 );
buf ( n90496 , n31655 );
buf ( n90497 , n30987 );
and ( n90498 , n32973 , n58397 );
xor ( n90499 , n33071 , n90498 );
and ( n90500 , n90499 , n33201 );
not ( n90501 , n41576 );
and ( n90502 , n90501 , n33071 );
buf ( n90503 , n90502 );
and ( n90504 , n90503 , n33189 );
and ( n90505 , n33071 , n41592 );
or ( n90506 , n90500 , n90504 , n90505 );
and ( n90507 , n90506 , n33208 );
and ( n90508 , n33071 , n39805 );
or ( n90509 , C0 , n90507 , n90508 );
buf ( n90510 , n90509 );
buf ( n90511 , n90510 );
buf ( n90512 , n30987 );
buf ( n90513 , n31655 );
not ( n90514 , n50828 );
not ( n90515 , n50834 );
and ( n90516 , n90515 , n40357 );
and ( n90517 , n73129 , n50834 );
or ( n90518 , n90516 , n90517 );
and ( n90519 , n90514 , n90518 );
and ( n90520 , n63218 , n50828 );
or ( n90521 , n90519 , n90520 );
buf ( n90522 , n90521 );
buf ( n90523 , n90522 );
buf ( n90524 , n31655 );
not ( n90525 , n46356 );
and ( n90526 , n90525 , n31208 );
not ( n90527 , n47831 );
and ( n90528 , n90527 , n31208 );
and ( n90529 , n31238 , n47831 );
or ( n90530 , n90528 , n90529 );
and ( n90531 , n90530 , n46356 );
or ( n90532 , n90526 , n90531 );
and ( n90533 , n90532 , n31649 );
not ( n90534 , n47839 );
not ( n90535 , n47831 );
and ( n90536 , n90535 , n31208 );
and ( n90537 , n49901 , n47831 );
or ( n90538 , n90536 , n90537 );
and ( n90539 , n90534 , n90538 );
and ( n90540 , n49901 , n47839 );
or ( n90541 , n90539 , n90540 );
and ( n90542 , n90541 , n31643 );
not ( n90543 , n31452 );
not ( n90544 , n47839 );
not ( n90545 , n47831 );
and ( n90546 , n90545 , n31208 );
and ( n90547 , n49901 , n47831 );
or ( n90548 , n90546 , n90547 );
and ( n90549 , n90544 , n90548 );
and ( n90550 , n49901 , n47839 );
or ( n90551 , n90549 , n90550 );
and ( n90552 , n90543 , n90551 );
not ( n90553 , n47866 );
not ( n90554 , n47868 );
and ( n90555 , n90554 , n90551 );
and ( n90556 , n49925 , n47868 );
or ( n90557 , n90555 , n90556 );
and ( n90558 , n90553 , n90557 );
and ( n90559 , n49933 , n47866 );
or ( n90560 , n90558 , n90559 );
and ( n90561 , n90560 , n31452 );
or ( n90562 , n90552 , n90561 );
and ( n90563 , n90562 , n31638 );
and ( n90564 , n31208 , n47277 );
or ( n90565 , C0 , n90533 , n90542 , n90563 , n90564 );
buf ( n90566 , n90565 );
buf ( n90567 , n90566 );
buf ( n90568 , n30987 );
not ( n90569 , n35278 );
and ( n90570 , n90569 , n69391 );
and ( n90571 , n69399 , n35278 );
or ( n90572 , n90570 , n90571 );
and ( n90573 , n90572 , n32417 );
not ( n90574 , n47912 );
and ( n90575 , n90574 , n69391 );
and ( n90576 , n83919 , n47912 );
or ( n90577 , n90575 , n90576 );
and ( n90578 , n90577 , n32415 );
and ( n90579 , n69391 , n48133 );
or ( n90580 , n90573 , n90578 , n90579 );
and ( n90581 , n90580 , n32456 );
and ( n90582 , n69391 , n47409 );
or ( n90583 , C0 , n90581 , n90582 );
buf ( n90584 , n90583 );
buf ( n90585 , n90584 );
buf ( n90586 , n31655 );
xor ( n90587 , n54146 , n78380 );
and ( n90588 , n90587 , n33199 );
not ( n90589 , n48648 );
and ( n90590 , n90589 , n54146 );
and ( n90591 , n34431 , n48648 );
or ( n90592 , n90590 , n90591 );
and ( n90593 , n90592 , n32924 );
not ( n90594 , n48660 );
and ( n90595 , n90594 , n54146 );
and ( n90596 , n64043 , n48660 );
or ( n90597 , n90595 , n90596 );
and ( n90598 , n90597 , n33172 );
not ( n90599 , n48730 );
and ( n90600 , n90599 , n54146 );
xor ( n90601 , n58574 , n58591 );
and ( n90602 , n90601 , n48730 );
or ( n90603 , n90600 , n90602 );
and ( n90604 , n90603 , n33187 );
and ( n90605 , n54146 , n54713 );
or ( n90606 , n90588 , n90593 , n90598 , n90604 , n90605 );
and ( n90607 , n90606 , n33208 );
and ( n90608 , n54146 , n39805 );
or ( n90609 , C0 , n90607 , n90608 );
buf ( n90610 , n90609 );
buf ( n90611 , n90610 );
buf ( n90612 , n30987 );
buf ( n90613 , n31655 );
buf ( n90614 , n30987 );
buf ( n90615 , n31655 );
not ( n90616 , n41532 );
and ( n90617 , n90616 , n34365 );
and ( n90618 , n78185 , n41532 );
or ( n90619 , n90617 , n90618 );
buf ( n90620 , n90619 );
buf ( n90621 , n90620 );
buf ( n90622 , n31655 );
and ( n90623 , n84892 , n31645 );
not ( n90624 , n45274 );
and ( n90625 , n90624 , n74194 );
not ( n90626 , n41809 );
and ( n90627 , n90626 , n41727 );
xor ( n90628 , n53295 , n53296 );
and ( n90629 , n90628 , n41809 );
or ( n90630 , n90627 , n90629 );
and ( n90631 , n90630 , n45274 );
or ( n90632 , n90625 , n90631 );
and ( n90633 , n90632 , n31373 );
not ( n90634 , n45280 );
and ( n90635 , n90634 , n74194 );
and ( n90636 , n90630 , n45280 );
or ( n90637 , n90635 , n90636 );
and ( n90638 , n90637 , n31468 );
and ( n90639 , n74194 , n45802 );
or ( n90640 , n90633 , n90638 , n90639 );
and ( n90641 , n90640 , n31557 );
and ( n90642 , n74194 , n45808 );
or ( n90643 , C0 , n90623 , n90641 , n90642 );
buf ( n90644 , n90643 );
buf ( n90645 , n90644 );
not ( n90646 , n40163 );
and ( n90647 , n90646 , n31867 );
not ( n90648 , n53227 );
and ( n90649 , n90648 , n31867 );
and ( n90650 , n32218 , n53227 );
or ( n90651 , n90649 , n90650 );
and ( n90652 , n90651 , n40163 );
or ( n90653 , n90647 , n90652 );
and ( n90654 , n90653 , n32498 );
not ( n90655 , n53235 );
not ( n90656 , n53227 );
and ( n90657 , n90656 , n31867 );
and ( n90658 , n42255 , n53227 );
or ( n90659 , n90657 , n90658 );
and ( n90660 , n90655 , n90659 );
and ( n90661 , n42255 , n53235 );
or ( n90662 , n90660 , n90661 );
and ( n90663 , n90662 , n32473 );
not ( n90664 , n32475 );
not ( n90665 , n53235 );
not ( n90666 , n53227 );
and ( n90667 , n90666 , n31867 );
and ( n90668 , n42255 , n53227 );
or ( n90669 , n90667 , n90668 );
and ( n90670 , n90665 , n90669 );
and ( n90671 , n42255 , n53235 );
or ( n90672 , n90670 , n90671 );
and ( n90673 , n90664 , n90672 );
not ( n90674 , n53260 );
not ( n90675 , n53262 );
and ( n90676 , n90675 , n90672 );
and ( n90677 , n42283 , n53262 );
or ( n90678 , n90676 , n90677 );
and ( n90679 , n90674 , n90678 );
and ( n90680 , n42291 , n53260 );
or ( n90681 , n90679 , n90680 );
and ( n90682 , n90681 , n32475 );
or ( n90683 , n90673 , n90682 );
and ( n90684 , n90683 , n32486 );
and ( n90685 , n31867 , n41278 );
or ( n90686 , C0 , n90654 , n90663 , n90684 , n90685 );
buf ( n90687 , n90686 );
buf ( n90688 , n90687 );
buf ( n90689 , n30987 );
buf ( n90690 , n30987 );
buf ( n90691 , n30987 );
not ( n90692 , n34150 );
and ( n90693 , n90692 , n32854 );
not ( n90694 , n56239 );
and ( n90695 , n90694 , n32854 );
and ( n90696 , n32856 , n56239 );
or ( n90697 , n90695 , n90696 );
and ( n90698 , n90697 , n34150 );
or ( n90699 , n90693 , n90698 );
and ( n90700 , n90699 , n33381 );
not ( n90701 , n56247 );
not ( n90702 , n56239 );
and ( n90703 , n90702 , n32854 );
and ( n90704 , n48160 , n56239 );
or ( n90705 , n90703 , n90704 );
and ( n90706 , n90701 , n90705 );
and ( n90707 , n48160 , n56247 );
or ( n90708 , n90706 , n90707 );
and ( n90709 , n90708 , n33375 );
not ( n90710 , n32968 );
not ( n90711 , n56247 );
not ( n90712 , n56239 );
and ( n90713 , n90712 , n32854 );
and ( n90714 , n48160 , n56239 );
or ( n90715 , n90713 , n90714 );
and ( n90716 , n90711 , n90715 );
and ( n90717 , n48160 , n56247 );
or ( n90718 , n90716 , n90717 );
and ( n90719 , n90710 , n90718 );
not ( n90720 , n56267 );
not ( n90721 , n56269 );
and ( n90722 , n90721 , n90718 );
and ( n90723 , n48186 , n56269 );
or ( n90724 , n90722 , n90723 );
and ( n90725 , n90720 , n90724 );
and ( n90726 , n48196 , n56267 );
or ( n90727 , n90725 , n90726 );
and ( n90728 , n90727 , n32968 );
or ( n90729 , n90719 , n90728 );
and ( n90730 , n90729 , n33370 );
and ( n90731 , n32854 , n35062 );
or ( n90732 , C0 , n90700 , n90709 , n90730 , n90731 );
buf ( n90733 , n90732 );
buf ( n90734 , n90733 );
not ( n90735 , n34150 );
and ( n90736 , n90735 , n32679 );
not ( n90737 , n56192 );
and ( n90738 , n90737 , n32679 );
and ( n90739 , n32689 , n56192 );
or ( n90740 , n90738 , n90739 );
and ( n90741 , n90740 , n34150 );
or ( n90742 , n90736 , n90741 );
and ( n90743 , n90742 , n33381 );
not ( n90744 , n56200 );
not ( n90745 , n56192 );
and ( n90746 , n90745 , n32679 );
and ( n90747 , n50682 , n56192 );
or ( n90748 , n90746 , n90747 );
and ( n90749 , n90744 , n90748 );
and ( n90750 , n50682 , n56200 );
or ( n90751 , n90749 , n90750 );
and ( n90752 , n90751 , n33375 );
not ( n90753 , n32968 );
not ( n90754 , n56200 );
not ( n90755 , n56192 );
and ( n90756 , n90755 , n32679 );
and ( n90757 , n50682 , n56192 );
or ( n90758 , n90756 , n90757 );
and ( n90759 , n90754 , n90758 );
and ( n90760 , n50682 , n56200 );
or ( n90761 , n90759 , n90760 );
and ( n90762 , n90753 , n90761 );
not ( n90763 , n56220 );
not ( n90764 , n56222 );
and ( n90765 , n90764 , n90761 );
and ( n90766 , n50706 , n56222 );
or ( n90767 , n90765 , n90766 );
and ( n90768 , n90763 , n90767 );
and ( n90769 , n50714 , n56220 );
or ( n90770 , n90768 , n90769 );
and ( n90771 , n90770 , n32968 );
or ( n90772 , n90762 , n90771 );
and ( n90773 , n90772 , n33370 );
and ( n90774 , n32679 , n35062 );
or ( n90775 , C0 , n90743 , n90752 , n90773 , n90774 );
buf ( n90776 , n90775 );
buf ( n90777 , n90776 );
buf ( n90778 , n31655 );
buf ( n90779 , n31655 );
buf ( n90780 , n30987 );
and ( n90781 , n81347 , n48639 );
not ( n90782 , n48642 );
and ( n90783 , n90782 , n56473 );
and ( n90784 , n81347 , n48642 );
or ( n90785 , n90783 , n90784 );
and ( n90786 , n90785 , n32890 );
not ( n90787 , n48648 );
and ( n90788 , n90787 , n56473 );
and ( n90789 , n81347 , n48648 );
or ( n90790 , n90788 , n90789 );
and ( n90791 , n90790 , n32924 );
not ( n90792 , n48654 );
and ( n90793 , n90792 , n56473 );
and ( n90794 , n81347 , n48654 );
or ( n90795 , n90793 , n90794 );
and ( n90796 , n90795 , n33038 );
not ( n90797 , n48660 );
and ( n90798 , n90797 , n56473 );
and ( n90799 , n81347 , n48660 );
or ( n90800 , n90798 , n90799 );
and ( n90801 , n90800 , n33172 );
not ( n90802 , n41576 );
and ( n90803 , n90802 , n56473 );
and ( n90804 , n81337 , n41576 );
or ( n90805 , n90803 , n90804 );
and ( n90806 , n90805 , n33189 );
not ( n90807 , n48730 );
and ( n90808 , n90807 , n56473 );
and ( n90809 , n81337 , n48730 );
or ( n90810 , n90808 , n90809 );
and ( n90811 , n90810 , n33187 );
not ( n90812 , n48765 );
and ( n90813 , n90812 , n56473 );
and ( n90814 , n81339 , n48765 );
or ( n90815 , n90813 , n90814 );
and ( n90816 , n90815 , n33180 );
not ( n90817 , n49054 );
and ( n90818 , n90817 , n56473 );
and ( n90819 , n81356 , n49054 );
or ( n90820 , n90818 , n90819 );
and ( n90821 , n90820 , n33178 );
and ( n90822 , n81352 , n49275 );
or ( n90823 , n90781 , n90786 , n90791 , n90796 , n90801 , n90806 , n90811 , n90816 , n90821 , n90822 );
and ( n90824 , n90823 , n33208 );
and ( n90825 , n32600 , n35056 );
and ( n90826 , n56473 , n49286 );
or ( n90827 , C0 , n90824 , n90825 , n90826 );
buf ( n90828 , n90827 );
buf ( n90829 , n90828 );
buf ( n90830 , n30987 );
buf ( n90831 , n31655 );
buf ( n90832 , n31655 );
buf ( n90833 , n31655 );
not ( n90834 , n46356 );
and ( n90835 , n90834 , n31266 );
not ( n90836 , n47423 );
and ( n90837 , n90836 , n31266 );
and ( n90838 , n31272 , n47423 );
or ( n90839 , n90837 , n90838 );
and ( n90840 , n90839 , n46356 );
or ( n90841 , n90835 , n90840 );
and ( n90842 , n90841 , n31649 );
not ( n90843 , n47431 );
not ( n90844 , n47423 );
and ( n90845 , n90844 , n31266 );
and ( n90846 , n49443 , n47423 );
or ( n90847 , n90845 , n90846 );
and ( n90848 , n90843 , n90847 );
and ( n90849 , n49443 , n47431 );
or ( n90850 , n90848 , n90849 );
and ( n90851 , n90850 , n31643 );
not ( n90852 , n31452 );
not ( n90853 , n47431 );
not ( n90854 , n47423 );
and ( n90855 , n90854 , n31266 );
and ( n90856 , n49443 , n47423 );
or ( n90857 , n90855 , n90856 );
and ( n90858 , n90853 , n90857 );
and ( n90859 , n49443 , n47431 );
or ( n90860 , n90858 , n90859 );
and ( n90861 , n90852 , n90860 );
not ( n90862 , n47466 );
not ( n90863 , n47468 );
and ( n90864 , n90863 , n90860 );
and ( n90865 , n49469 , n47468 );
or ( n90866 , n90864 , n90865 );
and ( n90867 , n90862 , n90866 );
and ( n90868 , n49477 , n47466 );
or ( n90869 , n90867 , n90868 );
and ( n90870 , n90869 , n31452 );
or ( n90871 , n90861 , n90870 );
and ( n90872 , n90871 , n31638 );
and ( n90873 , n31266 , n47277 );
or ( n90874 , C0 , n90842 , n90851 , n90872 , n90873 );
buf ( n90875 , n90874 );
buf ( n90876 , n90875 );
not ( n90877 , n35542 );
and ( n90878 , n90877 , n41840 );
and ( n90879 , n85624 , n35542 );
or ( n90880 , n90878 , n90879 );
buf ( n90881 , n90880 );
buf ( n90882 , n90881 );
buf ( n90883 , n30987 );
xor ( n90884 , n49597 , n60307 );
and ( n90885 , n90884 , n32433 );
not ( n90886 , n47331 );
and ( n90887 , n90886 , n49597 );
and ( n90888 , n73274 , n47331 );
or ( n90889 , n90887 , n90888 );
and ( n90890 , n90889 , n32413 );
and ( n90891 , n49597 , n47402 );
or ( n90892 , n90885 , n90890 , n90891 );
and ( n90893 , n90892 , n32456 );
and ( n90894 , n49597 , n47409 );
or ( n90895 , C0 , n90893 , n90894 );
buf ( n90896 , n90895 );
buf ( n90897 , n90896 );
buf ( n90898 , n31655 );
and ( n90899 , n49081 , n48639 );
not ( n90900 , n48642 );
and ( n90901 , n90900 , n48605 );
and ( n90902 , n49081 , n48642 );
or ( n90903 , n90901 , n90902 );
and ( n90904 , n90903 , n32890 );
not ( n90905 , n48648 );
and ( n90906 , n90905 , n48605 );
and ( n90907 , n49081 , n48648 );
or ( n90908 , n90906 , n90907 );
and ( n90909 , n90908 , n32924 );
not ( n90910 , n48654 );
and ( n90911 , n90910 , n48605 );
and ( n90912 , n49081 , n48654 );
or ( n90913 , n90911 , n90912 );
and ( n90914 , n90913 , n33038 );
not ( n90915 , n48660 );
and ( n90916 , n90915 , n48605 );
and ( n90917 , n49081 , n48660 );
or ( n90918 , n90916 , n90917 );
and ( n90919 , n90918 , n33172 );
not ( n90920 , n41576 );
and ( n90921 , n90920 , n48605 );
and ( n90922 , n48847 , n41576 );
or ( n90923 , n90921 , n90922 );
and ( n90924 , n90923 , n33189 );
not ( n90925 , n48730 );
and ( n90926 , n90925 , n48605 );
and ( n90927 , n48847 , n48730 );
or ( n90928 , n90926 , n90927 );
and ( n90929 , n90928 , n33187 );
not ( n90930 , n48765 );
and ( n90931 , n90930 , n48605 );
and ( n90932 , n66903 , n48765 );
or ( n90933 , n90931 , n90932 );
and ( n90934 , n90933 , n33180 );
not ( n90935 , n49054 );
and ( n90936 , n90935 , n48605 );
and ( n90937 , n66916 , n49054 );
or ( n90938 , n90936 , n90937 );
and ( n90939 , n90938 , n33178 );
and ( n90940 , n49192 , n49275 );
or ( n90941 , n90899 , n90904 , n90909 , n90914 , n90919 , n90924 , n90929 , n90934 , n90939 , n90940 );
and ( n90942 , n90941 , n33208 );
and ( n90943 , n32998 , n35056 );
and ( n90944 , n48605 , n49286 );
or ( n90945 , C0 , n90942 , n90943 , n90944 );
buf ( n90946 , n90945 );
buf ( n90947 , n90946 );
buf ( n90948 , n30987 );
buf ( n90949 , n30987 );
buf ( n90950 , n31655 );
buf ( n90951 , n31655 );
not ( n90952 , n46356 );
and ( n90953 , n90952 , n31168 );
not ( n90954 , n61975 );
and ( n90955 , n90954 , n31168 );
and ( n90956 , n31172 , n61975 );
or ( n90957 , n90955 , n90956 );
and ( n90958 , n90957 , n46356 );
or ( n90959 , n90953 , n90958 );
and ( n90960 , n90959 , n31649 );
not ( n90961 , n61983 );
not ( n90962 , n61975 );
and ( n90963 , n90962 , n31168 );
and ( n90964 , n46495 , n61975 );
or ( n90965 , n90963 , n90964 );
and ( n90966 , n90961 , n90965 );
and ( n90967 , n46495 , n61983 );
or ( n90968 , n90966 , n90967 );
and ( n90969 , n90968 , n31643 );
not ( n90970 , n31452 );
not ( n90971 , n61983 );
not ( n90972 , n61975 );
and ( n90973 , n90972 , n31168 );
and ( n90974 , n46495 , n61975 );
or ( n90975 , n90973 , n90974 );
and ( n90976 , n90971 , n90975 );
and ( n90977 , n46495 , n61983 );
or ( n90978 , n90976 , n90977 );
and ( n90979 , n90970 , n90978 );
not ( n90980 , n62003 );
not ( n90981 , n62005 );
and ( n90982 , n90981 , n90978 );
and ( n90983 , n46984 , n62005 );
or ( n90984 , n90982 , n90983 );
and ( n90985 , n90980 , n90984 );
and ( n90986 , n47267 , n62003 );
or ( n90987 , n90985 , n90986 );
and ( n90988 , n90987 , n31452 );
or ( n90989 , n90979 , n90988 );
and ( n90990 , n90989 , n31638 );
and ( n90991 , n31168 , n47277 );
or ( n90992 , C0 , n90960 , n90969 , n90990 , n90991 );
buf ( n90993 , n90992 );
buf ( n90994 , n90993 );
buf ( n90995 , n31655 );
buf ( n90996 , n30987 );
buf ( n90997 , n30987 );
xor ( n90998 , n49575 , n60318 );
and ( n90999 , n90998 , n32433 );
not ( n91000 , n47331 );
and ( n91001 , n91000 , n49575 );
xor ( n91002 , n60484 , n60542 );
and ( n91003 , n91002 , n47331 );
or ( n91004 , n91001 , n91003 );
and ( n91005 , n91004 , n32413 );
and ( n91006 , n49575 , n47402 );
or ( n91007 , n90999 , n91005 , n91006 );
and ( n91008 , n91007 , n32456 );
and ( n91009 , n49575 , n47409 );
or ( n91010 , C0 , n91008 , n91009 );
buf ( n91011 , n91010 );
buf ( n91012 , n91011 );
buf ( n91013 , n31655 );
not ( n91014 , n46356 );
and ( n91015 , n91014 , n31256 );
not ( n91016 , n55263 );
and ( n91017 , n91016 , n31256 );
and ( n91018 , n31272 , n55263 );
or ( n91019 , n91017 , n91018 );
and ( n91020 , n91019 , n46356 );
or ( n91021 , n91015 , n91020 );
and ( n91022 , n91021 , n31649 );
not ( n91023 , n55271 );
not ( n91024 , n55263 );
and ( n91025 , n91024 , n31256 );
and ( n91026 , n49443 , n55263 );
or ( n91027 , n91025 , n91026 );
and ( n91028 , n91023 , n91027 );
and ( n91029 , n49443 , n55271 );
or ( n91030 , n91028 , n91029 );
and ( n91031 , n91030 , n31643 );
not ( n91032 , n31452 );
not ( n91033 , n55271 );
not ( n91034 , n55263 );
and ( n91035 , n91034 , n31256 );
and ( n91036 , n49443 , n55263 );
or ( n91037 , n91035 , n91036 );
and ( n91038 , n91033 , n91037 );
and ( n91039 , n49443 , n55271 );
or ( n91040 , n91038 , n91039 );
and ( n91041 , n91032 , n91040 );
not ( n91042 , n55291 );
not ( n91043 , n55293 );
and ( n91044 , n91043 , n91040 );
and ( n91045 , n49469 , n55293 );
or ( n91046 , n91044 , n91045 );
and ( n91047 , n91042 , n91046 );
and ( n91048 , n49477 , n55291 );
or ( n91049 , n91047 , n91048 );
and ( n91050 , n91049 , n31452 );
or ( n91051 , n91041 , n91050 );
and ( n91052 , n91051 , n31638 );
and ( n91053 , n31256 , n47277 );
or ( n91054 , C0 , n91022 , n91031 , n91052 , n91053 );
buf ( n91055 , n91054 );
buf ( n91056 , n91055 );
buf ( n91057 , n31655 );
buf ( n91058 , n30987 );
xor ( n91059 , n46133 , n49989 );
and ( n91060 , n91059 , n32431 );
not ( n91061 , n50002 );
and ( n91062 , n91061 , n46133 );
and ( n91063 , n40305 , n50002 );
or ( n91064 , n91062 , n91063 );
and ( n91065 , n91064 , n32419 );
not ( n91066 , n50008 );
and ( n91067 , n91066 , n46133 );
not ( n91068 , n47910 );
and ( n91069 , n91068 , n55447 );
not ( n91070 , n48101 );
and ( n91071 , n91070 , n47965 );
xor ( n91072 , n48107 , n48115 );
and ( n91073 , n91072 , n48101 );
or ( n91074 , n91071 , n91073 );
and ( n91075 , n91074 , n47910 );
or ( n91076 , n91069 , n91075 );
and ( n91077 , n91076 , n50008 );
or ( n91078 , n91067 , n91077 );
and ( n91079 , n91078 , n32415 );
not ( n91080 , n50067 );
and ( n91081 , n91080 , n46133 );
and ( n91082 , n31928 , n50067 );
or ( n91083 , n91081 , n91082 );
and ( n91084 , n91083 , n32411 );
and ( n91085 , n46133 , n50098 );
or ( n91086 , n91060 , n91065 , n91079 , n91084 , n91085 );
and ( n91087 , n91086 , n32456 );
and ( n91088 , n46133 , n47409 );
or ( n91089 , C0 , n91087 , n91088 );
buf ( n91090 , n91089 );
buf ( n91091 , n91090 );
buf ( n91092 , n31655 );
buf ( n91093 , n30987 );
not ( n91094 , n34150 );
and ( n91095 , n91094 , n32875 );
not ( n91096 , n56836 );
and ( n91097 , n91096 , n32875 );
and ( n91098 , n32889 , n56836 );
or ( n91099 , n91097 , n91098 );
and ( n91100 , n91099 , n34150 );
or ( n91101 , n91095 , n91100 );
and ( n91102 , n91101 , n33381 );
not ( n91103 , n56844 );
not ( n91104 , n56836 );
and ( n91105 , n91104 , n32875 );
and ( n91106 , n52819 , n56836 );
or ( n91107 , n91105 , n91106 );
and ( n91108 , n91103 , n91107 );
and ( n91109 , n52819 , n56844 );
or ( n91110 , n91108 , n91109 );
and ( n91111 , n91110 , n33375 );
not ( n91112 , n32968 );
not ( n91113 , n56844 );
not ( n91114 , n56836 );
and ( n91115 , n91114 , n32875 );
and ( n91116 , n52819 , n56836 );
or ( n91117 , n91115 , n91116 );
and ( n91118 , n91113 , n91117 );
and ( n91119 , n52819 , n56844 );
or ( n91120 , n91118 , n91119 );
and ( n91121 , n91112 , n91120 );
not ( n91122 , n56864 );
not ( n91123 , n56866 );
and ( n91124 , n91123 , n91120 );
and ( n91125 , n52845 , n56866 );
or ( n91126 , n91124 , n91125 );
and ( n91127 , n91122 , n91126 );
and ( n91128 , n52855 , n56864 );
or ( n91129 , n91127 , n91128 );
and ( n91130 , n91129 , n32968 );
or ( n91131 , n91121 , n91130 );
and ( n91132 , n91131 , n33370 );
and ( n91133 , n32875 , n35062 );
or ( n91134 , C0 , n91102 , n91111 , n91132 , n91133 );
buf ( n91135 , n91134 );
buf ( n91136 , n91135 );
buf ( n91137 , n40200 );
buf ( n91138 , n30987 );
buf ( n91139 , n31655 );
buf ( n91140 , n31655 );
buf ( n91141 , n30987 );
buf ( n91142 , n31655 );
xor ( n91143 , n54158 , n54980 );
and ( n91144 , n91143 , n33199 );
not ( n91145 , n48648 );
and ( n91146 , n91145 , n54158 );
and ( n91147 , n34443 , n48648 );
or ( n91148 , n91146 , n91147 );
and ( n91149 , n91148 , n32924 );
not ( n91150 , n48660 );
and ( n91151 , n91150 , n54158 );
and ( n91152 , n83194 , n48660 );
or ( n91153 , n91151 , n91152 );
and ( n91154 , n91153 , n33172 );
not ( n91155 , n48730 );
and ( n91156 , n91155 , n54158 );
and ( n91157 , n32657 , n55215 );
and ( n91158 , n32659 , n55217 );
and ( n91159 , n32661 , n55219 );
and ( n91160 , n32663 , n55221 );
and ( n91161 , n32665 , n55223 );
and ( n91162 , n32667 , n55225 );
and ( n91163 , n32669 , n55227 );
and ( n91164 , n32671 , n55229 );
and ( n91165 , n32673 , n55231 );
and ( n91166 , n32675 , n55233 );
and ( n91167 , n32677 , n55235 );
and ( n91168 , n32679 , n55237 );
and ( n91169 , n32681 , n55239 );
and ( n91170 , n32683 , n55241 );
and ( n91171 , n32685 , n55243 );
and ( n91172 , n32687 , n55245 );
or ( n91173 , n91157 , n91158 , n91159 , n91160 , n91161 , n91162 , n91163 , n91164 , n91165 , n91166 , n91167 , n91168 , n91169 , n91170 , n91171 , n91172 );
and ( n91174 , n91173 , n48730 );
or ( n91175 , n91156 , n91174 );
and ( n91176 , n91175 , n33187 );
and ( n91177 , n54158 , n54713 );
or ( n91178 , n91144 , n91149 , n91154 , n91176 , n91177 );
and ( n91179 , n91178 , n33208 );
and ( n91180 , n54158 , n39805 );
or ( n91181 , C0 , n91179 , n91180 );
buf ( n91182 , n91181 );
buf ( n91183 , n91182 );
buf ( n91184 , n30987 );
buf ( n91185 , n31655 );
not ( n91186 , n41532 );
and ( n91187 , n91186 , n34435 );
buf ( n91188 , RI15b53d30_725);
and ( n91189 , n91188 , n41532 );
or ( n91190 , n91187 , n91189 );
buf ( n91191 , n91190 );
buf ( n91192 , n91191 );
and ( n91193 , n33220 , n32528 );
not ( n91194 , n32598 );
and ( n91195 , n91194 , n32983 );
buf ( n91196 , n91195 );
and ( n91197 , n91196 , n32890 );
not ( n91198 , n32919 );
and ( n91199 , n91198 , n32983 );
buf ( n91200 , n91199 );
and ( n91201 , n91200 , n32924 );
not ( n91202 , n32953 );
and ( n91203 , n91202 , n32983 );
not ( n91204 , n32971 );
and ( n91205 , n91204 , n33091 );
xor ( n91206 , n32983 , n33022 );
and ( n91207 , n91206 , n32971 );
or ( n91208 , n91205 , n91207 );
and ( n91209 , n91208 , n32953 );
or ( n91210 , n91203 , n91209 );
and ( n91211 , n91210 , n33038 );
not ( n91212 , n33067 );
and ( n91213 , n91212 , n32983 );
not ( n91214 , n32970 );
not ( n91215 , n33071 );
and ( n91216 , n91215 , n33091 );
xor ( n91217 , n33092 , n33154 );
and ( n91218 , n91217 , n33071 );
or ( n91219 , n91216 , n91218 );
and ( n91220 , n91214 , n91219 );
and ( n91221 , n91206 , n32970 );
or ( n91222 , n91220 , n91221 );
and ( n91223 , n91222 , n33067 );
or ( n91224 , n91213 , n91223 );
and ( n91225 , n91224 , n33172 );
and ( n91226 , n32983 , n33204 );
or ( n91227 , n91197 , n91201 , n91211 , n91225 , n91226 );
and ( n91228 , n91227 , n33208 );
not ( n91229 , n32968 );
not ( n91230 , n33270 );
and ( n91231 , n91230 , n33291 );
xor ( n91232 , n33292 , n33354 );
and ( n91233 , n91232 , n33270 );
or ( n91234 , n91231 , n91233 );
and ( n91235 , n91229 , n91234 );
and ( n91236 , n32983 , n32968 );
or ( n91237 , n91235 , n91236 );
and ( n91238 , n91237 , n33370 );
and ( n91239 , n32983 , n33382 );
or ( n91240 , C0 , n91193 , n91228 , n91238 , C0 , n91239 );
buf ( n91241 , n91240 );
buf ( n91242 , n91241 );
buf ( n91243 , n30987 );
buf ( n91244 , n31655 );
buf ( n91245 , n30987 );
buf ( n91246 , n31655 );
not ( n91247 , n31728 );
and ( n91248 , n91247 , n46030 );
and ( n91249 , n89822 , n31728 );
or ( n91250 , n91248 , n91249 );
and ( n91251 , n91250 , n32253 );
not ( n91252 , n32283 );
and ( n91253 , n91252 , n46030 );
and ( n91254 , n89833 , n32283 );
or ( n91255 , n91253 , n91254 );
and ( n91256 , n91255 , n32398 );
and ( n91257 , n46030 , n32436 );
or ( n91258 , n91251 , n91256 , n91257 );
and ( n91259 , n91258 , n32456 );
and ( n91260 , n49677 , n32473 );
not ( n91261 , n32475 );
and ( n91262 , n91261 , n49677 );
xor ( n91263 , n46030 , n47756 );
and ( n91264 , n91263 , n32475 );
or ( n91265 , n91262 , n91264 );
and ( n91266 , n91265 , n32486 );
and ( n91267 , n37557 , n32489 );
and ( n91268 , n46030 , n32501 );
or ( n91269 , C0 , n91259 , n91260 , n91266 , n91267 , n91268 );
buf ( n91270 , n91269 );
buf ( n91271 , n91270 );
buf ( n91272 , n30987 );
not ( n91273 , n48765 );
and ( n91274 , n91273 , n33231 );
and ( n91275 , n70548 , n48765 );
or ( n91276 , n91274 , n91275 );
and ( n91277 , n91276 , n33180 );
not ( n91278 , n49054 );
and ( n91279 , n91278 , n33231 );
and ( n91280 , n70559 , n49054 );
or ( n91281 , n91279 , n91280 );
and ( n91282 , n91281 , n33178 );
and ( n91283 , n33231 , n49774 );
or ( n91284 , n91277 , n91282 , n91283 );
and ( n91285 , n91284 , n33208 );
and ( n91286 , n33313 , n33375 );
not ( n91287 , n32968 );
and ( n91288 , n91287 , n33313 );
xor ( n91289 , n33231 , n53898 );
and ( n91290 , n91289 , n32968 );
or ( n91291 , n91288 , n91290 );
and ( n91292 , n91291 , n33370 );
and ( n91293 , n32994 , n35056 );
and ( n91294 , n33231 , n49794 );
or ( n91295 , C0 , n91285 , n91286 , n91292 , n91293 , n91294 );
buf ( n91296 , n91295 );
buf ( n91297 , n91296 );
buf ( n91298 , n31655 );
buf ( n91299 , n30987 );
buf ( n91300 , n31655 );
and ( n91301 , n46019 , n32500 );
not ( n91302 , n35211 );
and ( n91303 , n91302 , n37535 );
buf ( n91304 , n91303 );
and ( n91305 , n91304 , n32421 );
not ( n91306 , n35245 );
and ( n91307 , n91306 , n37535 );
buf ( n91308 , n91307 );
and ( n91309 , n91308 , n32419 );
not ( n91310 , n35278 );
and ( n91311 , n91310 , n37535 );
not ( n91312 , n35295 );
and ( n91313 , n91312 , n49565 );
xor ( n91314 , n37535 , n49548 );
and ( n91315 , n91314 , n35295 );
or ( n91316 , n91313 , n91315 );
and ( n91317 , n91316 , n35278 );
or ( n91318 , n91311 , n91317 );
and ( n91319 , n91318 , n32417 );
not ( n91320 , n35331 );
and ( n91321 , n91320 , n37535 );
not ( n91322 , n35294 );
not ( n91323 , n45995 );
and ( n91324 , n91323 , n49565 );
xor ( n91325 , n49566 , n49634 );
and ( n91326 , n91325 , n45995 );
or ( n91327 , n91324 , n91326 );
and ( n91328 , n91322 , n91327 );
and ( n91329 , n91314 , n35294 );
or ( n91330 , n91328 , n91329 );
and ( n91331 , n91330 , n35331 );
or ( n91332 , n91321 , n91331 );
and ( n91333 , n91332 , n32415 );
and ( n91334 , n37535 , n35354 );
or ( n91335 , n91305 , n91309 , n91319 , n91333 , n91334 );
and ( n91336 , n91335 , n32456 );
not ( n91337 , n32475 );
not ( n91338 , n46060 );
and ( n91339 , n91338 , n49656 );
xor ( n91340 , n49657 , n49728 );
and ( n91341 , n91340 , n46060 );
or ( n91342 , n91339 , n91341 );
and ( n91343 , n91337 , n91342 );
and ( n91344 , n37535 , n32475 );
or ( n91345 , n91343 , n91344 );
and ( n91346 , n91345 , n32486 );
and ( n91347 , n37535 , n35367 );
or ( n91348 , C0 , n91301 , n91336 , n91346 , C0 , n91347 );
buf ( n91349 , n91348 );
buf ( n91350 , n91349 );
not ( n91351 , n46356 );
and ( n91352 , n91351 , n31142 );
not ( n91353 , n47831 );
and ( n91354 , n91353 , n31142 );
and ( n91355 , n31172 , n47831 );
or ( n91356 , n91354 , n91355 );
and ( n91357 , n91356 , n46356 );
or ( n91358 , n91352 , n91357 );
and ( n91359 , n91358 , n31649 );
not ( n91360 , n47839 );
not ( n91361 , n47831 );
and ( n91362 , n91361 , n31142 );
and ( n91363 , n46495 , n47831 );
or ( n91364 , n91362 , n91363 );
and ( n91365 , n91360 , n91364 );
and ( n91366 , n46495 , n47839 );
or ( n91367 , n91365 , n91366 );
and ( n91368 , n91367 , n31643 );
not ( n91369 , n31452 );
not ( n91370 , n47839 );
not ( n91371 , n47831 );
and ( n91372 , n91371 , n31142 );
and ( n91373 , n46495 , n47831 );
or ( n91374 , n91372 , n91373 );
and ( n91375 , n91370 , n91374 );
and ( n91376 , n46495 , n47839 );
or ( n91377 , n91375 , n91376 );
and ( n91378 , n91369 , n91377 );
not ( n91379 , n47866 );
not ( n91380 , n47868 );
and ( n91381 , n91380 , n91377 );
and ( n91382 , n46984 , n47868 );
or ( n91383 , n91381 , n91382 );
and ( n91384 , n91379 , n91383 );
and ( n91385 , n47267 , n47866 );
or ( n91386 , n91384 , n91385 );
and ( n91387 , n91386 , n31452 );
or ( n91388 , n91378 , n91387 );
and ( n91389 , n91388 , n31638 );
and ( n91390 , n31142 , n47277 );
or ( n91391 , C0 , n91359 , n91368 , n91389 , n91390 );
buf ( n91392 , n91391 );
buf ( n91393 , n91392 );
buf ( n91394 , n31655 );
buf ( n91395 , n30987 );
not ( n91396 , n35278 );
and ( n91397 , n91396 , n46081 );
and ( n91398 , n46322 , n35278 );
or ( n91399 , n91397 , n91398 );
and ( n91400 , n91399 , n32417 );
not ( n91401 , n47912 );
and ( n91402 , n91401 , n46081 );
and ( n91403 , n63362 , n47912 );
or ( n91404 , n91402 , n91403 );
and ( n91405 , n91404 , n32415 );
and ( n91406 , n46081 , n48133 );
or ( n91407 , n91400 , n91405 , n91406 );
and ( n91408 , n91407 , n32456 );
and ( n91409 , n46081 , n47409 );
or ( n91410 , C0 , n91408 , n91409 );
buf ( n91411 , n91410 );
buf ( n91412 , n91411 );
buf ( n91413 , n31655 );
buf ( n91414 , n30987 );
not ( n91415 , n32953 );
and ( n91416 , n91415 , n55411 );
and ( n91417 , n81150 , n32953 );
or ( n91418 , n91416 , n91417 );
and ( n91419 , n91418 , n33038 );
not ( n91420 , n39586 );
and ( n91421 , n91420 , n55411 );
and ( n91422 , n55417 , n39586 );
or ( n91423 , n91421 , n91422 );
and ( n91424 , n91423 , n33172 );
and ( n91425 , n55411 , n39795 );
or ( n91426 , n91419 , n91424 , n91425 );
and ( n91427 , n91426 , n33208 );
and ( n91428 , n55411 , n39805 );
or ( n91429 , C0 , n91427 , n91428 );
buf ( n91430 , n91429 );
buf ( n91431 , n91430 );
buf ( n91432 , n31655 );
buf ( n91433 , n30987 );
buf ( n91434 , n31655 );
buf ( n91435 , n31655 );
xor ( n91436 , n41730 , n44785 );
and ( n91437 , n91436 , n31548 );
not ( n91438 , n44807 );
and ( n91439 , n91438 , n41730 );
and ( n91440 , n42030 , n44807 );
or ( n91441 , n91439 , n91440 );
and ( n91442 , n91441 , n31408 );
not ( n91443 , n44817 );
and ( n91444 , n91443 , n41730 );
not ( n91445 , n41835 );
and ( n91446 , n91445 , n53287 );
and ( n91447 , n89339 , n41835 );
or ( n91448 , n91446 , n91447 );
and ( n91449 , n91448 , n44817 );
or ( n91450 , n91444 , n91449 );
and ( n91451 , n91450 , n31521 );
not ( n91452 , n45059 );
and ( n91453 , n91452 , n41730 );
and ( n91454 , n60067 , n45059 );
or ( n91455 , n91453 , n91454 );
and ( n91456 , n91455 , n31536 );
and ( n91457 , n41730 , n45148 );
or ( n91458 , n91437 , n91442 , n91451 , n91456 , n91457 );
and ( n91459 , n91458 , n31557 );
and ( n91460 , n41730 , n40154 );
or ( n91461 , C0 , n91459 , n91460 );
buf ( n91462 , n91461 );
buf ( n91463 , n91462 );
not ( n91464 , n40163 );
and ( n91465 , n91464 , n31844 );
not ( n91466 , n49298 );
and ( n91467 , n91466 , n31844 );
and ( n91468 , n32235 , n49298 );
or ( n91469 , n91467 , n91468 );
and ( n91470 , n91469 , n40163 );
or ( n91471 , n91465 , n91470 );
and ( n91472 , n91471 , n32498 );
not ( n91473 , n49306 );
not ( n91474 , n49298 );
and ( n91475 , n91474 , n31844 );
and ( n91476 , n42188 , n49298 );
or ( n91477 , n91475 , n91476 );
and ( n91478 , n91473 , n91477 );
and ( n91479 , n42188 , n49306 );
or ( n91480 , n91478 , n91479 );
and ( n91481 , n91480 , n32473 );
not ( n91482 , n32475 );
not ( n91483 , n49306 );
not ( n91484 , n49298 );
and ( n91485 , n91484 , n31844 );
and ( n91486 , n42188 , n49298 );
or ( n91487 , n91485 , n91486 );
and ( n91488 , n91483 , n91487 );
and ( n91489 , n42188 , n49306 );
or ( n91490 , n91488 , n91489 );
and ( n91491 , n91482 , n91490 );
not ( n91492 , n49331 );
not ( n91493 , n49333 );
and ( n91494 , n91493 , n91490 );
and ( n91495 , n42216 , n49333 );
or ( n91496 , n91494 , n91495 );
and ( n91497 , n91492 , n91496 );
and ( n91498 , n42224 , n49331 );
or ( n91499 , n91497 , n91498 );
and ( n91500 , n91499 , n32475 );
or ( n91501 , n91491 , n91500 );
and ( n91502 , n91501 , n32486 );
and ( n91503 , n31844 , n41278 );
or ( n91504 , C0 , n91472 , n91481 , n91502 , n91503 );
buf ( n91505 , n91504 );
buf ( n91506 , n91505 );
buf ( n91507 , n30987 );
buf ( n91508 , n30987 );
buf ( n91509 , n31655 );
buf ( n91510 , n72718 );
xor ( n91511 , n35435 , n39946 );
and ( n91512 , n91511 , n31550 );
not ( n91513 , n39979 );
and ( n91514 , n91513 , n35435 );
xor ( n91515 , n40052 , n40128 );
and ( n91516 , n91515 , n39979 );
or ( n91517 , n91514 , n91516 );
and ( n91518 , n91517 , n31538 );
and ( n91519 , n35435 , n40143 );
or ( n91520 , n91512 , n91518 , n91519 );
and ( n91521 , n91520 , n31557 );
and ( n91522 , n35435 , n40154 );
or ( n91523 , C0 , n91521 , n91522 );
buf ( n91524 , n91523 );
buf ( n91525 , n91524 );
not ( n91526 , n40163 );
and ( n91527 , n91526 , n32064 );
not ( n91528 , n75905 );
and ( n91529 , n91528 , n32064 );
and ( n91530 , n32130 , n75905 );
or ( n91531 , n91529 , n91530 );
and ( n91532 , n91531 , n40163 );
or ( n91533 , n91527 , n91532 );
and ( n91534 , n91533 , n32498 );
not ( n91535 , n75913 );
not ( n91536 , n75905 );
and ( n91537 , n91536 , n32064 );
and ( n91538 , n45833 , n75905 );
or ( n91539 , n91537 , n91538 );
and ( n91540 , n91535 , n91539 );
and ( n91541 , n45833 , n75913 );
or ( n91542 , n91540 , n91541 );
and ( n91543 , n91542 , n32473 );
not ( n91544 , n32475 );
not ( n91545 , n75913 );
not ( n91546 , n75905 );
and ( n91547 , n91546 , n32064 );
and ( n91548 , n45833 , n75905 );
or ( n91549 , n91547 , n91548 );
and ( n91550 , n91545 , n91549 );
and ( n91551 , n45833 , n75913 );
or ( n91552 , n91550 , n91551 );
and ( n91553 , n91544 , n91552 );
not ( n91554 , n75933 );
not ( n91555 , n75935 );
and ( n91556 , n91555 , n91552 );
and ( n91557 , n45857 , n75935 );
or ( n91558 , n91556 , n91557 );
and ( n91559 , n91554 , n91558 );
and ( n91560 , n45865 , n75933 );
or ( n91561 , n91559 , n91560 );
and ( n91562 , n91561 , n32475 );
or ( n91563 , n91553 , n91562 );
and ( n91564 , n91563 , n32486 );
and ( n91565 , n32064 , n41278 );
or ( n91566 , C0 , n91534 , n91543 , n91564 , n91565 );
buf ( n91567 , n91566 );
buf ( n91568 , n91567 );
buf ( n91569 , n30987 );
buf ( n91570 , n30987 );
and ( n91571 , n33757 , n48455 );
not ( n91572 , n48457 );
and ( n91573 , n91572 , n33422 );
and ( n91574 , n33757 , n48457 );
or ( n91575 , n91573 , n91574 );
and ( n91576 , n91575 , n31373 );
not ( n91577 , n44807 );
and ( n91578 , n91577 , n33422 );
and ( n91579 , n33757 , n44807 );
or ( n91580 , n91578 , n91579 );
and ( n91581 , n91580 , n31408 );
not ( n91582 , n48468 );
and ( n91583 , n91582 , n33422 );
and ( n91584 , n33757 , n48468 );
or ( n91585 , n91583 , n91584 );
and ( n91586 , n91585 , n31468 );
not ( n91587 , n44817 );
and ( n91588 , n91587 , n33422 );
and ( n91589 , n33757 , n44817 );
or ( n91590 , n91588 , n91589 );
and ( n91591 , n91590 , n31521 );
not ( n91592 , n39979 );
and ( n91593 , n91592 , n33422 );
and ( n91594 , n33464 , n39979 );
or ( n91595 , n91593 , n91594 );
and ( n91596 , n91595 , n31538 );
not ( n91597 , n45059 );
and ( n91598 , n91597 , n33422 );
and ( n91599 , n33464 , n45059 );
or ( n91600 , n91598 , n91599 );
and ( n91601 , n91600 , n31536 );
not ( n91602 , n33419 );
and ( n91603 , n91602 , n33422 );
and ( n91604 , n33702 , n33419 );
or ( n91605 , n91603 , n91604 );
and ( n91606 , n91605 , n31529 );
not ( n91607 , n33734 );
and ( n91608 , n91607 , n33422 );
and ( n91609 , n33924 , n33734 );
or ( n91610 , n91608 , n91609 );
and ( n91611 , n91610 , n31527 );
and ( n91612 , n33842 , n48513 );
or ( n91613 , n91571 , n91576 , n91581 , n91586 , n91591 , n91596 , n91601 , n91606 , n91611 , n91612 );
and ( n91614 , n91613 , n31557 );
and ( n91615 , n33972 , n33973 );
and ( n91616 , n33422 , n48524 );
or ( n91617 , C0 , n91614 , n91615 , n91616 );
buf ( n91618 , n91617 );
buf ( n91619 , n91618 );
buf ( n91620 , n31655 );
buf ( n91621 , n30987 );
not ( n91622 , n38443 );
and ( n91623 , n91622 , n38388 );
xor ( n91624 , n69918 , n69919 );
and ( n91625 , n91624 , n38443 );
or ( n91626 , n91623 , n91625 );
and ( n91627 , n91626 , n38450 );
not ( n91628 , n39339 );
and ( n91629 , n91628 , n39288 );
xor ( n91630 , n69932 , n69933 );
and ( n91631 , n91630 , n39339 );
or ( n91632 , n91629 , n91631 );
and ( n91633 , n91632 , n39346 );
and ( n91634 , n40225 , n39359 );
or ( n91635 , n91627 , n91633 , n91634 );
buf ( n91636 , n91635 );
buf ( n91637 , n91636 );
buf ( n91638 , n31655 );
buf ( n91639 , n31655 );
not ( n91640 , n33419 );
and ( n91641 , n91640 , n31580 );
xor ( n91642 , n33474 , n33691 );
and ( n91643 , n91642 , n33419 );
or ( n91644 , n91641 , n91643 );
and ( n91645 , n91644 , n31529 );
not ( n91646 , n33734 );
and ( n91647 , n91646 , n31580 );
not ( n91648 , n33533 );
xor ( n91649 , n33767 , n33809 );
and ( n91650 , n91648 , n91649 );
xnor ( n91651 , n33852 , n33911 );
and ( n91652 , n91651 , n33533 );
or ( n91653 , n91650 , n91652 );
and ( n91654 , n91653 , n33734 );
or ( n91655 , n91647 , n91654 );
and ( n91656 , n91655 , n31527 );
and ( n91657 , n31580 , n33942 );
or ( n91658 , n91645 , n91656 , n91657 );
and ( n91659 , n91658 , n31557 );
and ( n91660 , n34105 , n31643 );
not ( n91661 , n31452 );
and ( n91662 , n91661 , n34105 );
xor ( n91663 , n31580 , n33957 );
and ( n91664 , n91663 , n31452 );
or ( n91665 , n91662 , n91664 );
and ( n91666 , n91665 , n31638 );
and ( n91667 , n34004 , n33973 );
and ( n91668 , n31580 , n33978 );
or ( n91669 , C0 , n91659 , n91660 , n91666 , n91667 , n91668 );
buf ( n91670 , n91669 );
buf ( n91671 , n91670 );
and ( n91672 , n31564 , n31007 );
not ( n91673 , n31077 );
and ( n91674 , n91673 , n35390 );
buf ( n91675 , n91674 );
and ( n91676 , n91675 , n31373 );
not ( n91677 , n31402 );
and ( n91678 , n91677 , n35390 );
buf ( n91679 , n91678 );
and ( n91680 , n91679 , n31408 );
not ( n91681 , n31437 );
and ( n91682 , n91681 , n35390 );
not ( n91683 , n31455 );
and ( n91684 , n91683 , n35429 );
xor ( n91685 , n35390 , n35408 );
and ( n91686 , n91685 , n31455 );
or ( n91687 , n91684 , n91686 );
and ( n91688 , n91687 , n31437 );
or ( n91689 , n91682 , n91688 );
and ( n91690 , n91689 , n31468 );
not ( n91691 , n31497 );
and ( n91692 , n91691 , n35390 );
not ( n91693 , n31454 );
not ( n91694 , n31501 );
and ( n91695 , n91694 , n35429 );
xor ( n91696 , n35430 , n35458 );
and ( n91697 , n91696 , n31501 );
or ( n91698 , n91695 , n91697 );
and ( n91699 , n91693 , n91698 );
and ( n91700 , n91685 , n31454 );
or ( n91701 , n91699 , n91700 );
and ( n91702 , n91701 , n31497 );
or ( n91703 , n91692 , n91702 );
and ( n91704 , n91703 , n31521 );
and ( n91705 , n35390 , n31553 );
or ( n91706 , n91676 , n91680 , n91690 , n91704 , n91705 );
and ( n91707 , n91706 , n31557 );
not ( n91708 , n31452 );
not ( n91709 , n31619 );
and ( n91710 , n91709 , n35484 );
xor ( n91711 , n35485 , n35512 );
and ( n91712 , n91711 , n31619 );
or ( n91713 , n91710 , n91712 );
and ( n91714 , n91708 , n91713 );
and ( n91715 , n35390 , n31452 );
or ( n91716 , n91714 , n91715 );
and ( n91717 , n91716 , n31638 );
and ( n91718 , n35390 , n31650 );
or ( n91719 , C0 , n91672 , n91707 , n91717 , C0 , n91718 );
buf ( n91720 , n91719 );
buf ( n91721 , n91720 );
buf ( n91722 , n30987 );
buf ( n91723 , n30987 );
buf ( n91724 , n30987 );
buf ( n91725 , n30987 );
not ( n91726 , n34150 );
and ( n91727 , n91726 , n32652 );
not ( n91728 , n56239 );
and ( n91729 , n91728 , n32652 );
and ( n91730 , n32655 , n56239 );
or ( n91731 , n91729 , n91730 );
and ( n91732 , n91731 , n34150 );
or ( n91733 , n91727 , n91732 );
and ( n91734 , n91733 , n33381 );
not ( n91735 , n56247 );
not ( n91736 , n56239 );
and ( n91737 , n91736 , n32652 );
and ( n91738 , n56044 , n56239 );
or ( n91739 , n91737 , n91738 );
and ( n91740 , n91735 , n91739 );
and ( n91741 , n56044 , n56247 );
or ( n91742 , n91740 , n91741 );
and ( n91743 , n91742 , n33375 );
not ( n91744 , n32968 );
not ( n91745 , n56247 );
not ( n91746 , n56239 );
and ( n91747 , n91746 , n32652 );
and ( n91748 , n56044 , n56239 );
or ( n91749 , n91747 , n91748 );
and ( n91750 , n91745 , n91749 );
and ( n91751 , n56044 , n56247 );
or ( n91752 , n91750 , n91751 );
and ( n91753 , n91744 , n91752 );
not ( n91754 , n56267 );
not ( n91755 , n56269 );
and ( n91756 , n91755 , n91752 );
and ( n91757 , n56068 , n56269 );
or ( n91758 , n91756 , n91757 );
and ( n91759 , n91754 , n91758 );
and ( n91760 , n56076 , n56267 );
or ( n91761 , n91759 , n91760 );
and ( n91762 , n91761 , n32968 );
or ( n91763 , n91753 , n91762 );
and ( n91764 , n91763 , n33370 );
and ( n91765 , n32652 , n35062 );
or ( n91766 , C0 , n91734 , n91743 , n91764 , n91765 );
buf ( n91767 , n91766 );
buf ( n91768 , n91767 );
not ( n91769 , n34150 );
and ( n91770 , n91769 , n32879 );
not ( n91771 , n56192 );
and ( n91772 , n91771 , n32879 );
and ( n91773 , n32889 , n56192 );
or ( n91774 , n91772 , n91773 );
and ( n91775 , n91774 , n34150 );
or ( n91776 , n91770 , n91775 );
and ( n91777 , n91776 , n33381 );
not ( n91778 , n56200 );
not ( n91779 , n56192 );
and ( n91780 , n91779 , n32879 );
and ( n91781 , n52819 , n56192 );
xor ( n91782 , n91780 , n91781 );
and ( n91783 , n91778 , n91782 );
and ( n91784 , n52819 , n56200 );
xor ( n91785 , n91783 , n91784 );
and ( n91786 , n91785 , n33375 );
not ( n91787 , n32968 );
not ( n91788 , n56200 );
not ( n91789 , n56192 );
and ( n91790 , n91789 , n32879 );
and ( n91791 , n52819 , n56192 );
or ( n91792 , n91790 , n91791 );
and ( n91793 , n91788 , n91792 );
and ( n91794 , n52819 , n56200 );
or ( n91795 , n91793 , n91794 );
and ( n91796 , n91787 , n91795 );
not ( n91797 , n56220 );
not ( n91798 , n56222 );
and ( n91799 , n91798 , n91795 );
and ( n91800 , n52845 , n56222 );
or ( n91801 , n91799 , n91800 );
and ( n91802 , n91797 , n91801 );
and ( n91803 , n52855 , n56220 );
or ( n91804 , n91802 , n91803 );
and ( n91805 , n91804 , n32968 );
or ( n91806 , n91796 , n91805 );
and ( n91807 , n91806 , n33370 );
and ( n91808 , n32879 , n35062 );
or ( n91809 , C0 , n91777 , n91786 , n91807 , n91808 );
buf ( n91810 , n91809 );
buf ( n91811 , n91810 );
buf ( n91812 , n31655 );
buf ( n91813 , n31655 );
buf ( n91814 , n31655 );
not ( n91815 , n36587 );
and ( n91816 , n91815 , n36464 );
xor ( n91817 , n50173 , n50214 );
and ( n91818 , n91817 , n36587 );
or ( n91819 , n91816 , n91818 );
and ( n91820 , n91819 , n36596 );
not ( n91821 , n37485 );
and ( n91822 , n91821 , n37366 );
xor ( n91823 , n50223 , n50264 );
and ( n91824 , n91823 , n37485 );
or ( n91825 , n91822 , n91824 );
and ( n91826 , n91825 , n37494 );
and ( n91827 , n41861 , n37506 );
or ( n91828 , n91820 , n91826 , n91827 );
buf ( n91829 , n91828 );
buf ( n91830 , n91829 );
and ( n91831 , n47654 , n50275 );
not ( n91832 , n50278 );
and ( n91833 , n91832 , n47567 );
and ( n91834 , n47654 , n50278 );
or ( n91835 , n91833 , n91834 );
and ( n91836 , n91835 , n32421 );
not ( n91837 , n50002 );
and ( n91838 , n91837 , n47567 );
and ( n91839 , n47654 , n50002 );
or ( n91840 , n91838 , n91839 );
and ( n91841 , n91840 , n32419 );
not ( n91842 , n50289 );
and ( n91843 , n91842 , n47567 );
and ( n91844 , n47654 , n50289 );
or ( n91845 , n91843 , n91844 );
and ( n91846 , n91845 , n32417 );
not ( n91847 , n50008 );
and ( n91848 , n91847 , n47567 );
and ( n91849 , n47654 , n50008 );
or ( n91850 , n91848 , n91849 );
and ( n91851 , n91850 , n32415 );
not ( n91852 , n47331 );
and ( n91853 , n91852 , n47567 );
and ( n91854 , n47599 , n47331 );
or ( n91855 , n91853 , n91854 );
and ( n91856 , n91855 , n32413 );
not ( n91857 , n50067 );
and ( n91858 , n91857 , n47567 );
and ( n91859 , n47599 , n50067 );
or ( n91860 , n91858 , n91859 );
and ( n91861 , n91860 , n32411 );
not ( n91862 , n31728 );
and ( n91863 , n91862 , n47567 );
and ( n91864 , n47631 , n31728 );
or ( n91865 , n91863 , n91864 );
and ( n91866 , n91865 , n32253 );
not ( n91867 , n32283 );
and ( n91868 , n91867 , n47567 );
and ( n91869 , n47738 , n32283 );
or ( n91870 , n91868 , n91869 );
and ( n91871 , n91870 , n32398 );
and ( n91872 , n47704 , n50334 );
or ( n91873 , n91831 , n91836 , n91841 , n91846 , n91851 , n91856 , n91861 , n91866 , n91871 , n91872 );
and ( n91874 , n91873 , n32456 );
and ( n91875 , n37541 , n32489 );
and ( n91876 , n47567 , n50345 );
or ( n91877 , C0 , n91874 , n91875 , n91876 );
buf ( n91878 , n91877 );
buf ( n91879 , n91878 );
buf ( n91880 , n30987 );
buf ( n91881 , n31655 );
not ( n91882 , n46356 );
and ( n91883 , n91882 , n31158 );
not ( n91884 , n50109 );
and ( n91885 , n91884 , n31158 );
and ( n91886 , n31172 , n50109 );
or ( n91887 , n91885 , n91886 );
and ( n91888 , n91887 , n46356 );
or ( n91889 , n91883 , n91888 );
and ( n91890 , n91889 , n31649 );
not ( n91891 , n50117 );
not ( n91892 , n50109 );
and ( n91893 , n91892 , n31158 );
and ( n91894 , n46495 , n50109 );
or ( n91895 , n91893 , n91894 );
and ( n91896 , n91891 , n91895 );
and ( n91897 , n46495 , n50117 );
or ( n91898 , n91896 , n91897 );
and ( n91899 , n91898 , n31643 );
not ( n91900 , n31452 );
not ( n91901 , n50117 );
not ( n91902 , n50109 );
and ( n91903 , n91902 , n31158 );
and ( n91904 , n46495 , n50109 );
or ( n91905 , n91903 , n91904 );
and ( n91906 , n91901 , n91905 );
and ( n91907 , n46495 , n50117 );
or ( n91908 , n91906 , n91907 );
and ( n91909 , n91900 , n91908 );
not ( n91910 , n50142 );
not ( n91911 , n50144 );
and ( n91912 , n91911 , n91908 );
and ( n91913 , n46984 , n50144 );
or ( n91914 , n91912 , n91913 );
and ( n91915 , n91910 , n91914 );
and ( n91916 , n47267 , n50142 );
or ( n91917 , n91915 , n91916 );
and ( n91918 , n91917 , n31452 );
or ( n91919 , n91909 , n91918 );
and ( n91920 , n91919 , n31638 );
and ( n91921 , n31158 , n47277 );
or ( n91922 , C0 , n91890 , n91899 , n91920 , n91921 );
buf ( n91923 , n91922 );
buf ( n91924 , n91923 );
buf ( n91925 , n30987 );
xor ( n91926 , n46276 , n64708 );
and ( n91927 , n91926 , n32431 );
not ( n91928 , n50002 );
and ( n91929 , n91928 , n46276 );
and ( n91930 , n40465 , n50002 );
or ( n91931 , n91929 , n91930 );
and ( n91932 , n91931 , n32419 );
not ( n91933 , n50008 );
and ( n91934 , n91933 , n46276 );
not ( n91935 , n47910 );
and ( n91936 , n91935 , n88732 );
not ( n91937 , n48101 );
and ( n91938 , n91937 , n48097 );
xor ( n91939 , n48097 , n40244 );
and ( n91940 , n50016 , n50029 );
xor ( n91941 , n91939 , n91940 );
and ( n91942 , n91941 , n48101 );
or ( n91943 , n91938 , n91942 );
and ( n91944 , n91943 , n47910 );
or ( n91945 , n91936 , n91944 );
and ( n91946 , n91945 , n50008 );
or ( n91947 , n91934 , n91946 );
and ( n91948 , n91947 , n32415 );
not ( n91949 , n50067 );
and ( n91950 , n91949 , n46276 );
and ( n91951 , n64111 , n50067 );
or ( n91952 , n91950 , n91951 );
and ( n91953 , n91952 , n32411 );
and ( n91954 , n46276 , n50098 );
or ( n91955 , n91927 , n91932 , n91948 , n91953 , n91954 );
and ( n91956 , n91955 , n32456 );
and ( n91957 , n46276 , n47409 );
or ( n91958 , C0 , n91956 , n91957 );
buf ( n91959 , n91958 );
buf ( n91960 , n91959 );
buf ( n91961 , n31655 );
buf ( n91962 , n30987 );
not ( n91963 , n34150 );
and ( n91964 , n91963 , n32700 );
not ( n91965 , n58762 );
and ( n91966 , n91965 , n32700 );
and ( n91967 , n32722 , n58762 );
or ( n91968 , n91966 , n91967 );
and ( n91969 , n91968 , n34150 );
or ( n91970 , n91964 , n91969 );
and ( n91971 , n91970 , n33381 );
not ( n91972 , n58770 );
not ( n91973 , n58762 );
and ( n91974 , n91973 , n32700 );
and ( n91975 , n42565 , n58762 );
or ( n91976 , n91974 , n91975 );
and ( n91977 , n91972 , n91976 );
and ( n91978 , n42565 , n58770 );
or ( n91979 , n91977 , n91978 );
and ( n91980 , n91979 , n33375 );
not ( n91981 , n32968 );
not ( n91982 , n58770 );
not ( n91983 , n58762 );
and ( n91984 , n91983 , n32700 );
and ( n91985 , n42565 , n58762 );
or ( n91986 , n91984 , n91985 );
and ( n91987 , n91982 , n91986 );
and ( n91988 , n42565 , n58770 );
or ( n91989 , n91987 , n91988 );
and ( n91990 , n91981 , n91989 );
not ( n91991 , n58790 );
not ( n91992 , n58792 );
and ( n91993 , n91992 , n91989 );
and ( n91994 , n42589 , n58792 );
or ( n91995 , n91993 , n91994 );
and ( n91996 , n91991 , n91995 );
and ( n91997 , n42597 , n58790 );
or ( n91998 , n91996 , n91997 );
and ( n91999 , n91998 , n32968 );
or ( n92000 , n91990 , n91999 );
and ( n92001 , n92000 , n33370 );
and ( n92002 , n32700 , n35062 );
or ( n92003 , C0 , n91971 , n91980 , n92001 , n92002 );
buf ( n92004 , n92003 );
buf ( n92005 , n92004 );
buf ( n92006 , n30987 );
buf ( n92007 , n31655 );
buf ( n92008 , n31655 );
not ( n92009 , n34150 );
and ( n92010 , n92009 , n32675 );
not ( n92011 , n56836 );
and ( n92012 , n92011 , n32675 );
and ( n92013 , n32689 , n56836 );
or ( n92014 , n92012 , n92013 );
and ( n92015 , n92014 , n34150 );
or ( n92016 , n92010 , n92015 );
and ( n92017 , n92016 , n33381 );
not ( n92018 , n56844 );
not ( n92019 , n56836 );
and ( n92020 , n92019 , n32675 );
and ( n92021 , n50682 , n56836 );
or ( n92022 , n92020 , n92021 );
and ( n92023 , n92018 , n92022 );
and ( n92024 , n50682 , n56844 );
or ( n92025 , n92023 , n92024 );
and ( n92026 , n92025 , n33375 );
not ( n92027 , n32968 );
not ( n92028 , n56844 );
not ( n92029 , n56836 );
and ( n92030 , n92029 , n32675 );
and ( n92031 , n50682 , n56836 );
or ( n92032 , n92030 , n92031 );
and ( n92033 , n92028 , n92032 );
and ( n92034 , n50682 , n56844 );
or ( n92035 , n92033 , n92034 );
and ( n92036 , n92027 , n92035 );
not ( n92037 , n56864 );
not ( n92038 , n56866 );
and ( n92039 , n92038 , n92035 );
and ( n92040 , n50706 , n56866 );
or ( n92041 , n92039 , n92040 );
and ( n92042 , n92037 , n92041 );
and ( n92043 , n50714 , n56864 );
or ( n92044 , n92042 , n92043 );
and ( n92045 , n92044 , n32968 );
or ( n92046 , n92036 , n92045 );
and ( n92047 , n92046 , n33370 );
and ( n92048 , n32675 , n35062 );
or ( n92049 , C0 , n92017 , n92026 , n92047 , n92048 );
buf ( n92050 , n92049 );
buf ( n92051 , n92050 );
buf ( n92052 , n30987 );
buf ( n92053 , n30987 );
not ( n92054 , n35542 );
and ( n92055 , n92054 , n41846 );
and ( n92056 , n67353 , n35542 );
or ( n92057 , n92055 , n92056 );
buf ( n92058 , n92057 );
buf ( n92059 , n92058 );
buf ( n92060 , n31655 );
buf ( n92061 , n31655 );
buf ( n92062 , n31655 );
and ( n92063 , n54004 , n31645 );
not ( n92064 , n45274 );
and ( n92065 , n92064 , n41535 );
not ( n92066 , n41809 );
and ( n92067 , n92066 , n41649 );
xor ( n92068 , n41817 , n41823 );
and ( n92069 , n92068 , n41809 );
or ( n92070 , n92067 , n92069 );
and ( n92071 , n92070 , n45274 );
or ( n92072 , n92065 , n92071 );
and ( n92073 , n92072 , n31373 );
not ( n92074 , n45280 );
and ( n92075 , n92074 , n41535 );
and ( n92076 , n92070 , n45280 );
or ( n92077 , n92075 , n92076 );
and ( n92078 , n92077 , n31468 );
and ( n92079 , n41535 , n45802 );
or ( n92080 , n92073 , n92078 , n92079 );
and ( n92081 , n92080 , n31557 );
and ( n92082 , n41535 , n45808 );
or ( n92083 , C0 , n92063 , n92081 , n92082 );
buf ( n92084 , n92083 );
buf ( n92085 , n92084 );
not ( n92086 , n40163 );
and ( n92087 , n92086 , n31935 );
not ( n92088 , n56287 );
and ( n92089 , n92088 , n31935 );
and ( n92090 , n32183 , n56287 );
or ( n92091 , n92089 , n92090 );
and ( n92092 , n92091 , n40163 );
or ( n92093 , n92087 , n92092 );
and ( n92094 , n92093 , n32498 );
not ( n92095 , n56295 );
not ( n92096 , n56287 );
and ( n92097 , n92096 , n31935 );
and ( n92098 , n45178 , n56287 );
or ( n92099 , n92097 , n92098 );
and ( n92100 , n92095 , n92099 );
and ( n92101 , n45178 , n56295 );
or ( n92102 , n92100 , n92101 );
and ( n92103 , n92102 , n32473 );
not ( n92104 , n32475 );
not ( n92105 , n56295 );
not ( n92106 , n56287 );
and ( n92107 , n92106 , n31935 );
and ( n92108 , n45178 , n56287 );
or ( n92109 , n92107 , n92108 );
and ( n92110 , n92105 , n92109 );
and ( n92111 , n45178 , n56295 );
or ( n92112 , n92110 , n92111 );
and ( n92113 , n92104 , n92112 );
not ( n92114 , n56315 );
not ( n92115 , n56317 );
and ( n92116 , n92115 , n92112 );
and ( n92117 , n45206 , n56317 );
or ( n92118 , n92116 , n92117 );
and ( n92119 , n92114 , n92118 );
and ( n92120 , n45214 , n56315 );
or ( n92121 , n92119 , n92120 );
and ( n92122 , n92121 , n32475 );
or ( n92123 , n92113 , n92122 );
and ( n92124 , n92123 , n32486 );
and ( n92125 , n31935 , n41278 );
or ( n92126 , C0 , n92094 , n92103 , n92124 , n92125 );
buf ( n92127 , n92126 );
buf ( n92128 , n92127 );
buf ( n92129 , n30987 );
buf ( n92130 , n31655 );
xor ( n92131 , n34046 , n39934 );
and ( n92132 , n92131 , n31550 );
not ( n92133 , n39979 );
and ( n92134 , n92133 , n34046 );
and ( n92135 , n65656 , n39979 );
or ( n92136 , n92134 , n92135 );
and ( n92137 , n92136 , n31538 );
and ( n92138 , n34046 , n40143 );
or ( n92139 , n92132 , n92137 , n92138 );
and ( n92140 , n92139 , n31557 );
and ( n92141 , n34046 , n40154 );
or ( n92142 , C0 , n92140 , n92141 );
buf ( n92143 , n92142 );
buf ( n92144 , n92143 );
not ( n92145 , n40163 );
and ( n92146 , n92145 , n31922 );
not ( n92147 , n42238 );
and ( n92148 , n92147 , n31922 );
and ( n92149 , n32200 , n42238 );
or ( n92150 , n92148 , n92149 );
and ( n92151 , n92150 , n40163 );
or ( n92152 , n92146 , n92151 );
and ( n92153 , n92152 , n32498 );
not ( n92154 , n42247 );
not ( n92155 , n42238 );
and ( n92156 , n92155 , n31922 );
and ( n92157 , n53243 , n42238 );
or ( n92158 , n92156 , n92157 );
and ( n92159 , n92154 , n92158 );
and ( n92160 , n53243 , n42247 );
or ( n92161 , n92159 , n92160 );
and ( n92162 , n92161 , n32473 );
not ( n92163 , n32475 );
not ( n92164 , n42247 );
not ( n92165 , n42238 );
and ( n92166 , n92165 , n31922 );
and ( n92167 , n53243 , n42238 );
or ( n92168 , n92166 , n92167 );
and ( n92169 , n92164 , n92168 );
and ( n92170 , n53243 , n42247 );
or ( n92171 , n92169 , n92170 );
and ( n92172 , n92163 , n92171 );
not ( n92173 , n42273 );
not ( n92174 , n42276 );
and ( n92175 , n92174 , n92171 );
and ( n92176 , n53269 , n42276 );
or ( n92177 , n92175 , n92176 );
and ( n92178 , n92173 , n92177 );
and ( n92179 , n53277 , n42273 );
or ( n92180 , n92178 , n92179 );
and ( n92181 , n92180 , n32475 );
or ( n92182 , n92172 , n92181 );
and ( n92183 , n92182 , n32486 );
and ( n92184 , n31922 , n41278 );
or ( n92185 , C0 , n92153 , n92162 , n92183 , n92184 );
buf ( n92186 , n92185 );
buf ( n92187 , n92186 );
buf ( n92188 , n30987 );
buf ( n92189 , n30987 );
buf ( n92190 , n31655 );
or ( n92191 , n37497 , n37499 );
or ( n92192 , n92191 , n37501 );
buf ( n92193 , n92192 );
or ( n92194 , n37496 , n37503 );
or ( n92195 , n92194 , n37505 );
and ( n92196 , n41517 , n92195 );
or ( n92197 , C0 , n92193 , n92196 );
buf ( n92198 , n92197 );
buf ( n92199 , n92198 );
and ( n92200 , n47665 , n50275 );
not ( n92201 , n50278 );
and ( n92202 , n92201 , n47578 );
and ( n92203 , n47665 , n50278 );
or ( n92204 , n92202 , n92203 );
and ( n92205 , n92204 , n32421 );
not ( n92206 , n50002 );
and ( n92207 , n92206 , n47578 );
and ( n92208 , n47665 , n50002 );
or ( n92209 , n92207 , n92208 );
and ( n92210 , n92209 , n32419 );
not ( n92211 , n50289 );
and ( n92212 , n92211 , n47578 );
and ( n92213 , n47665 , n50289 );
or ( n92214 , n92212 , n92213 );
and ( n92215 , n92214 , n32417 );
not ( n92216 , n50008 );
and ( n92217 , n92216 , n47578 );
and ( n92218 , n47665 , n50008 );
or ( n92219 , n92217 , n92218 );
and ( n92220 , n92219 , n32415 );
not ( n92221 , n47331 );
and ( n92222 , n92221 , n47578 );
and ( n92223 , n47610 , n47331 );
or ( n92224 , n92222 , n92223 );
and ( n92225 , n92224 , n32413 );
not ( n92226 , n50067 );
and ( n92227 , n92226 , n47578 );
and ( n92228 , n47610 , n50067 );
or ( n92229 , n92227 , n92228 );
and ( n92230 , n92229 , n32411 );
not ( n92231 , n31728 );
and ( n92232 , n92231 , n47578 );
and ( n92233 , n71180 , n31728 );
or ( n92234 , n92232 , n92233 );
and ( n92235 , n92234 , n32253 );
not ( n92236 , n32283 );
and ( n92237 , n92236 , n47578 );
and ( n92238 , n71191 , n32283 );
or ( n92239 , n92237 , n92238 );
and ( n92240 , n92239 , n32398 );
and ( n92241 , n47715 , n50334 );
or ( n92242 , n92200 , n92205 , n92210 , n92215 , n92220 , n92225 , n92230 , n92235 , n92240 , n92241 );
and ( n92243 , n92242 , n32456 );
and ( n92244 , n37563 , n32489 );
and ( n92245 , n47578 , n50345 );
or ( n92246 , C0 , n92243 , n92244 , n92245 );
buf ( n92247 , n92246 );
buf ( n92248 , n92247 );
buf ( n92249 , n30987 );
and ( n92250 , n49064 , n48639 );
not ( n92251 , n48642 );
and ( n92252 , n92251 , n48589 );
and ( n92253 , n49064 , n48642 );
or ( n92254 , n92252 , n92253 );
and ( n92255 , n92254 , n32890 );
not ( n92256 , n48648 );
and ( n92257 , n92256 , n48589 );
and ( n92258 , n49064 , n48648 );
or ( n92259 , n92257 , n92258 );
and ( n92260 , n92259 , n32924 );
not ( n92261 , n48654 );
and ( n92262 , n92261 , n48589 );
and ( n92263 , n49064 , n48654 );
or ( n92264 , n92262 , n92263 );
and ( n92265 , n92264 , n33038 );
not ( n92266 , n48660 );
and ( n92267 , n92266 , n48589 );
and ( n92268 , n49064 , n48660 );
or ( n92269 , n92267 , n92268 );
and ( n92270 , n92269 , n33172 );
not ( n92271 , n41576 );
and ( n92272 , n92271 , n48589 );
and ( n92273 , n48774 , n41576 );
or ( n92274 , n92272 , n92273 );
and ( n92275 , n92274 , n33189 );
not ( n92276 , n48730 );
and ( n92277 , n92276 , n48589 );
and ( n92278 , n48774 , n48730 );
or ( n92279 , n92277 , n92278 );
and ( n92280 , n92279 , n33187 );
not ( n92281 , n48765 );
and ( n92282 , n92281 , n48589 );
and ( n92283 , n77459 , n48765 );
or ( n92284 , n92282 , n92283 );
and ( n92285 , n92284 , n33180 );
not ( n92286 , n49054 );
and ( n92287 , n92286 , n48589 );
and ( n92288 , n77470 , n49054 );
or ( n92289 , n92287 , n92288 );
and ( n92290 , n92289 , n33178 );
and ( n92291 , n49173 , n49275 );
or ( n92292 , n92250 , n92255 , n92260 , n92265 , n92270 , n92275 , n92280 , n92285 , n92290 , n92291 );
and ( n92293 , n92292 , n33208 );
and ( n92294 , n32982 , n35056 );
and ( n92295 , n48589 , n49286 );
or ( n92296 , C0 , n92293 , n92294 , n92295 );
buf ( n92297 , n92296 );
buf ( n92298 , n92297 );
buf ( n92299 , n30987 );
buf ( n92300 , n30987 );
buf ( n92301 , n31655 );
buf ( n92302 , n31655 );
and ( n92303 , n33767 , n48455 );
not ( n92304 , n48457 );
and ( n92305 , n92304 , n33432 );
and ( n92306 , n33767 , n48457 );
or ( n92307 , n92305 , n92306 );
and ( n92308 , n92307 , n31373 );
not ( n92309 , n44807 );
and ( n92310 , n92309 , n33432 );
and ( n92311 , n33767 , n44807 );
or ( n92312 , n92310 , n92311 );
and ( n92313 , n92312 , n31408 );
not ( n92314 , n48468 );
and ( n92315 , n92314 , n33432 );
and ( n92316 , n33767 , n48468 );
or ( n92317 , n92315 , n92316 );
and ( n92318 , n92317 , n31468 );
not ( n92319 , n44817 );
and ( n92320 , n92319 , n33432 );
and ( n92321 , n33767 , n44817 );
or ( n92322 , n92320 , n92321 );
and ( n92323 , n92322 , n31521 );
not ( n92324 , n39979 );
and ( n92325 , n92324 , n33432 );
and ( n92326 , n33474 , n39979 );
or ( n92327 , n92325 , n92326 );
and ( n92328 , n92327 , n31538 );
not ( n92329 , n45059 );
and ( n92330 , n92329 , n33432 );
and ( n92331 , n33474 , n45059 );
or ( n92332 , n92330 , n92331 );
and ( n92333 , n92332 , n31536 );
not ( n92334 , n33419 );
and ( n92335 , n92334 , n33432 );
and ( n92336 , n91642 , n33419 );
or ( n92337 , n92335 , n92336 );
and ( n92338 , n92337 , n31529 );
not ( n92339 , n33734 );
and ( n92340 , n92339 , n33432 );
and ( n92341 , n91653 , n33734 );
or ( n92342 , n92340 , n92341 );
and ( n92343 , n92342 , n31527 );
and ( n92344 , n33852 , n48513 );
or ( n92345 , n92303 , n92308 , n92313 , n92318 , n92323 , n92328 , n92333 , n92338 , n92343 , n92344 );
and ( n92346 , n92345 , n31557 );
and ( n92347 , n34004 , n33973 );
and ( n92348 , n33432 , n48524 );
or ( n92349 , C0 , n92346 , n92347 , n92348 );
buf ( n92350 , n92349 );
buf ( n92351 , n92350 );
buf ( n92352 , n31655 );
buf ( n92353 , n30987 );
not ( n92354 , n35278 );
and ( n92355 , n92354 , n80196 );
and ( n92356 , n80208 , n35278 );
or ( n92357 , n92355 , n92356 );
and ( n92358 , n92357 , n32417 );
not ( n92359 , n50008 );
and ( n92360 , n92359 , n80196 );
and ( n92361 , n75150 , n50008 );
or ( n92362 , n92360 , n92361 );
and ( n92363 , n92362 , n32415 );
and ( n92364 , n80196 , n48133 );
or ( n92365 , n92358 , n92363 , n92364 );
and ( n92366 , n92365 , n32456 );
and ( n92367 , n80196 , n47409 );
or ( n92368 , C0 , n92366 , n92367 );
buf ( n92369 , n92368 );
buf ( n92370 , n92369 );
xor ( n92371 , n33129 , n41542 );
and ( n92372 , n92371 , n33201 );
not ( n92373 , n41576 );
and ( n92374 , n92373 , n33129 );
buf ( n92375 , n32720 );
and ( n92376 , n92375 , n41576 );
or ( n92377 , n92374 , n92376 );
and ( n92378 , n92377 , n33189 );
and ( n92379 , n33129 , n41592 );
or ( n92380 , n92372 , n92378 , n92379 );
and ( n92381 , n92380 , n33208 );
and ( n92382 , n33129 , n39805 );
or ( n92383 , C0 , n92381 , n92382 );
buf ( n92384 , n92383 );
buf ( n92385 , n92384 );
buf ( n92386 , n31655 );
buf ( n92387 , n30987 );
buf ( n92388 , n30987 );
buf ( n92389 , n31655 );
not ( n92390 , n41532 );
and ( n92391 , n92390 , n34234 );
and ( n92392 , n50837 , n41532 );
or ( n92393 , n92391 , n92392 );
buf ( n92394 , n92393 );
buf ( n92395 , n92394 );
not ( n92396 , n52719 );
not ( n92397 , n92396 );
not ( n92398 , n92397 );
and ( n92399 , n92398 , n90343 );
and ( n92400 , n42739 , n62377 );
or ( n92401 , n92399 , C0 , n92400 );
buf ( n92402 , n92401 );
buf ( n92403 , n92402 );
buf ( n92404 , n30987 );
buf ( n92405 , n31655 );
buf ( n92406 , n30987 );
buf ( n92407 , n31655 );
buf ( n92408 , n30987 );
not ( n92409 , n43755 );
and ( n92410 , n92409 , n43275 );
xor ( n92411 , n43763 , n43765 );
and ( n92412 , n92411 , n43755 );
or ( n92413 , n92410 , n92412 );
and ( n92414 , n92413 , n43774 );
not ( n92415 , n44663 );
and ( n92416 , n92415 , n44187 );
xor ( n92417 , n44671 , n44673 );
and ( n92418 , n92417 , n44663 );
or ( n92419 , n92416 , n92418 );
and ( n92420 , n92419 , n44682 );
and ( n92421 , n35546 , n44695 );
or ( n92422 , n92414 , n92420 , n92421 );
buf ( n92423 , n92422 );
buf ( n92424 , n92423 );
buf ( n92425 , n30987 );
buf ( n92426 , n31655 );
buf ( n92427 , n31655 );
buf ( n92428 , n31655 );
not ( n92429 , n46356 );
and ( n92430 , n92429 , n31173 );
not ( n92431 , n63024 );
and ( n92432 , n92431 , n31173 );
and ( n92433 , n31205 , n63024 );
or ( n92434 , n92432 , n92433 );
and ( n92435 , n92434 , n46356 );
or ( n92436 , n92430 , n92435 );
and ( n92437 , n92436 , n31649 );
not ( n92438 , n63032 );
not ( n92439 , n63024 );
and ( n92440 , n92439 , n31173 );
and ( n92441 , n50125 , n63024 );
or ( n92442 , n92440 , n92441 );
and ( n92443 , n92438 , n92442 );
and ( n92444 , n50125 , n63032 );
or ( n92445 , n92443 , n92444 );
and ( n92446 , n92445 , n31643 );
not ( n92447 , n31452 );
not ( n92448 , n63032 );
not ( n92449 , n63024 );
and ( n92450 , n92449 , n31173 );
and ( n92451 , n50125 , n63024 );
or ( n92452 , n92450 , n92451 );
and ( n92453 , n92448 , n92452 );
and ( n92454 , n50125 , n63032 );
or ( n92455 , n92453 , n92454 );
and ( n92456 , n92447 , n92455 );
not ( n92457 , n63052 );
not ( n92458 , n63054 );
and ( n92459 , n92458 , n92455 );
and ( n92460 , n50151 , n63054 );
or ( n92461 , n92459 , n92460 );
and ( n92462 , n92457 , n92461 );
and ( n92463 , n50159 , n63052 );
or ( n92464 , n92462 , n92463 );
and ( n92465 , n92464 , n31452 );
or ( n92466 , n92456 , n92465 );
and ( n92467 , n92466 , n31638 );
and ( n92468 , n31173 , n47277 );
or ( n92469 , C0 , n92437 , n92446 , n92467 , n92468 );
buf ( n92470 , n92469 );
buf ( n92471 , n92470 );
buf ( n92472 , n30987 );
not ( n92473 , n35278 );
and ( n92474 , n92473 , n55447 );
and ( n92475 , n55455 , n35278 );
or ( n92476 , n92474 , n92475 );
and ( n92477 , n92476 , n32417 );
not ( n92478 , n47912 );
and ( n92479 , n92478 , n55447 );
and ( n92480 , n91074 , n47912 );
or ( n92481 , n92479 , n92480 );
and ( n92482 , n92481 , n32415 );
and ( n92483 , n55447 , n48133 );
or ( n92484 , n92477 , n92482 , n92483 );
and ( n92485 , n92484 , n32456 );
and ( n92486 , n55447 , n47409 );
or ( n92487 , C0 , n92485 , n92486 );
buf ( n92488 , n92487 );
buf ( n92489 , n92488 );
buf ( n92490 , n31655 );
not ( n92491 , n31437 );
and ( n92492 , n92491 , n54004 );
and ( n92493 , n92070 , n31437 );
or ( n92494 , n92492 , n92493 );
and ( n92495 , n92494 , n31468 );
not ( n92496 , n41837 );
and ( n92497 , n92496 , n54004 );
and ( n92498 , n54010 , n41837 );
or ( n92499 , n92497 , n92498 );
and ( n92500 , n92499 , n31521 );
and ( n92501 , n54004 , n42158 );
or ( n92502 , n92495 , n92500 , n92501 );
and ( n92503 , n92502 , n31557 );
and ( n92504 , n54004 , n40154 );
or ( n92505 , C0 , n92503 , n92504 );
buf ( n92506 , n92505 );
buf ( n92507 , n92506 );
not ( n92508 , n40163 );
and ( n92509 , n92508 , n31931 );
not ( n92510 , n56988 );
and ( n92511 , n92510 , n31931 );
and ( n92512 , n32183 , n56988 );
or ( n92513 , n92511 , n92512 );
and ( n92514 , n92513 , n40163 );
or ( n92515 , n92509 , n92514 );
and ( n92516 , n92515 , n32498 );
not ( n92517 , n56996 );
not ( n92518 , n56988 );
and ( n92519 , n92518 , n31931 );
and ( n92520 , n45178 , n56988 );
or ( n92521 , n92519 , n92520 );
and ( n92522 , n92517 , n92521 );
and ( n92523 , n45178 , n56996 );
or ( n92524 , n92522 , n92523 );
and ( n92525 , n92524 , n32473 );
not ( n92526 , n32475 );
not ( n92527 , n56996 );
not ( n92528 , n56988 );
and ( n92529 , n92528 , n31931 );
and ( n92530 , n45178 , n56988 );
or ( n92531 , n92529 , n92530 );
and ( n92532 , n92527 , n92531 );
and ( n92533 , n45178 , n56996 );
or ( n92534 , n92532 , n92533 );
and ( n92535 , n92526 , n92534 );
not ( n92536 , n57016 );
not ( n92537 , n57018 );
and ( n92538 , n92537 , n92534 );
and ( n92539 , n45206 , n57018 );
or ( n92540 , n92538 , n92539 );
and ( n92541 , n92536 , n92540 );
and ( n92542 , n45214 , n57016 );
or ( n92543 , n92541 , n92542 );
and ( n92544 , n92543 , n32475 );
or ( n92545 , n92535 , n92544 );
and ( n92546 , n92545 , n32486 );
and ( n92547 , n31931 , n41278 );
or ( n92548 , C0 , n92516 , n92525 , n92546 , n92547 );
buf ( n92549 , n92548 );
buf ( n92550 , n92549 );
buf ( n92551 , n30987 );
buf ( n92552 , n31655 );
and ( n92553 , n33766 , n48455 );
not ( n92554 , n48457 );
and ( n92555 , n92554 , n33431 );
and ( n92556 , n33766 , n48457 );
or ( n92557 , n92555 , n92556 );
and ( n92558 , n92557 , n31373 );
not ( n92559 , n44807 );
and ( n92560 , n92559 , n33431 );
and ( n92561 , n33766 , n44807 );
or ( n92562 , n92560 , n92561 );
and ( n92563 , n92562 , n31408 );
not ( n92564 , n48468 );
and ( n92565 , n92564 , n33431 );
and ( n92566 , n33766 , n48468 );
or ( n92567 , n92565 , n92566 );
and ( n92568 , n92567 , n31468 );
not ( n92569 , n44817 );
and ( n92570 , n92569 , n33431 );
and ( n92571 , n33766 , n44817 );
or ( n92572 , n92570 , n92571 );
and ( n92573 , n92572 , n31521 );
not ( n92574 , n39979 );
and ( n92575 , n92574 , n33431 );
and ( n92576 , n33473 , n39979 );
or ( n92577 , n92575 , n92576 );
and ( n92578 , n92577 , n31538 );
not ( n92579 , n45059 );
and ( n92580 , n92579 , n33431 );
and ( n92581 , n33473 , n45059 );
or ( n92582 , n92580 , n92581 );
and ( n92583 , n92582 , n31536 );
not ( n92584 , n33419 );
and ( n92585 , n92584 , n33431 );
and ( n92586 , n71429 , n33419 );
or ( n92587 , n92585 , n92586 );
and ( n92588 , n92587 , n31529 );
not ( n92589 , n33734 );
and ( n92590 , n92589 , n33431 );
and ( n92591 , n71440 , n33734 );
or ( n92592 , n92590 , n92591 );
and ( n92593 , n92592 , n31527 );
and ( n92594 , n33851 , n48513 );
or ( n92595 , n92553 , n92558 , n92563 , n92568 , n92573 , n92578 , n92583 , n92588 , n92593 , n92594 );
and ( n92596 , n92595 , n31557 );
and ( n92597 , n34003 , n33973 );
and ( n92598 , n33431 , n48524 );
or ( n92599 , C0 , n92596 , n92597 , n92598 );
buf ( n92600 , n92599 );
buf ( n92601 , n92600 );
buf ( n92602 , n30987 );
not ( n92603 , n35278 );
and ( n92604 , n92603 , n82377 );
and ( n92605 , n82390 , n35278 );
or ( n92606 , n92604 , n92605 );
and ( n92607 , n92606 , n32417 );
not ( n92608 , n50008 );
and ( n92609 , n92608 , n82377 );
and ( n92610 , n80579 , n50008 );
or ( n92611 , n92609 , n92610 );
and ( n92612 , n92611 , n32415 );
and ( n92613 , n82377 , n48133 );
or ( n92614 , n92607 , n92612 , n92613 );
and ( n92615 , n92614 , n32456 );
and ( n92616 , n82377 , n47409 );
or ( n92617 , C0 , n92615 , n92616 );
buf ( n92618 , n92617 );
buf ( n92619 , n92618 );
buf ( n92620 , n31655 );
buf ( n92621 , n53756 );
buf ( n92622 , n92621 );
and ( n92623 , n92622 , n53793 );
buf ( n92624 , n53756 );
buf ( n92625 , n53832 );
or ( n92626 , C0 , n92624 , C0 , C0 , n92625 );
and ( n92627 , n92626 , n53828 );
buf ( n92628 , n53756 );
buf ( n92629 , n67277 );
buf ( n92630 , n53832 );
or ( n92631 , C0 , n92628 , C0 , n92629 , n92630 );
and ( n92632 , n92631 , n53864 );
or ( n92633 , C0 , n92623 , n92627 , n92632 );
buf ( n92634 , n92633 );
buf ( n92635 , n92634 );
not ( n92636 , n40163 );
and ( n92637 , n92636 , n32048 );
not ( n92638 , n52903 );
and ( n92639 , n92638 , n32048 );
and ( n92640 , n32130 , n52903 );
or ( n92641 , n92639 , n92640 );
and ( n92642 , n92641 , n40163 );
or ( n92643 , n92637 , n92642 );
and ( n92644 , n92643 , n32498 );
not ( n92645 , n52911 );
not ( n92646 , n52903 );
and ( n92647 , n92646 , n32048 );
and ( n92648 , n45833 , n52903 );
or ( n92649 , n92647 , n92648 );
and ( n92650 , n92645 , n92649 );
and ( n92651 , n45833 , n52911 );
or ( n92652 , n92650 , n92651 );
and ( n92653 , n92652 , n32473 );
not ( n92654 , n32475 );
not ( n92655 , n52911 );
not ( n92656 , n52903 );
and ( n92657 , n92656 , n32048 );
and ( n92658 , n45833 , n52903 );
or ( n92659 , n92657 , n92658 );
and ( n92660 , n92655 , n92659 );
and ( n92661 , n45833 , n52911 );
or ( n92662 , n92660 , n92661 );
and ( n92663 , n92654 , n92662 );
not ( n92664 , n52931 );
not ( n92665 , n52933 );
and ( n92666 , n92665 , n92662 );
and ( n92667 , n45857 , n52933 );
or ( n92668 , n92666 , n92667 );
and ( n92669 , n92664 , n92668 );
and ( n92670 , n45865 , n52931 );
or ( n92671 , n92669 , n92670 );
and ( n92672 , n92671 , n32475 );
or ( n92673 , n92663 , n92672 );
and ( n92674 , n92673 , n32486 );
and ( n92675 , n32048 , n41278 );
or ( n92676 , C0 , n92644 , n92653 , n92674 , n92675 );
buf ( n92677 , n92676 );
buf ( n92678 , n92677 );
buf ( n92679 , n30987 );
buf ( n92680 , n30987 );
buf ( n92681 , n30987 );
buf ( n92682 , n30987 );
not ( n92683 , n43755 );
and ( n92684 , n92683 , n43496 );
xor ( n92685 , n52313 , n52316 );
and ( n92686 , n92685 , n43755 );
or ( n92687 , n92684 , n92686 );
and ( n92688 , n92687 , n43774 );
not ( n92689 , n44663 );
and ( n92690 , n92689 , n44408 );
xor ( n92691 , n52351 , n52354 );
and ( n92692 , n92691 , n44663 );
or ( n92693 , n92690 , n92692 );
and ( n92694 , n92693 , n44682 );
buf ( n92695 , RI15b45708_234);
and ( n92696 , n92695 , n44695 );
or ( n92697 , n92688 , n92694 , n92696 );
buf ( n92698 , n92697 );
buf ( n92699 , n92698 );
buf ( n92700 , n31655 );
buf ( n92701 , n31655 );
buf ( n92702 , n31655 );
buf ( n92703 , n31655 );
not ( n92704 , n33419 );
and ( n92705 , n92704 , n31582 );
xor ( n92706 , n33476 , n33689 );
and ( n92707 , n92706 , n33419 );
or ( n92708 , n92705 , n92707 );
and ( n92709 , n92708 , n31529 );
not ( n92710 , n33734 );
and ( n92711 , n92710 , n31582 );
not ( n92712 , n33533 );
xor ( n92713 , n33769 , n33807 );
and ( n92714 , n92712 , n92713 );
xnor ( n92715 , n33854 , n33909 );
and ( n92716 , n92715 , n33533 );
or ( n92717 , n92714 , n92716 );
and ( n92718 , n92717 , n33734 );
or ( n92719 , n92711 , n92718 );
and ( n92720 , n92719 , n31527 );
and ( n92721 , n31582 , n33942 );
or ( n92722 , n92709 , n92720 , n92721 );
and ( n92723 , n92722 , n31557 );
and ( n92724 , n34109 , n31643 );
not ( n92725 , n31452 );
and ( n92726 , n92725 , n34109 );
xor ( n92727 , n31582 , n33955 );
and ( n92728 , n92727 , n31452 );
or ( n92729 , n92726 , n92728 );
and ( n92730 , n92729 , n31638 );
and ( n92731 , n34006 , n33973 );
and ( n92732 , n31582 , n33978 );
or ( n92733 , C0 , n92723 , n92724 , n92730 , n92731 , n92732 );
buf ( n92734 , n92733 );
buf ( n92735 , n92734 );
and ( n92736 , n31562 , n31007 );
not ( n92737 , n31077 );
and ( n92738 , n92737 , n35388 );
buf ( n92739 , n92738 );
and ( n92740 , n92739 , n31373 );
not ( n92741 , n31402 );
and ( n92742 , n92741 , n35388 );
buf ( n92743 , n92742 );
and ( n92744 , n92743 , n31408 );
not ( n92745 , n31437 );
and ( n92746 , n92745 , n35388 );
not ( n92747 , n31455 );
and ( n92748 , n92747 , n35425 );
xor ( n92749 , n35388 , n35410 );
and ( n92750 , n92749 , n31455 );
or ( n92751 , n92748 , n92750 );
and ( n92752 , n92751 , n31437 );
or ( n92753 , n92746 , n92752 );
and ( n92754 , n92753 , n31468 );
not ( n92755 , n31497 );
and ( n92756 , n92755 , n35388 );
not ( n92757 , n31454 );
not ( n92758 , n31501 );
and ( n92759 , n92758 , n35425 );
xor ( n92760 , n35426 , n35460 );
and ( n92761 , n92760 , n31501 );
or ( n92762 , n92759 , n92761 );
and ( n92763 , n92757 , n92762 );
and ( n92764 , n92749 , n31454 );
or ( n92765 , n92763 , n92764 );
and ( n92766 , n92765 , n31497 );
or ( n92767 , n92756 , n92766 );
and ( n92768 , n92767 , n31521 );
and ( n92769 , n35388 , n31553 );
or ( n92770 , n92740 , n92744 , n92754 , n92768 , n92769 );
and ( n92771 , n92770 , n31557 );
not ( n92772 , n31452 );
not ( n92773 , n31619 );
and ( n92774 , n92773 , n35480 );
xor ( n92775 , n35481 , n35514 );
and ( n92776 , n92775 , n31619 );
or ( n92777 , n92774 , n92776 );
and ( n92778 , n92772 , n92777 );
and ( n92779 , n35388 , n31452 );
or ( n92780 , n92778 , n92779 );
and ( n92781 , n92780 , n31638 );
and ( n92782 , n35388 , n31650 );
or ( n92783 , C0 , n92736 , n92771 , n92781 , C0 , n92782 );
buf ( n92784 , n92783 );
buf ( n92785 , n92784 );
buf ( n92786 , n30987 );
buf ( n92787 , n30987 );
buf ( n92788 , n31655 );
not ( n92789 , n46356 );
and ( n92790 , n92789 , n31276 );
not ( n92791 , n47831 );
and ( n92792 , n92791 , n31276 );
and ( n92793 , n31306 , n47831 );
or ( n92794 , n92792 , n92793 );
and ( n92795 , n92794 , n46356 );
or ( n92796 , n92790 , n92795 );
and ( n92797 , n92796 , n31649 );
not ( n92798 , n47839 );
not ( n92799 , n47831 );
and ( n92800 , n92799 , n31276 );
and ( n92801 , n58061 , n47831 );
or ( n92802 , n92800 , n92801 );
and ( n92803 , n92798 , n92802 );
and ( n92804 , n58061 , n47839 );
or ( n92805 , n92803 , n92804 );
and ( n92806 , n92805 , n31643 );
not ( n92807 , n31452 );
not ( n92808 , n47839 );
not ( n92809 , n47831 );
and ( n92810 , n92809 , n31276 );
and ( n92811 , n58061 , n47831 );
or ( n92812 , n92810 , n92811 );
and ( n92813 , n92808 , n92812 );
and ( n92814 , n58061 , n47839 );
or ( n92815 , n92813 , n92814 );
and ( n92816 , n92807 , n92815 );
not ( n92817 , n47866 );
not ( n92818 , n47868 );
and ( n92819 , n92818 , n92815 );
and ( n92820 , n58085 , n47868 );
or ( n92821 , n92819 , n92820 );
and ( n92822 , n92817 , n92821 );
and ( n92823 , n58093 , n47866 );
or ( n92824 , n92822 , n92823 );
and ( n92825 , n92824 , n31452 );
or ( n92826 , n92816 , n92825 );
and ( n92827 , n92826 , n31638 );
and ( n92828 , n31276 , n47277 );
or ( n92829 , C0 , n92797 , n92806 , n92827 , n92828 );
buf ( n92830 , n92829 );
buf ( n92831 , n92830 );
buf ( n92832 , n30987 );
not ( n92833 , n35278 );
and ( n92834 , n92833 , n61466 );
and ( n92835 , n86773 , n35278 );
or ( n92836 , n92834 , n92835 );
and ( n92837 , n92836 , n32417 );
not ( n92838 , n47912 );
and ( n92839 , n92838 , n61466 );
and ( n92840 , n61472 , n47912 );
or ( n92841 , n92839 , n92840 );
and ( n92842 , n92841 , n32415 );
and ( n92843 , n61466 , n48133 );
or ( n92844 , n92837 , n92842 , n92843 );
and ( n92845 , n92844 , n32456 );
and ( n92846 , n61466 , n47409 );
or ( n92847 , C0 , n92845 , n92846 );
buf ( n92848 , n92847 );
buf ( n92849 , n92848 );
and ( n92850 , n33768 , n48455 );
not ( n92851 , n48457 );
and ( n92852 , n92851 , n33433 );
and ( n92853 , n33768 , n48457 );
or ( n92854 , n92852 , n92853 );
and ( n92855 , n92854 , n31373 );
not ( n92856 , n44807 );
and ( n92857 , n92856 , n33433 );
and ( n92858 , n33768 , n44807 );
or ( n92859 , n92857 , n92858 );
and ( n92860 , n92859 , n31408 );
not ( n92861 , n48468 );
and ( n92862 , n92861 , n33433 );
and ( n92863 , n33768 , n48468 );
or ( n92864 , n92862 , n92863 );
and ( n92865 , n92864 , n31468 );
not ( n92866 , n44817 );
and ( n92867 , n92866 , n33433 );
and ( n92868 , n33768 , n44817 );
or ( n92869 , n92867 , n92868 );
and ( n92870 , n92869 , n31521 );
not ( n92871 , n39979 );
and ( n92872 , n92871 , n33433 );
and ( n92873 , n33475 , n39979 );
or ( n92874 , n92872 , n92873 );
and ( n92875 , n92874 , n31538 );
not ( n92876 , n45059 );
and ( n92877 , n92876 , n33433 );
and ( n92878 , n33475 , n45059 );
or ( n92879 , n92877 , n92878 );
and ( n92880 , n92879 , n31536 );
not ( n92881 , n33419 );
and ( n92882 , n92881 , n33433 );
and ( n92883 , n70627 , n33419 );
or ( n92884 , n92882 , n92883 );
and ( n92885 , n92884 , n31529 );
not ( n92886 , n33734 );
and ( n92887 , n92886 , n33433 );
and ( n92888 , n70638 , n33734 );
or ( n92889 , n92887 , n92888 );
and ( n92890 , n92889 , n31527 );
and ( n92891 , n33853 , n48513 );
or ( n92892 , n92850 , n92855 , n92860 , n92865 , n92870 , n92875 , n92880 , n92885 , n92890 , n92891 );
and ( n92893 , n92892 , n31557 );
and ( n92894 , n34005 , n33973 );
and ( n92895 , n33433 , n48524 );
or ( n92896 , C0 , n92893 , n92894 , n92895 );
buf ( n92897 , n92896 );
buf ( n92898 , n92897 );
buf ( n92899 , n31655 );
buf ( n92900 , n30987 );
not ( n92901 , n35278 );
and ( n92902 , n92901 , n78755 );
and ( n92903 , n78768 , n35278 );
or ( n92904 , n92902 , n92903 );
and ( n92905 , n92904 , n32417 );
not ( n92906 , n50008 );
and ( n92907 , n92906 , n78755 );
and ( n92908 , n71746 , n50008 );
or ( n92909 , n92907 , n92908 );
and ( n92910 , n92909 , n32415 );
and ( n92911 , n78755 , n48133 );
or ( n92912 , n92905 , n92910 , n92911 );
and ( n92913 , n92912 , n32456 );
and ( n92914 , n78755 , n47409 );
or ( n92915 , C0 , n92913 , n92914 );
buf ( n92916 , n92915 );
buf ( n92917 , n92916 );
buf ( n92918 , n31655 );
buf ( n92919 , RI15b54528_742);
and ( n92920 , n92919 , n58921 );
and ( n92921 , n41529 , n37506 );
or ( n92922 , n92920 , n92921 );
buf ( n92923 , n92922 );
buf ( n92924 , n92923 );
buf ( n92925 , n30987 );
not ( n92926 , n38443 );
and ( n92927 , n92926 , n37997 );
xor ( n92928 , n53482 , n53487 );
and ( n92929 , n92928 , n38443 );
or ( n92930 , n92927 , n92929 );
and ( n92931 , n92930 , n38450 );
not ( n92932 , n39339 );
and ( n92933 , n92932 , n38897 );
xor ( n92934 , n53538 , n53543 );
and ( n92935 , n92934 , n39339 );
or ( n92936 , n92933 , n92935 );
and ( n92937 , n92936 , n39346 );
and ( n92938 , n40202 , n39359 );
or ( n92939 , n92931 , n92937 , n92938 );
buf ( n92940 , n92939 );
buf ( n92941 , n92940 );
buf ( n92942 , n31655 );
not ( n92943 , n31437 );
and ( n92944 , n92943 , n84892 );
and ( n92945 , n90630 , n31437 );
or ( n92946 , n92944 , n92945 );
and ( n92947 , n92946 , n31468 );
not ( n92948 , n41837 );
and ( n92949 , n92948 , n84892 );
and ( n92950 , n84898 , n41837 );
or ( n92951 , n92949 , n92950 );
and ( n92952 , n92951 , n31521 );
and ( n92953 , n84892 , n42158 );
or ( n92954 , n92947 , n92952 , n92953 );
and ( n92955 , n92954 , n31557 );
and ( n92956 , n84892 , n40154 );
or ( n92957 , C0 , n92955 , n92956 );
buf ( n92958 , n92957 );
buf ( n92959 , n92958 );
not ( n92960 , n40163 );
and ( n92961 , n92960 , n31863 );
not ( n92962 , n42171 );
and ( n92963 , n92962 , n31863 );
and ( n92964 , n32218 , n42171 );
or ( n92965 , n92963 , n92964 );
and ( n92966 , n92965 , n40163 );
or ( n92967 , n92961 , n92966 );
and ( n92968 , n92967 , n32498 );
not ( n92969 , n42180 );
not ( n92970 , n42171 );
and ( n92971 , n92970 , n31863 );
and ( n92972 , n42255 , n42171 );
or ( n92973 , n92971 , n92972 );
and ( n92974 , n92969 , n92973 );
and ( n92975 , n42255 , n42180 );
or ( n92976 , n92974 , n92975 );
and ( n92977 , n92976 , n32473 );
not ( n92978 , n32475 );
not ( n92979 , n42180 );
not ( n92980 , n42171 );
and ( n92981 , n92980 , n31863 );
and ( n92982 , n42255 , n42171 );
or ( n92983 , n92981 , n92982 );
and ( n92984 , n92979 , n92983 );
and ( n92985 , n42255 , n42180 );
or ( n92986 , n92984 , n92985 );
and ( n92987 , n92978 , n92986 );
not ( n92988 , n42206 );
not ( n92989 , n42209 );
and ( n92990 , n92989 , n92986 );
and ( n92991 , n42283 , n42209 );
or ( n92992 , n92990 , n92991 );
and ( n92993 , n92988 , n92992 );
and ( n92994 , n42291 , n42206 );
or ( n92995 , n92993 , n92994 );
and ( n92996 , n92995 , n32475 );
or ( n92997 , n92987 , n92996 );
and ( n92998 , n92997 , n32486 );
and ( n92999 , n31863 , n41278 );
or ( n93000 , C0 , n92968 , n92977 , n92998 , n92999 );
buf ( n93001 , n93000 );
buf ( n93002 , n93001 );
buf ( n93003 , n30987 );
buf ( n93004 , n30987 );
buf ( n93005 , n30987 );
not ( n93006 , n34150 );
and ( n93007 , n93006 , n32611 );
not ( n93008 , n60126 );
and ( n93009 , n93008 , n32611 );
and ( n93010 , n32655 , n60126 );
or ( n93011 , n93009 , n93010 );
and ( n93012 , n93011 , n34150 );
or ( n93013 , n93007 , n93012 );
and ( n93014 , n93013 , n33381 );
not ( n93015 , n60134 );
not ( n93016 , n60126 );
and ( n93017 , n93016 , n32611 );
and ( n93018 , n56044 , n60126 );
or ( n93019 , n93017 , n93018 );
and ( n93020 , n93015 , n93019 );
and ( n93021 , n56044 , n60134 );
or ( n93022 , n93020 , n93021 );
and ( n93023 , n93022 , n33375 );
not ( n93024 , n32968 );
not ( n93025 , n60134 );
not ( n93026 , n60126 );
and ( n93027 , n93026 , n32611 );
and ( n93028 , n56044 , n60126 );
or ( n93029 , n93027 , n93028 );
and ( n93030 , n93025 , n93029 );
and ( n93031 , n56044 , n60134 );
or ( n93032 , n93030 , n93031 );
and ( n93033 , n93024 , n93032 );
not ( n93034 , n60154 );
not ( n93035 , n60156 );
and ( n93036 , n93035 , n93032 );
and ( n93037 , n56068 , n60156 );
or ( n93038 , n93036 , n93037 );
and ( n93039 , n93034 , n93038 );
and ( n93040 , n56076 , n60154 );
or ( n93041 , n93039 , n93040 );
and ( n93042 , n93041 , n32968 );
or ( n93043 , n93033 , n93042 );
and ( n93044 , n93043 , n33370 );
and ( n93045 , n32611 , n35062 );
or ( n93046 , C0 , n93014 , n93023 , n93044 , n93045 );
buf ( n93047 , n93046 );
buf ( n93048 , n93047 );
buf ( n93049 , n31655 );
buf ( n93050 , n31655 );
buf ( n93051 , n30987 );
buf ( n93052 , n88433 );
buf ( n93053 , n31655 );
not ( n93054 , n48765 );
and ( n93055 , n93054 , n33224 );
and ( n93056 , n89647 , n48765 );
or ( n93057 , n93055 , n93056 );
and ( n93058 , n93057 , n33180 );
not ( n93059 , n49054 );
and ( n93060 , n93059 , n33224 );
and ( n93061 , n89658 , n49054 );
or ( n93062 , n93060 , n93061 );
and ( n93063 , n93062 , n33178 );
and ( n93064 , n33224 , n49774 );
or ( n93065 , n93058 , n93063 , n93064 );
and ( n93066 , n93065 , n33208 );
and ( n93067 , n33299 , n33375 );
not ( n93068 , n32968 );
and ( n93069 , n93068 , n33299 );
xor ( n93070 , n33224 , n53905 );
and ( n93071 , n93070 , n32968 );
or ( n93072 , n93069 , n93071 );
and ( n93073 , n93072 , n33370 );
and ( n93074 , n32987 , n35056 );
and ( n93075 , n33224 , n49794 );
or ( n93076 , C0 , n93066 , n93067 , n93073 , n93074 , n93075 );
buf ( n93077 , n93076 );
buf ( n93078 , n93077 );
buf ( n93079 , n30987 );
buf ( n93080 , n31655 );
and ( n93081 , n46026 , n32500 );
not ( n93082 , n35211 );
and ( n93083 , n93082 , n37549 );
buf ( n93084 , n93083 );
and ( n93085 , n93084 , n32421 );
not ( n93086 , n35245 );
and ( n93087 , n93086 , n37549 );
buf ( n93088 , n93087 );
and ( n93089 , n93088 , n32419 );
not ( n93090 , n35278 );
and ( n93091 , n93090 , n37549 );
not ( n93092 , n35295 );
and ( n93093 , n93092 , n49579 );
xor ( n93094 , n37549 , n49541 );
and ( n93095 , n93094 , n35295 );
or ( n93096 , n93093 , n93095 );
and ( n93097 , n93096 , n35278 );
or ( n93098 , n93091 , n93097 );
and ( n93099 , n93098 , n32417 );
not ( n93100 , n35331 );
and ( n93101 , n93100 , n37549 );
not ( n93102 , n35294 );
not ( n93103 , n45995 );
and ( n93104 , n93103 , n49579 );
xor ( n93105 , n49580 , n49627 );
and ( n93106 , n93105 , n45995 );
or ( n93107 , n93104 , n93106 );
and ( n93108 , n93102 , n93107 );
and ( n93109 , n93094 , n35294 );
or ( n93110 , n93108 , n93109 );
and ( n93111 , n93110 , n35331 );
or ( n93112 , n93101 , n93111 );
and ( n93113 , n93112 , n32415 );
and ( n93114 , n37549 , n35354 );
or ( n93115 , n93085 , n93089 , n93099 , n93113 , n93114 );
and ( n93116 , n93115 , n32456 );
not ( n93117 , n32475 );
not ( n93118 , n46060 );
and ( n93119 , n93118 , n49669 );
xor ( n93120 , n49670 , n49721 );
and ( n93121 , n93120 , n46060 );
or ( n93122 , n93119 , n93121 );
and ( n93123 , n93117 , n93122 );
and ( n93124 , n37549 , n32475 );
or ( n93125 , n93123 , n93124 );
and ( n93126 , n93125 , n32486 );
and ( n93127 , n37549 , n35367 );
or ( n93128 , C0 , n93081 , n93116 , n93126 , C0 , n93127 );
buf ( n93129 , n93128 );
buf ( n93130 , n93129 );
not ( n93131 , n46356 );
and ( n93132 , n93131 , n31098 );
not ( n93133 , n46362 );
and ( n93134 , n93133 , n31098 );
and ( n93135 , n31138 , n46362 );
or ( n93136 , n93134 , n93135 );
and ( n93137 , n93136 , n46356 );
or ( n93138 , n93132 , n93137 );
and ( n93139 , n93138 , n31649 );
not ( n93140 , n46393 );
not ( n93141 , n46362 );
and ( n93142 , n93141 , n31098 );
and ( n93143 , n56920 , n46362 );
or ( n93144 , n93142 , n93143 );
and ( n93145 , n93140 , n93144 );
and ( n93146 , n56920 , n46393 );
or ( n93147 , n93145 , n93146 );
and ( n93148 , n93147 , n31643 );
not ( n93149 , n31452 );
not ( n93150 , n46393 );
not ( n93151 , n46362 );
and ( n93152 , n93151 , n31098 );
and ( n93153 , n56920 , n46362 );
or ( n93154 , n93152 , n93153 );
and ( n93155 , n93150 , n93154 );
and ( n93156 , n56920 , n46393 );
or ( n93157 , n93155 , n93156 );
and ( n93158 , n93149 , n93157 );
not ( n93159 , n46550 );
not ( n93160 , n46554 );
and ( n93161 , n93160 , n93157 );
and ( n93162 , n56946 , n46554 );
or ( n93163 , n93161 , n93162 );
and ( n93164 , n93159 , n93163 );
and ( n93165 , n56954 , n46550 );
or ( n93166 , n93164 , n93165 );
and ( n93167 , n93166 , n31452 );
or ( n93168 , n93158 , n93167 );
and ( n93169 , n93168 , n31638 );
and ( n93170 , n31098 , n47277 );
or ( n93171 , C0 , n93139 , n93148 , n93169 , n93170 );
buf ( n93172 , n93171 );
buf ( n93173 , n93172 );
buf ( n93174 , n31655 );
buf ( n93175 , n30987 );
and ( n93176 , n50012 , n32494 );
not ( n93177 , n46083 );
and ( n93178 , n93177 , n70742 );
and ( n93179 , n72082 , n46083 );
or ( n93180 , n93178 , n93179 );
and ( n93181 , n93180 , n32421 );
not ( n93182 , n46326 );
and ( n93183 , n93182 , n70742 );
and ( n93184 , n72082 , n46326 );
or ( n93185 , n93183 , n93184 );
and ( n93186 , n93185 , n32417 );
and ( n93187 , n70742 , n46340 );
or ( n93188 , n93181 , n93186 , n93187 );
and ( n93189 , n93188 , n32456 );
and ( n93190 , n70742 , n46349 );
or ( n93191 , C0 , n93176 , n93189 , n93190 );
buf ( n93192 , n93191 );
buf ( n93193 , n93192 );
buf ( n93194 , n31655 );
buf ( n93195 , n31655 );
and ( n93196 , n76107 , n31645 );
not ( n93197 , n45274 );
and ( n93198 , n93197 , n83507 );
and ( n93199 , n82670 , n45274 );
or ( n93200 , n93198 , n93199 );
and ( n93201 , n93200 , n31373 );
not ( n93202 , n45280 );
and ( n93203 , n93202 , n83507 );
and ( n93204 , n82670 , n45280 );
or ( n93205 , n93203 , n93204 );
and ( n93206 , n93205 , n31468 );
and ( n93207 , n83507 , n45802 );
or ( n93208 , n93201 , n93206 , n93207 );
and ( n93209 , n93208 , n31557 );
and ( n93210 , n83507 , n45808 );
or ( n93211 , C0 , n93196 , n93209 , n93210 );
buf ( n93212 , n93211 );
buf ( n93213 , n93212 );
not ( n93214 , n40163 );
and ( n93215 , n93214 , n32007 );
not ( n93216 , n53227 );
and ( n93217 , n93216 , n32007 );
and ( n93218 , n32147 , n53227 );
or ( n93219 , n93217 , n93218 );
and ( n93220 , n93219 , n40163 );
or ( n93221 , n93215 , n93220 );
and ( n93222 , n93221 , n32498 );
not ( n93223 , n53235 );
not ( n93224 , n53227 );
and ( n93225 , n93224 , n32007 );
and ( n93226 , n49314 , n53227 );
or ( n93227 , n93225 , n93226 );
and ( n93228 , n93223 , n93227 );
and ( n93229 , n49314 , n53235 );
or ( n93230 , n93228 , n93229 );
and ( n93231 , n93230 , n32473 );
not ( n93232 , n32475 );
not ( n93233 , n53235 );
not ( n93234 , n53227 );
and ( n93235 , n93234 , n32007 );
and ( n93236 , n49314 , n53227 );
or ( n93237 , n93235 , n93236 );
and ( n93238 , n93233 , n93237 );
and ( n93239 , n49314 , n53235 );
or ( n93240 , n93238 , n93239 );
and ( n93241 , n93232 , n93240 );
not ( n93242 , n53260 );
not ( n93243 , n53262 );
and ( n93244 , n93243 , n93240 );
and ( n93245 , n49340 , n53262 );
or ( n93246 , n93244 , n93245 );
and ( n93247 , n93242 , n93246 );
and ( n93248 , n49348 , n53260 );
or ( n93249 , n93247 , n93248 );
and ( n93250 , n93249 , n32475 );
or ( n93251 , n93241 , n93250 );
and ( n93252 , n93251 , n32486 );
and ( n93253 , n32007 , n41278 );
or ( n93254 , C0 , n93222 , n93231 , n93252 , n93253 );
buf ( n93255 , n93254 );
buf ( n93256 , n93255 );
buf ( n93257 , n30987 );
buf ( n93258 , n30987 );
buf ( n93259 , n30987 );
not ( n93260 , n34150 );
and ( n93261 , n93260 , n32618 );
not ( n93262 , n59105 );
and ( n93263 , n93262 , n32618 );
and ( n93264 , n32655 , n59105 );
or ( n93265 , n93263 , n93264 );
and ( n93266 , n93265 , n34150 );
or ( n93267 , n93261 , n93266 );
and ( n93268 , n93267 , n33381 );
not ( n93269 , n59113 );
not ( n93270 , n59105 );
and ( n93271 , n93270 , n32618 );
and ( n93272 , n56044 , n59105 );
or ( n93273 , n93271 , n93272 );
and ( n93274 , n93269 , n93273 );
and ( n93275 , n56044 , n59113 );
or ( n93276 , n93274 , n93275 );
and ( n93277 , n93276 , n33375 );
not ( n93278 , n32968 );
not ( n93279 , n59113 );
not ( n93280 , n59105 );
and ( n93281 , n93280 , n32618 );
and ( n93282 , n56044 , n59105 );
or ( n93283 , n93281 , n93282 );
and ( n93284 , n93279 , n93283 );
and ( n93285 , n56044 , n59113 );
or ( n93286 , n93284 , n93285 );
and ( n93287 , n93278 , n93286 );
not ( n93288 , n59133 );
not ( n93289 , n59135 );
and ( n93290 , n93289 , n93286 );
and ( n93291 , n56068 , n59135 );
or ( n93292 , n93290 , n93291 );
and ( n93293 , n93288 , n93292 );
and ( n93294 , n56076 , n59133 );
or ( n93295 , n93293 , n93294 );
and ( n93296 , n93295 , n32968 );
or ( n93297 , n93287 , n93296 );
and ( n93298 , n93297 , n33370 );
and ( n93299 , n32618 , n35062 );
or ( n93300 , C0 , n93268 , n93277 , n93298 , n93299 );
buf ( n93301 , n93300 );
buf ( n93302 , n93301 );
buf ( n93303 , n31655 );
buf ( n93304 , n31655 );
and ( n93305 , n59411 , n48455 );
not ( n93306 , n48457 );
and ( n93307 , n93306 , n52394 );
and ( n93308 , n59411 , n48457 );
or ( n93309 , n93307 , n93308 );
and ( n93310 , n93309 , n31373 );
not ( n93311 , n44807 );
and ( n93312 , n93311 , n52394 );
and ( n93313 , n59411 , n44807 );
or ( n93314 , n93312 , n93313 );
and ( n93315 , n93314 , n31408 );
not ( n93316 , n48468 );
and ( n93317 , n93316 , n52394 );
and ( n93318 , n59411 , n48468 );
or ( n93319 , n93317 , n93318 );
and ( n93320 , n93319 , n31468 );
not ( n93321 , n44817 );
and ( n93322 , n93321 , n52394 );
and ( n93323 , n59411 , n44817 );
or ( n93324 , n93322 , n93323 );
and ( n93325 , n93324 , n31521 );
not ( n93326 , n39979 );
and ( n93327 , n93326 , n52394 );
and ( n93328 , n59398 , n39979 );
or ( n93329 , n93327 , n93328 );
and ( n93330 , n93329 , n31538 );
not ( n93331 , n45059 );
and ( n93332 , n93331 , n52394 );
and ( n93333 , n59398 , n45059 );
or ( n93334 , n93332 , n93333 );
and ( n93335 , n93334 , n31536 );
not ( n93336 , n33419 );
and ( n93337 , n93336 , n52394 );
and ( n93338 , n59402 , n33419 );
or ( n93339 , n93337 , n93338 );
and ( n93340 , n93339 , n31529 );
not ( n93341 , n33734 );
and ( n93342 , n93341 , n52394 );
and ( n93343 , n59425 , n33734 );
or ( n93344 , n93342 , n93343 );
and ( n93345 , n93344 , n31527 );
and ( n93346 , n59419 , n48513 );
or ( n93347 , n93305 , n93310 , n93315 , n93320 , n93325 , n93330 , n93335 , n93340 , n93345 , n93346 );
and ( n93348 , n93347 , n31557 );
and ( n93349 , n35375 , n33973 );
and ( n93350 , n52394 , n48524 );
or ( n93351 , C0 , n93348 , n93349 , n93350 );
buf ( n93352 , n93351 );
buf ( n93353 , n93352 );
buf ( n93354 , n31655 );
buf ( n93355 , n30987 );
not ( n93356 , n38443 );
and ( n93357 , n93356 , n38218 );
xor ( n93358 , n53469 , n53500 );
and ( n93359 , n93358 , n38443 );
or ( n93360 , n93357 , n93359 );
and ( n93361 , n93360 , n38450 );
not ( n93362 , n39339 );
and ( n93363 , n93362 , n39118 );
xor ( n93364 , n53525 , n53556 );
and ( n93365 , n93364 , n39339 );
or ( n93366 , n93363 , n93365 );
and ( n93367 , n93366 , n39346 );
and ( n93368 , n40215 , n39359 );
or ( n93369 , n93361 , n93367 , n93368 );
buf ( n93370 , n93369 );
buf ( n93371 , n93370 );
buf ( n93372 , n31655 );
xor ( n93373 , n44767 , n44800 );
and ( n93374 , n93373 , n31548 );
not ( n93375 , n44807 );
and ( n93376 , n93375 , n44767 );
and ( n93377 , n46632 , n44807 );
or ( n93378 , n93376 , n93377 );
and ( n93379 , n93378 , n31408 );
not ( n93380 , n44817 );
and ( n93381 , n93380 , n44767 );
and ( n93382 , n87046 , n44817 );
or ( n93383 , n93381 , n93382 );
and ( n93384 , n93383 , n31521 );
not ( n93385 , n45059 );
and ( n93386 , n93385 , n44767 );
xor ( n93387 , n40035 , n45131 );
and ( n93388 , n93387 , n45059 );
or ( n93389 , n93386 , n93388 );
and ( n93390 , n93389 , n31536 );
and ( n93391 , n44767 , n45148 );
or ( n93392 , n93374 , n93379 , n93384 , n93390 , n93391 );
and ( n93393 , n93392 , n31557 );
and ( n93394 , n44767 , n40154 );
or ( n93395 , C0 , n93393 , n93394 );
buf ( n93396 , n93395 );
buf ( n93397 , n93396 );
not ( n93398 , n40163 );
and ( n93399 , n93398 , n31808 );
not ( n93400 , n45161 );
and ( n93401 , n93400 , n31808 );
and ( n93402 , n32252 , n45161 );
or ( n93403 , n93401 , n93402 );
and ( n93404 , n93403 , n40163 );
or ( n93405 , n93399 , n93404 );
and ( n93406 , n93405 , n32498 );
not ( n93407 , n45170 );
not ( n93408 , n45161 );
and ( n93409 , n93408 , n31808 );
and ( n93410 , n40393 , n45161 );
or ( n93411 , n93409 , n93410 );
and ( n93412 , n93407 , n93411 );
and ( n93413 , n40393 , n45170 );
or ( n93414 , n93412 , n93413 );
and ( n93415 , n93414 , n32473 );
not ( n93416 , n32475 );
not ( n93417 , n45170 );
not ( n93418 , n45161 );
and ( n93419 , n93418 , n31808 );
and ( n93420 , n40393 , n45161 );
or ( n93421 , n93419 , n93420 );
and ( n93422 , n93417 , n93421 );
and ( n93423 , n40393 , n45170 );
or ( n93424 , n93422 , n93423 );
and ( n93425 , n93416 , n93424 );
not ( n93426 , n45196 );
not ( n93427 , n45199 );
and ( n93428 , n93427 , n93424 );
and ( n93429 , n40972 , n45199 );
or ( n93430 , n93428 , n93429 );
and ( n93431 , n93426 , n93430 );
and ( n93432 , n41267 , n45196 );
or ( n93433 , n93431 , n93432 );
and ( n93434 , n93433 , n32475 );
or ( n93435 , n93425 , n93434 );
and ( n93436 , n93435 , n32486 );
and ( n93437 , n31808 , n41278 );
or ( n93438 , C0 , n93406 , n93415 , n93436 , n93437 );
buf ( n93439 , n93438 );
buf ( n93440 , n93439 );
buf ( n93441 , n30987 );
buf ( n93442 , n30987 );
buf ( n93443 , n31655 );
and ( n93444 , n65494 , n31645 );
not ( n93445 , n45274 );
and ( n93446 , n93445 , n66712 );
and ( n93447 , n78189 , n78190 );
buf ( n93448 , n93447 );
and ( n93449 , n93448 , n41809 );
buf ( n93450 , n93449 );
and ( n93451 , n93450 , n45274 );
or ( n93452 , n93446 , n93451 );
and ( n93453 , n93452 , n31373 );
not ( n93454 , n45280 );
and ( n93455 , n93454 , n66712 );
and ( n93456 , n65500 , n45280 );
or ( n93457 , n93455 , n93456 );
and ( n93458 , n93457 , n31468 );
and ( n93459 , n66712 , n45802 );
or ( n93460 , n93453 , n93458 , n93459 );
and ( n93461 , n93460 , n31557 );
and ( n93462 , n66712 , n45808 );
or ( n93463 , C0 , n93444 , n93461 , n93462 );
buf ( n93464 , n93463 );
buf ( n93465 , n93464 );
not ( n93466 , n40163 );
and ( n93467 , n93466 , n31834 );
not ( n93468 , n54629 );
and ( n93469 , n93468 , n31834 );
and ( n93470 , n32235 , n54629 );
or ( n93471 , n93469 , n93470 );
and ( n93472 , n93471 , n40163 );
or ( n93473 , n93467 , n93472 );
and ( n93474 , n93473 , n32498 );
not ( n93475 , n54637 );
not ( n93476 , n54629 );
and ( n93477 , n93476 , n31834 );
and ( n93478 , n42188 , n54629 );
or ( n93479 , n93477 , n93478 );
and ( n93480 , n93475 , n93479 );
and ( n93481 , n42188 , n54637 );
or ( n93482 , n93480 , n93481 );
and ( n93483 , n93482 , n32473 );
not ( n93484 , n32475 );
not ( n93485 , n54637 );
not ( n93486 , n54629 );
and ( n93487 , n93486 , n31834 );
and ( n93488 , n42188 , n54629 );
or ( n93489 , n93487 , n93488 );
and ( n93490 , n93485 , n93489 );
and ( n93491 , n42188 , n54637 );
or ( n93492 , n93490 , n93491 );
and ( n93493 , n93484 , n93492 );
not ( n93494 , n54657 );
not ( n93495 , n54659 );
and ( n93496 , n93495 , n93492 );
and ( n93497 , n42216 , n54659 );
or ( n93498 , n93496 , n93497 );
and ( n93499 , n93494 , n93498 );
and ( n93500 , n42224 , n54657 );
or ( n93501 , n93499 , n93500 );
and ( n93502 , n93501 , n32475 );
or ( n93503 , n93493 , n93502 );
and ( n93504 , n93503 , n32486 );
and ( n93505 , n31834 , n41278 );
or ( n93506 , C0 , n93474 , n93483 , n93504 , n93505 );
buf ( n93507 , n93506 );
buf ( n93508 , n93507 );
buf ( n93509 , n30987 );
not ( n93510 , n43755 );
and ( n93511 , n93510 , n43598 );
xor ( n93512 , n52307 , n52322 );
and ( n93513 , n93512 , n43755 );
or ( n93514 , n93511 , n93513 );
and ( n93515 , n93514 , n43774 );
not ( n93516 , n44663 );
and ( n93517 , n93516 , n44510 );
xor ( n93518 , n52345 , n52360 );
and ( n93519 , n93518 , n44663 );
or ( n93520 , n93517 , n93519 );
and ( n93521 , n93520 , n44682 );
buf ( n93522 , RI15b459d8_240);
and ( n93523 , n93522 , n44695 );
or ( n93524 , n93515 , n93521 , n93523 );
buf ( n93525 , n93524 );
buf ( n93526 , n93525 );
buf ( n93527 , n30987 );
buf ( n93528 , n30987 );
buf ( n93529 , n31655 );
buf ( n93530 , n31655 );
buf ( n93531 , n31655 );
not ( n93532 , n46356 );
and ( n93533 , n93532 , n31218 );
not ( n93534 , n52734 );
and ( n93535 , n93534 , n31218 );
and ( n93536 , n31238 , n52734 );
or ( n93537 , n93535 , n93536 );
and ( n93538 , n93537 , n46356 );
or ( n93539 , n93533 , n93538 );
and ( n93540 , n93539 , n31649 );
not ( n93541 , n52742 );
not ( n93542 , n52734 );
and ( n93543 , n93542 , n31218 );
and ( n93544 , n49901 , n52734 );
or ( n93545 , n93543 , n93544 );
and ( n93546 , n93541 , n93545 );
and ( n93547 , n49901 , n52742 );
or ( n93548 , n93546 , n93547 );
and ( n93549 , n93548 , n31643 );
not ( n93550 , n31452 );
not ( n93551 , n52742 );
not ( n93552 , n52734 );
and ( n93553 , n93552 , n31218 );
and ( n93554 , n49901 , n52734 );
or ( n93555 , n93553 , n93554 );
and ( n93556 , n93551 , n93555 );
and ( n93557 , n49901 , n52742 );
or ( n93558 , n93556 , n93557 );
and ( n93559 , n93550 , n93558 );
not ( n93560 , n52762 );
not ( n93561 , n52764 );
and ( n93562 , n93561 , n93558 );
and ( n93563 , n49925 , n52764 );
or ( n93564 , n93562 , n93563 );
and ( n93565 , n93560 , n93564 );
and ( n93566 , n49933 , n52762 );
or ( n93567 , n93565 , n93566 );
and ( n93568 , n93567 , n31452 );
or ( n93569 , n93559 , n93568 );
and ( n93570 , n93569 , n31638 );
and ( n93571 , n31218 , n47277 );
or ( n93572 , C0 , n93540 , n93549 , n93570 , n93571 );
buf ( n93573 , n93572 );
buf ( n93574 , n93573 );
buf ( n93575 , n30987 );
not ( n93576 , n35211 );
and ( n93577 , n48530 , n93576 );
and ( n93578 , n93577 , n32421 );
not ( n93579 , n35245 );
and ( n93580 , n48530 , n93579 );
and ( n93581 , n93580 , n32419 );
not ( n93582 , n35278 );
and ( n93583 , n93582 , n48530 );
buf ( n93584 , n35278 );
or ( n93585 , n93583 , n93584 );
and ( n93586 , n93585 , n32417 );
not ( n93587 , n35331 );
and ( n93588 , n93587 , n48530 );
buf ( n93589 , n35331 );
or ( n93590 , n93588 , n93589 );
and ( n93591 , n93590 , n32415 );
and ( n93592 , n48530 , n35354 );
or ( n93593 , n93578 , n93581 , n93586 , n93591 , n93592 );
and ( n93594 , n93593 , n32456 );
and ( n93595 , n48530 , n81226 );
buf ( n93596 , n68574 );
or ( n93597 , C0 , n93594 , n93595 , n93596 );
buf ( n93598 , n93597 );
buf ( n93599 , n93598 );
buf ( n93600 , n31655 );
buf ( n93601 , n30987 );
buf ( n93602 , n30987 );
not ( n93603 , n34150 );
and ( n93604 , n93603 , n32696 );
not ( n93605 , n59574 );
and ( n93606 , n93605 , n32696 );
and ( n93607 , n32722 , n59574 );
or ( n93608 , n93606 , n93607 );
and ( n93609 , n93608 , n34150 );
or ( n93610 , n93604 , n93609 );
and ( n93611 , n93610 , n33381 );
not ( n93612 , n59582 );
not ( n93613 , n59574 );
and ( n93614 , n93613 , n32696 );
and ( n93615 , n42565 , n59574 );
or ( n93616 , n93614 , n93615 );
and ( n93617 , n93612 , n93616 );
and ( n93618 , n42565 , n59582 );
or ( n93619 , n93617 , n93618 );
and ( n93620 , n93619 , n33375 );
not ( n93621 , n32968 );
not ( n93622 , n59582 );
not ( n93623 , n59574 );
and ( n93624 , n93623 , n32696 );
and ( n93625 , n42565 , n59574 );
or ( n93626 , n93624 , n93625 );
and ( n93627 , n93622 , n93626 );
and ( n93628 , n42565 , n59582 );
or ( n93629 , n93627 , n93628 );
and ( n93630 , n93621 , n93629 );
not ( n93631 , n59602 );
not ( n93632 , n59604 );
and ( n93633 , n93632 , n93629 );
and ( n93634 , n42589 , n59604 );
or ( n93635 , n93633 , n93634 );
and ( n93636 , n93631 , n93635 );
and ( n93637 , n42597 , n59602 );
or ( n93638 , n93636 , n93637 );
and ( n93639 , n93638 , n32968 );
or ( n93640 , n93630 , n93639 );
and ( n93641 , n93640 , n33370 );
and ( n93642 , n32696 , n35062 );
or ( n93643 , C0 , n93611 , n93620 , n93641 , n93642 );
buf ( n93644 , n93643 );
buf ( n93645 , n93644 );
buf ( n93646 , n31655 );
buf ( n93647 , n31655 );
buf ( n93648 , n30987 );
buf ( n93649 , n30987 );
not ( n93650 , n34150 );
and ( n93651 , n93650 , n32718 );
not ( n93652 , n56140 );
and ( n93653 , n93652 , n32718 );
and ( n93654 , n32722 , n56140 );
or ( n93655 , n93653 , n93654 );
and ( n93656 , n93655 , n34150 );
or ( n93657 , n93651 , n93656 );
and ( n93658 , n93657 , n33381 );
not ( n93659 , n56148 );
not ( n93660 , n56140 );
and ( n93661 , n93660 , n32718 );
and ( n93662 , n42565 , n56140 );
or ( n93663 , n93661 , n93662 );
and ( n93664 , n93659 , n93663 );
and ( n93665 , n42565 , n56148 );
or ( n93666 , n93664 , n93665 );
and ( n93667 , n93666 , n33375 );
not ( n93668 , n32968 );
not ( n93669 , n56148 );
not ( n93670 , n56140 );
and ( n93671 , n93670 , n32718 );
and ( n93672 , n42565 , n56140 );
or ( n93673 , n93671 , n93672 );
and ( n93674 , n93669 , n93673 );
and ( n93675 , n42565 , n56148 );
or ( n93676 , n93674 , n93675 );
and ( n93677 , n93668 , n93676 );
not ( n93678 , n56168 );
not ( n93679 , n56170 );
and ( n93680 , n93679 , n93676 );
and ( n93681 , n42589 , n56170 );
or ( n93682 , n93680 , n93681 );
and ( n93683 , n93678 , n93682 );
and ( n93684 , n42597 , n56168 );
or ( n93685 , n93683 , n93684 );
and ( n93686 , n93685 , n32968 );
or ( n93687 , n93677 , n93686 );
and ( n93688 , n93687 , n33370 );
and ( n93689 , n32718 , n35062 );
or ( n93690 , C0 , n93658 , n93667 , n93688 , n93689 );
buf ( n93691 , n93690 );
buf ( n93692 , n93691 );
not ( n93693 , n34150 );
and ( n93694 , n93693 , n32815 );
not ( n93695 , n56093 );
and ( n93696 , n93695 , n32815 );
and ( n93697 , n32823 , n56093 );
or ( n93698 , n93696 , n93697 );
and ( n93699 , n93698 , n34150 );
or ( n93700 , n93694 , n93699 );
and ( n93701 , n93700 , n33381 );
not ( n93702 , n56101 );
not ( n93703 , n56093 );
and ( n93704 , n93703 , n32815 );
and ( n93705 , n41464 , n56093 );
or ( n93706 , n93704 , n93705 );
and ( n93707 , n93702 , n93706 );
and ( n93708 , n41464 , n56101 );
or ( n93709 , n93707 , n93708 );
and ( n93710 , n93709 , n33375 );
not ( n93711 , n32968 );
not ( n93712 , n56101 );
not ( n93713 , n56093 );
and ( n93714 , n93713 , n32815 );
and ( n93715 , n41464 , n56093 );
or ( n93716 , n93714 , n93715 );
and ( n93717 , n93712 , n93716 );
and ( n93718 , n41464 , n56101 );
or ( n93719 , n93717 , n93718 );
and ( n93720 , n93711 , n93719 );
not ( n93721 , n56121 );
not ( n93722 , n56123 );
and ( n93723 , n93722 , n93719 );
and ( n93724 , n41490 , n56123 );
or ( n93725 , n93723 , n93724 );
and ( n93726 , n93721 , n93725 );
and ( n93727 , n41500 , n56121 );
or ( n93728 , n93726 , n93727 );
and ( n93729 , n93728 , n32968 );
or ( n93730 , n93720 , n93729 );
and ( n93731 , n93730 , n33370 );
and ( n93732 , n32815 , n35062 );
or ( n93733 , C0 , n93701 , n93710 , n93731 , n93732 );
buf ( n93734 , n93733 );
buf ( n93735 , n93734 );
buf ( n93736 , n31655 );
buf ( n93737 , n31655 );
not ( n93738 , n36587 );
and ( n93739 , n93738 , n36192 );
xor ( n93740 , n50189 , n50198 );
and ( n93741 , n93740 , n36587 );
or ( n93742 , n93739 , n93741 );
and ( n93743 , n93742 , n36596 );
not ( n93744 , n37485 );
and ( n93745 , n93744 , n37094 );
xor ( n93746 , n50239 , n50248 );
and ( n93747 , n93746 , n37485 );
or ( n93748 , n93745 , n93747 );
and ( n93749 , n93748 , n37494 );
and ( n93750 , n41845 , n37506 );
or ( n93751 , n93743 , n93749 , n93750 );
buf ( n93752 , n93751 );
buf ( n93753 , n93752 );
buf ( n93754 , n31655 );
buf ( n93755 , n30987 );
buf ( n93756 , n32498 );
buf ( n93757 , n32496 );
not ( n93758 , n76230 );
not ( n93759 , n76232 );
and ( n93760 , n93759 , n32440 );
buf ( n93761 , n93760 );
and ( n93762 , n93761 , n32417 );
and ( n93763 , n32440 , n76244 );
or ( n93764 , n93762 , n93763 );
and ( n93765 , n93758 , n93764 );
buf ( n93766 , n93765 );
and ( n93767 , n93766 , n32456 );
or ( n93768 , C0 , n93756 , n93757 , C0 , n93767 , C0 , C0 , C0 , C0 , C0 );
buf ( n93769 , n93768 );
buf ( n93770 , n93769 );
buf ( n93771 , n31655 );
and ( n93772 , n33765 , n48455 );
not ( n93773 , n48457 );
and ( n93774 , n93773 , n33430 );
and ( n93775 , n33765 , n48457 );
or ( n93776 , n93774 , n93775 );
and ( n93777 , n93776 , n31373 );
not ( n93778 , n44807 );
and ( n93779 , n93778 , n33430 );
and ( n93780 , n33765 , n44807 );
or ( n93781 , n93779 , n93780 );
and ( n93782 , n93781 , n31408 );
not ( n93783 , n48468 );
and ( n93784 , n93783 , n33430 );
and ( n93785 , n33765 , n48468 );
or ( n93786 , n93784 , n93785 );
and ( n93787 , n93786 , n31468 );
not ( n93788 , n44817 );
and ( n93789 , n93788 , n33430 );
and ( n93790 , n33765 , n44817 );
or ( n93791 , n93789 , n93790 );
and ( n93792 , n93791 , n31521 );
not ( n93793 , n39979 );
and ( n93794 , n93793 , n33430 );
and ( n93795 , n33472 , n39979 );
or ( n93796 , n93794 , n93795 );
and ( n93797 , n93796 , n31538 );
not ( n93798 , n45059 );
and ( n93799 , n93798 , n33430 );
and ( n93800 , n33472 , n45059 );
or ( n93801 , n93799 , n93800 );
and ( n93802 , n93801 , n31536 );
not ( n93803 , n33419 );
and ( n93804 , n93803 , n33430 );
xor ( n93805 , n33472 , n33693 );
and ( n93806 , n93805 , n33419 );
or ( n93807 , n93804 , n93806 );
and ( n93808 , n93807 , n31529 );
not ( n93809 , n33734 );
and ( n93810 , n93809 , n33430 );
not ( n93811 , n33533 );
xor ( n93812 , n33765 , n33811 );
and ( n93813 , n93811 , n93812 );
xnor ( n93814 , n33850 , n33913 );
and ( n93815 , n93814 , n33533 );
or ( n93816 , n93813 , n93815 );
and ( n93817 , n93816 , n33734 );
or ( n93818 , n93810 , n93817 );
and ( n93819 , n93818 , n31527 );
and ( n93820 , n33850 , n48513 );
or ( n93821 , n93772 , n93777 , n93782 , n93787 , n93792 , n93797 , n93802 , n93808 , n93819 , n93820 );
and ( n93822 , n93821 , n31557 );
and ( n93823 , n34002 , n33973 );
and ( n93824 , n33430 , n48524 );
or ( n93825 , C0 , n93822 , n93823 , n93824 );
buf ( n93826 , n93825 );
buf ( n93827 , n93826 );
buf ( n93828 , n30987 );
not ( n93829 , n35278 );
and ( n93830 , n93829 , n85029 );
and ( n93831 , n85048 , n35278 );
or ( n93832 , n93830 , n93831 );
and ( n93833 , n93832 , n32417 );
not ( n93834 , n50008 );
and ( n93835 , n93834 , n85029 );
and ( n93836 , n85959 , n50008 );
or ( n93837 , n93835 , n93836 );
and ( n93838 , n93837 , n32415 );
and ( n93839 , n85029 , n48133 );
or ( n93840 , n93833 , n93838 , n93839 );
and ( n93841 , n93840 , n32456 );
and ( n93842 , n85029 , n47409 );
or ( n93843 , C0 , n93841 , n93842 );
buf ( n93844 , n93843 );
buf ( n93845 , n93844 );
not ( n93846 , n46356 );
and ( n93847 , n93846 , n31337 );
not ( n93848 , n60564 );
and ( n93849 , n93848 , n31337 );
and ( n93850 , n31339 , n60564 );
or ( n93851 , n93849 , n93850 );
and ( n93852 , n93851 , n46356 );
or ( n93853 , n93847 , n93852 );
and ( n93854 , n93853 , n31649 );
not ( n93855 , n60572 );
not ( n93856 , n60564 );
and ( n93857 , n93856 , n31337 );
and ( n93858 , n47449 , n60564 );
or ( n93859 , n93857 , n93858 );
and ( n93860 , n93855 , n93859 );
and ( n93861 , n47449 , n60572 );
or ( n93862 , n93860 , n93861 );
and ( n93863 , n93862 , n31643 );
not ( n93864 , n31452 );
not ( n93865 , n60572 );
not ( n93866 , n60564 );
and ( n93867 , n93866 , n31337 );
and ( n93868 , n47449 , n60564 );
or ( n93869 , n93867 , n93868 );
and ( n93870 , n93865 , n93869 );
and ( n93871 , n47449 , n60572 );
or ( n93872 , n93870 , n93871 );
and ( n93873 , n93864 , n93872 );
not ( n93874 , n60592 );
not ( n93875 , n60594 );
and ( n93876 , n93875 , n93872 );
and ( n93877 , n47485 , n60594 );
or ( n93878 , n93876 , n93877 );
and ( n93879 , n93874 , n93878 );
and ( n93880 , n47503 , n60592 );
or ( n93881 , n93879 , n93880 );
and ( n93882 , n93881 , n31452 );
or ( n93883 , n93873 , n93882 );
and ( n93884 , n93883 , n31638 );
and ( n93885 , n31337 , n47277 );
or ( n93886 , C0 , n93854 , n93863 , n93884 , n93885 );
buf ( n93887 , n93886 );
buf ( n93888 , n93887 );
buf ( n93889 , n31655 );
buf ( n93890 , n30987 );
buf ( n93891 , n30987 );
xor ( n93892 , n49569 , n60321 );
and ( n93893 , n93892 , n32433 );
not ( n93894 , n47331 );
and ( n93895 , n93894 , n49569 );
xor ( n93896 , n60433 , n60545 );
and ( n93897 , n93896 , n47331 );
or ( n93898 , n93895 , n93897 );
and ( n93899 , n93898 , n32413 );
and ( n93900 , n49569 , n47402 );
or ( n93901 , n93893 , n93899 , n93900 );
and ( n93902 , n93901 , n32456 );
and ( n93903 , n49569 , n47409 );
or ( n93904 , C0 , n93902 , n93903 );
buf ( n93905 , n93904 );
buf ( n93906 , n93905 );
buf ( n93907 , n31655 );
buf ( n93908 , n30987 );
not ( n93909 , n34150 );
and ( n93910 , n93909 , n32739 );
not ( n93911 , n57038 );
and ( n93912 , n93911 , n32739 );
and ( n93913 , n32755 , n57038 );
or ( n93914 , n93912 , n93913 );
and ( n93915 , n93914 , n34150 );
or ( n93916 , n93910 , n93915 );
and ( n93917 , n93916 , n33381 );
not ( n93918 , n57046 );
not ( n93919 , n57038 );
and ( n93920 , n93919 , n32739 );
and ( n93921 , n35083 , n57038 );
or ( n93922 , n93920 , n93921 );
and ( n93923 , n93918 , n93922 );
and ( n93924 , n35083 , n57046 );
or ( n93925 , n93923 , n93924 );
and ( n93926 , n93925 , n33375 );
not ( n93927 , n32968 );
not ( n93928 , n57046 );
not ( n93929 , n57038 );
and ( n93930 , n93929 , n32739 );
and ( n93931 , n35083 , n57038 );
or ( n93932 , n93930 , n93931 );
and ( n93933 , n93928 , n93932 );
and ( n93934 , n35083 , n57046 );
or ( n93935 , n93933 , n93934 );
and ( n93936 , n93927 , n93935 );
not ( n93937 , n57066 );
not ( n93938 , n57068 );
and ( n93939 , n93938 , n93935 );
and ( n93940 , n35107 , n57068 );
or ( n93941 , n93939 , n93940 );
and ( n93942 , n93937 , n93941 );
and ( n93943 , n35115 , n57066 );
or ( n93944 , n93942 , n93943 );
and ( n93945 , n93944 , n32968 );
or ( n93946 , n93936 , n93945 );
and ( n93947 , n93946 , n33370 );
and ( n93948 , n32739 , n35062 );
or ( n93949 , C0 , n93917 , n93926 , n93947 , n93948 );
buf ( n93950 , n93949 );
buf ( n93951 , n93950 );
buf ( n93952 , n40216 );
buf ( n93953 , n30987 );
buf ( n93954 , n31655 );
buf ( n93955 , n31655 );
buf ( n93956 , n31655 );
xor ( n93957 , n44765 , n44802 );
and ( n93958 , n93957 , n31548 );
not ( n93959 , n44807 );
and ( n93960 , n93959 , n44765 );
and ( n93961 , n46622 , n44807 );
or ( n93962 , n93960 , n93961 );
and ( n93963 , n93962 , n31408 );
not ( n93964 , n44817 );
and ( n93965 , n93964 , n44765 );
not ( n93966 , n44994 );
and ( n93967 , n93966 , n44954 );
xor ( n93968 , n44999 , n45021 );
and ( n93969 , n93968 , n44994 );
or ( n93970 , n93967 , n93969 );
and ( n93971 , n93970 , n44817 );
or ( n93972 , n93965 , n93971 );
and ( n93973 , n93972 , n31521 );
not ( n93974 , n45059 );
and ( n93975 , n93974 , n44765 );
xor ( n93976 , n45112 , n45133 );
and ( n93977 , n93976 , n45059 );
or ( n93978 , n93975 , n93977 );
and ( n93979 , n93978 , n31536 );
and ( n93980 , n44765 , n45148 );
or ( n93981 , n93958 , n93963 , n93973 , n93979 , n93980 );
and ( n93982 , n93981 , n31557 );
and ( n93983 , n44765 , n40154 );
or ( n93984 , C0 , n93982 , n93983 );
buf ( n93985 , n93984 );
buf ( n93986 , n93985 );
not ( n93987 , n40163 );
and ( n93988 , n93987 , n31883 );
not ( n93989 , n45161 );
and ( n93990 , n93989 , n31883 );
and ( n93991 , n32218 , n45161 );
or ( n93992 , n93990 , n93991 );
and ( n93993 , n93992 , n40163 );
or ( n93994 , n93988 , n93993 );
and ( n93995 , n93994 , n32498 );
not ( n93996 , n45170 );
not ( n93997 , n45161 );
and ( n93998 , n93997 , n31883 );
and ( n93999 , n42255 , n45161 );
or ( n94000 , n93998 , n93999 );
and ( n94001 , n93996 , n94000 );
and ( n94002 , n42255 , n45170 );
or ( n94003 , n94001 , n94002 );
and ( n94004 , n94003 , n32473 );
not ( n94005 , n32475 );
not ( n94006 , n45170 );
not ( n94007 , n45161 );
and ( n94008 , n94007 , n31883 );
and ( n94009 , n42255 , n45161 );
or ( n94010 , n94008 , n94009 );
and ( n94011 , n94006 , n94010 );
and ( n94012 , n42255 , n45170 );
or ( n94013 , n94011 , n94012 );
and ( n94014 , n94005 , n94013 );
not ( n94015 , n45196 );
not ( n94016 , n45199 );
and ( n94017 , n94016 , n94013 );
and ( n94018 , n42283 , n45199 );
or ( n94019 , n94017 , n94018 );
and ( n94020 , n94015 , n94019 );
and ( n94021 , n42291 , n45196 );
or ( n94022 , n94020 , n94021 );
and ( n94023 , n94022 , n32475 );
or ( n94024 , n94014 , n94023 );
and ( n94025 , n94024 , n32486 );
and ( n94026 , n31883 , n41278 );
or ( n94027 , C0 , n93995 , n94004 , n94025 , n94026 );
buf ( n94028 , n94027 );
buf ( n94029 , n94028 );
buf ( n94030 , n30987 );
buf ( n94031 , n30987 );
xor ( n94032 , n33099 , n58384 );
and ( n94033 , n94032 , n33201 );
not ( n94034 , n41576 );
and ( n94035 , n94034 , n33099 );
and ( n94036 , n91173 , n41576 );
or ( n94037 , n94035 , n94036 );
and ( n94038 , n94037 , n33189 );
and ( n94039 , n33099 , n41592 );
or ( n94040 , n94033 , n94038 , n94039 );
and ( n94041 , n94040 , n33208 );
and ( n94042 , n33099 , n39805 );
or ( n94043 , C0 , n94041 , n94042 );
buf ( n94044 , n94043 );
buf ( n94045 , n94044 );
buf ( n94046 , n31655 );
buf ( n94047 , n30987 );
buf ( n94048 , n30987 );
buf ( n94049 , n31655 );
not ( n94050 , n50828 );
not ( n94051 , n50834 );
and ( n94052 , n94051 , n40618 );
and ( n94053 , n91188 , n50834 );
or ( n94054 , n94052 , n94053 );
and ( n94055 , n94050 , n94054 );
and ( n94056 , n79208 , n50828 );
or ( n94057 , n94055 , n94056 );
buf ( n94058 , n94057 );
buf ( n94059 , n94058 );
not ( n94060 , n46356 );
and ( n94061 , n94060 , n31325 );
not ( n94062 , n50109 );
and ( n94063 , n94062 , n31325 );
and ( n94064 , n31339 , n50109 );
or ( n94065 , n94063 , n94064 );
and ( n94066 , n94065 , n46356 );
or ( n94067 , n94061 , n94066 );
and ( n94068 , n94067 , n31649 );
not ( n94069 , n50117 );
not ( n94070 , n50109 );
and ( n94071 , n94070 , n31325 );
and ( n94072 , n47449 , n50109 );
or ( n94073 , n94071 , n94072 );
and ( n94074 , n94069 , n94073 );
and ( n94075 , n47449 , n50117 );
or ( n94076 , n94074 , n94075 );
and ( n94077 , n94076 , n31643 );
not ( n94078 , n31452 );
not ( n94079 , n50117 );
not ( n94080 , n50109 );
and ( n94081 , n94080 , n31325 );
and ( n94082 , n47449 , n50109 );
or ( n94083 , n94081 , n94082 );
and ( n94084 , n94079 , n94083 );
and ( n94085 , n47449 , n50117 );
or ( n94086 , n94084 , n94085 );
and ( n94087 , n94078 , n94086 );
not ( n94088 , n50142 );
not ( n94089 , n50144 );
and ( n94090 , n94089 , n94086 );
and ( n94091 , n47485 , n50144 );
or ( n94092 , n94090 , n94091 );
and ( n94093 , n94088 , n94092 );
and ( n94094 , n47503 , n50142 );
or ( n94095 , n94093 , n94094 );
and ( n94096 , n94095 , n31452 );
or ( n94097 , n94087 , n94096 );
and ( n94098 , n94097 , n31638 );
and ( n94099 , n31325 , n47277 );
or ( n94100 , C0 , n94068 , n94077 , n94098 , n94099 );
buf ( n94101 , n94100 );
buf ( n94102 , n94101 );
buf ( n94103 , n31655 );
buf ( n94104 , n30987 );
xor ( n94105 , n46211 , n49995 );
and ( n94106 , n94105 , n32431 );
not ( n94107 , n50002 );
and ( n94108 , n94107 , n46211 );
and ( n94109 , n40500 , n50002 );
or ( n94110 , n94108 , n94109 );
and ( n94111 , n94110 , n32419 );
not ( n94112 , n50008 );
and ( n94113 , n94112 , n46211 );
not ( n94114 , n47910 );
and ( n94115 , n94114 , n69733 );
and ( n94116 , n69749 , n47910 );
or ( n94117 , n94115 , n94116 );
and ( n94118 , n94117 , n50008 );
or ( n94119 , n94113 , n94118 );
and ( n94120 , n94119 , n32415 );
not ( n94121 , n50067 );
and ( n94122 , n94121 , n46211 );
and ( n94123 , n47389 , n50067 );
or ( n94124 , n94122 , n94123 );
and ( n94125 , n94124 , n32411 );
and ( n94126 , n46211 , n50098 );
or ( n94127 , n94106 , n94111 , n94120 , n94125 , n94126 );
and ( n94128 , n94127 , n32456 );
and ( n94129 , n46211 , n47409 );
or ( n94130 , C0 , n94128 , n94129 );
buf ( n94131 , n94130 );
buf ( n94132 , n94131 );
buf ( n94133 , n31655 );
buf ( n94134 , n31655 );
not ( n94135 , n46356 );
and ( n94136 , n94135 , n31274 );
not ( n94137 , n63024 );
and ( n94138 , n94137 , n31274 );
and ( n94139 , n31306 , n63024 );
or ( n94140 , n94138 , n94139 );
and ( n94141 , n94140 , n46356 );
or ( n94142 , n94136 , n94141 );
and ( n94143 , n94142 , n31649 );
not ( n94144 , n63032 );
not ( n94145 , n63024 );
and ( n94146 , n94145 , n31274 );
and ( n94147 , n58061 , n63024 );
or ( n94148 , n94146 , n94147 );
and ( n94149 , n94144 , n94148 );
and ( n94150 , n58061 , n63032 );
or ( n94151 , n94149 , n94150 );
and ( n94152 , n94151 , n31643 );
not ( n94153 , n31452 );
not ( n94154 , n63032 );
not ( n94155 , n63024 );
and ( n94156 , n94155 , n31274 );
and ( n94157 , n58061 , n63024 );
or ( n94158 , n94156 , n94157 );
and ( n94159 , n94154 , n94158 );
and ( n94160 , n58061 , n63032 );
or ( n94161 , n94159 , n94160 );
and ( n94162 , n94153 , n94161 );
not ( n94163 , n63052 );
not ( n94164 , n63054 );
and ( n94165 , n94164 , n94161 );
and ( n94166 , n58085 , n63054 );
or ( n94167 , n94165 , n94166 );
and ( n94168 , n94163 , n94167 );
and ( n94169 , n58093 , n63052 );
or ( n94170 , n94168 , n94169 );
and ( n94171 , n94170 , n31452 );
or ( n94172 , n94162 , n94171 );
and ( n94173 , n94172 , n31638 );
and ( n94174 , n31274 , n47277 );
or ( n94175 , C0 , n94143 , n94152 , n94173 , n94174 );
buf ( n94176 , n94175 );
buf ( n94177 , n94176 );
buf ( n94178 , n30987 );
not ( n94179 , n35278 );
and ( n94180 , n94179 , n55319 );
and ( n94181 , n60224 , n35278 );
or ( n94182 , n94180 , n94181 );
and ( n94183 , n94182 , n32417 );
not ( n94184 , n47912 );
and ( n94185 , n94184 , n55319 );
and ( n94186 , n55325 , n47912 );
or ( n94187 , n94185 , n94186 );
and ( n94188 , n94187 , n32415 );
and ( n94189 , n55319 , n48133 );
or ( n94190 , n94183 , n94188 , n94189 );
and ( n94191 , n94190 , n32456 );
and ( n94192 , n55319 , n47409 );
or ( n94193 , C0 , n94191 , n94192 );
buf ( n94194 , n94193 );
buf ( n94195 , n94194 );
and ( n94196 , n33769 , n48455 );
not ( n94197 , n48457 );
and ( n94198 , n94197 , n33434 );
and ( n94199 , n33769 , n48457 );
or ( n94200 , n94198 , n94199 );
and ( n94201 , n94200 , n31373 );
not ( n94202 , n44807 );
and ( n94203 , n94202 , n33434 );
and ( n94204 , n33769 , n44807 );
or ( n94205 , n94203 , n94204 );
and ( n94206 , n94205 , n31408 );
not ( n94207 , n48468 );
and ( n94208 , n94207 , n33434 );
and ( n94209 , n33769 , n48468 );
or ( n94210 , n94208 , n94209 );
and ( n94211 , n94210 , n31468 );
not ( n94212 , n44817 );
and ( n94213 , n94212 , n33434 );
and ( n94214 , n33769 , n44817 );
or ( n94215 , n94213 , n94214 );
and ( n94216 , n94215 , n31521 );
not ( n94217 , n39979 );
and ( n94218 , n94217 , n33434 );
and ( n94219 , n33476 , n39979 );
or ( n94220 , n94218 , n94219 );
and ( n94221 , n94220 , n31538 );
not ( n94222 , n45059 );
and ( n94223 , n94222 , n33434 );
and ( n94224 , n33476 , n45059 );
or ( n94225 , n94223 , n94224 );
and ( n94226 , n94225 , n31536 );
not ( n94227 , n33419 );
and ( n94228 , n94227 , n33434 );
and ( n94229 , n92706 , n33419 );
or ( n94230 , n94228 , n94229 );
and ( n94231 , n94230 , n31529 );
not ( n94232 , n33734 );
and ( n94233 , n94232 , n33434 );
and ( n94234 , n92717 , n33734 );
or ( n94235 , n94233 , n94234 );
and ( n94236 , n94235 , n31527 );
and ( n94237 , n33854 , n48513 );
or ( n94238 , n94196 , n94201 , n94206 , n94211 , n94216 , n94221 , n94226 , n94231 , n94236 , n94237 );
and ( n94239 , n94238 , n31557 );
and ( n94240 , n34006 , n33973 );
and ( n94241 , n33434 , n48524 );
or ( n94242 , C0 , n94239 , n94240 , n94241 );
buf ( n94243 , n94242 );
buf ( n94244 , n94243 );
buf ( n94245 , n31655 );
buf ( n94246 , n30987 );
not ( n94247 , n35278 );
and ( n94248 , n94247 , n78296 );
and ( n94249 , n78308 , n35278 );
or ( n94250 , n94248 , n94249 );
and ( n94251 , n94250 , n32417 );
not ( n94252 , n50008 );
and ( n94253 , n94252 , n78296 );
and ( n94254 , n68940 , n50008 );
or ( n94255 , n94253 , n94254 );
and ( n94256 , n94255 , n32415 );
and ( n94257 , n78296 , n48133 );
or ( n94258 , n94251 , n94256 , n94257 );
and ( n94259 , n94258 , n32456 );
and ( n94260 , n78296 , n47409 );
or ( n94261 , C0 , n94259 , n94260 );
buf ( n94262 , n94261 );
buf ( n94263 , n94262 );
not ( n94264 , n48765 );
and ( n94265 , n94264 , n33217 );
and ( n94266 , n64430 , n48765 );
or ( n94267 , n94265 , n94266 );
and ( n94268 , n94267 , n33180 );
not ( n94269 , n49054 );
and ( n94270 , n94269 , n33217 );
and ( n94271 , n64441 , n49054 );
or ( n94272 , n94270 , n94271 );
and ( n94273 , n94272 , n33178 );
and ( n94274 , n33217 , n49774 );
or ( n94275 , n94268 , n94273 , n94274 );
and ( n94276 , n94275 , n33208 );
and ( n94277 , n33285 , n33375 );
not ( n94278 , n32968 );
and ( n94279 , n94278 , n33285 );
xor ( n94280 , n33217 , n59701 );
and ( n94281 , n94280 , n32968 );
or ( n94282 , n94279 , n94281 );
and ( n94283 , n94282 , n33370 );
and ( n94284 , n32980 , n35056 );
and ( n94285 , n33217 , n49794 );
or ( n94286 , C0 , n94276 , n94277 , n94283 , n94284 , n94285 );
buf ( n94287 , n94286 );
buf ( n94288 , n94287 );
buf ( n94289 , n30987 );
buf ( n94290 , n40211 );
buf ( n94291 , n31655 );
buf ( n94292 , n30987 );
buf ( n94293 , n31655 );
and ( n94294 , n46033 , n32500 );
not ( n94295 , n35211 );
and ( n94296 , n94295 , n37563 );
buf ( n94297 , n94296 );
and ( n94298 , n94297 , n32421 );
not ( n94299 , n35245 );
and ( n94300 , n94299 , n37563 );
buf ( n94301 , n94300 );
and ( n94302 , n94301 , n32419 );
not ( n94303 , n35278 );
and ( n94304 , n94303 , n37563 );
not ( n94305 , n35295 );
and ( n94306 , n94305 , n49593 );
xor ( n94307 , n37563 , n49534 );
and ( n94308 , n94307 , n35295 );
or ( n94309 , n94306 , n94308 );
and ( n94310 , n94309 , n35278 );
or ( n94311 , n94304 , n94310 );
and ( n94312 , n94311 , n32417 );
not ( n94313 , n35331 );
and ( n94314 , n94313 , n37563 );
not ( n94315 , n35294 );
not ( n94316 , n45995 );
and ( n94317 , n94316 , n49593 );
xor ( n94318 , n49594 , n49620 );
and ( n94319 , n94318 , n45995 );
or ( n94320 , n94317 , n94319 );
and ( n94321 , n94315 , n94320 );
and ( n94322 , n94307 , n35294 );
or ( n94323 , n94321 , n94322 );
and ( n94324 , n94323 , n35331 );
or ( n94325 , n94314 , n94324 );
and ( n94326 , n94325 , n32415 );
and ( n94327 , n37563 , n35354 );
or ( n94328 , n94298 , n94302 , n94312 , n94326 , n94327 );
and ( n94329 , n94328 , n32456 );
not ( n94330 , n32475 );
not ( n94331 , n46060 );
and ( n94332 , n94331 , n49683 );
xor ( n94333 , n49684 , n49714 );
and ( n94334 , n94333 , n46060 );
or ( n94335 , n94332 , n94334 );
and ( n94336 , n94330 , n94335 );
and ( n94337 , n37563 , n32475 );
or ( n94338 , n94336 , n94337 );
and ( n94339 , n94338 , n32486 );
buf ( n94340 , n32489 );
and ( n94341 , n37563 , n35367 );
or ( n94342 , C0 , n94294 , n94329 , n94339 , n94340 , n94341 );
buf ( n94343 , n94342 );
buf ( n94344 , n94343 );
buf ( n94345 , n31655 );
not ( n94346 , n46356 );
and ( n94347 , n94346 , n31108 );
not ( n94348 , n52734 );
and ( n94349 , n94348 , n31108 );
and ( n94350 , n31138 , n52734 );
or ( n94351 , n94349 , n94350 );
and ( n94352 , n94351 , n46356 );
or ( n94353 , n94347 , n94352 );
and ( n94354 , n94353 , n31649 );
not ( n94355 , n52742 );
not ( n94356 , n52734 );
and ( n94357 , n94356 , n31108 );
and ( n94358 , n56920 , n52734 );
or ( n94359 , n94357 , n94358 );
and ( n94360 , n94355 , n94359 );
and ( n94361 , n56920 , n52742 );
or ( n94362 , n94360 , n94361 );
and ( n94363 , n94362 , n31643 );
not ( n94364 , n31452 );
not ( n94365 , n52742 );
not ( n94366 , n52734 );
and ( n94367 , n94366 , n31108 );
and ( n94368 , n56920 , n52734 );
or ( n94369 , n94367 , n94368 );
and ( n94370 , n94365 , n94369 );
and ( n94371 , n56920 , n52742 );
or ( n94372 , n94370 , n94371 );
and ( n94373 , n94364 , n94372 );
not ( n94374 , n52762 );
not ( n94375 , n52764 );
and ( n94376 , n94375 , n94372 );
and ( n94377 , n56946 , n52764 );
or ( n94378 , n94376 , n94377 );
and ( n94379 , n94374 , n94378 );
and ( n94380 , n56954 , n52762 );
or ( n94381 , n94379 , n94380 );
and ( n94382 , n94381 , n31452 );
or ( n94383 , n94373 , n94382 );
and ( n94384 , n94383 , n31638 );
and ( n94385 , n31108 , n47277 );
or ( n94386 , C0 , n94354 , n94363 , n94384 , n94385 );
buf ( n94387 , n94386 );
buf ( n94388 , n94387 );
buf ( n94389 , n30987 );
buf ( n94390 , n67631 );
buf ( n94391 , n79276 );
or ( n94392 , n94390 , n94391 , C0 , C0 );
and ( n94393 , n94392 , n67665 );
buf ( n94394 , n67631 );
buf ( n94395 , n79276 );
or ( n94396 , C0 , n94394 , n94395 , C0 , C0 );
and ( n94397 , n94396 , n67701 );
buf ( n94398 , n67631 );
buf ( n94399 , n79276 );
buf ( n94400 , n67668 );
or ( n94401 , C0 , n94398 , n94399 , C0 , n94400 );
and ( n94402 , n94401 , n67737 );
or ( n94403 , C0 , n94393 , n94397 , n94402 );
buf ( n94404 , n94403 );
buf ( n94405 , n94404 );
buf ( n94406 , n31655 );
and ( n94407 , n49087 , n48639 );
not ( n94408 , n48642 );
and ( n94409 , n94408 , n48608 );
and ( n94410 , n49087 , n48642 );
or ( n94411 , n94409 , n94410 );
and ( n94412 , n94411 , n32890 );
not ( n94413 , n48648 );
and ( n94414 , n94413 , n48608 );
and ( n94415 , n49087 , n48648 );
or ( n94416 , n94414 , n94415 );
and ( n94417 , n94416 , n32924 );
not ( n94418 , n48654 );
and ( n94419 , n94418 , n48608 );
and ( n94420 , n49087 , n48654 );
or ( n94421 , n94419 , n94420 );
and ( n94422 , n94421 , n33038 );
not ( n94423 , n48660 );
and ( n94424 , n94423 , n48608 );
and ( n94425 , n49087 , n48660 );
or ( n94426 , n94424 , n94425 );
and ( n94427 , n94426 , n33172 );
not ( n94428 , n41576 );
and ( n94429 , n94428 , n48608 );
and ( n94430 , n48904 , n41576 );
or ( n94431 , n94429 , n94430 );
and ( n94432 , n94431 , n33189 );
not ( n94433 , n48730 );
and ( n94434 , n94433 , n48608 );
and ( n94435 , n48904 , n48730 );
or ( n94436 , n94434 , n94435 );
and ( n94437 , n94436 , n33187 );
not ( n94438 , n48765 );
and ( n94439 , n94438 , n48608 );
and ( n94440 , n90384 , n48765 );
or ( n94441 , n94439 , n94440 );
and ( n94442 , n94441 , n33180 );
not ( n94443 , n49054 );
and ( n94444 , n94443 , n48608 );
and ( n94445 , n90397 , n49054 );
or ( n94446 , n94444 , n94445 );
and ( n94447 , n94446 , n33178 );
and ( n94448 , n49204 , n49275 );
or ( n94449 , n94407 , n94412 , n94417 , n94422 , n94427 , n94432 , n94437 , n94442 , n94447 , n94448 );
and ( n94450 , n94449 , n33208 );
and ( n94451 , n33001 , n35056 );
and ( n94452 , n48608 , n49286 );
or ( n94453 , C0 , n94450 , n94451 , n94452 );
buf ( n94454 , n94453 );
buf ( n94455 , n94454 );
buf ( n94456 , n30987 );
buf ( n94457 , n30987 );
buf ( n94458 , n31655 );
buf ( n94459 , n31655 );
and ( n94460 , n77648 , n33377 );
not ( n94461 , n48545 );
and ( n94462 , n94461 , n88453 );
buf ( n94463 , n94462 );
and ( n94464 , n94463 , n32890 );
not ( n94465 , n48557 );
and ( n94466 , n94465 , n88453 );
and ( n94467 , n77654 , n48557 );
or ( n94468 , n94466 , n94467 );
and ( n94469 , n94468 , n33038 );
and ( n94470 , n88453 , n48571 );
or ( n94471 , n94464 , n94469 , n94470 );
and ( n94472 , n94471 , n33208 );
and ( n94473 , n88453 , n48577 );
or ( n94474 , C0 , n94460 , n94472 , n94473 );
buf ( n94475 , n94474 );
buf ( n94476 , n94475 );
buf ( n94477 , n31655 );
buf ( n94478 , n30987 );
buf ( n94479 , n30987 );
buf ( n94480 , n31655 );
buf ( n94481 , n31655 );
buf ( n94482 , n31655 );
not ( n94483 , n33419 );
and ( n94484 , n94483 , n31578 );
and ( n94485 , n93805 , n33419 );
or ( n94486 , n94484 , n94485 );
and ( n94487 , n94486 , n31529 );
not ( n94488 , n33734 );
and ( n94489 , n94488 , n31578 );
and ( n94490 , n93816 , n33734 );
or ( n94491 , n94489 , n94490 );
and ( n94492 , n94491 , n31527 );
and ( n94493 , n31578 , n33942 );
or ( n94494 , n94487 , n94492 , n94493 );
and ( n94495 , n94494 , n31557 );
and ( n94496 , n34101 , n31643 );
not ( n94497 , n31452 );
and ( n94498 , n94497 , n34101 );
xor ( n94499 , n31578 , n33959 );
and ( n94500 , n94499 , n31452 );
or ( n94501 , n94498 , n94500 );
and ( n94502 , n94501 , n31638 );
and ( n94503 , n34002 , n33973 );
and ( n94504 , n31578 , n33978 );
or ( n94505 , C0 , n94495 , n94496 , n94502 , n94503 , n94504 );
buf ( n94506 , n94505 );
buf ( n94507 , n94506 );
and ( n94508 , n31566 , n31007 );
not ( n94509 , n31077 );
and ( n94510 , n94509 , n35392 );
buf ( n94511 , n94510 );
and ( n94512 , n94511 , n31373 );
not ( n94513 , n31402 );
and ( n94514 , n94513 , n35392 );
buf ( n94515 , n94514 );
and ( n94516 , n94515 , n31408 );
not ( n94517 , n31437 );
and ( n94518 , n94517 , n35392 );
not ( n94519 , n31455 );
and ( n94520 , n94519 , n35433 );
xor ( n94521 , n35392 , n35406 );
and ( n94522 , n94521 , n31455 );
xor ( n94523 , n94520 , n94522 );
and ( n94524 , n94523 , n31437 );
xor ( n94525 , n94518 , n94524 );
and ( n94526 , n94525 , n31468 );
not ( n94527 , n31497 );
and ( n94528 , n94527 , n35392 );
not ( n94529 , n31454 );
not ( n94530 , n31501 );
and ( n94531 , n94530 , n35433 );
xor ( n94532 , n35434 , n35456 );
and ( n94533 , n94532 , n31501 );
or ( n94534 , n94531 , n94533 );
and ( n94535 , n94529 , n94534 );
and ( n94536 , n94521 , n31454 );
or ( n94537 , n94535 , n94536 );
and ( n94538 , n94537 , n31497 );
or ( n94539 , n94528 , n94538 );
and ( n94540 , n94539 , n31521 );
and ( n94541 , n35392 , n31553 );
or ( n94542 , n94512 , n94516 , n94526 , n94540 , n94541 );
and ( n94543 , n94542 , n31557 );
not ( n94544 , n31452 );
not ( n94545 , n31619 );
and ( n94546 , n94545 , n35488 );
xor ( n94547 , n35489 , n35510 );
and ( n94548 , n94547 , n31619 );
or ( n94549 , n94546 , n94548 );
and ( n94550 , n94544 , n94549 );
and ( n94551 , n35392 , n31452 );
or ( n94552 , n94550 , n94551 );
and ( n94553 , n94552 , n31638 );
and ( n94554 , n35392 , n31650 );
or ( n94555 , C0 , n94508 , n94543 , n94553 , C0 , n94554 );
buf ( n94556 , n94555 );
buf ( n94557 , n94556 );
buf ( n94558 , n30987 );
buf ( n94559 , n30987 );
buf ( n94560 , n31655 );
not ( n94561 , n36587 );
and ( n94562 , n94561 , n36549 );
xor ( n94563 , n61939 , n61946 );
and ( n94564 , n94563 , n36587 );
or ( n94565 , n94562 , n94564 );
and ( n94566 , n94565 , n36596 );
not ( n94567 , n37485 );
and ( n94568 , n94567 , n37451 );
xor ( n94569 , n61955 , n61962 );
and ( n94570 , n94569 , n37485 );
or ( n94571 , n94568 , n94570 );
and ( n94572 , n94571 , n37494 );
and ( n94573 , n41866 , n37506 );
or ( n94574 , n94566 , n94572 , n94573 );
buf ( n94575 , n94574 );
buf ( n94576 , n94575 );
and ( n94577 , n47659 , n50275 );
not ( n94578 , n50278 );
and ( n94579 , n94578 , n47572 );
and ( n94580 , n47659 , n50278 );
or ( n94581 , n94579 , n94580 );
and ( n94582 , n94581 , n32421 );
not ( n94583 , n50002 );
and ( n94584 , n94583 , n47572 );
and ( n94585 , n47659 , n50002 );
or ( n94586 , n94584 , n94585 );
and ( n94587 , n94586 , n32419 );
not ( n94588 , n50289 );
and ( n94589 , n94588 , n47572 );
and ( n94590 , n47659 , n50289 );
or ( n94591 , n94589 , n94590 );
and ( n94592 , n94591 , n32417 );
not ( n94593 , n50008 );
and ( n94594 , n94593 , n47572 );
and ( n94595 , n47659 , n50008 );
or ( n94596 , n94594 , n94595 );
and ( n94597 , n94596 , n32415 );
not ( n94598 , n47331 );
and ( n94599 , n94598 , n47572 );
and ( n94600 , n47604 , n47331 );
or ( n94601 , n94599 , n94600 );
and ( n94602 , n94601 , n32413 );
not ( n94603 , n50067 );
and ( n94604 , n94603 , n47572 );
and ( n94605 , n47604 , n50067 );
or ( n94606 , n94604 , n94605 );
and ( n94607 , n94606 , n32411 );
not ( n94608 , n31728 );
and ( n94609 , n94608 , n47572 );
and ( n94610 , n76883 , n31728 );
or ( n94611 , n94609 , n94610 );
and ( n94612 , n94611 , n32253 );
not ( n94613 , n32283 );
and ( n94614 , n94613 , n47572 );
and ( n94615 , n76894 , n32283 );
or ( n94616 , n94614 , n94615 );
and ( n94617 , n94616 , n32398 );
and ( n94618 , n47709 , n50334 );
or ( n94619 , n94577 , n94582 , n94587 , n94592 , n94597 , n94602 , n94607 , n94612 , n94617 , n94618 );
and ( n94620 , n94619 , n32456 );
and ( n94621 , n37551 , n32489 );
and ( n94622 , n47572 , n50345 );
or ( n94623 , C0 , n94620 , n94621 , n94622 );
buf ( n94624 , n94623 );
buf ( n94625 , n94624 );
buf ( n94626 , n30987 );
buf ( n94627 , n30987 );
not ( n94628 , n34150 );
and ( n94629 , n94628 , n32836 );
not ( n94630 , n57872 );
and ( n94631 , n94630 , n32836 );
and ( n94632 , n32856 , n57872 );
or ( n94633 , n94631 , n94632 );
and ( n94634 , n94633 , n34150 );
or ( n94635 , n94629 , n94634 );
and ( n94636 , n94635 , n33381 );
not ( n94637 , n57880 );
not ( n94638 , n57872 );
and ( n94639 , n94638 , n32836 );
and ( n94640 , n48160 , n57872 );
or ( n94641 , n94639 , n94640 );
and ( n94642 , n94637 , n94641 );
and ( n94643 , n48160 , n57880 );
or ( n94644 , n94642 , n94643 );
and ( n94645 , n94644 , n33375 );
not ( n94646 , n32968 );
not ( n94647 , n57880 );
not ( n94648 , n57872 );
and ( n94649 , n94648 , n32836 );
and ( n94650 , n48160 , n57872 );
or ( n94651 , n94649 , n94650 );
and ( n94652 , n94647 , n94651 );
and ( n94653 , n48160 , n57880 );
or ( n94654 , n94652 , n94653 );
and ( n94655 , n94646 , n94654 );
not ( n94656 , n57900 );
not ( n94657 , n57902 );
and ( n94658 , n94657 , n94654 );
and ( n94659 , n48186 , n57902 );
or ( n94660 , n94658 , n94659 );
and ( n94661 , n94656 , n94660 );
and ( n94662 , n48196 , n57900 );
or ( n94663 , n94661 , n94662 );
and ( n94664 , n94663 , n32968 );
or ( n94665 , n94655 , n94664 );
and ( n94666 , n94665 , n33370 );
and ( n94667 , n32836 , n35062 );
or ( n94668 , C0 , n94636 , n94645 , n94666 , n94667 );
buf ( n94669 , n94668 );
buf ( n94670 , n94669 );
buf ( n94671 , n30987 );
buf ( n94672 , n31655 );
buf ( n94673 , n31655 );
buf ( n94674 , n31655 );
and ( n94675 , n33783 , n48455 );
not ( n94676 , n48457 );
and ( n94677 , n94676 , n33442 );
and ( n94678 , n33783 , n48457 );
or ( n94679 , n94677 , n94678 );
and ( n94680 , n94679 , n31373 );
not ( n94681 , n44807 );
and ( n94682 , n94681 , n33442 );
and ( n94683 , n33783 , n44807 );
or ( n94684 , n94682 , n94683 );
and ( n94685 , n94684 , n31408 );
not ( n94686 , n48468 );
and ( n94687 , n94686 , n33442 );
and ( n94688 , n33783 , n48468 );
or ( n94689 , n94687 , n94688 );
and ( n94690 , n94689 , n31468 );
not ( n94691 , n44817 );
and ( n94692 , n94691 , n33442 );
and ( n94693 , n33783 , n44817 );
or ( n94694 , n94692 , n94693 );
and ( n94695 , n94694 , n31521 );
not ( n94696 , n39979 );
and ( n94697 , n94696 , n33442 );
and ( n94698 , n33630 , n39979 );
or ( n94699 , n94697 , n94698 );
and ( n94700 , n94699 , n31538 );
not ( n94701 , n45059 );
and ( n94702 , n94701 , n33442 );
and ( n94703 , n33630 , n45059 );
or ( n94704 , n94702 , n94703 );
and ( n94705 , n94704 , n31536 );
not ( n94706 , n33419 );
and ( n94707 , n94706 , n33442 );
and ( n94708 , n88918 , n33419 );
or ( n94709 , n94707 , n94708 );
and ( n94710 , n94709 , n31529 );
not ( n94711 , n33734 );
and ( n94712 , n94711 , n33442 );
and ( n94713 , n88931 , n33734 );
or ( n94714 , n94712 , n94713 );
and ( n94715 , n94714 , n31527 );
and ( n94716 , n33880 , n48513 );
or ( n94717 , n94675 , n94680 , n94685 , n94690 , n94695 , n94700 , n94705 , n94710 , n94715 , n94716 );
and ( n94718 , n94717 , n31557 );
and ( n94719 , n31460 , n33973 );
and ( n94720 , n33442 , n48524 );
or ( n94721 , C0 , n94718 , n94719 , n94720 );
buf ( n94722 , n94721 );
buf ( n94723 , n94722 );
buf ( n94724 , n30987 );
not ( n94725 , n35278 );
and ( n94726 , n94725 , n63555 );
and ( n94727 , n63568 , n35278 );
or ( n94728 , n94726 , n94727 );
and ( n94729 , n94728 , n32417 );
not ( n94730 , n50008 );
and ( n94731 , n94730 , n63555 );
and ( n94732 , n77583 , n50008 );
or ( n94733 , n94731 , n94732 );
and ( n94734 , n94733 , n32415 );
and ( n94735 , n63555 , n48133 );
or ( n94736 , n94729 , n94734 , n94735 );
and ( n94737 , n94736 , n32456 );
and ( n94738 , n63555 , n47409 );
or ( n94739 , C0 , n94737 , n94738 );
buf ( n94740 , n94739 );
buf ( n94741 , n94740 );
buf ( n94742 , n30987 );
not ( n94743 , n68284 );
not ( n94744 , n68286 );
not ( n94745 , n68289 );
and ( n94746 , n94745 , n68293 );
buf ( n94747 , n68289 );
or ( n94748 , n94746 , n94747 );
and ( n94749 , n94744 , n94748 );
buf ( n94750 , n94749 );
and ( n94751 , n94743 , n94750 );
buf ( n94752 , n68284 );
or ( n94753 , n94751 , n94752 );
and ( n94754 , n94753 , n44694 );
and ( n94755 , n57860 , n43774 );
and ( n94756 , n68304 , n44692 );
not ( n94757 , n68313 );
not ( n94758 , n68316 );
and ( n94759 , n94758 , n48294 );
buf ( n94760 , n68316 );
or ( n94761 , n94759 , n94760 );
and ( n94762 , n94757 , n94761 );
buf ( n94763 , n68313 );
or ( n94764 , n94762 , n94763 );
and ( n94765 , n94764 , n44690 );
not ( n94766 , n68289 );
not ( n94767 , n68327 );
not ( n94768 , n68331 );
not ( n94769 , n68334 );
not ( n94770 , n68336 );
not ( n94771 , n68338 );
and ( n94772 , n94770 , n94771 );
buf ( n94773 , n94772 );
and ( n94774 , n94769 , n94773 );
buf ( n94775 , n68334 );
or ( n94776 , n94774 , n94775 );
and ( n94777 , n94768 , n94776 );
buf ( n94778 , n68331 );
or ( n94779 , n94777 , n94778 );
and ( n94780 , n94767 , n94779 );
and ( n94781 , n32957 , n68327 );
or ( n94782 , n94780 , n94781 );
and ( n94783 , n94766 , n94782 );
buf ( n94784 , n68289 );
or ( n94785 , n94783 , n94784 );
and ( n94786 , n94785 , n44688 );
buf ( n94787 , n44682 );
and ( n94788 , n68281 , n44685 );
or ( n94789 , n94754 , n94755 , n94756 , n94765 , n94786 , n94787 , n94788 , C0 );
buf ( n94790 , n94789 );
buf ( n94791 , n94790 );
buf ( n94792 , n31655 );
buf ( n94793 , n30987 );
buf ( n94794 , n31655 );
buf ( n94795 , n31655 );
buf ( n94796 , n30987 );
and ( n94797 , n79986 , n33377 );
not ( n94798 , n48545 );
and ( n94799 , n94798 , n80472 );
and ( n94800 , n79992 , n48545 );
or ( n94801 , n94799 , n94800 );
and ( n94802 , n94801 , n32890 );
not ( n94803 , n48557 );
and ( n94804 , n94803 , n80472 );
and ( n94805 , n79992 , n48557 );
or ( n94806 , n94804 , n94805 );
and ( n94807 , n94806 , n33038 );
and ( n94808 , n80472 , n48571 );
or ( n94809 , n94802 , n94807 , n94808 );
and ( n94810 , n94809 , n33208 );
and ( n94811 , n80472 , n48577 );
or ( n94812 , C0 , n94797 , n94810 , n94811 );
buf ( n94813 , n94812 );
buf ( n94814 , n94813 );
buf ( n94815 , n30987 );
buf ( n94816 , n31655 );
buf ( n94817 , n30987 );
and ( n94818 , n86492 , n33377 );
not ( n94819 , n48545 );
and ( n94820 , n94819 , n83086 );
and ( n94821 , n90362 , n48545 );
or ( n94822 , n94820 , n94821 );
and ( n94823 , n94822 , n32890 );
not ( n94824 , n48557 );
and ( n94825 , n94824 , n83086 );
and ( n94826 , n90362 , n48557 );
or ( n94827 , n94825 , n94826 );
and ( n94828 , n94827 , n33038 );
and ( n94829 , n83086 , n48571 );
or ( n94830 , n94823 , n94828 , n94829 );
and ( n94831 , n94830 , n33208 );
and ( n94832 , n83086 , n48577 );
or ( n94833 , C0 , n94818 , n94831 , n94832 );
buf ( n94834 , n94833 );
buf ( n94835 , n94834 );
buf ( n94836 , n31655 );
buf ( n94837 , n30987 );
buf ( n94838 , n31655 );
buf ( n94839 , n31655 );
buf ( n94840 , n31655 );
not ( n94841 , n33419 );
and ( n94842 , n94841 , n31573 );
and ( n94843 , n69979 , n33419 );
or ( n94844 , n94842 , n94843 );
and ( n94845 , n94844 , n31529 );
not ( n94846 , n33734 );
and ( n94847 , n94846 , n31573 );
and ( n94848 , n69990 , n33734 );
or ( n94849 , n94847 , n94848 );
and ( n94850 , n94849 , n31527 );
and ( n94851 , n31573 , n33942 );
or ( n94852 , n94845 , n94850 , n94851 );
and ( n94853 , n94852 , n31557 );
and ( n94854 , n35501 , n31643 );
not ( n94855 , n31452 );
and ( n94856 , n94855 , n35501 );
or ( n94857 , n31573 , n33964 );
and ( n94858 , n94857 , n31452 );
or ( n94859 , n94856 , n94858 );
and ( n94860 , n94859 , n31638 );
and ( n94861 , n35398 , n33973 );
and ( n94862 , n31573 , n33978 );
or ( n94863 , C0 , n94853 , n94854 , n94860 , n94861 , n94862 );
buf ( n94864 , n94863 );
buf ( n94865 , n94864 );
and ( n94866 , n31571 , n31007 );
not ( n94867 , n31077 );
and ( n94868 , n94867 , n35396 );
buf ( n94869 , n94868 );
and ( n94870 , n94869 , n31373 );
not ( n94871 , n31402 );
and ( n94872 , n94871 , n35396 );
buf ( n94873 , n94872 );
and ( n94874 , n94873 , n31408 );
not ( n94875 , n31437 );
and ( n94876 , n94875 , n35396 );
not ( n94877 , n31455 );
and ( n94878 , n94877 , n35443 );
xor ( n94879 , n35396 , n35401 );
and ( n94880 , n94879 , n31455 );
or ( n94881 , n94878 , n94880 );
and ( n94882 , n94881 , n31437 );
or ( n94883 , n94876 , n94882 );
and ( n94884 , n94883 , n31468 );
not ( n94885 , n31497 );
and ( n94886 , n94885 , n35396 );
not ( n94887 , n31454 );
not ( n94888 , n31501 );
and ( n94889 , n94888 , n35443 );
xor ( n94890 , n35444 , n35451 );
and ( n94891 , n94890 , n31501 );
or ( n94892 , n94889 , n94891 );
and ( n94893 , n94887 , n94892 );
and ( n94894 , n94879 , n31454 );
or ( n94895 , n94893 , n94894 );
and ( n94896 , n94895 , n31497 );
or ( n94897 , n94886 , n94896 );
and ( n94898 , n94897 , n31521 );
and ( n94899 , n35396 , n31553 );
or ( n94900 , n94870 , n94874 , n94884 , n94898 , n94899 );
and ( n94901 , n94900 , n31557 );
not ( n94902 , n31452 );
not ( n94903 , n31619 );
and ( n94904 , n94903 , n35497 );
xor ( n94905 , n35498 , n35505 );
and ( n94906 , n94905 , n31619 );
or ( n94907 , n94904 , n94906 );
and ( n94908 , n94902 , n94907 );
and ( n94909 , n35396 , n31452 );
or ( n94910 , n94908 , n94909 );
and ( n94911 , n94910 , n31638 );
and ( n94912 , n35396 , n31650 );
or ( n94913 , C0 , n94866 , n94901 , n94911 , C0 , n94912 );
buf ( n94914 , n94913 );
buf ( n94915 , n94914 );
buf ( n94916 , n30987 );
buf ( n94917 , n30987 );
buf ( n94918 , n31655 );
not ( n94919 , n35542 );
and ( n94920 , n94919 , n41859 );
and ( n94921 , n93522 , n35542 );
or ( n94922 , n94920 , n94921 );
buf ( n94923 , n94922 );
buf ( n94924 , n94923 );
not ( n94925 , n46356 );
and ( n94926 , n94925 , n31164 );
not ( n94927 , n49427 );
and ( n94928 , n94927 , n31164 );
and ( n94929 , n31172 , n49427 );
or ( n94930 , n94928 , n94929 );
and ( n94931 , n94930 , n46356 );
or ( n94932 , n94926 , n94931 );
and ( n94933 , n94932 , n31649 );
not ( n94934 , n49435 );
not ( n94935 , n49427 );
and ( n94936 , n94935 , n31164 );
and ( n94937 , n46495 , n49427 );
or ( n94938 , n94936 , n94937 );
and ( n94939 , n94934 , n94938 );
and ( n94940 , n46495 , n49435 );
or ( n94941 , n94939 , n94940 );
and ( n94942 , n94941 , n31643 );
not ( n94943 , n31452 );
not ( n94944 , n49435 );
not ( n94945 , n49427 );
and ( n94946 , n94945 , n31164 );
and ( n94947 , n46495 , n49427 );
or ( n94948 , n94946 , n94947 );
and ( n94949 , n94944 , n94948 );
and ( n94950 , n46495 , n49435 );
or ( n94951 , n94949 , n94950 );
and ( n94952 , n94943 , n94951 );
not ( n94953 , n49460 );
not ( n94954 , n49462 );
and ( n94955 , n94954 , n94951 );
and ( n94956 , n46984 , n49462 );
or ( n94957 , n94955 , n94956 );
and ( n94958 , n94953 , n94957 );
and ( n94959 , n47267 , n49460 );
or ( n94960 , n94958 , n94959 );
and ( n94961 , n94960 , n31452 );
or ( n94962 , n94952 , n94961 );
and ( n94963 , n94962 , n31638 );
and ( n94964 , n31164 , n47277 );
or ( n94965 , C0 , n94933 , n94942 , n94963 , n94964 );
buf ( n94966 , n94965 );
buf ( n94967 , n94966 );
buf ( n94968 , n30987 );
xor ( n94969 , n47286 , n47296 );
and ( n94970 , n94969 , n32433 );
not ( n94971 , n47331 );
and ( n94972 , n94971 , n47286 );
buf ( n94973 , n31820 );
and ( n94974 , n94973 , n47331 );
or ( n94975 , n94972 , n94974 );
and ( n94976 , n94975 , n32413 );
and ( n94977 , n47286 , n47402 );
or ( n94978 , n94970 , n94976 , n94977 );
and ( n94979 , n94978 , n32456 );
and ( n94980 , n47286 , n47409 );
or ( n94981 , C0 , n94979 , n94980 );
buf ( n94982 , n94981 );
buf ( n94983 , n94982 );
buf ( n94984 , n31655 );
buf ( n94985 , n30987 );
buf ( n94986 , n30987 );
not ( n94987 , n43755 );
and ( n94988 , n94987 , n43411 );
xor ( n94989 , n50500 , n50505 );
and ( n94990 , n94989 , n43755 );
or ( n94991 , n94988 , n94990 );
and ( n94992 , n94991 , n43774 );
not ( n94993 , n44663 );
and ( n94994 , n94993 , n44323 );
xor ( n94995 , n50518 , n50523 );
and ( n94996 , n94995 , n44663 );
or ( n94997 , n94994 , n94996 );
and ( n94998 , n94997 , n44682 );
and ( n94999 , n61073 , n44695 );
or ( n95000 , n94992 , n94998 , n94999 );
buf ( n95001 , n95000 );
buf ( n95002 , n95001 );
buf ( n95003 , n31655 );
buf ( n95004 , n31655 );
buf ( n95005 , n31655 );
buf ( n95006 , n30987 );
not ( n95007 , n48765 );
and ( n95008 , n95007 , n33232 );
xor ( n95009 , n48787 , n49001 );
and ( n95010 , n95009 , n48765 );
or ( n95011 , n95008 , n95010 );
and ( n95012 , n95011 , n33180 );
not ( n95013 , n49054 );
and ( n95014 , n95013 , n33232 );
not ( n95015 , n48845 );
xor ( n95016 , n49077 , n49115 );
and ( n95017 , n95015 , n95016 );
xnor ( n95018 , n49186 , n49241 );
and ( n95019 , n95018 , n48845 );
or ( n95020 , n95017 , n95019 );
and ( n95021 , n95020 , n49054 );
or ( n95022 , n95014 , n95021 );
and ( n95023 , n95022 , n33178 );
and ( n95024 , n33232 , n49774 );
or ( n95025 , n95012 , n95023 , n95024 );
and ( n95026 , n95025 , n33208 );
and ( n95027 , n33315 , n33375 );
not ( n95028 , n32968 );
and ( n95029 , n95028 , n33315 );
xor ( n95030 , n33232 , n53897 );
and ( n95031 , n95030 , n32968 );
or ( n95032 , n95029 , n95031 );
and ( n95033 , n95032 , n33370 );
and ( n95034 , n32995 , n35056 );
and ( n95035 , n33232 , n49794 );
or ( n95036 , C0 , n95026 , n95027 , n95033 , n95034 , n95035 );
buf ( n95037 , n95036 );
buf ( n95038 , n95037 );
buf ( n95039 , n30987 );
buf ( n95040 , n31655 );
and ( n95041 , n46018 , n32500 );
not ( n95042 , n35211 );
and ( n95043 , n95042 , n37533 );
buf ( n95044 , n95043 );
and ( n95045 , n95044 , n32421 );
not ( n95046 , n35245 );
and ( n95047 , n95046 , n37533 );
buf ( n95048 , n95047 );
and ( n95049 , n95048 , n32419 );
not ( n95050 , n35278 );
and ( n95051 , n95050 , n37533 );
not ( n95052 , n35295 );
and ( n95053 , n95052 , n49563 );
xor ( n95054 , n37533 , n49549 );
and ( n95055 , n95054 , n35295 );
or ( n95056 , n95053 , n95055 );
and ( n95057 , n95056 , n35278 );
or ( n95058 , n95051 , n95057 );
and ( n95059 , n95058 , n32417 );
not ( n95060 , n35331 );
and ( n95061 , n95060 , n37533 );
not ( n95062 , n35294 );
not ( n95063 , n45995 );
and ( n95064 , n95063 , n49563 );
xor ( n95065 , n49564 , n49635 );
and ( n95066 , n95065 , n45995 );
or ( n95067 , n95064 , n95066 );
and ( n95068 , n95062 , n95067 );
and ( n95069 , n95054 , n35294 );
or ( n95070 , n95068 , n95069 );
and ( n95071 , n95070 , n35331 );
or ( n95072 , n95061 , n95071 );
and ( n95073 , n95072 , n32415 );
and ( n95074 , n37533 , n35354 );
or ( n95075 , n95045 , n95049 , n95059 , n95073 , n95074 );
and ( n95076 , n95075 , n32456 );
not ( n95077 , n32475 );
not ( n95078 , n46060 );
and ( n95079 , n95078 , n49654 );
xor ( n95080 , n49655 , n49729 );
and ( n95081 , n95080 , n46060 );
or ( n95082 , n95079 , n95081 );
and ( n95083 , n95077 , n95082 );
and ( n95084 , n37533 , n32475 );
or ( n95085 , n95083 , n95084 );
and ( n95086 , n95085 , n32486 );
and ( n95087 , n37533 , n35367 );
or ( n95088 , C0 , n95041 , n95076 , n95086 , C0 , n95087 );
buf ( n95089 , n95088 );
buf ( n95090 , n95089 );
buf ( n95091 , n31655 );
not ( n95092 , n46356 );
and ( n95093 , n95092 , n31250 );
not ( n95094 , n53353 );
and ( n95095 , n95094 , n31250 );
and ( n95096 , n31272 , n53353 );
or ( n95097 , n95095 , n95096 );
and ( n95098 , n95097 , n46356 );
or ( n95099 , n95093 , n95098 );
and ( n95100 , n95099 , n31649 );
not ( n95101 , n53361 );
not ( n95102 , n53353 );
and ( n95103 , n95102 , n31250 );
and ( n95104 , n49443 , n53353 );
or ( n95105 , n95103 , n95104 );
and ( n95106 , n95101 , n95105 );
and ( n95107 , n49443 , n53361 );
or ( n95108 , n95106 , n95107 );
and ( n95109 , n95108 , n31643 );
not ( n95110 , n31452 );
not ( n95111 , n53361 );
not ( n95112 , n53353 );
and ( n95113 , n95112 , n31250 );
and ( n95114 , n49443 , n53353 );
or ( n95115 , n95113 , n95114 );
and ( n95116 , n95111 , n95115 );
and ( n95117 , n49443 , n53361 );
or ( n95118 , n95116 , n95117 );
and ( n95119 , n95110 , n95118 );
not ( n95120 , n53381 );
not ( n95121 , n53383 );
and ( n95122 , n95121 , n95118 );
and ( n95123 , n49469 , n53383 );
or ( n95124 , n95122 , n95123 );
and ( n95125 , n95120 , n95124 );
and ( n95126 , n49477 , n53381 );
or ( n95127 , n95125 , n95126 );
and ( n95128 , n95127 , n31452 );
or ( n95129 , n95119 , n95128 );
and ( n95130 , n95129 , n31638 );
and ( n95131 , n31250 , n47277 );
or ( n95132 , C0 , n95100 , n95109 , n95130 , n95131 );
buf ( n95133 , n95132 );
buf ( n95134 , n95133 );
buf ( n95135 , n30987 );
and ( n95136 , n78780 , n32494 );
not ( n95137 , n46083 );
and ( n95138 , n95137 , n52211 );
buf ( n95139 , n95138 );
and ( n95140 , n95139 , n32421 );
not ( n95141 , n46326 );
and ( n95142 , n95141 , n52211 );
and ( n95143 , n78786 , n46326 );
or ( n95144 , n95142 , n95143 );
and ( n95145 , n95144 , n32417 );
and ( n95146 , n52211 , n46340 );
or ( n95147 , n95140 , n95145 , n95146 );
and ( n95148 , n95147 , n32456 );
and ( n95149 , n52211 , n46349 );
or ( n95150 , C0 , n95136 , n95148 , n95149 );
buf ( n95151 , n95150 );
buf ( n95152 , n95151 );
buf ( n95153 , n31655 );
buf ( n95154 , n30987 );
buf ( n95155 , n31655 );
and ( n95156 , n61232 , n33377 );
not ( n95157 , n48545 );
and ( n95158 , n95157 , n53870 );
and ( n95159 , n61238 , n48545 );
or ( n95160 , n95158 , n95159 );
and ( n95161 , n95160 , n32890 );
not ( n95162 , n48557 );
and ( n95163 , n95162 , n53870 );
and ( n95164 , n61238 , n48557 );
or ( n95165 , n95163 , n95164 );
and ( n95166 , n95165 , n33038 );
and ( n95167 , n53870 , n48571 );
or ( n95168 , n95161 , n95166 , n95167 );
and ( n95169 , n95168 , n33208 );
and ( n95170 , n53870 , n48577 );
or ( n95171 , C0 , n95156 , n95169 , n95170 );
buf ( n95172 , n95171 );
buf ( n95173 , n95172 );
buf ( n95174 , n30987 );
buf ( n95175 , n31655 );
buf ( n95176 , n31655 );
buf ( n95177 , n40221 );
not ( n95178 , n46356 );
and ( n95179 , n95178 , n31162 );
not ( n95180 , n56904 );
and ( n95181 , n95180 , n31162 );
and ( n95182 , n31172 , n56904 );
or ( n95183 , n95181 , n95182 );
and ( n95184 , n95183 , n46356 );
or ( n95185 , n95179 , n95184 );
and ( n95186 , n95185 , n31649 );
not ( n95187 , n56912 );
not ( n95188 , n56904 );
and ( n95189 , n95188 , n31162 );
and ( n95190 , n46495 , n56904 );
or ( n95191 , n95189 , n95190 );
and ( n95192 , n95187 , n95191 );
and ( n95193 , n46495 , n56912 );
or ( n95194 , n95192 , n95193 );
and ( n95195 , n95194 , n31643 );
not ( n95196 , n31452 );
not ( n95197 , n56912 );
not ( n95198 , n56904 );
and ( n95199 , n95198 , n31162 );
and ( n95200 , n46495 , n56904 );
or ( n95201 , n95199 , n95200 );
and ( n95202 , n95197 , n95201 );
and ( n95203 , n46495 , n56912 );
or ( n95204 , n95202 , n95203 );
and ( n95205 , n95196 , n95204 );
not ( n95206 , n56937 );
not ( n95207 , n56939 );
and ( n95208 , n95207 , n95204 );
and ( n95209 , n46984 , n56939 );
or ( n95210 , n95208 , n95209 );
and ( n95211 , n95206 , n95210 );
and ( n95212 , n47267 , n56937 );
or ( n95213 , n95211 , n95212 );
and ( n95214 , n95213 , n31452 );
or ( n95215 , n95205 , n95214 );
and ( n95216 , n95215 , n31638 );
and ( n95217 , n31162 , n47277 );
or ( n95218 , C0 , n95186 , n95195 , n95216 , n95217 );
buf ( n95219 , n95218 );
buf ( n95220 , n95219 );
buf ( n95221 , n30987 );
and ( n95222 , n50947 , n88642 );
xor ( n95223 , n46092 , n95222 );
and ( n95224 , n95223 , n32431 );
not ( n95225 , n50002 );
and ( n95226 , n95225 , n46092 );
and ( n95227 , n40244 , n50002 );
or ( n95228 , n95226 , n95227 );
and ( n95229 , n95228 , n32419 );
not ( n95230 , n50008 );
and ( n95231 , n95230 , n46092 );
buf ( n95232 , n95231 );
and ( n95233 , n95232 , n32415 );
not ( n95234 , n50067 );
and ( n95235 , n95234 , n46092 );
buf ( n95236 , n95235 );
and ( n95237 , n95236 , n32411 );
and ( n95238 , n46092 , n50098 );
or ( n95239 , n95224 , n95229 , n95233 , n95237 , n95238 );
and ( n95240 , n95239 , n32456 );
and ( n95241 , n46092 , n47409 );
or ( n95242 , C0 , n95240 , n95241 );
buf ( n95243 , n95242 );
buf ( n95244 , n95243 );
buf ( n95245 , n31655 );
buf ( n95246 , n30987 );
buf ( n95247 , n31655 );
xor ( n95248 , n39532 , n54976 );
and ( n95249 , n95248 , n33199 );
not ( n95250 , n48648 );
and ( n95251 , n95250 , n39532 );
and ( n95252 , n34369 , n48648 );
or ( n95253 , n95251 , n95252 );
and ( n95254 , n95253 , n32924 );
not ( n95255 , n48660 );
and ( n95256 , n95255 , n39532 );
not ( n95257 , n39584 );
and ( n95258 , n95257 , n79986 );
and ( n95259 , n80002 , n39584 );
or ( n95260 , n95258 , n95259 );
and ( n95261 , n95260 , n48660 );
or ( n95262 , n95256 , n95261 );
and ( n95263 , n95262 , n33172 );
not ( n95264 , n48730 );
and ( n95265 , n95264 , n39532 );
and ( n95266 , n71584 , n48730 );
or ( n95267 , n95265 , n95266 );
and ( n95268 , n95267 , n33187 );
and ( n95269 , n39532 , n54713 );
or ( n95270 , n95249 , n95254 , n95263 , n95268 , n95269 );
and ( n95271 , n95270 , n33208 );
and ( n95272 , n39532 , n39805 );
or ( n95273 , C0 , n95271 , n95272 );
buf ( n95274 , n95273 );
buf ( n95275 , n95274 );
buf ( n95276 , n30987 );
buf ( n95277 , n31655 );
not ( n95278 , n41532 );
and ( n95279 , n95278 , n34427 );
and ( n95280 , n45276 , n41532 );
or ( n95281 , n95279 , n95280 );
buf ( n95282 , n95281 );
buf ( n95283 , n95282 );
xor ( n95284 , n33117 , n52220 );
and ( n95285 , n95284 , n33201 );
not ( n95286 , n41576 );
and ( n95287 , n95286 , n33117 );
and ( n95288 , n87692 , n41576 );
or ( n95289 , n95287 , n95288 );
and ( n95290 , n95289 , n33189 );
and ( n95291 , n33117 , n41592 );
or ( n95292 , n95285 , n95290 , n95291 );
and ( n95293 , n95292 , n33208 );
and ( n95294 , n33117 , n39805 );
nor ( n95295 , C0 , n95293 , n95294 );
buf ( n95296 , n95295 );
buf ( n95297 , n95296 );
buf ( n95298 , n31655 );
buf ( n95299 , n30987 );
buf ( n95300 , n30987 );
buf ( n95301 , n31655 );
not ( n95302 , n50828 );
not ( n95303 , n50834 );
and ( n95304 , n95303 , n40555 );
and ( n95305 , n35533 , n50834 );
or ( n95306 , n95304 , n95305 );
and ( n95307 , n95302 , n95306 );
and ( n95308 , n35529 , n50828 );
or ( n95309 , n95307 , n95308 );
buf ( n95310 , n95309 );
buf ( n95311 , n95310 );
buf ( n95312 , n31655 );
xor ( n95313 , n33083 , n58392 );
and ( n95314 , n95313 , n33201 );
not ( n95315 , n41576 );
and ( n95316 , n95315 , n33083 );
xor ( n95317 , n58540 , n58593 );
and ( n95318 , n95317 , n41576 );
or ( n95319 , n95316 , n95318 );
and ( n95320 , n95319 , n33189 );
and ( n95321 , n33083 , n41592 );
or ( n95322 , n95314 , n95320 , n95321 );
and ( n95323 , n95322 , n33208 );
and ( n95324 , n33083 , n39805 );
or ( n95325 , C0 , n95323 , n95324 );
buf ( n95326 , n95325 );
buf ( n95327 , n95326 );
buf ( n95328 , n30987 );
buf ( n95329 , n30987 );
buf ( n95330 , n31655 );
not ( n95331 , n50828 );
not ( n95332 , n50834 );
and ( n95333 , n95332 , n40477 );
and ( n95334 , n83507 , n50834 );
or ( n95335 , n95333 , n95334 );
and ( n95336 , n95331 , n95335 );
and ( n95337 , n46085 , n50828 );
or ( n95338 , n95336 , n95337 );
buf ( n95339 , n95338 );
buf ( n95340 , n95339 );
buf ( n95341 , n30987 );
or ( n95342 , n44686 , n44688 );
or ( n95343 , n95342 , n44690 );
buf ( n95344 , n95343 );
or ( n95345 , n44685 , n44692 );
or ( n95346 , n95345 , n44694 );
and ( n95347 , n54724 , n95346 );
or ( n95348 , C0 , n95344 , n95347 );
buf ( n95349 , n95348 );
buf ( n95350 , n95349 );
buf ( n95351 , n30987 );
buf ( n95352 , n31655 );
buf ( n95353 , n31655 );
buf ( n95354 , n31655 );
not ( n95355 , n31437 );
and ( n95356 , n95355 , n45875 );
and ( n95357 , n45897 , n31437 );
or ( n95358 , n95356 , n95357 );
and ( n95359 , n95358 , n31468 );
not ( n95360 , n44817 );
and ( n95361 , n95360 , n45875 );
and ( n95362 , n80887 , n44817 );
or ( n95363 , n95361 , n95362 );
and ( n95364 , n95363 , n31521 );
and ( n95365 , n45875 , n42158 );
or ( n95366 , n95359 , n95364 , n95365 );
and ( n95367 , n95366 , n31557 );
and ( n95368 , n45875 , n40154 );
or ( n95369 , C0 , n95367 , n95368 );
buf ( n95370 , n95369 );
buf ( n95371 , n95370 );
not ( n95372 , n40163 );
and ( n95373 , n95372 , n31750 );
not ( n95374 , n56988 );
and ( n95375 , n95374 , n31750 );
and ( n95376 , n32252 , n56988 );
or ( n95377 , n95375 , n95376 );
and ( n95378 , n95377 , n40163 );
or ( n95379 , n95373 , n95378 );
and ( n95380 , n95379 , n32498 );
not ( n95381 , n56996 );
not ( n95382 , n56988 );
and ( n95383 , n95382 , n31750 );
and ( n95384 , n40393 , n56988 );
or ( n95385 , n95383 , n95384 );
and ( n95386 , n95381 , n95385 );
and ( n95387 , n40393 , n56996 );
or ( n95388 , n95386 , n95387 );
and ( n95389 , n95388 , n32473 );
not ( n95390 , n32475 );
not ( n95391 , n56996 );
not ( n95392 , n56988 );
and ( n95393 , n95392 , n31750 );
and ( n95394 , n40393 , n56988 );
or ( n95395 , n95393 , n95394 );
and ( n95396 , n95391 , n95395 );
and ( n95397 , n40393 , n56996 );
or ( n95398 , n95396 , n95397 );
and ( n95399 , n95390 , n95398 );
not ( n95400 , n57016 );
not ( n95401 , n57018 );
and ( n95402 , n95401 , n95398 );
and ( n95403 , n40972 , n57018 );
or ( n95404 , n95402 , n95403 );
and ( n95405 , n95400 , n95404 );
and ( n95406 , n41267 , n57016 );
or ( n95407 , n95405 , n95406 );
and ( n95408 , n95407 , n32475 );
or ( n95409 , n95399 , n95408 );
and ( n95410 , n95409 , n32486 );
and ( n95411 , n31750 , n41278 );
or ( n95412 , C0 , n95380 , n95389 , n95410 , n95411 );
buf ( n95413 , n95412 );
buf ( n95414 , n95413 );
buf ( n95415 , n30987 );
buf ( n95416 , n30987 );
buf ( n95417 , n31655 );
xor ( n95418 , n54148 , n78379 );
and ( n95419 , n95418 , n33199 );
not ( n95420 , n48648 );
and ( n95421 , n95420 , n54148 );
and ( n95422 , n34433 , n48648 );
or ( n95423 , n95421 , n95422 );
and ( n95424 , n95423 , n32924 );
not ( n95425 , n48660 );
and ( n95426 , n95425 , n54148 );
and ( n95427 , n64930 , n48660 );
or ( n95428 , n95426 , n95427 );
and ( n95429 , n95428 , n33172 );
not ( n95430 , n48730 );
and ( n95431 , n95430 , n54148 );
and ( n95432 , n66743 , n48730 );
or ( n95433 , n95431 , n95432 );
and ( n95434 , n95433 , n33187 );
and ( n95435 , n54148 , n54713 );
or ( n95436 , n95419 , n95424 , n95429 , n95434 , n95435 );
and ( n95437 , n95436 , n33208 );
and ( n95438 , n54148 , n39805 );
or ( n95439 , C0 , n95437 , n95438 );
buf ( n95440 , n95439 );
buf ( n95441 , n95440 );
buf ( n95442 , n30987 );
buf ( n95443 , n31655 );
not ( n95444 , n41532 );
and ( n95445 , n95444 , n34362 );
and ( n95446 , n66712 , n41532 );
or ( n95447 , n95445 , n95446 );
buf ( n95448 , n95447 );
buf ( n95449 , n95448 );
and ( n95450 , n49077 , n48639 );
not ( n95451 , n48642 );
and ( n95452 , n95451 , n48602 );
and ( n95453 , n49077 , n48642 );
or ( n95454 , n95452 , n95453 );
and ( n95455 , n95454 , n32890 );
not ( n95456 , n48648 );
and ( n95457 , n95456 , n48602 );
and ( n95458 , n49077 , n48648 );
or ( n95459 , n95457 , n95458 );
and ( n95460 , n95459 , n32924 );
not ( n95461 , n48654 );
and ( n95462 , n95461 , n48602 );
and ( n95463 , n49077 , n48654 );
or ( n95464 , n95462 , n95463 );
and ( n95465 , n95464 , n33038 );
not ( n95466 , n48660 );
and ( n95467 , n95466 , n48602 );
and ( n95468 , n49077 , n48660 );
or ( n95469 , n95467 , n95468 );
and ( n95470 , n95469 , n33172 );
not ( n95471 , n41576 );
and ( n95472 , n95471 , n48602 );
and ( n95473 , n48787 , n41576 );
or ( n95474 , n95472 , n95473 );
and ( n95475 , n95474 , n33189 );
not ( n95476 , n48730 );
and ( n95477 , n95476 , n48602 );
and ( n95478 , n48787 , n48730 );
or ( n95479 , n95477 , n95478 );
and ( n95480 , n95479 , n33187 );
not ( n95481 , n48765 );
and ( n95482 , n95481 , n48602 );
and ( n95483 , n95009 , n48765 );
or ( n95484 , n95482 , n95483 );
and ( n95485 , n95484 , n33180 );
not ( n95486 , n49054 );
and ( n95487 , n95486 , n48602 );
and ( n95488 , n95020 , n49054 );
or ( n95489 , n95487 , n95488 );
and ( n95490 , n95489 , n33178 );
and ( n95491 , n49186 , n49275 );
or ( n95492 , n95450 , n95455 , n95460 , n95465 , n95470 , n95475 , n95480 , n95485 , n95490 , n95491 );
and ( n95493 , n95492 , n33208 );
and ( n95494 , n32995 , n35056 );
and ( n95495 , n48602 , n49286 );
or ( n95496 , C0 , n95493 , n95494 , n95495 );
buf ( n95497 , n95496 );
buf ( n95498 , n95497 );
buf ( n95499 , n30987 );
buf ( n95500 , n30987 );
buf ( n95501 , n31655 );
buf ( n95502 , n31655 );
not ( n95503 , n46356 );
and ( n95504 , n95503 , n31203 );
not ( n95505 , n60564 );
and ( n95506 , n95505 , n31203 );
and ( n95507 , n31205 , n60564 );
or ( n95508 , n95506 , n95507 );
and ( n95509 , n95508 , n46356 );
or ( n95510 , n95504 , n95509 );
and ( n95511 , n95510 , n31649 );
not ( n95512 , n60572 );
not ( n95513 , n60564 );
and ( n95514 , n95513 , n31203 );
and ( n95515 , n50125 , n60564 );
or ( n95516 , n95514 , n95515 );
and ( n95517 , n95512 , n95516 );
and ( n95518 , n50125 , n60572 );
or ( n95519 , n95517 , n95518 );
and ( n95520 , n95519 , n31643 );
not ( n95521 , n31452 );
not ( n95522 , n60572 );
not ( n95523 , n60564 );
and ( n95524 , n95523 , n31203 );
and ( n95525 , n50125 , n60564 );
or ( n95526 , n95524 , n95525 );
and ( n95527 , n95522 , n95526 );
and ( n95528 , n50125 , n60572 );
or ( n95529 , n95527 , n95528 );
and ( n95530 , n95521 , n95529 );
not ( n95531 , n60592 );
not ( n95532 , n60594 );
and ( n95533 , n95532 , n95529 );
and ( n95534 , n50151 , n60594 );
or ( n95535 , n95533 , n95534 );
and ( n95536 , n95531 , n95535 );
and ( n95537 , n50159 , n60592 );
or ( n95538 , n95536 , n95537 );
and ( n95539 , n95538 , n31452 );
or ( n95540 , n95530 , n95539 );
and ( n95541 , n95540 , n31638 );
and ( n95542 , n31203 , n47277 );
or ( n95543 , C0 , n95511 , n95520 , n95541 , n95542 );
buf ( n95544 , n95543 );
buf ( n95545 , n95544 );
buf ( n95546 , n31655 );
buf ( n95547 , n30987 );
buf ( n95548 , n30987 );
xor ( n95549 , n49521 , n87870 );
and ( n95550 , n95549 , n32433 );
not ( n95551 , n47331 );
and ( n95552 , n95551 , n49521 );
and ( n95553 , n60382 , n60548 );
xor ( n95554 , n88673 , n95553 );
and ( n95555 , n95554 , n47331 );
or ( n95556 , n95552 , n95555 );
and ( n95557 , n95556 , n32413 );
and ( n95558 , n49521 , n47402 );
or ( n95559 , n95550 , n95557 , n95558 );
and ( n95560 , n95559 , n32456 );
and ( n95561 , n49521 , n47409 );
or ( n95562 , C0 , n95560 , n95561 );
buf ( n95563 , n95562 );
buf ( n95564 , n95563 );
buf ( n95565 , n31655 );
buf ( n95566 , n30987 );
not ( n95567 , n48765 );
and ( n95568 , n95567 , n33211 );
and ( n95569 , n84806 , n48765 );
or ( n95570 , n95568 , n95569 );
and ( n95571 , n95570 , n33180 );
not ( n95572 , n49054 );
and ( n95573 , n95572 , n33211 );
and ( n95574 , n84821 , n49054 );
or ( n95575 , n95573 , n95574 );
and ( n95576 , n95575 , n33178 );
and ( n95577 , n33211 , n49774 );
or ( n95578 , n95571 , n95576 , n95577 );
and ( n95579 , n95578 , n33208 );
and ( n95580 , n33270 , n33375 );
not ( n95581 , n32968 );
and ( n95582 , n95581 , n33270 );
and ( n95583 , n32510 , n81366 );
xor ( n95584 , n33211 , n95583 );
and ( n95585 , n95584 , n32968 );
or ( n95586 , n95582 , n95585 );
and ( n95587 , n95586 , n33370 );
and ( n95588 , n35592 , n35056 );
and ( n95589 , n33211 , n49794 );
or ( n95590 , C0 , n95579 , n95580 , n95587 , n95588 , n95589 );
buf ( n95591 , n95590 );
buf ( n95592 , n95591 );
buf ( n95593 , n31655 );
not ( n95594 , n35542 );
and ( n95595 , n95594 , n41853 );
and ( n95596 , n92695 , n35542 );
or ( n95597 , n95595 , n95596 );
buf ( n95598 , n95597 );
buf ( n95599 , n95598 );
buf ( n95600 , n30987 );
buf ( n95601 , n31655 );
and ( n95602 , n32458 , n32500 );
not ( n95603 , n35211 );
and ( n95604 , n95603 , n35677 );
buf ( n95605 , n95604 );
and ( n95606 , n95605 , n32421 );
not ( n95607 , n35245 );
and ( n95608 , n95607 , n35677 );
buf ( n95609 , n95608 );
and ( n95610 , n95609 , n32419 );
not ( n95611 , n35278 );
and ( n95612 , n95611 , n35677 );
not ( n95613 , n35295 );
and ( n95614 , n95613 , n47286 );
xor ( n95615 , n35677 , n49527 );
and ( n95616 , n95615 , n35295 );
or ( n95617 , n95614 , n95616 );
and ( n95618 , n95617 , n35278 );
or ( n95619 , n95612 , n95618 );
and ( n95620 , n95619 , n32417 );
not ( n95621 , n35331 );
and ( n95622 , n95621 , n35677 );
not ( n95623 , n35294 );
not ( n95624 , n45995 );
and ( n95625 , n95624 , n47286 );
xor ( n95626 , n49604 , n49613 );
and ( n95627 , n95626 , n45995 );
or ( n95628 , n95625 , n95627 );
and ( n95629 , n95623 , n95628 );
and ( n95630 , n95615 , n35294 );
or ( n95631 , n95629 , n95630 );
and ( n95632 , n95631 , n35331 );
or ( n95633 , n95622 , n95632 );
and ( n95634 , n95633 , n32415 );
and ( n95635 , n35677 , n35354 );
or ( n95636 , n95606 , n95610 , n95620 , n95634 , n95635 );
and ( n95637 , n95636 , n32456 );
not ( n95638 , n32475 );
not ( n95639 , n46060 );
and ( n95640 , n95639 , n35669 );
xor ( n95641 , n49695 , n49707 );
and ( n95642 , n95641 , n46060 );
or ( n95643 , n95640 , n95642 );
and ( n95644 , n95638 , n95643 );
and ( n95645 , n35677 , n32475 );
or ( n95646 , n95644 , n95645 );
and ( n95647 , n95646 , n32486 );
buf ( n95648 , n32489 );
and ( n95649 , n35677 , n35367 );
or ( n95650 , C0 , n95602 , n95637 , n95647 , n95648 , n95649 );
buf ( n95651 , n95650 );
buf ( n95652 , n95651 );
buf ( n95653 , n30987 );
buf ( n95654 , n30987 );
not ( n95655 , n34150 );
and ( n95656 , n95655 , n32761 );
not ( n95657 , n60126 );
and ( n95658 , n95657 , n32761 );
and ( n95659 , n32789 , n60126 );
or ( n95660 , n95658 , n95659 );
and ( n95661 , n95660 , n34150 );
or ( n95662 , n95656 , n95661 );
and ( n95663 , n95662 , n33381 );
not ( n95664 , n60134 );
not ( n95665 , n60126 );
and ( n95666 , n95665 , n32761 );
and ( n95667 , n34301 , n60126 );
or ( n95668 , n95666 , n95667 );
and ( n95669 , n95664 , n95668 );
and ( n95670 , n34301 , n60134 );
or ( n95671 , n95669 , n95670 );
and ( n95672 , n95671 , n33375 );
not ( n95673 , n32968 );
not ( n95674 , n60134 );
not ( n95675 , n60126 );
and ( n95676 , n95675 , n32761 );
and ( n95677 , n34301 , n60126 );
or ( n95678 , n95676 , n95677 );
and ( n95679 , n95674 , n95678 );
and ( n95680 , n34301 , n60134 );
or ( n95681 , n95679 , n95680 );
and ( n95682 , n95673 , n95681 );
not ( n95683 , n60154 );
not ( n95684 , n60156 );
and ( n95685 , n95684 , n95681 );
and ( n95686 , n34761 , n60156 );
or ( n95687 , n95685 , n95686 );
and ( n95688 , n95683 , n95687 );
and ( n95689 , n35050 , n60154 );
or ( n95690 , n95688 , n95689 );
and ( n95691 , n95690 , n32968 );
or ( n95692 , n95682 , n95691 );
and ( n95693 , n95692 , n33370 );
and ( n95694 , n32761 , n35062 );
or ( n95695 , C0 , n95663 , n95672 , n95693 , n95694 );
buf ( n95696 , n95695 );
buf ( n95697 , n95696 );
buf ( n95698 , n31655 );
buf ( n95699 , n31655 );
not ( n95700 , n31655 );
and ( n95701 , n33764 , n48455 );
not ( n95702 , n48457 );
and ( n95703 , n95702 , n33429 );
and ( n95704 , n33764 , n48457 );
or ( n95705 , n95703 , n95704 );
and ( n95706 , n95705 , n31373 );
not ( n95707 , n44807 );
and ( n95708 , n95707 , n33429 );
and ( n95709 , n33764 , n44807 );
or ( n95710 , n95708 , n95709 );
and ( n95711 , n95710 , n31408 );
not ( n95712 , n48468 );
and ( n95713 , n95712 , n33429 );
and ( n95714 , n33764 , n48468 );
or ( n95715 , n95713 , n95714 );
and ( n95716 , n95715 , n31468 );
not ( n95717 , n44817 );
and ( n95718 , n95717 , n33429 );
and ( n95719 , n33764 , n44817 );
or ( n95720 , n95718 , n95719 );
and ( n95721 , n95720 , n31521 );
not ( n95722 , n39979 );
and ( n95723 , n95722 , n33429 );
and ( n95724 , n33471 , n39979 );
or ( n95725 , n95723 , n95724 );
and ( n95726 , n95725 , n31538 );
not ( n95727 , n45059 );
and ( n95728 , n95727 , n33429 );
and ( n95729 , n33471 , n45059 );
or ( n95730 , n95728 , n95729 );
and ( n95731 , n95730 , n31536 );
not ( n95732 , n33419 );
and ( n95733 , n95732 , n33429 );
and ( n95734 , n75416 , n33419 );
or ( n95735 , n95733 , n95734 );
and ( n95736 , n95735 , n31529 );
not ( n95737 , n33734 );
and ( n95738 , n95737 , n33429 );
and ( n95739 , n75427 , n33734 );
or ( n95740 , n95738 , n95739 );
and ( n95741 , n95740 , n31527 );
and ( n95742 , n33849 , n48513 );
or ( n95743 , n95701 , n95706 , n95711 , n95716 , n95721 , n95726 , n95731 , n95736 , n95741 , n95742 );
and ( n95744 , n95743 , n31557 );
and ( n95745 , n34001 , n33973 );
and ( n95746 , n33429 , n48524 );
or ( n95747 , C0 , n95744 , n95745 , n95746 );
buf ( n95748 , n95747 );
buf ( n95749 , n95748 );
buf ( n95750 , n30987 );
or ( n95751 , n39350 , n39352 );
or ( n95752 , n95751 , n39354 );
buf ( n95753 , n95752 );
or ( n95754 , n39349 , n39356 );
or ( n95755 , n95754 , n39358 );
and ( n95756 , n50814 , n95755 );
or ( n95757 , C0 , n95753 , n95756 );
buf ( n95758 , n95757 );
buf ( n95759 , n95758 );
buf ( n95760 , n31655 );
and ( n95761 , n81697 , n31645 );
not ( n95762 , n45274 );
and ( n95763 , n95762 , n56397 );
buf ( n95764 , n95763 );
and ( n95765 , n95764 , n31373 );
not ( n95766 , n45280 );
and ( n95767 , n95766 , n56397 );
and ( n95768 , n81703 , n45280 );
or ( n95769 , n95767 , n95768 );
and ( n95770 , n95769 , n31468 );
and ( n95771 , n56397 , n45802 );
or ( n95772 , n95765 , n95770 , n95771 );
and ( n95773 , n95772 , n31557 );
and ( n95774 , n56397 , n45808 );
or ( n95775 , C0 , n95761 , n95773 , n95774 );
buf ( n95776 , n95775 );
buf ( n95777 , n95776 );
not ( n95778 , n40163 );
and ( n95779 , n95778 , n31790 );
not ( n95780 , n45227 );
and ( n95781 , n95780 , n31790 );
and ( n95782 , n32252 , n45227 );
or ( n95783 , n95781 , n95782 );
and ( n95784 , n95783 , n40163 );
or ( n95785 , n95779 , n95784 );
and ( n95786 , n95785 , n32498 );
not ( n95787 , n45235 );
not ( n95788 , n45227 );
and ( n95789 , n95788 , n31790 );
and ( n95790 , n40393 , n45227 );
or ( n95791 , n95789 , n95790 );
and ( n95792 , n95787 , n95791 );
and ( n95793 , n40393 , n45235 );
or ( n95794 , n95792 , n95793 );
and ( n95795 , n95794 , n32473 );
not ( n95796 , n32475 );
not ( n95797 , n45235 );
not ( n95798 , n45227 );
and ( n95799 , n95798 , n31790 );
and ( n95800 , n40393 , n45227 );
or ( n95801 , n95799 , n95800 );
and ( n95802 , n95797 , n95801 );
and ( n95803 , n40393 , n45235 );
or ( n95804 , n95802 , n95803 );
and ( n95805 , n95796 , n95804 );
not ( n95806 , n45255 );
not ( n95807 , n45257 );
and ( n95808 , n95807 , n95804 );
and ( n95809 , n40972 , n45257 );
or ( n95810 , n95808 , n95809 );
and ( n95811 , n95806 , n95810 );
and ( n95812 , n41267 , n45255 );
or ( n95813 , n95811 , n95812 );
and ( n95814 , n95813 , n32475 );
or ( n95815 , n95805 , n95814 );
and ( n95816 , n95815 , n32486 );
and ( n95817 , n31790 , n41278 );
or ( n95818 , C0 , n95786 , n95795 , n95816 , n95817 );
buf ( n95819 , n95818 );
buf ( n95820 , n95819 );
buf ( n95821 , n30987 );
buf ( n95822 , n30987 );
buf ( n95823 , n30987 );
and ( n95824 , n49061 , n48639 );
not ( n95825 , n48642 );
and ( n95826 , n95825 , n48586 );
and ( n95827 , n49061 , n48642 );
or ( n95828 , n95826 , n95827 );
and ( n95829 , n95828 , n32890 );
not ( n95830 , n48648 );
and ( n95831 , n95830 , n48586 );
and ( n95832 , n49061 , n48648 );
or ( n95833 , n95831 , n95832 );
and ( n95834 , n95833 , n32924 );
not ( n95835 , n48654 );
and ( n95836 , n95835 , n48586 );
and ( n95837 , n49061 , n48654 );
or ( n95838 , n95836 , n95837 );
and ( n95839 , n95838 , n33038 );
not ( n95840 , n48660 );
and ( n95841 , n95840 , n48586 );
and ( n95842 , n49061 , n48660 );
or ( n95843 , n95841 , n95842 );
and ( n95844 , n95843 , n33172 );
not ( n95845 , n41576 );
and ( n95846 , n95845 , n48586 );
nand ( n95847 , n48771 , n41576 );
nor ( n95848 , n95846 , n95847 );
and ( n95849 , n95848 , n33189 );
not ( n95850 , n48730 );
and ( n95851 , n95850 , n48586 );
and ( n95852 , n48771 , n48730 );
or ( n95853 , n95851 , n95852 );
and ( n95854 , n95853 , n33187 );
not ( n95855 , n48765 );
and ( n95856 , n95855 , n48586 );
and ( n95857 , n59676 , n48765 );
or ( n95858 , n95856 , n95857 );
and ( n95859 , n95858 , n33180 );
not ( n95860 , n49054 );
and ( n95861 , n95860 , n48586 );
and ( n95862 , n59687 , n49054 );
or ( n95863 , n95861 , n95862 );
and ( n95864 , n95863 , n33178 );
and ( n95865 , n49170 , n49275 );
or ( n95866 , n95824 , n95829 , n95834 , n95839 , n95844 , n95849 , n95854 , n95859 , n95864 , n95865 );
and ( n95867 , n95866 , n33208 );
and ( n95868 , n32979 , n35056 );
and ( n95869 , n48586 , n49286 );
or ( n95870 , C0 , n95867 , n95868 , n95869 );
buf ( n95871 , n95870 );
buf ( n95872 , n95871 );
buf ( n95873 , n30987 );
buf ( n95874 , n31655 );
buf ( n95875 , n31655 );
buf ( n95876 , n31655 );
xor ( n95877 , n44769 , n44798 );
and ( n95878 , n95877 , n31548 );
not ( n95879 , n44807 );
and ( n95880 , n95879 , n44769 );
and ( n95881 , n46642 , n44807 );
or ( n95882 , n95880 , n95881 );
and ( n95883 , n95882 , n31408 );
not ( n95884 , n44817 );
and ( n95885 , n95884 , n44769 );
and ( n95886 , n81713 , n44817 );
or ( n95887 , n95885 , n95886 );
and ( n95888 , n95887 , n31521 );
not ( n95889 , n45059 );
and ( n95890 , n95889 , n44769 );
xor ( n95891 , n40069 , n40127 );
and ( n95892 , n95891 , n45059 );
or ( n95893 , n95890 , n95892 );
and ( n95894 , n95893 , n31536 );
and ( n95895 , n44769 , n45148 );
or ( n95896 , n95878 , n95883 , n95888 , n95894 , n95895 );
and ( n95897 , n95896 , n31557 );
and ( n95898 , n44769 , n40154 );
or ( n95899 , C0 , n95897 , n95898 );
buf ( n95900 , n95899 );
buf ( n95901 , n95900 );
not ( n95902 , n40163 );
and ( n95903 , n95902 , n32021 );
not ( n95904 , n55888 );
and ( n95905 , n95904 , n32021 );
and ( n95906 , n32147 , n55888 );
or ( n95907 , n95905 , n95906 );
and ( n95908 , n95907 , n40163 );
or ( n95909 , n95903 , n95908 );
and ( n95910 , n95909 , n32498 );
not ( n95911 , n55896 );
not ( n95912 , n55888 );
and ( n95913 , n95912 , n32021 );
and ( n95914 , n49314 , n55888 );
or ( n95915 , n95913 , n95914 );
and ( n95916 , n95911 , n95915 );
and ( n95917 , n49314 , n55896 );
or ( n95918 , n95916 , n95917 );
and ( n95919 , n95918 , n32473 );
not ( n95920 , n32475 );
not ( n95921 , n55896 );
not ( n95922 , n55888 );
and ( n95923 , n95922 , n32021 );
and ( n95924 , n49314 , n55888 );
or ( n95925 , n95923 , n95924 );
and ( n95926 , n95921 , n95925 );
and ( n95927 , n49314 , n55896 );
or ( n95928 , n95926 , n95927 );
and ( n95929 , n95920 , n95928 );
not ( n95930 , n55916 );
not ( n95931 , n55918 );
and ( n95932 , n95931 , n95928 );
and ( n95933 , n49340 , n55918 );
or ( n95934 , n95932 , n95933 );
and ( n95935 , n95930 , n95934 );
and ( n95936 , n49348 , n55916 );
or ( n95937 , n95935 , n95936 );
and ( n95938 , n95937 , n32475 );
or ( n95939 , n95929 , n95938 );
and ( n95940 , n95939 , n32486 );
and ( n95941 , n32021 , n41278 );
or ( n95942 , C1 , n95910 , n95919 , n95940 , n95941 );
buf ( n95943 , n95942 );
buf ( n95944 , n95943 );
buf ( n95945 , n30987 );
buf ( n95946 , n30987 );
not ( n95947 , n48765 );
and ( n95948 , n95947 , n33213 );
and ( n95949 , n63532 , n48765 );
or ( n95950 , n95948 , n95949 );
and ( n95951 , n95950 , n33180 );
not ( n95952 , n49054 );
and ( n95953 , n95952 , n33213 );
and ( n95954 , n63543 , n49054 );
or ( n95955 , n95953 , n95954 );
and ( n95956 , n95955 , n33178 );
and ( n95957 , n33213 , n49774 );
or ( n95958 , n95951 , n95956 , n95957 );
and ( n95959 , n95958 , n33208 );
and ( n95960 , n33277 , n33375 );
not ( n95961 , n32968 );
and ( n95962 , n95961 , n33277 );
xor ( n95963 , n33213 , n66022 );
and ( n95964 , n95963 , n32968 );
or ( n95965 , n95962 , n95964 );
and ( n95966 , n95965 , n33370 );
and ( n95967 , n32976 , n35056 );
and ( n95968 , n33213 , n49794 );
or ( n95969 , C0 , n95959 , n95960 , n95966 , n95967 , n95968 );
buf ( n95970 , n95969 );
buf ( n95971 , n95970 );
buf ( n95972 , n30987 );
not ( n95973 , n35542 );
and ( n95974 , n95973 , n41865 );
and ( n95975 , n83173 , n35542 );
or ( n95976 , n95974 , n95975 );
buf ( n95977 , n95976 );
buf ( n95978 , n95977 );
buf ( n95979 , n31655 );
buf ( n95980 , n30987 );
buf ( n95981 , n31655 );
and ( n95982 , n46037 , n32500 );
not ( n95983 , n35211 );
and ( n95984 , n95983 , n37571 );
buf ( n95985 , n95984 );
and ( n95986 , n95985 , n32421 );
not ( n95987 , n35245 );
and ( n95988 , n95987 , n37571 );
buf ( n95989 , n95988 );
and ( n95990 , n95989 , n32419 );
not ( n95991 , n35278 );
and ( n95992 , n95991 , n37571 );
not ( n95993 , n35295 );
and ( n95994 , n95993 , n47283 );
xor ( n95995 , n37571 , n49530 );
and ( n95996 , n95995 , n35295 );
or ( n95997 , n95994 , n95996 );
and ( n95998 , n95997 , n35278 );
or ( n95999 , n95992 , n95998 );
and ( n96000 , n95999 , n32417 );
not ( n96001 , n35331 );
and ( n96002 , n96001 , n37571 );
not ( n96003 , n35294 );
not ( n96004 , n45995 );
and ( n96005 , n96004 , n47283 );
xor ( n96006 , n49601 , n49616 );
and ( n96007 , n96006 , n45995 );
or ( n96008 , n96005 , n96007 );
and ( n96009 , n96003 , n96008 );
and ( n96010 , n95995 , n35294 );
or ( n96011 , n96009 , n96010 );
and ( n96012 , n96011 , n35331 );
or ( n96013 , n96002 , n96012 );
and ( n96014 , n96013 , n32415 );
and ( n96015 , n37571 , n35354 );
or ( n96016 , n95986 , n95990 , n96000 , n96014 , n96015 );
and ( n96017 , n96016 , n32456 );
not ( n96018 , n32475 );
not ( n96019 , n46060 );
and ( n96020 , n96019 , n49691 );
xor ( n96021 , n49692 , n49710 );
and ( n96022 , n96021 , n46060 );
or ( n96023 , n96020 , n96022 );
and ( n96024 , n96018 , n96023 );
and ( n96025 , n37571 , n32475 );
or ( n96026 , n96024 , n96025 );
and ( n96027 , n96026 , n32486 );
buf ( n96028 , n32489 );
and ( n96029 , n37571 , n35367 );
or ( n96030 , C0 , n95982 , n96017 , n96027 , n96028 , n96029 );
buf ( n96031 , n96030 );
buf ( n96032 , n96031 );
buf ( n96033 , n31655 );
buf ( n96034 , n40206 );
xor ( n96035 , n35423 , n62857 );
and ( n96036 , n96035 , n31550 );
not ( n96037 , n39979 );
and ( n96038 , n96037 , n35423 );
and ( n96039 , n45078 , n86357 );
xor ( n96040 , n80909 , n96039 );
and ( n96041 , n96040 , n39979 );
or ( n96042 , n96038 , n96041 );
and ( n96043 , n96042 , n31538 );
and ( n96044 , n35423 , n40143 );
or ( n96045 , n96036 , n96043 , n96044 );
and ( n96046 , n96045 , n31557 );
and ( n96047 , n35423 , n40154 );
or ( n96048 , C0 , n96046 , n96047 );
buf ( n96049 , n96048 );
buf ( n96050 , n96049 );
not ( n96051 , n40163 );
and ( n96052 , n96051 , n31996 );
not ( n96053 , n40166 );
and ( n96054 , n96053 , n31996 );
and ( n96055 , n32165 , n40166 );
or ( n96056 , n96054 , n96055 );
and ( n96057 , n96056 , n40163 );
or ( n96058 , n96052 , n96057 );
and ( n96059 , n96058 , n32498 );
not ( n96060 , n40195 );
not ( n96061 , n40166 );
and ( n96062 , n96061 , n31996 );
and ( n96063 , n59005 , n40166 );
or ( n96064 , n96062 , n96063 );
and ( n96065 , n96060 , n96064 );
and ( n96066 , n59005 , n40195 );
or ( n96067 , n96065 , n96066 );
and ( n96068 , n96067 , n32473 );
not ( n96069 , n32475 );
not ( n96070 , n40195 );
not ( n96071 , n40166 );
and ( n96072 , n96071 , n31996 );
and ( n96073 , n59005 , n40166 );
or ( n96074 , n96072 , n96073 );
and ( n96075 , n96070 , n96074 );
and ( n96076 , n59005 , n40195 );
or ( n96077 , n96075 , n96076 );
and ( n96078 , n96069 , n96077 );
not ( n96079 , n40446 );
not ( n96080 , n40448 );
and ( n96081 , n96080 , n96077 );
and ( n96082 , n59029 , n40448 );
or ( n96083 , n96081 , n96082 );
and ( n96084 , n96079 , n96083 );
and ( n96085 , n59037 , n40446 );
or ( n96086 , n96084 , n96085 );
and ( n96087 , n96086 , n32475 );
or ( n96088 , n96078 , n96087 );
and ( n96089 , n96088 , n32486 );
and ( n96090 , n31996 , n41278 );
or ( n96091 , C0 , n96059 , n96068 , n96089 , n96090 );
buf ( n96092 , n96091 );
buf ( n96093 , n96092 );
buf ( n96094 , n30987 );
buf ( n96095 , n30987 );
not ( n96096 , n46356 );
and ( n96097 , n96096 , n31268 );
not ( n96098 , n61975 );
and ( n96099 , n96098 , n31268 );
and ( n96100 , n31272 , n61975 );
or ( n96101 , n96099 , n96100 );
and ( n96102 , n96101 , n46356 );
or ( n96103 , n96097 , n96102 );
and ( n96104 , n96103 , n31649 );
not ( n96105 , n61983 );
not ( n96106 , n61975 );
and ( n96107 , n96106 , n31268 );
and ( n96108 , n49443 , n61975 );
or ( n96109 , n96107 , n96108 );
and ( n96110 , n96105 , n96109 );
and ( n96111 , n49443 , n61983 );
or ( n96112 , n96110 , n96111 );
and ( n96113 , n96112 , n31643 );
not ( n96114 , n31452 );
not ( n96115 , n61983 );
not ( n96116 , n61975 );
and ( n96117 , n96116 , n31268 );
and ( n96118 , n49443 , n61975 );
or ( n96119 , n96117 , n96118 );
and ( n96120 , n96115 , n96119 );
and ( n96121 , n49443 , n61983 );
or ( n96122 , n96120 , n96121 );
and ( n96123 , n96114 , n96122 );
not ( n96124 , n62003 );
not ( n96125 , n62005 );
and ( n96126 , n96125 , n96122 );
and ( n96127 , n49469 , n62005 );
or ( n96128 , n96126 , n96127 );
and ( n96129 , n96124 , n96128 );
and ( n96130 , n49477 , n62003 );
or ( n96131 , n96129 , n96130 );
and ( n96132 , n96131 , n31452 );
or ( n96133 , n96123 , n96132 );
and ( n96134 , n96133 , n31638 );
and ( n96135 , n31268 , n47277 );
or ( n96136 , n96104 , n96113 , n96134 , n96135 );
buf ( n96137 , n96136 );
buf ( n96138 , n96137 );
buf ( n96139 , n31655 );
buf ( n96140 , n30987 );
buf ( n96141 , n30987 );
xor ( n96142 , n49581 , n60315 );
and ( n96143 , n96142 , n32433 );
not ( n96144 , n47331 );
and ( n96145 , n96144 , n49581 );
and ( n96146 , n68962 , n47331 );
or ( n96147 , n96145 , n96146 );
and ( n96148 , n96147 , n32413 );
and ( n96149 , n49581 , n47402 );
or ( n96150 , n96143 , n96148 , n96149 );
and ( n96151 , n96150 , n32456 );
and ( n96152 , n49581 , n47409 );
or ( n96153 , n96151 , n96152 );
buf ( n96154 , n96153 );
buf ( n96155 , n96154 );
buf ( n96156 , n31655 );
buf ( n96157 , n31655 );
not ( n96158 , n31437 );
and ( n96159 , n96158 , n59975 );
and ( n96160 , n59988 , n31437 );
or ( n96161 , n96159 , n96160 );
and ( n96162 , n96161 , n31468 );
not ( n96163 , n44817 );
and ( n96164 , n96163 , n59975 );
and ( n96165 , n93970 , n44817 );
or ( n96166 , n96164 , n96165 );
and ( n96167 , n96166 , n31521 );
and ( n96168 , n59975 , n42158 );
or ( n96169 , n96162 , n96167 , n96168 );
and ( n96170 , n96169 , n31557 );
and ( n96171 , n59975 , n40154 );
nor ( n96172 , n96170 , n96171 );
not ( n96173 , n96172 );
buf ( n96174 , n96173 );
and ( n96175 , n32304 , n50275 );
not ( n96176 , n50278 );
and ( n96177 , n96176 , n31738 );
and ( n96178 , n32304 , n50278 );
or ( n96179 , n96177 , n96178 );
and ( n96180 , n96179 , n32421 );
not ( n96181 , n50002 );
and ( n96182 , n96181 , n31738 );
and ( n96183 , n32304 , n50002 );
or ( n96184 , n96182 , n96183 );
and ( n96185 , n96184 , n32419 );
not ( n96186 , n50289 );
and ( n96187 , n96186 , n31738 );
and ( n96188 , n32304 , n50289 );
or ( n96189 , n96187 , n96188 );
and ( n96190 , n96189 , n32417 );
not ( n96191 , n50008 );
and ( n96192 , n96191 , n31738 );
and ( n96193 , n32304 , n50008 );
or ( n96194 , n96192 , n96193 );
and ( n96195 , n96194 , n32415 );
not ( n96196 , n47331 );
and ( n96197 , n96196 , n31738 );
and ( n96198 , n31965 , n47331 );
or ( n96199 , n96197 , n96198 );
and ( n96200 , n96199 , n32413 );
not ( n96201 , n50067 );
and ( n96202 , n96201 , n31738 );
and ( n96203 , n31965 , n50067 );
or ( n96204 , n96202 , n96203 );
and ( n96205 , n96204 , n32411 );
not ( n96206 , n31728 );
and ( n96207 , n96206 , n31738 );
and ( n96208 , n68458 , n31728 );
or ( n96209 , n96207 , n96208 );
and ( n96210 , n96209 , n32253 );
not ( n96211 , n32283 );
and ( n96212 , n96211 , n31738 );
and ( n96213 , n68471 , n32283 );
or ( n96214 , n96212 , n96213 );
and ( n96215 , n96214 , n32398 );
and ( n96216 , n32360 , n50334 );
or ( n96217 , n96175 , n96180 , n96185 , n96190 , n96195 , n96200 , n96205 , n96210 , n96215 , n96216 );
and ( n96218 , n96217 , n32456 );
and ( n96219 , n37585 , n32489 );
and ( n96220 , n31738 , n50345 );
or ( n96221 , n96218 , n96219 , n96220 );
buf ( n96222 , n96221 );
buf ( n96223 , n96222 );
buf ( n96224 , n30987 );
buf ( n96225 , n31655 );
buf ( n96226 , n31649 );
buf ( n96227 , n31647 );
not ( n96228 , n63845 );
not ( n96229 , n63847 );
and ( n96230 , n96229 , n30992 );
buf ( n96231 , n96230 );
and ( n96232 , n96231 , n31468 );
and ( n96233 , n30992 , n63859 );
or ( n96234 , n96232 , n96233 );
and ( n96235 , n96228 , n96234 );
buf ( n96236 , n96235 );
and ( n96237 , n96236 , n31557 );
or ( n96238 , n96226 , n96227 , n96237 );
buf ( n96239 , n96238 );
buf ( n96240 , n96239 );
buf ( n96241 , n30987 );
not ( n96242 , n38443 );
and ( n96243 , n96242 , n38048 );
xor ( n96244 , n53479 , n53490 );
and ( n96245 , n96244 , n38443 );
or ( n96246 , n96243 , n96245 );
and ( n96247 , n96246 , n38450 );
not ( n96248 , n39339 );
and ( n96249 , n96248 , n38948 );
xor ( n96250 , n53535 , n53546 );
and ( n96251 , n96250 , n39339 );
or ( n96252 , n96249 , n96251 );
and ( n96253 , n96252 , n39346 );
and ( n96254 , n40205 , n39359 );
or ( n96255 , n96247 , n96253 , n96254 );
buf ( n96256 , n96255 );
buf ( n96257 , n96256 );
not ( n96258 , n46356 );
and ( n96259 , n96258 , n31344 );
not ( n96260 , n55473 );
and ( n96261 , n96260 , n31344 );
and ( n96262 , n31372 , n55473 );
or ( n96263 , n96261 , n96262 );
and ( n96264 , n96263 , n46356 );
or ( n96265 , n96259 , n96264 );
and ( n96266 , n96265 , n31649 );
not ( n96267 , n55481 );
not ( n96268 , n55473 );
and ( n96269 , n96268 , n31344 );
and ( n96270 , n47849 , n55473 );
or ( n96271 , n96269 , n96270 );
and ( n96272 , n96267 , n96271 );
and ( n96273 , n47849 , n55481 );
or ( n96274 , n96272 , n96273 );
and ( n96275 , n96274 , n31643 );
not ( n96276 , n31452 );
not ( n96277 , n55481 );
not ( n96278 , n55473 );
and ( n96279 , n96278 , n31344 );
and ( n96280 , n47849 , n55473 );
or ( n96281 , n96279 , n96280 );
and ( n96282 , n96277 , n96281 );
and ( n96283 , n47849 , n55481 );
or ( n96284 , n96282 , n96283 );
and ( n96285 , n96276 , n96284 );
not ( n96286 , n55501 );
not ( n96287 , n55503 );
and ( n96288 , n96287 , n96284 );
and ( n96289 , n47877 , n55503 );
or ( n96290 , n96288 , n96289 );
and ( n96291 , n96286 , n96290 );
and ( n96292 , n47887 , n55501 );
or ( n96293 , n96291 , n96292 );
and ( n96294 , n96293 , n31452 );
or ( n96295 , n96285 , n96294 );
and ( n96296 , n96295 , n31638 );
and ( n96297 , n31344 , n47277 );
or ( n96298 , n96266 , n96275 , n96296 , n96297 );
buf ( n96299 , n96298 );
buf ( n96300 , n96299 );
buf ( n96301 , n31655 );
buf ( n96302 , n30987 );
not ( n96303 , n35278 );
and ( n96304 , n96303 , n88732 );
or ( n96305 , n88741 , n35278 );
or ( n96306 , n96304 , n96305 );
or ( n96307 , n96306 , n32417 );
not ( n96308 , n47912 );
and ( n96309 , n96308 , n88732 );
and ( n96310 , n91943 , n47912 );
or ( n96311 , n96309 , n96310 );
and ( n96312 , n96311 , n32415 );
and ( n96313 , n88732 , n48133 );
or ( n96314 , n96307 , n96312 , n96313 );
and ( n96315 , n96314 , n32456 );
and ( n96316 , n88732 , n47409 );
or ( n96317 , n96315 , n96316 );
buf ( n96318 , n96317 );
buf ( n96319 , n96318 );
buf ( n96320 , n31655 );
and ( n96321 , n49067 , n48639 );
not ( n96322 , n48642 );
and ( n96323 , n96322 , n48592 );
and ( n96324 , n49067 , n48642 );
or ( n96325 , n96323 , n96324 );
and ( n96326 , n96325 , n32890 );
not ( n96327 , n48648 );
and ( n96328 , n96327 , n48592 );
and ( n96329 , n49067 , n48648 );
or ( n96330 , n96328 , n96329 );
and ( n96331 , n96330 , n32924 );
not ( n96332 , n48654 );
and ( n96333 , n96332 , n48592 );
and ( n96334 , n49067 , n48654 );
or ( n96335 , n96333 , n96334 );
and ( n96336 , n96335 , n33038 );
not ( n96337 , n48660 );
and ( n96338 , n96337 , n48592 );
and ( n96339 , n49067 , n48660 );
or ( n96340 , n96338 , n96339 );
and ( n96341 , n96340 , n33172 );
not ( n96342 , n41576 );
and ( n96343 , n96342 , n48592 );
and ( n96344 , n48777 , n41576 );
or ( n96345 , n96343 , n96344 );
and ( n96346 , n96345 , n33189 );
not ( n96347 , n48730 );
and ( n96348 , n96347 , n48592 );
and ( n96349 , n48777 , n48730 );
or ( n96350 , n96348 , n96349 );
and ( n96351 , n96350 , n33187 );
not ( n96352 , n48765 );
and ( n96353 , n96352 , n48592 );
and ( n96354 , n53876 , n48765 );
or ( n96355 , n96353 , n96354 );
and ( n96356 , n96355 , n33180 );
not ( n96357 , n49054 );
and ( n96358 , n96357 , n48592 );
and ( n96359 , n53887 , n49054 );
or ( n96360 , n96358 , n96359 );
and ( n96361 , n96360 , n33178 );
and ( n96362 , n49176 , n49275 );
or ( n96363 , n96321 , n96326 , n96331 , n96336 , n96341 , n96346 , n96351 , n96356 , n96361 , n96362 );
and ( n96364 , n96363 , n33208 );
and ( n96365 , n32985 , n35056 );
and ( n96366 , n48592 , n49286 );
or ( n96367 , n96364 , n96365 , n96366 );
buf ( n96368 , n96367 );
buf ( n96369 , n96368 );
buf ( n96370 , n30987 );
buf ( n96371 , n30987 );
buf ( n96372 , n31655 );
buf ( n96373 , n31655 );
buf ( n96374 , n30987 );
buf ( n96375 , n31655 );
xor ( n96376 , n39493 , n54973 );
and ( n96377 , n96376 , n33199 );
not ( n96378 , n48648 );
and ( n96379 , n96378 , n39493 );
and ( n96380 , n34375 , n48648 );
or ( n96381 , n96379 , n96380 );
and ( n96382 , n96381 , n32924 );
not ( n96383 , n48660 );
and ( n96384 , n96383 , n39493 );
not ( n96385 , n39584 );
and ( n96386 , n96385 , n72102 );
and ( n96387 , n72118 , n39584 );
or ( n96388 , n96386 , n96387 );
and ( n96389 , n96388 , n48660 );
or ( n96390 , n96384 , n96389 );
and ( n96391 , n96390 , n33172 );
not ( n96392 , n48730 );
and ( n96393 , n96392 , n39493 );
and ( n96394 , n74257 , n48730 );
or ( n96395 , n96393 , n96394 );
and ( n96396 , n96395 , n33187 );
and ( n96397 , n39493 , n54713 );
or ( n96398 , n96377 , n96382 , n96391 , n96396 , n96397 );
and ( n96399 , n96398 , n33208 );
and ( n96400 , n39493 , n39805 );
or ( n96401 , n96399 , n96400 );
buf ( n96402 , n96401 );
buf ( n96403 , n96402 );
buf ( n96404 , n30987 );
buf ( n96405 , n31655 );
not ( n96406 , n41532 );
and ( n96407 , n96406 , n34421 );
and ( n96408 , n74228 , n41532 );
or ( n96409 , n96407 , n96408 );
buf ( n96410 , n96409 );
buf ( n96411 , n96410 );
not ( n96412 , n46356 );
and ( n96413 , n96412 , n31313 );
not ( n96414 , n46362 );
and ( n96415 , n96414 , n31313 );
and ( n96416 , n31339 , n46362 );
or ( n96417 , n96415 , n96416 );
and ( n96418 , n96417 , n46356 );
or ( n96419 , n96413 , n96418 );
and ( n96420 , n96419 , n31649 );
not ( n96421 , n46393 );
not ( n96422 , n46362 );
and ( n96423 , n96422 , n31313 );
and ( n96424 , n47449 , n46362 );
or ( n96425 , n96423 , n96424 );
and ( n96426 , n96421 , n96425 );
and ( n96427 , n47449 , n46393 );
or ( n96428 , n96426 , n96427 );
and ( n96429 , n96428 , n31643 );
not ( n96430 , n31452 );
not ( n96431 , n46393 );
not ( n96432 , n46362 );
and ( n96433 , n96432 , n31313 );
and ( n96434 , n47449 , n46362 );
or ( n96435 , n96433 , n96434 );
and ( n96436 , n96431 , n96435 );
and ( n96437 , n47449 , n46393 );
or ( n96438 , n96436 , n96437 );
and ( n96439 , n96430 , n96438 );
not ( n96440 , n46550 );
not ( n96441 , n46554 );
and ( n96442 , n96441 , n96438 );
and ( n96443 , n47485 , n46554 );
or ( n96444 , n96442 , n96443 );
and ( n96445 , n96440 , n96444 );
and ( n96446 , n47503 , n46550 );
or ( n96447 , n96445 , n96446 );
and ( n96448 , n96447 , n31452 );
or ( n96449 , n96439 , n96448 );
and ( n96450 , n96449 , n31638 );
and ( n96451 , n31313 , n47277 );
or ( n96452 , n96420 , n96429 , n96450 , n96451 );
buf ( n96453 , n96452 );
buf ( n96454 , n96453 );
buf ( n96455 , n31655 );
buf ( n96456 , n30987 );
and ( n96457 , n73740 , n32494 );
not ( n96458 , n46083 );
and ( n96459 , n96458 , n58618 );
and ( n96460 , n73746 , n46083 );
or ( n96461 , n96459 , n96460 );
and ( n96462 , n96461 , n32421 );
not ( n96463 , n46326 );
and ( n96464 , n96463 , n58618 );
and ( n96465 , n73746 , n46326 );
or ( n96466 , n96464 , n96465 );
and ( n96467 , n96466 , n32417 );
and ( n96468 , n58618 , n46340 );
or ( n96469 , n96462 , n96467 , n96468 );
and ( n96470 , n96469 , n32456 );
and ( n96471 , n58618 , n46349 );
or ( n96472 , n96457 , n96470 , n96471 );
buf ( n96473 , n96472 );
buf ( n96474 , n96473 );
buf ( n96475 , n31655 );
buf ( n96476 , n30987 );
not ( n96477 , n43755 );
and ( n96478 , n96477 , n43683 );
xor ( n96479 , n52302 , n52327 );
and ( n96480 , n96479 , n43755 );
or ( n96481 , n96478 , n96480 );
and ( n96482 , n96481 , n43774 );
not ( n96483 , n44663 );
and ( n96484 , n96483 , n44595 );
xor ( n96485 , n52340 , n52365 );
and ( n96486 , n96485 , n44663 );
or ( n96487 , n96484 , n96486 );
and ( n96488 , n96487 , n44682 );
and ( n96489 , n88909 , n44695 );
or ( n96490 , n96482 , n96488 , n96489 );
buf ( n96491 , n96490 );
buf ( n96492 , n96491 );
buf ( n96493 , n30987 );
buf ( n96494 , n31655 );
buf ( n96495 , n31655 );
buf ( n96496 , n31655 );
or ( n96497 , n33379 , n33381 );
or ( n96498 , n96497 , n32528 );
and ( n96499 , n68281 , n96498 );
not ( n96500 , n32967 );
and ( n96501 , n68281 , n96500 );
and ( n96502 , n96501 , n33377 );
not ( n96503 , n32598 );
and ( n96504 , n96503 , n68281 );
not ( n96505 , n32963 );
buf ( n96506 , n96505 );
and ( n96507 , n32966 , n32963 );
or ( n96508 , n96506 , n96507 );
and ( n96509 , n96508 , n32598 );
or ( n96510 , n96504 , n96509 );
and ( n96511 , n96510 , n32890 );
not ( n96512 , n32919 );
and ( n96513 , n96512 , n68281 );
and ( n96514 , n32966 , n32919 );
or ( n96515 , n96513 , n96514 );
and ( n96516 , n96515 , n32924 );
not ( n96517 , n32953 );
and ( n96518 , n96517 , n68281 );
not ( n96519 , n48641 );
buf ( n96520 , n96519 );
and ( n96521 , n32969 , n48641 );
or ( n96522 , n96520 , n96521 );
and ( n96523 , n96522 , n32953 );
or ( n96524 , n96518 , n96523 );
and ( n96525 , n96524 , n33038 );
not ( n96526 , n33067 );
and ( n96527 , n96526 , n68281 );
not ( n96528 , n32967 );
buf ( n96529 , n96528 );
not ( n96530 , n96529 );
and ( n96531 , n96530 , n33067 );
or ( n96532 , n96527 , n96531 );
and ( n96533 , n96532 , n33172 );
and ( n96534 , n68281 , n33204 );
nor ( n96535 , n96511 , n96516 , n96525 , n96533 , n96534 );
nand ( n96536 , n96535 , n33208 );
or ( n96537 , n58910 , n33373 );
buf ( n96538 , n96537 );
or ( n96539 , n96499 , n96502 , n96536 , n96538 );
buf ( n96540 , n96539 );
buf ( n96541 , n96540 );
buf ( n96542 , n30987 );
buf ( n96543 , n30987 );
buf ( n96544 , n31655 );
buf ( n96545 , n31655 );
xor ( n96546 , n44774 , n44793 );
and ( n96547 , n96546 , n31548 );
not ( n96548 , n44807 );
and ( n96549 , n96548 , n44774 );
and ( n96550 , n46667 , n44807 );
or ( n96551 , n96549 , n96550 );
and ( n96552 , n96551 , n31408 );
not ( n96553 , n44817 );
and ( n96554 , n96553 , n44774 );
and ( n96555 , n57106 , n44817 );
or ( n96556 , n96554 , n96555 );
and ( n96557 , n96556 , n31521 );
not ( n96558 , n45059 );
and ( n96559 , n96558 , n44774 );
and ( n96560 , n75970 , n45059 );
or ( n96561 , n96559 , n96560 );
and ( n96562 , n96561 , n31536 );
and ( n96563 , n44774 , n45148 );
or ( n96564 , n96547 , n96552 , n96557 , n96562 , n96563 );
and ( n96565 , n96564 , n31557 );
and ( n96566 , n44774 , n40154 );
or ( n96567 , n96565 , n96566 );
buf ( n96568 , n96567 );
buf ( n96569 , n96568 );
not ( n96570 , n40163 );
and ( n96571 , n96570 , n31846 );
not ( n96572 , n55888 );
and ( n96573 , n96572 , n31846 );
and ( n96574 , n32235 , n55888 );
or ( n96575 , n96573 , n96574 );
and ( n96576 , n96575 , n40163 );
or ( n96577 , n96571 , n96576 );
and ( n96578 , n96577 , n32498 );
not ( n96579 , n55896 );
not ( n96580 , n55888 );
and ( n96581 , n96580 , n31846 );
and ( n96582 , n42188 , n55888 );
or ( n96583 , n96581 , n96582 );
and ( n96584 , n96579 , n96583 );
and ( n96585 , n42188 , n55896 );
or ( n96586 , n96584 , n96585 );
and ( n96587 , n96586 , n32473 );
not ( n96588 , n32475 );
not ( n96589 , n55896 );
not ( n96590 , n55888 );
and ( n96591 , n96590 , n31846 );
and ( n96592 , n42188 , n55888 );
or ( n96593 , n96591 , n96592 );
and ( n96594 , n96589 , n96593 );
and ( n96595 , n42188 , n55896 );
or ( n96596 , n96594 , n96595 );
and ( n96597 , n96588 , n96596 );
not ( n96598 , n55916 );
not ( n96599 , n55918 );
and ( n96600 , n96599 , n96596 );
and ( n96601 , n42216 , n55918 );
or ( n96602 , n96600 , n96601 );
and ( n96603 , n96598 , n96602 );
and ( n96604 , n42224 , n55916 );
or ( n96605 , n96603 , n96604 );
and ( n96606 , n96605 , n32475 );
or ( n96607 , n96597 , n96606 );
and ( n96608 , n96607 , n32486 );
and ( n96609 , n31846 , n41278 );
or ( n96610 , n96578 , n96587 , n96608 , n96609 );
buf ( n96611 , n96610 );
buf ( n96612 , n96611 );
buf ( n96613 , n30987 );
buf ( n96614 , n30987 );
and ( n96615 , n33770 , n48455 );
not ( n96616 , n48457 );
and ( n96617 , n96616 , n33435 );
and ( n96618 , n33770 , n48457 );
or ( n96619 , n96617 , n96618 );
and ( n96620 , n96619 , n31373 );
not ( n96621 , n44807 );
and ( n96622 , n96621 , n33435 );
and ( n96623 , n33770 , n44807 );
or ( n96624 , n96622 , n96623 );
and ( n96625 , n96624 , n31408 );
not ( n96626 , n48468 );
and ( n96627 , n96626 , n33435 );
and ( n96628 , n33770 , n48468 );
or ( n96629 , n96627 , n96628 );
and ( n96630 , n96629 , n31468 );
not ( n96631 , n44817 );
and ( n96632 , n96631 , n33435 );
and ( n96633 , n33770 , n44817 );
or ( n96634 , n96632 , n96633 );
and ( n96635 , n96634 , n31521 );
not ( n96636 , n39979 );
and ( n96637 , n96636 , n33435 );
and ( n96638 , n33477 , n39979 );
or ( n96639 , n96637 , n96638 );
and ( n96640 , n96639 , n31538 );
not ( n96641 , n45059 );
and ( n96642 , n96641 , n33435 );
and ( n96643 , n33477 , n45059 );
or ( n96644 , n96642 , n96643 );
and ( n96645 , n96644 , n31536 );
not ( n96646 , n33419 );
and ( n96647 , n96646 , n33435 );
and ( n96648 , n72842 , n33419 );
or ( n96649 , n96647 , n96648 );
and ( n96650 , n96649 , n31529 );
not ( n96651 , n33734 );
and ( n96652 , n96651 , n33435 );
and ( n96653 , n72853 , n33734 );
or ( n96654 , n96652 , n96653 );
and ( n96655 , n96654 , n31527 );
and ( n96656 , n33855 , n48513 );
or ( n96657 , n96615 , n96620 , n96625 , n96630 , n96635 , n96640 , n96645 , n96650 , n96655 , n96656 );
and ( n96658 , n96657 , n31557 );
and ( n96659 , n34007 , n33973 );
and ( n96660 , n33435 , n48524 );
or ( n96661 , n96658 , n96659 , n96660 );
buf ( n96662 , n96661 );
buf ( n96663 , n96662 );
buf ( n96664 , n31655 );
buf ( n96665 , n30987 );
not ( n96666 , n35278 );
and ( n96667 , n96666 , n79205 );
and ( n96668 , n79218 , n35278 );
or ( n96669 , n96667 , n96668 );
and ( n96670 , n96669 , n32417 );
not ( n96671 , n50008 );
and ( n96672 , n96671 , n79205 );
and ( n96673 , n66674 , n50008 );
or ( n96674 , n96672 , n96673 );
and ( n96675 , n96674 , n32415 );
and ( n96676 , n79205 , n48133 );
or ( n96677 , n96670 , n96675 , n96676 );
and ( n96678 , n96677 , n32456 );
and ( n96679 , n79205 , n47409 );
or ( n96680 , n96678 , n96679 );
buf ( n96681 , n96680 );
buf ( n96682 , n96681 );
not ( n96683 , n48765 );
and ( n96684 , n96683 , n33223 );
and ( n96685 , n70890 , n48765 );
or ( n96686 , n96684 , n96685 );
and ( n96687 , n96686 , n33180 );
not ( n96688 , n49054 );
and ( n96689 , n96688 , n33223 );
and ( n96690 , n70901 , n49054 );
or ( n96691 , n96689 , n96690 );
and ( n96692 , n96691 , n33178 );
and ( n96693 , n33223 , n49774 );
or ( n96694 , n96687 , n96692 , n96693 );
and ( n96695 , n96694 , n33208 );
and ( n96696 , n33297 , n33375 );
not ( n96697 , n32968 );
and ( n96698 , n96697 , n33297 );
xor ( n96699 , n33223 , n53906 );
and ( n96700 , n96699 , n32968 );
or ( n96701 , n96698 , n96700 );
and ( n96702 , n96701 , n33370 );
and ( n96703 , n32986 , n35056 );
and ( n96704 , n33223 , n49794 );
or ( n96705 , n96695 , n96696 , n96702 , n96703 , n96704 );
buf ( n96706 , n96705 );
buf ( n96707 , n96706 );
buf ( n96708 , n30987 );
buf ( n96709 , n61736 );
buf ( n96710 , n31655 );
buf ( n96711 , n30987 );
buf ( n96712 , n31655 );
and ( n96713 , n46027 , n32500 );
not ( n96714 , n35211 );
and ( n96715 , n96714 , n37551 );
buf ( n96716 , n96715 );
and ( n96717 , n96716 , n32421 );
not ( n96718 , n35245 );
and ( n96719 , n96718 , n37551 );
buf ( n96720 , n96719 );
and ( n96721 , n96720 , n32419 );
not ( n96722 , n35278 );
and ( n96723 , n96722 , n37551 );
not ( n96724 , n35295 );
and ( n96725 , n96724 , n49581 );
xor ( n96726 , n37551 , n49540 );
and ( n96727 , n96726 , n35295 );
or ( n96728 , n96725 , n96727 );
and ( n96729 , n96728 , n35278 );
or ( n96730 , n96723 , n96729 );
and ( n96731 , n96730 , n32417 );
not ( n96732 , n35331 );
and ( n96733 , n96732 , n37551 );
not ( n96734 , n35294 );
not ( n96735 , n45995 );
and ( n96736 , n96735 , n49581 );
xor ( n96737 , n49582 , n49626 );
and ( n96738 , n96737 , n45995 );
or ( n96739 , n96736 , n96738 );
and ( n96740 , n96734 , n96739 );
and ( n96741 , n96726 , n35294 );
or ( n96742 , n96740 , n96741 );
and ( n96743 , n96742 , n35331 );
or ( n96744 , n96733 , n96743 );
and ( n96745 , n96744 , n32415 );
and ( n96746 , n37551 , n35354 );
or ( n96747 , n96717 , n96721 , n96731 , n96745 , n96746 );
and ( n96748 , n96747 , n32456 );
not ( n96749 , n32475 );
not ( n96750 , n46060 );
and ( n96751 , n96750 , n49671 );
xor ( n96752 , n49672 , n49720 );
and ( n96753 , n96752 , n46060 );
xor ( n96754 , n96751 , n96753 );
and ( n96755 , n96749 , n96754 );
and ( n96756 , n37551 , n32475 );
xor ( n96757 , n96755 , n96756 );
nand ( n96758 , n96757 , n32486 );
and ( n96759 , n37551 , n35367 );
nor ( n96760 , n96713 , n96748 , n96758 , n96759 );
buf ( n96761 , n96760 );
buf ( n96762 , n96761 );
buf ( n96763 , n31655 );
xor ( n96764 , n34058 , n39928 );
and ( n96765 , n96764 , n31550 );
not ( n96766 , n39979 );
and ( n96767 , n96766 , n34058 );
buf ( n96768 , n31337 );
and ( n96769 , n96768 , n39979 );
or ( n96770 , n96767 , n96769 );
and ( n96771 , n96770 , n31538 );
and ( n96772 , n34058 , n40143 );
or ( n96773 , n96765 , n96771 , n96772 );
and ( n96774 , n96773 , n31557 );
and ( n96775 , n34058 , n40154 );
or ( n96776 , n96774 , n96775 );
buf ( n96777 , n96776 );
buf ( n96778 , n96777 );
not ( n96779 , n40163 );
and ( n96780 , n96779 , n31990 );
not ( n96781 , n57233 );
and ( n96782 , n96781 , n31990 );
and ( n96783 , n32165 , n57233 );
or ( n96784 , n96782 , n96783 );
and ( n96785 , n96784 , n40163 );
or ( n96786 , n96780 , n96785 );
and ( n96787 , n96786 , n32498 );
not ( n96788 , n57241 );
not ( n96789 , n57233 );
and ( n96790 , n96789 , n31990 );
and ( n96791 , n59005 , n57233 );
or ( n96792 , n96790 , n96791 );
and ( n96793 , n96788 , n96792 );
and ( n96794 , n59005 , n57241 );
or ( n96795 , n96793 , n96794 );
and ( n96796 , n96795 , n32473 );
not ( n96797 , n32475 );
not ( n96798 , n57241 );
not ( n96799 , n57233 );
and ( n96800 , n96799 , n31990 );
and ( n96801 , n59005 , n57233 );
or ( n96802 , n96800 , n96801 );
and ( n96803 , n96798 , n96802 );
and ( n96804 , n59005 , n57241 );
or ( n96805 , n96803 , n96804 );
and ( n96806 , n96797 , n96805 );
not ( n96807 , n57261 );
not ( n96808 , n57263 );
and ( n96809 , n96808 , n96805 );
and ( n96810 , n59029 , n57263 );
or ( n96811 , n96809 , n96810 );
and ( n96812 , n96807 , n96811 );
and ( n96813 , n59037 , n57261 );
or ( n96814 , n96812 , n96813 );
and ( n96815 , n96814 , n32475 );
or ( n96816 , n96806 , n96815 );
and ( n96817 , n96816 , n32486 );
and ( n96818 , n31990 , n41278 );
or ( n96819 , n96787 , n96796 , n96817 , n96818 );
buf ( n96820 , n96819 );
buf ( n96821 , n96820 );
buf ( n96822 , n30987 );
buf ( n96823 , n30987 );
not ( n96824 , n34150 );
and ( n96825 , n96824 , n32857 );
not ( n96826 , n56708 );
and ( n96827 , n96826 , n32857 );
and ( n96828 , n32889 , n56708 );
or ( n96829 , n96827 , n96828 );
and ( n96830 , n96829 , n34150 );
or ( n96831 , n96825 , n96830 );
and ( n96832 , n96831 , n33381 );
not ( n96833 , n56716 );
not ( n96834 , n56708 );
and ( n96835 , n96834 , n32857 );
and ( n96836 , n52819 , n56708 );
or ( n96837 , n96835 , n96836 );
and ( n96838 , n96833 , n96837 );
and ( n96839 , n52819 , n56716 );
or ( n96840 , n96838 , n96839 );
and ( n96841 , n96840 , n33375 );
not ( n96842 , n32968 );
not ( n96843 , n56716 );
not ( n96844 , n56708 );
and ( n96845 , n96844 , n32857 );
and ( n96846 , n52819 , n56708 );
or ( n96847 , n96845 , n96846 );
and ( n96848 , n96843 , n96847 );
and ( n96849 , n52819 , n56716 );
or ( n96850 , n96848 , n96849 );
and ( n96851 , n96842 , n96850 );
not ( n96852 , n56736 );
not ( n96853 , n56738 );
and ( n96854 , n96853 , n96850 );
and ( n96855 , n52845 , n56738 );
or ( n96856 , n96854 , n96855 );
and ( n96857 , n96852 , n96856 );
and ( n96858 , n52855 , n56736 );
or ( n96859 , n96857 , n96858 );
and ( n96860 , n96859 , n32968 );
or ( n96861 , n96851 , n96860 );
and ( n96862 , n96861 , n33370 );
and ( n96863 , n32857 , n35062 );
or ( n96864 , n96832 , n96841 , n96862 , n96863 );
buf ( n96865 , n96864 );
buf ( n96866 , n96865 );
buf ( n96867 , n30987 );
buf ( n96868 , n30987 );
buf ( n96869 , n31655 );
buf ( n96870 , n31655 );
buf ( n96871 , n31655 );
and ( n96872 , n58634 , n31645 );
not ( n96873 , n45274 );
and ( n96874 , n96873 , n50837 );
and ( n96875 , n83745 , n45274 );
or ( n96876 , n96874 , n96875 );
and ( n96877 , n96876 , n31373 );
not ( n96878 , n45280 );
and ( n96879 , n96878 , n50837 );
and ( n96880 , n83745 , n45280 );
or ( n96881 , n96879 , n96880 );
and ( n96882 , n96881 , n31468 );
and ( n96883 , n50837 , n45802 );
or ( n96884 , n96877 , n96882 , n96883 );
and ( n96885 , n96884 , n31557 );
and ( n96886 , n50837 , n45808 );
or ( n96887 , n96872 , n96885 , n96886 );
buf ( n96888 , n96887 );
buf ( n96889 , n96888 );
not ( n96890 , n40163 );
and ( n96891 , n96890 , n31970 );
not ( n96892 , n56287 );
and ( n96893 , n96892 , n31970 );
and ( n96894 , n32165 , n56287 );
or ( n96895 , n96893 , n96894 );
and ( n96896 , n96895 , n40163 );
or ( n96897 , n96891 , n96896 );
and ( n96898 , n96897 , n32498 );
not ( n96899 , n56295 );
not ( n96900 , n56287 );
and ( n96901 , n96900 , n31970 );
and ( n96902 , n59005 , n56287 );
or ( n96903 , n96901 , n96902 );
and ( n96904 , n96899 , n96903 );
and ( n96905 , n59005 , n56295 );
or ( n96906 , n96904 , n96905 );
and ( n96907 , n96906 , n32473 );
not ( n96908 , n32475 );
not ( n96909 , n56295 );
not ( n96910 , n56287 );
and ( n96911 , n96910 , n31970 );
and ( n96912 , n59005 , n56287 );
or ( n96913 , n96911 , n96912 );
and ( n96914 , n96909 , n96913 );
and ( n96915 , n59005 , n56295 );
or ( n96916 , n96914 , n96915 );
and ( n96917 , n96908 , n96916 );
not ( n96918 , n56315 );
not ( n96919 , n56317 );
and ( n96920 , n96919 , n96916 );
and ( n96921 , n59029 , n56317 );
or ( n96922 , n96920 , n96921 );
and ( n96923 , n96918 , n96922 );
and ( n96924 , n59037 , n56315 );
or ( n96925 , n96923 , n96924 );
and ( n96926 , n96925 , n32475 );
or ( n96927 , n96917 , n96926 );
and ( n96928 , n96927 , n32486 );
and ( n96929 , n31970 , n41278 );
or ( n96930 , n96898 , n96907 , n96928 , n96929 );
buf ( n96931 , n96930 );
buf ( n96932 , n96931 );
buf ( n96933 , n30987 );
buf ( n96934 , n31655 );
and ( n96935 , n78686 , n31645 );
not ( n96936 , n45274 );
and ( n96937 , n96936 , n91188 );
buf ( n96938 , n96937 );
and ( n96939 , n96938 , n31373 );
not ( n96940 , n45280 );
and ( n96941 , n96940 , n91188 );
and ( n96942 , n78692 , n45280 );
or ( n96943 , n96941 , n96942 );
and ( n96944 , n96943 , n31468 );
and ( n96945 , n91188 , n45802 );
or ( n96946 , n96939 , n96944 , n96945 );
and ( n96947 , n96946 , n31557 );
and ( n96948 , n91188 , n45808 );
or ( n96949 , n96935 , n96947 , n96948 );
buf ( n96950 , n96949 );
buf ( n96951 , n96950 );
not ( n96952 , n40163 );
and ( n96953 , n96952 , n32009 );
not ( n96954 , n54629 );
and ( n96955 , n96954 , n32009 );
and ( n96956 , n32147 , n54629 );
or ( n96957 , n96955 , n96956 );
and ( n96958 , n96957 , n40163 );
or ( n96959 , n96953 , n96958 );
and ( n96960 , n96959 , n32498 );
not ( n96961 , n54637 );
not ( n96962 , n54629 );
and ( n96963 , n96962 , n32009 );
and ( n96964 , n49314 , n54629 );
or ( n96965 , n96963 , n96964 );
and ( n96966 , n96961 , n96965 );
and ( n96967 , n49314 , n54637 );
or ( n96968 , n96966 , n96967 );
and ( n96969 , n96968 , n32473 );
not ( n96970 , n32475 );
not ( n96971 , n54637 );
not ( n96972 , n54629 );
and ( n96973 , n96972 , n32009 );
and ( n96974 , n49314 , n54629 );
or ( n96975 , n96973 , n96974 );
and ( n96976 , n96971 , n96975 );
and ( n96977 , n49314 , n54637 );
or ( n96978 , n96976 , n96977 );
and ( n96979 , n96970 , n96978 );
not ( n96980 , n54657 );
not ( n96981 , n54659 );
and ( n96982 , n96981 , n96978 );
and ( n96983 , n49340 , n54659 );
or ( n96984 , n96982 , n96983 );
and ( n96985 , n96980 , n96984 );
and ( n96986 , n49348 , n54657 );
or ( n96987 , n96985 , n96986 );
and ( n96988 , n96987 , n32475 );
or ( n96989 , n96979 , n96988 );
and ( n96990 , n96989 , n32486 );
and ( n96991 , n32009 , n41278 );
or ( n96992 , n96960 , n96969 , n96990 , n96991 );
buf ( n96993 , n96992 );
buf ( n96994 , n96993 );
buf ( n96995 , n30987 );
and ( C0 , n31018 , n31019 );
and ( C1 , n31018 , n31019 );
endmodule

