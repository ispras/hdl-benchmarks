//NOTE: no-implementation module stub

module GTECH_MUX8 (
    input wire D0,
    input wire D1,
    input wire D2,
    input wire D3,
    input wire D4,
    input wire D5,
    input wire D6,
    input wire D7,
    input wire A,
    input wire B,
    input wire C,
    output wire Z
);

endmodule
