//NOTE: no-implementation module stub

module GtCLK_NAND3 (
    output Z,
    input A,
    input B,
    input C
);

endmodule
